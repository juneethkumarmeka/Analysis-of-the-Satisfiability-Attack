module basic_5000_50000_5000_10_levels_5xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,In_3000,In_3001,In_3002,In_3003,In_3004,In_3005,In_3006,In_3007,In_3008,In_3009,In_3010,In_3011,In_3012,In_3013,In_3014,In_3015,In_3016,In_3017,In_3018,In_3019,In_3020,In_3021,In_3022,In_3023,In_3024,In_3025,In_3026,In_3027,In_3028,In_3029,In_3030,In_3031,In_3032,In_3033,In_3034,In_3035,In_3036,In_3037,In_3038,In_3039,In_3040,In_3041,In_3042,In_3043,In_3044,In_3045,In_3046,In_3047,In_3048,In_3049,In_3050,In_3051,In_3052,In_3053,In_3054,In_3055,In_3056,In_3057,In_3058,In_3059,In_3060,In_3061,In_3062,In_3063,In_3064,In_3065,In_3066,In_3067,In_3068,In_3069,In_3070,In_3071,In_3072,In_3073,In_3074,In_3075,In_3076,In_3077,In_3078,In_3079,In_3080,In_3081,In_3082,In_3083,In_3084,In_3085,In_3086,In_3087,In_3088,In_3089,In_3090,In_3091,In_3092,In_3093,In_3094,In_3095,In_3096,In_3097,In_3098,In_3099,In_3100,In_3101,In_3102,In_3103,In_3104,In_3105,In_3106,In_3107,In_3108,In_3109,In_3110,In_3111,In_3112,In_3113,In_3114,In_3115,In_3116,In_3117,In_3118,In_3119,In_3120,In_3121,In_3122,In_3123,In_3124,In_3125,In_3126,In_3127,In_3128,In_3129,In_3130,In_3131,In_3132,In_3133,In_3134,In_3135,In_3136,In_3137,In_3138,In_3139,In_3140,In_3141,In_3142,In_3143,In_3144,In_3145,In_3146,In_3147,In_3148,In_3149,In_3150,In_3151,In_3152,In_3153,In_3154,In_3155,In_3156,In_3157,In_3158,In_3159,In_3160,In_3161,In_3162,In_3163,In_3164,In_3165,In_3166,In_3167,In_3168,In_3169,In_3170,In_3171,In_3172,In_3173,In_3174,In_3175,In_3176,In_3177,In_3178,In_3179,In_3180,In_3181,In_3182,In_3183,In_3184,In_3185,In_3186,In_3187,In_3188,In_3189,In_3190,In_3191,In_3192,In_3193,In_3194,In_3195,In_3196,In_3197,In_3198,In_3199,In_3200,In_3201,In_3202,In_3203,In_3204,In_3205,In_3206,In_3207,In_3208,In_3209,In_3210,In_3211,In_3212,In_3213,In_3214,In_3215,In_3216,In_3217,In_3218,In_3219,In_3220,In_3221,In_3222,In_3223,In_3224,In_3225,In_3226,In_3227,In_3228,In_3229,In_3230,In_3231,In_3232,In_3233,In_3234,In_3235,In_3236,In_3237,In_3238,In_3239,In_3240,In_3241,In_3242,In_3243,In_3244,In_3245,In_3246,In_3247,In_3248,In_3249,In_3250,In_3251,In_3252,In_3253,In_3254,In_3255,In_3256,In_3257,In_3258,In_3259,In_3260,In_3261,In_3262,In_3263,In_3264,In_3265,In_3266,In_3267,In_3268,In_3269,In_3270,In_3271,In_3272,In_3273,In_3274,In_3275,In_3276,In_3277,In_3278,In_3279,In_3280,In_3281,In_3282,In_3283,In_3284,In_3285,In_3286,In_3287,In_3288,In_3289,In_3290,In_3291,In_3292,In_3293,In_3294,In_3295,In_3296,In_3297,In_3298,In_3299,In_3300,In_3301,In_3302,In_3303,In_3304,In_3305,In_3306,In_3307,In_3308,In_3309,In_3310,In_3311,In_3312,In_3313,In_3314,In_3315,In_3316,In_3317,In_3318,In_3319,In_3320,In_3321,In_3322,In_3323,In_3324,In_3325,In_3326,In_3327,In_3328,In_3329,In_3330,In_3331,In_3332,In_3333,In_3334,In_3335,In_3336,In_3337,In_3338,In_3339,In_3340,In_3341,In_3342,In_3343,In_3344,In_3345,In_3346,In_3347,In_3348,In_3349,In_3350,In_3351,In_3352,In_3353,In_3354,In_3355,In_3356,In_3357,In_3358,In_3359,In_3360,In_3361,In_3362,In_3363,In_3364,In_3365,In_3366,In_3367,In_3368,In_3369,In_3370,In_3371,In_3372,In_3373,In_3374,In_3375,In_3376,In_3377,In_3378,In_3379,In_3380,In_3381,In_3382,In_3383,In_3384,In_3385,In_3386,In_3387,In_3388,In_3389,In_3390,In_3391,In_3392,In_3393,In_3394,In_3395,In_3396,In_3397,In_3398,In_3399,In_3400,In_3401,In_3402,In_3403,In_3404,In_3405,In_3406,In_3407,In_3408,In_3409,In_3410,In_3411,In_3412,In_3413,In_3414,In_3415,In_3416,In_3417,In_3418,In_3419,In_3420,In_3421,In_3422,In_3423,In_3424,In_3425,In_3426,In_3427,In_3428,In_3429,In_3430,In_3431,In_3432,In_3433,In_3434,In_3435,In_3436,In_3437,In_3438,In_3439,In_3440,In_3441,In_3442,In_3443,In_3444,In_3445,In_3446,In_3447,In_3448,In_3449,In_3450,In_3451,In_3452,In_3453,In_3454,In_3455,In_3456,In_3457,In_3458,In_3459,In_3460,In_3461,In_3462,In_3463,In_3464,In_3465,In_3466,In_3467,In_3468,In_3469,In_3470,In_3471,In_3472,In_3473,In_3474,In_3475,In_3476,In_3477,In_3478,In_3479,In_3480,In_3481,In_3482,In_3483,In_3484,In_3485,In_3486,In_3487,In_3488,In_3489,In_3490,In_3491,In_3492,In_3493,In_3494,In_3495,In_3496,In_3497,In_3498,In_3499,In_3500,In_3501,In_3502,In_3503,In_3504,In_3505,In_3506,In_3507,In_3508,In_3509,In_3510,In_3511,In_3512,In_3513,In_3514,In_3515,In_3516,In_3517,In_3518,In_3519,In_3520,In_3521,In_3522,In_3523,In_3524,In_3525,In_3526,In_3527,In_3528,In_3529,In_3530,In_3531,In_3532,In_3533,In_3534,In_3535,In_3536,In_3537,In_3538,In_3539,In_3540,In_3541,In_3542,In_3543,In_3544,In_3545,In_3546,In_3547,In_3548,In_3549,In_3550,In_3551,In_3552,In_3553,In_3554,In_3555,In_3556,In_3557,In_3558,In_3559,In_3560,In_3561,In_3562,In_3563,In_3564,In_3565,In_3566,In_3567,In_3568,In_3569,In_3570,In_3571,In_3572,In_3573,In_3574,In_3575,In_3576,In_3577,In_3578,In_3579,In_3580,In_3581,In_3582,In_3583,In_3584,In_3585,In_3586,In_3587,In_3588,In_3589,In_3590,In_3591,In_3592,In_3593,In_3594,In_3595,In_3596,In_3597,In_3598,In_3599,In_3600,In_3601,In_3602,In_3603,In_3604,In_3605,In_3606,In_3607,In_3608,In_3609,In_3610,In_3611,In_3612,In_3613,In_3614,In_3615,In_3616,In_3617,In_3618,In_3619,In_3620,In_3621,In_3622,In_3623,In_3624,In_3625,In_3626,In_3627,In_3628,In_3629,In_3630,In_3631,In_3632,In_3633,In_3634,In_3635,In_3636,In_3637,In_3638,In_3639,In_3640,In_3641,In_3642,In_3643,In_3644,In_3645,In_3646,In_3647,In_3648,In_3649,In_3650,In_3651,In_3652,In_3653,In_3654,In_3655,In_3656,In_3657,In_3658,In_3659,In_3660,In_3661,In_3662,In_3663,In_3664,In_3665,In_3666,In_3667,In_3668,In_3669,In_3670,In_3671,In_3672,In_3673,In_3674,In_3675,In_3676,In_3677,In_3678,In_3679,In_3680,In_3681,In_3682,In_3683,In_3684,In_3685,In_3686,In_3687,In_3688,In_3689,In_3690,In_3691,In_3692,In_3693,In_3694,In_3695,In_3696,In_3697,In_3698,In_3699,In_3700,In_3701,In_3702,In_3703,In_3704,In_3705,In_3706,In_3707,In_3708,In_3709,In_3710,In_3711,In_3712,In_3713,In_3714,In_3715,In_3716,In_3717,In_3718,In_3719,In_3720,In_3721,In_3722,In_3723,In_3724,In_3725,In_3726,In_3727,In_3728,In_3729,In_3730,In_3731,In_3732,In_3733,In_3734,In_3735,In_3736,In_3737,In_3738,In_3739,In_3740,In_3741,In_3742,In_3743,In_3744,In_3745,In_3746,In_3747,In_3748,In_3749,In_3750,In_3751,In_3752,In_3753,In_3754,In_3755,In_3756,In_3757,In_3758,In_3759,In_3760,In_3761,In_3762,In_3763,In_3764,In_3765,In_3766,In_3767,In_3768,In_3769,In_3770,In_3771,In_3772,In_3773,In_3774,In_3775,In_3776,In_3777,In_3778,In_3779,In_3780,In_3781,In_3782,In_3783,In_3784,In_3785,In_3786,In_3787,In_3788,In_3789,In_3790,In_3791,In_3792,In_3793,In_3794,In_3795,In_3796,In_3797,In_3798,In_3799,In_3800,In_3801,In_3802,In_3803,In_3804,In_3805,In_3806,In_3807,In_3808,In_3809,In_3810,In_3811,In_3812,In_3813,In_3814,In_3815,In_3816,In_3817,In_3818,In_3819,In_3820,In_3821,In_3822,In_3823,In_3824,In_3825,In_3826,In_3827,In_3828,In_3829,In_3830,In_3831,In_3832,In_3833,In_3834,In_3835,In_3836,In_3837,In_3838,In_3839,In_3840,In_3841,In_3842,In_3843,In_3844,In_3845,In_3846,In_3847,In_3848,In_3849,In_3850,In_3851,In_3852,In_3853,In_3854,In_3855,In_3856,In_3857,In_3858,In_3859,In_3860,In_3861,In_3862,In_3863,In_3864,In_3865,In_3866,In_3867,In_3868,In_3869,In_3870,In_3871,In_3872,In_3873,In_3874,In_3875,In_3876,In_3877,In_3878,In_3879,In_3880,In_3881,In_3882,In_3883,In_3884,In_3885,In_3886,In_3887,In_3888,In_3889,In_3890,In_3891,In_3892,In_3893,In_3894,In_3895,In_3896,In_3897,In_3898,In_3899,In_3900,In_3901,In_3902,In_3903,In_3904,In_3905,In_3906,In_3907,In_3908,In_3909,In_3910,In_3911,In_3912,In_3913,In_3914,In_3915,In_3916,In_3917,In_3918,In_3919,In_3920,In_3921,In_3922,In_3923,In_3924,In_3925,In_3926,In_3927,In_3928,In_3929,In_3930,In_3931,In_3932,In_3933,In_3934,In_3935,In_3936,In_3937,In_3938,In_3939,In_3940,In_3941,In_3942,In_3943,In_3944,In_3945,In_3946,In_3947,In_3948,In_3949,In_3950,In_3951,In_3952,In_3953,In_3954,In_3955,In_3956,In_3957,In_3958,In_3959,In_3960,In_3961,In_3962,In_3963,In_3964,In_3965,In_3966,In_3967,In_3968,In_3969,In_3970,In_3971,In_3972,In_3973,In_3974,In_3975,In_3976,In_3977,In_3978,In_3979,In_3980,In_3981,In_3982,In_3983,In_3984,In_3985,In_3986,In_3987,In_3988,In_3989,In_3990,In_3991,In_3992,In_3993,In_3994,In_3995,In_3996,In_3997,In_3998,In_3999,In_4000,In_4001,In_4002,In_4003,In_4004,In_4005,In_4006,In_4007,In_4008,In_4009,In_4010,In_4011,In_4012,In_4013,In_4014,In_4015,In_4016,In_4017,In_4018,In_4019,In_4020,In_4021,In_4022,In_4023,In_4024,In_4025,In_4026,In_4027,In_4028,In_4029,In_4030,In_4031,In_4032,In_4033,In_4034,In_4035,In_4036,In_4037,In_4038,In_4039,In_4040,In_4041,In_4042,In_4043,In_4044,In_4045,In_4046,In_4047,In_4048,In_4049,In_4050,In_4051,In_4052,In_4053,In_4054,In_4055,In_4056,In_4057,In_4058,In_4059,In_4060,In_4061,In_4062,In_4063,In_4064,In_4065,In_4066,In_4067,In_4068,In_4069,In_4070,In_4071,In_4072,In_4073,In_4074,In_4075,In_4076,In_4077,In_4078,In_4079,In_4080,In_4081,In_4082,In_4083,In_4084,In_4085,In_4086,In_4087,In_4088,In_4089,In_4090,In_4091,In_4092,In_4093,In_4094,In_4095,In_4096,In_4097,In_4098,In_4099,In_4100,In_4101,In_4102,In_4103,In_4104,In_4105,In_4106,In_4107,In_4108,In_4109,In_4110,In_4111,In_4112,In_4113,In_4114,In_4115,In_4116,In_4117,In_4118,In_4119,In_4120,In_4121,In_4122,In_4123,In_4124,In_4125,In_4126,In_4127,In_4128,In_4129,In_4130,In_4131,In_4132,In_4133,In_4134,In_4135,In_4136,In_4137,In_4138,In_4139,In_4140,In_4141,In_4142,In_4143,In_4144,In_4145,In_4146,In_4147,In_4148,In_4149,In_4150,In_4151,In_4152,In_4153,In_4154,In_4155,In_4156,In_4157,In_4158,In_4159,In_4160,In_4161,In_4162,In_4163,In_4164,In_4165,In_4166,In_4167,In_4168,In_4169,In_4170,In_4171,In_4172,In_4173,In_4174,In_4175,In_4176,In_4177,In_4178,In_4179,In_4180,In_4181,In_4182,In_4183,In_4184,In_4185,In_4186,In_4187,In_4188,In_4189,In_4190,In_4191,In_4192,In_4193,In_4194,In_4195,In_4196,In_4197,In_4198,In_4199,In_4200,In_4201,In_4202,In_4203,In_4204,In_4205,In_4206,In_4207,In_4208,In_4209,In_4210,In_4211,In_4212,In_4213,In_4214,In_4215,In_4216,In_4217,In_4218,In_4219,In_4220,In_4221,In_4222,In_4223,In_4224,In_4225,In_4226,In_4227,In_4228,In_4229,In_4230,In_4231,In_4232,In_4233,In_4234,In_4235,In_4236,In_4237,In_4238,In_4239,In_4240,In_4241,In_4242,In_4243,In_4244,In_4245,In_4246,In_4247,In_4248,In_4249,In_4250,In_4251,In_4252,In_4253,In_4254,In_4255,In_4256,In_4257,In_4258,In_4259,In_4260,In_4261,In_4262,In_4263,In_4264,In_4265,In_4266,In_4267,In_4268,In_4269,In_4270,In_4271,In_4272,In_4273,In_4274,In_4275,In_4276,In_4277,In_4278,In_4279,In_4280,In_4281,In_4282,In_4283,In_4284,In_4285,In_4286,In_4287,In_4288,In_4289,In_4290,In_4291,In_4292,In_4293,In_4294,In_4295,In_4296,In_4297,In_4298,In_4299,In_4300,In_4301,In_4302,In_4303,In_4304,In_4305,In_4306,In_4307,In_4308,In_4309,In_4310,In_4311,In_4312,In_4313,In_4314,In_4315,In_4316,In_4317,In_4318,In_4319,In_4320,In_4321,In_4322,In_4323,In_4324,In_4325,In_4326,In_4327,In_4328,In_4329,In_4330,In_4331,In_4332,In_4333,In_4334,In_4335,In_4336,In_4337,In_4338,In_4339,In_4340,In_4341,In_4342,In_4343,In_4344,In_4345,In_4346,In_4347,In_4348,In_4349,In_4350,In_4351,In_4352,In_4353,In_4354,In_4355,In_4356,In_4357,In_4358,In_4359,In_4360,In_4361,In_4362,In_4363,In_4364,In_4365,In_4366,In_4367,In_4368,In_4369,In_4370,In_4371,In_4372,In_4373,In_4374,In_4375,In_4376,In_4377,In_4378,In_4379,In_4380,In_4381,In_4382,In_4383,In_4384,In_4385,In_4386,In_4387,In_4388,In_4389,In_4390,In_4391,In_4392,In_4393,In_4394,In_4395,In_4396,In_4397,In_4398,In_4399,In_4400,In_4401,In_4402,In_4403,In_4404,In_4405,In_4406,In_4407,In_4408,In_4409,In_4410,In_4411,In_4412,In_4413,In_4414,In_4415,In_4416,In_4417,In_4418,In_4419,In_4420,In_4421,In_4422,In_4423,In_4424,In_4425,In_4426,In_4427,In_4428,In_4429,In_4430,In_4431,In_4432,In_4433,In_4434,In_4435,In_4436,In_4437,In_4438,In_4439,In_4440,In_4441,In_4442,In_4443,In_4444,In_4445,In_4446,In_4447,In_4448,In_4449,In_4450,In_4451,In_4452,In_4453,In_4454,In_4455,In_4456,In_4457,In_4458,In_4459,In_4460,In_4461,In_4462,In_4463,In_4464,In_4465,In_4466,In_4467,In_4468,In_4469,In_4470,In_4471,In_4472,In_4473,In_4474,In_4475,In_4476,In_4477,In_4478,In_4479,In_4480,In_4481,In_4482,In_4483,In_4484,In_4485,In_4486,In_4487,In_4488,In_4489,In_4490,In_4491,In_4492,In_4493,In_4494,In_4495,In_4496,In_4497,In_4498,In_4499,In_4500,In_4501,In_4502,In_4503,In_4504,In_4505,In_4506,In_4507,In_4508,In_4509,In_4510,In_4511,In_4512,In_4513,In_4514,In_4515,In_4516,In_4517,In_4518,In_4519,In_4520,In_4521,In_4522,In_4523,In_4524,In_4525,In_4526,In_4527,In_4528,In_4529,In_4530,In_4531,In_4532,In_4533,In_4534,In_4535,In_4536,In_4537,In_4538,In_4539,In_4540,In_4541,In_4542,In_4543,In_4544,In_4545,In_4546,In_4547,In_4548,In_4549,In_4550,In_4551,In_4552,In_4553,In_4554,In_4555,In_4556,In_4557,In_4558,In_4559,In_4560,In_4561,In_4562,In_4563,In_4564,In_4565,In_4566,In_4567,In_4568,In_4569,In_4570,In_4571,In_4572,In_4573,In_4574,In_4575,In_4576,In_4577,In_4578,In_4579,In_4580,In_4581,In_4582,In_4583,In_4584,In_4585,In_4586,In_4587,In_4588,In_4589,In_4590,In_4591,In_4592,In_4593,In_4594,In_4595,In_4596,In_4597,In_4598,In_4599,In_4600,In_4601,In_4602,In_4603,In_4604,In_4605,In_4606,In_4607,In_4608,In_4609,In_4610,In_4611,In_4612,In_4613,In_4614,In_4615,In_4616,In_4617,In_4618,In_4619,In_4620,In_4621,In_4622,In_4623,In_4624,In_4625,In_4626,In_4627,In_4628,In_4629,In_4630,In_4631,In_4632,In_4633,In_4634,In_4635,In_4636,In_4637,In_4638,In_4639,In_4640,In_4641,In_4642,In_4643,In_4644,In_4645,In_4646,In_4647,In_4648,In_4649,In_4650,In_4651,In_4652,In_4653,In_4654,In_4655,In_4656,In_4657,In_4658,In_4659,In_4660,In_4661,In_4662,In_4663,In_4664,In_4665,In_4666,In_4667,In_4668,In_4669,In_4670,In_4671,In_4672,In_4673,In_4674,In_4675,In_4676,In_4677,In_4678,In_4679,In_4680,In_4681,In_4682,In_4683,In_4684,In_4685,In_4686,In_4687,In_4688,In_4689,In_4690,In_4691,In_4692,In_4693,In_4694,In_4695,In_4696,In_4697,In_4698,In_4699,In_4700,In_4701,In_4702,In_4703,In_4704,In_4705,In_4706,In_4707,In_4708,In_4709,In_4710,In_4711,In_4712,In_4713,In_4714,In_4715,In_4716,In_4717,In_4718,In_4719,In_4720,In_4721,In_4722,In_4723,In_4724,In_4725,In_4726,In_4727,In_4728,In_4729,In_4730,In_4731,In_4732,In_4733,In_4734,In_4735,In_4736,In_4737,In_4738,In_4739,In_4740,In_4741,In_4742,In_4743,In_4744,In_4745,In_4746,In_4747,In_4748,In_4749,In_4750,In_4751,In_4752,In_4753,In_4754,In_4755,In_4756,In_4757,In_4758,In_4759,In_4760,In_4761,In_4762,In_4763,In_4764,In_4765,In_4766,In_4767,In_4768,In_4769,In_4770,In_4771,In_4772,In_4773,In_4774,In_4775,In_4776,In_4777,In_4778,In_4779,In_4780,In_4781,In_4782,In_4783,In_4784,In_4785,In_4786,In_4787,In_4788,In_4789,In_4790,In_4791,In_4792,In_4793,In_4794,In_4795,In_4796,In_4797,In_4798,In_4799,In_4800,In_4801,In_4802,In_4803,In_4804,In_4805,In_4806,In_4807,In_4808,In_4809,In_4810,In_4811,In_4812,In_4813,In_4814,In_4815,In_4816,In_4817,In_4818,In_4819,In_4820,In_4821,In_4822,In_4823,In_4824,In_4825,In_4826,In_4827,In_4828,In_4829,In_4830,In_4831,In_4832,In_4833,In_4834,In_4835,In_4836,In_4837,In_4838,In_4839,In_4840,In_4841,In_4842,In_4843,In_4844,In_4845,In_4846,In_4847,In_4848,In_4849,In_4850,In_4851,In_4852,In_4853,In_4854,In_4855,In_4856,In_4857,In_4858,In_4859,In_4860,In_4861,In_4862,In_4863,In_4864,In_4865,In_4866,In_4867,In_4868,In_4869,In_4870,In_4871,In_4872,In_4873,In_4874,In_4875,In_4876,In_4877,In_4878,In_4879,In_4880,In_4881,In_4882,In_4883,In_4884,In_4885,In_4886,In_4887,In_4888,In_4889,In_4890,In_4891,In_4892,In_4893,In_4894,In_4895,In_4896,In_4897,In_4898,In_4899,In_4900,In_4901,In_4902,In_4903,In_4904,In_4905,In_4906,In_4907,In_4908,In_4909,In_4910,In_4911,In_4912,In_4913,In_4914,In_4915,In_4916,In_4917,In_4918,In_4919,In_4920,In_4921,In_4922,In_4923,In_4924,In_4925,In_4926,In_4927,In_4928,In_4929,In_4930,In_4931,In_4932,In_4933,In_4934,In_4935,In_4936,In_4937,In_4938,In_4939,In_4940,In_4941,In_4942,In_4943,In_4944,In_4945,In_4946,In_4947,In_4948,In_4949,In_4950,In_4951,In_4952,In_4953,In_4954,In_4955,In_4956,In_4957,In_4958,In_4959,In_4960,In_4961,In_4962,In_4963,In_4964,In_4965,In_4966,In_4967,In_4968,In_4969,In_4970,In_4971,In_4972,In_4973,In_4974,In_4975,In_4976,In_4977,In_4978,In_4979,In_4980,In_4981,In_4982,In_4983,In_4984,In_4985,In_4986,In_4987,In_4988,In_4989,In_4990,In_4991,In_4992,In_4993,In_4994,In_4995,In_4996,In_4997,In_4998,In_4999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499,O_3500,O_3501,O_3502,O_3503,O_3504,O_3505,O_3506,O_3507,O_3508,O_3509,O_3510,O_3511,O_3512,O_3513,O_3514,O_3515,O_3516,O_3517,O_3518,O_3519,O_3520,O_3521,O_3522,O_3523,O_3524,O_3525,O_3526,O_3527,O_3528,O_3529,O_3530,O_3531,O_3532,O_3533,O_3534,O_3535,O_3536,O_3537,O_3538,O_3539,O_3540,O_3541,O_3542,O_3543,O_3544,O_3545,O_3546,O_3547,O_3548,O_3549,O_3550,O_3551,O_3552,O_3553,O_3554,O_3555,O_3556,O_3557,O_3558,O_3559,O_3560,O_3561,O_3562,O_3563,O_3564,O_3565,O_3566,O_3567,O_3568,O_3569,O_3570,O_3571,O_3572,O_3573,O_3574,O_3575,O_3576,O_3577,O_3578,O_3579,O_3580,O_3581,O_3582,O_3583,O_3584,O_3585,O_3586,O_3587,O_3588,O_3589,O_3590,O_3591,O_3592,O_3593,O_3594,O_3595,O_3596,O_3597,O_3598,O_3599,O_3600,O_3601,O_3602,O_3603,O_3604,O_3605,O_3606,O_3607,O_3608,O_3609,O_3610,O_3611,O_3612,O_3613,O_3614,O_3615,O_3616,O_3617,O_3618,O_3619,O_3620,O_3621,O_3622,O_3623,O_3624,O_3625,O_3626,O_3627,O_3628,O_3629,O_3630,O_3631,O_3632,O_3633,O_3634,O_3635,O_3636,O_3637,O_3638,O_3639,O_3640,O_3641,O_3642,O_3643,O_3644,O_3645,O_3646,O_3647,O_3648,O_3649,O_3650,O_3651,O_3652,O_3653,O_3654,O_3655,O_3656,O_3657,O_3658,O_3659,O_3660,O_3661,O_3662,O_3663,O_3664,O_3665,O_3666,O_3667,O_3668,O_3669,O_3670,O_3671,O_3672,O_3673,O_3674,O_3675,O_3676,O_3677,O_3678,O_3679,O_3680,O_3681,O_3682,O_3683,O_3684,O_3685,O_3686,O_3687,O_3688,O_3689,O_3690,O_3691,O_3692,O_3693,O_3694,O_3695,O_3696,O_3697,O_3698,O_3699,O_3700,O_3701,O_3702,O_3703,O_3704,O_3705,O_3706,O_3707,O_3708,O_3709,O_3710,O_3711,O_3712,O_3713,O_3714,O_3715,O_3716,O_3717,O_3718,O_3719,O_3720,O_3721,O_3722,O_3723,O_3724,O_3725,O_3726,O_3727,O_3728,O_3729,O_3730,O_3731,O_3732,O_3733,O_3734,O_3735,O_3736,O_3737,O_3738,O_3739,O_3740,O_3741,O_3742,O_3743,O_3744,O_3745,O_3746,O_3747,O_3748,O_3749,O_3750,O_3751,O_3752,O_3753,O_3754,O_3755,O_3756,O_3757,O_3758,O_3759,O_3760,O_3761,O_3762,O_3763,O_3764,O_3765,O_3766,O_3767,O_3768,O_3769,O_3770,O_3771,O_3772,O_3773,O_3774,O_3775,O_3776,O_3777,O_3778,O_3779,O_3780,O_3781,O_3782,O_3783,O_3784,O_3785,O_3786,O_3787,O_3788,O_3789,O_3790,O_3791,O_3792,O_3793,O_3794,O_3795,O_3796,O_3797,O_3798,O_3799,O_3800,O_3801,O_3802,O_3803,O_3804,O_3805,O_3806,O_3807,O_3808,O_3809,O_3810,O_3811,O_3812,O_3813,O_3814,O_3815,O_3816,O_3817,O_3818,O_3819,O_3820,O_3821,O_3822,O_3823,O_3824,O_3825,O_3826,O_3827,O_3828,O_3829,O_3830,O_3831,O_3832,O_3833,O_3834,O_3835,O_3836,O_3837,O_3838,O_3839,O_3840,O_3841,O_3842,O_3843,O_3844,O_3845,O_3846,O_3847,O_3848,O_3849,O_3850,O_3851,O_3852,O_3853,O_3854,O_3855,O_3856,O_3857,O_3858,O_3859,O_3860,O_3861,O_3862,O_3863,O_3864,O_3865,O_3866,O_3867,O_3868,O_3869,O_3870,O_3871,O_3872,O_3873,O_3874,O_3875,O_3876,O_3877,O_3878,O_3879,O_3880,O_3881,O_3882,O_3883,O_3884,O_3885,O_3886,O_3887,O_3888,O_3889,O_3890,O_3891,O_3892,O_3893,O_3894,O_3895,O_3896,O_3897,O_3898,O_3899,O_3900,O_3901,O_3902,O_3903,O_3904,O_3905,O_3906,O_3907,O_3908,O_3909,O_3910,O_3911,O_3912,O_3913,O_3914,O_3915,O_3916,O_3917,O_3918,O_3919,O_3920,O_3921,O_3922,O_3923,O_3924,O_3925,O_3926,O_3927,O_3928,O_3929,O_3930,O_3931,O_3932,O_3933,O_3934,O_3935,O_3936,O_3937,O_3938,O_3939,O_3940,O_3941,O_3942,O_3943,O_3944,O_3945,O_3946,O_3947,O_3948,O_3949,O_3950,O_3951,O_3952,O_3953,O_3954,O_3955,O_3956,O_3957,O_3958,O_3959,O_3960,O_3961,O_3962,O_3963,O_3964,O_3965,O_3966,O_3967,O_3968,O_3969,O_3970,O_3971,O_3972,O_3973,O_3974,O_3975,O_3976,O_3977,O_3978,O_3979,O_3980,O_3981,O_3982,O_3983,O_3984,O_3985,O_3986,O_3987,O_3988,O_3989,O_3990,O_3991,O_3992,O_3993,O_3994,O_3995,O_3996,O_3997,O_3998,O_3999,O_4000,O_4001,O_4002,O_4003,O_4004,O_4005,O_4006,O_4007,O_4008,O_4009,O_4010,O_4011,O_4012,O_4013,O_4014,O_4015,O_4016,O_4017,O_4018,O_4019,O_4020,O_4021,O_4022,O_4023,O_4024,O_4025,O_4026,O_4027,O_4028,O_4029,O_4030,O_4031,O_4032,O_4033,O_4034,O_4035,O_4036,O_4037,O_4038,O_4039,O_4040,O_4041,O_4042,O_4043,O_4044,O_4045,O_4046,O_4047,O_4048,O_4049,O_4050,O_4051,O_4052,O_4053,O_4054,O_4055,O_4056,O_4057,O_4058,O_4059,O_4060,O_4061,O_4062,O_4063,O_4064,O_4065,O_4066,O_4067,O_4068,O_4069,O_4070,O_4071,O_4072,O_4073,O_4074,O_4075,O_4076,O_4077,O_4078,O_4079,O_4080,O_4081,O_4082,O_4083,O_4084,O_4085,O_4086,O_4087,O_4088,O_4089,O_4090,O_4091,O_4092,O_4093,O_4094,O_4095,O_4096,O_4097,O_4098,O_4099,O_4100,O_4101,O_4102,O_4103,O_4104,O_4105,O_4106,O_4107,O_4108,O_4109,O_4110,O_4111,O_4112,O_4113,O_4114,O_4115,O_4116,O_4117,O_4118,O_4119,O_4120,O_4121,O_4122,O_4123,O_4124,O_4125,O_4126,O_4127,O_4128,O_4129,O_4130,O_4131,O_4132,O_4133,O_4134,O_4135,O_4136,O_4137,O_4138,O_4139,O_4140,O_4141,O_4142,O_4143,O_4144,O_4145,O_4146,O_4147,O_4148,O_4149,O_4150,O_4151,O_4152,O_4153,O_4154,O_4155,O_4156,O_4157,O_4158,O_4159,O_4160,O_4161,O_4162,O_4163,O_4164,O_4165,O_4166,O_4167,O_4168,O_4169,O_4170,O_4171,O_4172,O_4173,O_4174,O_4175,O_4176,O_4177,O_4178,O_4179,O_4180,O_4181,O_4182,O_4183,O_4184,O_4185,O_4186,O_4187,O_4188,O_4189,O_4190,O_4191,O_4192,O_4193,O_4194,O_4195,O_4196,O_4197,O_4198,O_4199,O_4200,O_4201,O_4202,O_4203,O_4204,O_4205,O_4206,O_4207,O_4208,O_4209,O_4210,O_4211,O_4212,O_4213,O_4214,O_4215,O_4216,O_4217,O_4218,O_4219,O_4220,O_4221,O_4222,O_4223,O_4224,O_4225,O_4226,O_4227,O_4228,O_4229,O_4230,O_4231,O_4232,O_4233,O_4234,O_4235,O_4236,O_4237,O_4238,O_4239,O_4240,O_4241,O_4242,O_4243,O_4244,O_4245,O_4246,O_4247,O_4248,O_4249,O_4250,O_4251,O_4252,O_4253,O_4254,O_4255,O_4256,O_4257,O_4258,O_4259,O_4260,O_4261,O_4262,O_4263,O_4264,O_4265,O_4266,O_4267,O_4268,O_4269,O_4270,O_4271,O_4272,O_4273,O_4274,O_4275,O_4276,O_4277,O_4278,O_4279,O_4280,O_4281,O_4282,O_4283,O_4284,O_4285,O_4286,O_4287,O_4288,O_4289,O_4290,O_4291,O_4292,O_4293,O_4294,O_4295,O_4296,O_4297,O_4298,O_4299,O_4300,O_4301,O_4302,O_4303,O_4304,O_4305,O_4306,O_4307,O_4308,O_4309,O_4310,O_4311,O_4312,O_4313,O_4314,O_4315,O_4316,O_4317,O_4318,O_4319,O_4320,O_4321,O_4322,O_4323,O_4324,O_4325,O_4326,O_4327,O_4328,O_4329,O_4330,O_4331,O_4332,O_4333,O_4334,O_4335,O_4336,O_4337,O_4338,O_4339,O_4340,O_4341,O_4342,O_4343,O_4344,O_4345,O_4346,O_4347,O_4348,O_4349,O_4350,O_4351,O_4352,O_4353,O_4354,O_4355,O_4356,O_4357,O_4358,O_4359,O_4360,O_4361,O_4362,O_4363,O_4364,O_4365,O_4366,O_4367,O_4368,O_4369,O_4370,O_4371,O_4372,O_4373,O_4374,O_4375,O_4376,O_4377,O_4378,O_4379,O_4380,O_4381,O_4382,O_4383,O_4384,O_4385,O_4386,O_4387,O_4388,O_4389,O_4390,O_4391,O_4392,O_4393,O_4394,O_4395,O_4396,O_4397,O_4398,O_4399,O_4400,O_4401,O_4402,O_4403,O_4404,O_4405,O_4406,O_4407,O_4408,O_4409,O_4410,O_4411,O_4412,O_4413,O_4414,O_4415,O_4416,O_4417,O_4418,O_4419,O_4420,O_4421,O_4422,O_4423,O_4424,O_4425,O_4426,O_4427,O_4428,O_4429,O_4430,O_4431,O_4432,O_4433,O_4434,O_4435,O_4436,O_4437,O_4438,O_4439,O_4440,O_4441,O_4442,O_4443,O_4444,O_4445,O_4446,O_4447,O_4448,O_4449,O_4450,O_4451,O_4452,O_4453,O_4454,O_4455,O_4456,O_4457,O_4458,O_4459,O_4460,O_4461,O_4462,O_4463,O_4464,O_4465,O_4466,O_4467,O_4468,O_4469,O_4470,O_4471,O_4472,O_4473,O_4474,O_4475,O_4476,O_4477,O_4478,O_4479,O_4480,O_4481,O_4482,O_4483,O_4484,O_4485,O_4486,O_4487,O_4488,O_4489,O_4490,O_4491,O_4492,O_4493,O_4494,O_4495,O_4496,O_4497,O_4498,O_4499,O_4500,O_4501,O_4502,O_4503,O_4504,O_4505,O_4506,O_4507,O_4508,O_4509,O_4510,O_4511,O_4512,O_4513,O_4514,O_4515,O_4516,O_4517,O_4518,O_4519,O_4520,O_4521,O_4522,O_4523,O_4524,O_4525,O_4526,O_4527,O_4528,O_4529,O_4530,O_4531,O_4532,O_4533,O_4534,O_4535,O_4536,O_4537,O_4538,O_4539,O_4540,O_4541,O_4542,O_4543,O_4544,O_4545,O_4546,O_4547,O_4548,O_4549,O_4550,O_4551,O_4552,O_4553,O_4554,O_4555,O_4556,O_4557,O_4558,O_4559,O_4560,O_4561,O_4562,O_4563,O_4564,O_4565,O_4566,O_4567,O_4568,O_4569,O_4570,O_4571,O_4572,O_4573,O_4574,O_4575,O_4576,O_4577,O_4578,O_4579,O_4580,O_4581,O_4582,O_4583,O_4584,O_4585,O_4586,O_4587,O_4588,O_4589,O_4590,O_4591,O_4592,O_4593,O_4594,O_4595,O_4596,O_4597,O_4598,O_4599,O_4600,O_4601,O_4602,O_4603,O_4604,O_4605,O_4606,O_4607,O_4608,O_4609,O_4610,O_4611,O_4612,O_4613,O_4614,O_4615,O_4616,O_4617,O_4618,O_4619,O_4620,O_4621,O_4622,O_4623,O_4624,O_4625,O_4626,O_4627,O_4628,O_4629,O_4630,O_4631,O_4632,O_4633,O_4634,O_4635,O_4636,O_4637,O_4638,O_4639,O_4640,O_4641,O_4642,O_4643,O_4644,O_4645,O_4646,O_4647,O_4648,O_4649,O_4650,O_4651,O_4652,O_4653,O_4654,O_4655,O_4656,O_4657,O_4658,O_4659,O_4660,O_4661,O_4662,O_4663,O_4664,O_4665,O_4666,O_4667,O_4668,O_4669,O_4670,O_4671,O_4672,O_4673,O_4674,O_4675,O_4676,O_4677,O_4678,O_4679,O_4680,O_4681,O_4682,O_4683,O_4684,O_4685,O_4686,O_4687,O_4688,O_4689,O_4690,O_4691,O_4692,O_4693,O_4694,O_4695,O_4696,O_4697,O_4698,O_4699,O_4700,O_4701,O_4702,O_4703,O_4704,O_4705,O_4706,O_4707,O_4708,O_4709,O_4710,O_4711,O_4712,O_4713,O_4714,O_4715,O_4716,O_4717,O_4718,O_4719,O_4720,O_4721,O_4722,O_4723,O_4724,O_4725,O_4726,O_4727,O_4728,O_4729,O_4730,O_4731,O_4732,O_4733,O_4734,O_4735,O_4736,O_4737,O_4738,O_4739,O_4740,O_4741,O_4742,O_4743,O_4744,O_4745,O_4746,O_4747,O_4748,O_4749,O_4750,O_4751,O_4752,O_4753,O_4754,O_4755,O_4756,O_4757,O_4758,O_4759,O_4760,O_4761,O_4762,O_4763,O_4764,O_4765,O_4766,O_4767,O_4768,O_4769,O_4770,O_4771,O_4772,O_4773,O_4774,O_4775,O_4776,O_4777,O_4778,O_4779,O_4780,O_4781,O_4782,O_4783,O_4784,O_4785,O_4786,O_4787,O_4788,O_4789,O_4790,O_4791,O_4792,O_4793,O_4794,O_4795,O_4796,O_4797,O_4798,O_4799,O_4800,O_4801,O_4802,O_4803,O_4804,O_4805,O_4806,O_4807,O_4808,O_4809,O_4810,O_4811,O_4812,O_4813,O_4814,O_4815,O_4816,O_4817,O_4818,O_4819,O_4820,O_4821,O_4822,O_4823,O_4824,O_4825,O_4826,O_4827,O_4828,O_4829,O_4830,O_4831,O_4832,O_4833,O_4834,O_4835,O_4836,O_4837,O_4838,O_4839,O_4840,O_4841,O_4842,O_4843,O_4844,O_4845,O_4846,O_4847,O_4848,O_4849,O_4850,O_4851,O_4852,O_4853,O_4854,O_4855,O_4856,O_4857,O_4858,O_4859,O_4860,O_4861,O_4862,O_4863,O_4864,O_4865,O_4866,O_4867,O_4868,O_4869,O_4870,O_4871,O_4872,O_4873,O_4874,O_4875,O_4876,O_4877,O_4878,O_4879,O_4880,O_4881,O_4882,O_4883,O_4884,O_4885,O_4886,O_4887,O_4888,O_4889,O_4890,O_4891,O_4892,O_4893,O_4894,O_4895,O_4896,O_4897,O_4898,O_4899,O_4900,O_4901,O_4902,O_4903,O_4904,O_4905,O_4906,O_4907,O_4908,O_4909,O_4910,O_4911,O_4912,O_4913,O_4914,O_4915,O_4916,O_4917,O_4918,O_4919,O_4920,O_4921,O_4922,O_4923,O_4924,O_4925,O_4926,O_4927,O_4928,O_4929,O_4930,O_4931,O_4932,O_4933,O_4934,O_4935,O_4936,O_4937,O_4938,O_4939,O_4940,O_4941,O_4942,O_4943,O_4944,O_4945,O_4946,O_4947,O_4948,O_4949,O_4950,O_4951,O_4952,O_4953,O_4954,O_4955,O_4956,O_4957,O_4958,O_4959,O_4960,O_4961,O_4962,O_4963,O_4964,O_4965,O_4966,O_4967,O_4968,O_4969,O_4970,O_4971,O_4972,O_4973,O_4974,O_4975,O_4976,O_4977,O_4978,O_4979,O_4980,O_4981,O_4982,O_4983,O_4984,O_4985,O_4986,O_4987,O_4988,O_4989,O_4990,O_4991,O_4992,O_4993,O_4994,O_4995,O_4996,O_4997,O_4998,O_4999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,In_3000,In_3001,In_3002,In_3003,In_3004,In_3005,In_3006,In_3007,In_3008,In_3009,In_3010,In_3011,In_3012,In_3013,In_3014,In_3015,In_3016,In_3017,In_3018,In_3019,In_3020,In_3021,In_3022,In_3023,In_3024,In_3025,In_3026,In_3027,In_3028,In_3029,In_3030,In_3031,In_3032,In_3033,In_3034,In_3035,In_3036,In_3037,In_3038,In_3039,In_3040,In_3041,In_3042,In_3043,In_3044,In_3045,In_3046,In_3047,In_3048,In_3049,In_3050,In_3051,In_3052,In_3053,In_3054,In_3055,In_3056,In_3057,In_3058,In_3059,In_3060,In_3061,In_3062,In_3063,In_3064,In_3065,In_3066,In_3067,In_3068,In_3069,In_3070,In_3071,In_3072,In_3073,In_3074,In_3075,In_3076,In_3077,In_3078,In_3079,In_3080,In_3081,In_3082,In_3083,In_3084,In_3085,In_3086,In_3087,In_3088,In_3089,In_3090,In_3091,In_3092,In_3093,In_3094,In_3095,In_3096,In_3097,In_3098,In_3099,In_3100,In_3101,In_3102,In_3103,In_3104,In_3105,In_3106,In_3107,In_3108,In_3109,In_3110,In_3111,In_3112,In_3113,In_3114,In_3115,In_3116,In_3117,In_3118,In_3119,In_3120,In_3121,In_3122,In_3123,In_3124,In_3125,In_3126,In_3127,In_3128,In_3129,In_3130,In_3131,In_3132,In_3133,In_3134,In_3135,In_3136,In_3137,In_3138,In_3139,In_3140,In_3141,In_3142,In_3143,In_3144,In_3145,In_3146,In_3147,In_3148,In_3149,In_3150,In_3151,In_3152,In_3153,In_3154,In_3155,In_3156,In_3157,In_3158,In_3159,In_3160,In_3161,In_3162,In_3163,In_3164,In_3165,In_3166,In_3167,In_3168,In_3169,In_3170,In_3171,In_3172,In_3173,In_3174,In_3175,In_3176,In_3177,In_3178,In_3179,In_3180,In_3181,In_3182,In_3183,In_3184,In_3185,In_3186,In_3187,In_3188,In_3189,In_3190,In_3191,In_3192,In_3193,In_3194,In_3195,In_3196,In_3197,In_3198,In_3199,In_3200,In_3201,In_3202,In_3203,In_3204,In_3205,In_3206,In_3207,In_3208,In_3209,In_3210,In_3211,In_3212,In_3213,In_3214,In_3215,In_3216,In_3217,In_3218,In_3219,In_3220,In_3221,In_3222,In_3223,In_3224,In_3225,In_3226,In_3227,In_3228,In_3229,In_3230,In_3231,In_3232,In_3233,In_3234,In_3235,In_3236,In_3237,In_3238,In_3239,In_3240,In_3241,In_3242,In_3243,In_3244,In_3245,In_3246,In_3247,In_3248,In_3249,In_3250,In_3251,In_3252,In_3253,In_3254,In_3255,In_3256,In_3257,In_3258,In_3259,In_3260,In_3261,In_3262,In_3263,In_3264,In_3265,In_3266,In_3267,In_3268,In_3269,In_3270,In_3271,In_3272,In_3273,In_3274,In_3275,In_3276,In_3277,In_3278,In_3279,In_3280,In_3281,In_3282,In_3283,In_3284,In_3285,In_3286,In_3287,In_3288,In_3289,In_3290,In_3291,In_3292,In_3293,In_3294,In_3295,In_3296,In_3297,In_3298,In_3299,In_3300,In_3301,In_3302,In_3303,In_3304,In_3305,In_3306,In_3307,In_3308,In_3309,In_3310,In_3311,In_3312,In_3313,In_3314,In_3315,In_3316,In_3317,In_3318,In_3319,In_3320,In_3321,In_3322,In_3323,In_3324,In_3325,In_3326,In_3327,In_3328,In_3329,In_3330,In_3331,In_3332,In_3333,In_3334,In_3335,In_3336,In_3337,In_3338,In_3339,In_3340,In_3341,In_3342,In_3343,In_3344,In_3345,In_3346,In_3347,In_3348,In_3349,In_3350,In_3351,In_3352,In_3353,In_3354,In_3355,In_3356,In_3357,In_3358,In_3359,In_3360,In_3361,In_3362,In_3363,In_3364,In_3365,In_3366,In_3367,In_3368,In_3369,In_3370,In_3371,In_3372,In_3373,In_3374,In_3375,In_3376,In_3377,In_3378,In_3379,In_3380,In_3381,In_3382,In_3383,In_3384,In_3385,In_3386,In_3387,In_3388,In_3389,In_3390,In_3391,In_3392,In_3393,In_3394,In_3395,In_3396,In_3397,In_3398,In_3399,In_3400,In_3401,In_3402,In_3403,In_3404,In_3405,In_3406,In_3407,In_3408,In_3409,In_3410,In_3411,In_3412,In_3413,In_3414,In_3415,In_3416,In_3417,In_3418,In_3419,In_3420,In_3421,In_3422,In_3423,In_3424,In_3425,In_3426,In_3427,In_3428,In_3429,In_3430,In_3431,In_3432,In_3433,In_3434,In_3435,In_3436,In_3437,In_3438,In_3439,In_3440,In_3441,In_3442,In_3443,In_3444,In_3445,In_3446,In_3447,In_3448,In_3449,In_3450,In_3451,In_3452,In_3453,In_3454,In_3455,In_3456,In_3457,In_3458,In_3459,In_3460,In_3461,In_3462,In_3463,In_3464,In_3465,In_3466,In_3467,In_3468,In_3469,In_3470,In_3471,In_3472,In_3473,In_3474,In_3475,In_3476,In_3477,In_3478,In_3479,In_3480,In_3481,In_3482,In_3483,In_3484,In_3485,In_3486,In_3487,In_3488,In_3489,In_3490,In_3491,In_3492,In_3493,In_3494,In_3495,In_3496,In_3497,In_3498,In_3499,In_3500,In_3501,In_3502,In_3503,In_3504,In_3505,In_3506,In_3507,In_3508,In_3509,In_3510,In_3511,In_3512,In_3513,In_3514,In_3515,In_3516,In_3517,In_3518,In_3519,In_3520,In_3521,In_3522,In_3523,In_3524,In_3525,In_3526,In_3527,In_3528,In_3529,In_3530,In_3531,In_3532,In_3533,In_3534,In_3535,In_3536,In_3537,In_3538,In_3539,In_3540,In_3541,In_3542,In_3543,In_3544,In_3545,In_3546,In_3547,In_3548,In_3549,In_3550,In_3551,In_3552,In_3553,In_3554,In_3555,In_3556,In_3557,In_3558,In_3559,In_3560,In_3561,In_3562,In_3563,In_3564,In_3565,In_3566,In_3567,In_3568,In_3569,In_3570,In_3571,In_3572,In_3573,In_3574,In_3575,In_3576,In_3577,In_3578,In_3579,In_3580,In_3581,In_3582,In_3583,In_3584,In_3585,In_3586,In_3587,In_3588,In_3589,In_3590,In_3591,In_3592,In_3593,In_3594,In_3595,In_3596,In_3597,In_3598,In_3599,In_3600,In_3601,In_3602,In_3603,In_3604,In_3605,In_3606,In_3607,In_3608,In_3609,In_3610,In_3611,In_3612,In_3613,In_3614,In_3615,In_3616,In_3617,In_3618,In_3619,In_3620,In_3621,In_3622,In_3623,In_3624,In_3625,In_3626,In_3627,In_3628,In_3629,In_3630,In_3631,In_3632,In_3633,In_3634,In_3635,In_3636,In_3637,In_3638,In_3639,In_3640,In_3641,In_3642,In_3643,In_3644,In_3645,In_3646,In_3647,In_3648,In_3649,In_3650,In_3651,In_3652,In_3653,In_3654,In_3655,In_3656,In_3657,In_3658,In_3659,In_3660,In_3661,In_3662,In_3663,In_3664,In_3665,In_3666,In_3667,In_3668,In_3669,In_3670,In_3671,In_3672,In_3673,In_3674,In_3675,In_3676,In_3677,In_3678,In_3679,In_3680,In_3681,In_3682,In_3683,In_3684,In_3685,In_3686,In_3687,In_3688,In_3689,In_3690,In_3691,In_3692,In_3693,In_3694,In_3695,In_3696,In_3697,In_3698,In_3699,In_3700,In_3701,In_3702,In_3703,In_3704,In_3705,In_3706,In_3707,In_3708,In_3709,In_3710,In_3711,In_3712,In_3713,In_3714,In_3715,In_3716,In_3717,In_3718,In_3719,In_3720,In_3721,In_3722,In_3723,In_3724,In_3725,In_3726,In_3727,In_3728,In_3729,In_3730,In_3731,In_3732,In_3733,In_3734,In_3735,In_3736,In_3737,In_3738,In_3739,In_3740,In_3741,In_3742,In_3743,In_3744,In_3745,In_3746,In_3747,In_3748,In_3749,In_3750,In_3751,In_3752,In_3753,In_3754,In_3755,In_3756,In_3757,In_3758,In_3759,In_3760,In_3761,In_3762,In_3763,In_3764,In_3765,In_3766,In_3767,In_3768,In_3769,In_3770,In_3771,In_3772,In_3773,In_3774,In_3775,In_3776,In_3777,In_3778,In_3779,In_3780,In_3781,In_3782,In_3783,In_3784,In_3785,In_3786,In_3787,In_3788,In_3789,In_3790,In_3791,In_3792,In_3793,In_3794,In_3795,In_3796,In_3797,In_3798,In_3799,In_3800,In_3801,In_3802,In_3803,In_3804,In_3805,In_3806,In_3807,In_3808,In_3809,In_3810,In_3811,In_3812,In_3813,In_3814,In_3815,In_3816,In_3817,In_3818,In_3819,In_3820,In_3821,In_3822,In_3823,In_3824,In_3825,In_3826,In_3827,In_3828,In_3829,In_3830,In_3831,In_3832,In_3833,In_3834,In_3835,In_3836,In_3837,In_3838,In_3839,In_3840,In_3841,In_3842,In_3843,In_3844,In_3845,In_3846,In_3847,In_3848,In_3849,In_3850,In_3851,In_3852,In_3853,In_3854,In_3855,In_3856,In_3857,In_3858,In_3859,In_3860,In_3861,In_3862,In_3863,In_3864,In_3865,In_3866,In_3867,In_3868,In_3869,In_3870,In_3871,In_3872,In_3873,In_3874,In_3875,In_3876,In_3877,In_3878,In_3879,In_3880,In_3881,In_3882,In_3883,In_3884,In_3885,In_3886,In_3887,In_3888,In_3889,In_3890,In_3891,In_3892,In_3893,In_3894,In_3895,In_3896,In_3897,In_3898,In_3899,In_3900,In_3901,In_3902,In_3903,In_3904,In_3905,In_3906,In_3907,In_3908,In_3909,In_3910,In_3911,In_3912,In_3913,In_3914,In_3915,In_3916,In_3917,In_3918,In_3919,In_3920,In_3921,In_3922,In_3923,In_3924,In_3925,In_3926,In_3927,In_3928,In_3929,In_3930,In_3931,In_3932,In_3933,In_3934,In_3935,In_3936,In_3937,In_3938,In_3939,In_3940,In_3941,In_3942,In_3943,In_3944,In_3945,In_3946,In_3947,In_3948,In_3949,In_3950,In_3951,In_3952,In_3953,In_3954,In_3955,In_3956,In_3957,In_3958,In_3959,In_3960,In_3961,In_3962,In_3963,In_3964,In_3965,In_3966,In_3967,In_3968,In_3969,In_3970,In_3971,In_3972,In_3973,In_3974,In_3975,In_3976,In_3977,In_3978,In_3979,In_3980,In_3981,In_3982,In_3983,In_3984,In_3985,In_3986,In_3987,In_3988,In_3989,In_3990,In_3991,In_3992,In_3993,In_3994,In_3995,In_3996,In_3997,In_3998,In_3999,In_4000,In_4001,In_4002,In_4003,In_4004,In_4005,In_4006,In_4007,In_4008,In_4009,In_4010,In_4011,In_4012,In_4013,In_4014,In_4015,In_4016,In_4017,In_4018,In_4019,In_4020,In_4021,In_4022,In_4023,In_4024,In_4025,In_4026,In_4027,In_4028,In_4029,In_4030,In_4031,In_4032,In_4033,In_4034,In_4035,In_4036,In_4037,In_4038,In_4039,In_4040,In_4041,In_4042,In_4043,In_4044,In_4045,In_4046,In_4047,In_4048,In_4049,In_4050,In_4051,In_4052,In_4053,In_4054,In_4055,In_4056,In_4057,In_4058,In_4059,In_4060,In_4061,In_4062,In_4063,In_4064,In_4065,In_4066,In_4067,In_4068,In_4069,In_4070,In_4071,In_4072,In_4073,In_4074,In_4075,In_4076,In_4077,In_4078,In_4079,In_4080,In_4081,In_4082,In_4083,In_4084,In_4085,In_4086,In_4087,In_4088,In_4089,In_4090,In_4091,In_4092,In_4093,In_4094,In_4095,In_4096,In_4097,In_4098,In_4099,In_4100,In_4101,In_4102,In_4103,In_4104,In_4105,In_4106,In_4107,In_4108,In_4109,In_4110,In_4111,In_4112,In_4113,In_4114,In_4115,In_4116,In_4117,In_4118,In_4119,In_4120,In_4121,In_4122,In_4123,In_4124,In_4125,In_4126,In_4127,In_4128,In_4129,In_4130,In_4131,In_4132,In_4133,In_4134,In_4135,In_4136,In_4137,In_4138,In_4139,In_4140,In_4141,In_4142,In_4143,In_4144,In_4145,In_4146,In_4147,In_4148,In_4149,In_4150,In_4151,In_4152,In_4153,In_4154,In_4155,In_4156,In_4157,In_4158,In_4159,In_4160,In_4161,In_4162,In_4163,In_4164,In_4165,In_4166,In_4167,In_4168,In_4169,In_4170,In_4171,In_4172,In_4173,In_4174,In_4175,In_4176,In_4177,In_4178,In_4179,In_4180,In_4181,In_4182,In_4183,In_4184,In_4185,In_4186,In_4187,In_4188,In_4189,In_4190,In_4191,In_4192,In_4193,In_4194,In_4195,In_4196,In_4197,In_4198,In_4199,In_4200,In_4201,In_4202,In_4203,In_4204,In_4205,In_4206,In_4207,In_4208,In_4209,In_4210,In_4211,In_4212,In_4213,In_4214,In_4215,In_4216,In_4217,In_4218,In_4219,In_4220,In_4221,In_4222,In_4223,In_4224,In_4225,In_4226,In_4227,In_4228,In_4229,In_4230,In_4231,In_4232,In_4233,In_4234,In_4235,In_4236,In_4237,In_4238,In_4239,In_4240,In_4241,In_4242,In_4243,In_4244,In_4245,In_4246,In_4247,In_4248,In_4249,In_4250,In_4251,In_4252,In_4253,In_4254,In_4255,In_4256,In_4257,In_4258,In_4259,In_4260,In_4261,In_4262,In_4263,In_4264,In_4265,In_4266,In_4267,In_4268,In_4269,In_4270,In_4271,In_4272,In_4273,In_4274,In_4275,In_4276,In_4277,In_4278,In_4279,In_4280,In_4281,In_4282,In_4283,In_4284,In_4285,In_4286,In_4287,In_4288,In_4289,In_4290,In_4291,In_4292,In_4293,In_4294,In_4295,In_4296,In_4297,In_4298,In_4299,In_4300,In_4301,In_4302,In_4303,In_4304,In_4305,In_4306,In_4307,In_4308,In_4309,In_4310,In_4311,In_4312,In_4313,In_4314,In_4315,In_4316,In_4317,In_4318,In_4319,In_4320,In_4321,In_4322,In_4323,In_4324,In_4325,In_4326,In_4327,In_4328,In_4329,In_4330,In_4331,In_4332,In_4333,In_4334,In_4335,In_4336,In_4337,In_4338,In_4339,In_4340,In_4341,In_4342,In_4343,In_4344,In_4345,In_4346,In_4347,In_4348,In_4349,In_4350,In_4351,In_4352,In_4353,In_4354,In_4355,In_4356,In_4357,In_4358,In_4359,In_4360,In_4361,In_4362,In_4363,In_4364,In_4365,In_4366,In_4367,In_4368,In_4369,In_4370,In_4371,In_4372,In_4373,In_4374,In_4375,In_4376,In_4377,In_4378,In_4379,In_4380,In_4381,In_4382,In_4383,In_4384,In_4385,In_4386,In_4387,In_4388,In_4389,In_4390,In_4391,In_4392,In_4393,In_4394,In_4395,In_4396,In_4397,In_4398,In_4399,In_4400,In_4401,In_4402,In_4403,In_4404,In_4405,In_4406,In_4407,In_4408,In_4409,In_4410,In_4411,In_4412,In_4413,In_4414,In_4415,In_4416,In_4417,In_4418,In_4419,In_4420,In_4421,In_4422,In_4423,In_4424,In_4425,In_4426,In_4427,In_4428,In_4429,In_4430,In_4431,In_4432,In_4433,In_4434,In_4435,In_4436,In_4437,In_4438,In_4439,In_4440,In_4441,In_4442,In_4443,In_4444,In_4445,In_4446,In_4447,In_4448,In_4449,In_4450,In_4451,In_4452,In_4453,In_4454,In_4455,In_4456,In_4457,In_4458,In_4459,In_4460,In_4461,In_4462,In_4463,In_4464,In_4465,In_4466,In_4467,In_4468,In_4469,In_4470,In_4471,In_4472,In_4473,In_4474,In_4475,In_4476,In_4477,In_4478,In_4479,In_4480,In_4481,In_4482,In_4483,In_4484,In_4485,In_4486,In_4487,In_4488,In_4489,In_4490,In_4491,In_4492,In_4493,In_4494,In_4495,In_4496,In_4497,In_4498,In_4499,In_4500,In_4501,In_4502,In_4503,In_4504,In_4505,In_4506,In_4507,In_4508,In_4509,In_4510,In_4511,In_4512,In_4513,In_4514,In_4515,In_4516,In_4517,In_4518,In_4519,In_4520,In_4521,In_4522,In_4523,In_4524,In_4525,In_4526,In_4527,In_4528,In_4529,In_4530,In_4531,In_4532,In_4533,In_4534,In_4535,In_4536,In_4537,In_4538,In_4539,In_4540,In_4541,In_4542,In_4543,In_4544,In_4545,In_4546,In_4547,In_4548,In_4549,In_4550,In_4551,In_4552,In_4553,In_4554,In_4555,In_4556,In_4557,In_4558,In_4559,In_4560,In_4561,In_4562,In_4563,In_4564,In_4565,In_4566,In_4567,In_4568,In_4569,In_4570,In_4571,In_4572,In_4573,In_4574,In_4575,In_4576,In_4577,In_4578,In_4579,In_4580,In_4581,In_4582,In_4583,In_4584,In_4585,In_4586,In_4587,In_4588,In_4589,In_4590,In_4591,In_4592,In_4593,In_4594,In_4595,In_4596,In_4597,In_4598,In_4599,In_4600,In_4601,In_4602,In_4603,In_4604,In_4605,In_4606,In_4607,In_4608,In_4609,In_4610,In_4611,In_4612,In_4613,In_4614,In_4615,In_4616,In_4617,In_4618,In_4619,In_4620,In_4621,In_4622,In_4623,In_4624,In_4625,In_4626,In_4627,In_4628,In_4629,In_4630,In_4631,In_4632,In_4633,In_4634,In_4635,In_4636,In_4637,In_4638,In_4639,In_4640,In_4641,In_4642,In_4643,In_4644,In_4645,In_4646,In_4647,In_4648,In_4649,In_4650,In_4651,In_4652,In_4653,In_4654,In_4655,In_4656,In_4657,In_4658,In_4659,In_4660,In_4661,In_4662,In_4663,In_4664,In_4665,In_4666,In_4667,In_4668,In_4669,In_4670,In_4671,In_4672,In_4673,In_4674,In_4675,In_4676,In_4677,In_4678,In_4679,In_4680,In_4681,In_4682,In_4683,In_4684,In_4685,In_4686,In_4687,In_4688,In_4689,In_4690,In_4691,In_4692,In_4693,In_4694,In_4695,In_4696,In_4697,In_4698,In_4699,In_4700,In_4701,In_4702,In_4703,In_4704,In_4705,In_4706,In_4707,In_4708,In_4709,In_4710,In_4711,In_4712,In_4713,In_4714,In_4715,In_4716,In_4717,In_4718,In_4719,In_4720,In_4721,In_4722,In_4723,In_4724,In_4725,In_4726,In_4727,In_4728,In_4729,In_4730,In_4731,In_4732,In_4733,In_4734,In_4735,In_4736,In_4737,In_4738,In_4739,In_4740,In_4741,In_4742,In_4743,In_4744,In_4745,In_4746,In_4747,In_4748,In_4749,In_4750,In_4751,In_4752,In_4753,In_4754,In_4755,In_4756,In_4757,In_4758,In_4759,In_4760,In_4761,In_4762,In_4763,In_4764,In_4765,In_4766,In_4767,In_4768,In_4769,In_4770,In_4771,In_4772,In_4773,In_4774,In_4775,In_4776,In_4777,In_4778,In_4779,In_4780,In_4781,In_4782,In_4783,In_4784,In_4785,In_4786,In_4787,In_4788,In_4789,In_4790,In_4791,In_4792,In_4793,In_4794,In_4795,In_4796,In_4797,In_4798,In_4799,In_4800,In_4801,In_4802,In_4803,In_4804,In_4805,In_4806,In_4807,In_4808,In_4809,In_4810,In_4811,In_4812,In_4813,In_4814,In_4815,In_4816,In_4817,In_4818,In_4819,In_4820,In_4821,In_4822,In_4823,In_4824,In_4825,In_4826,In_4827,In_4828,In_4829,In_4830,In_4831,In_4832,In_4833,In_4834,In_4835,In_4836,In_4837,In_4838,In_4839,In_4840,In_4841,In_4842,In_4843,In_4844,In_4845,In_4846,In_4847,In_4848,In_4849,In_4850,In_4851,In_4852,In_4853,In_4854,In_4855,In_4856,In_4857,In_4858,In_4859,In_4860,In_4861,In_4862,In_4863,In_4864,In_4865,In_4866,In_4867,In_4868,In_4869,In_4870,In_4871,In_4872,In_4873,In_4874,In_4875,In_4876,In_4877,In_4878,In_4879,In_4880,In_4881,In_4882,In_4883,In_4884,In_4885,In_4886,In_4887,In_4888,In_4889,In_4890,In_4891,In_4892,In_4893,In_4894,In_4895,In_4896,In_4897,In_4898,In_4899,In_4900,In_4901,In_4902,In_4903,In_4904,In_4905,In_4906,In_4907,In_4908,In_4909,In_4910,In_4911,In_4912,In_4913,In_4914,In_4915,In_4916,In_4917,In_4918,In_4919,In_4920,In_4921,In_4922,In_4923,In_4924,In_4925,In_4926,In_4927,In_4928,In_4929,In_4930,In_4931,In_4932,In_4933,In_4934,In_4935,In_4936,In_4937,In_4938,In_4939,In_4940,In_4941,In_4942,In_4943,In_4944,In_4945,In_4946,In_4947,In_4948,In_4949,In_4950,In_4951,In_4952,In_4953,In_4954,In_4955,In_4956,In_4957,In_4958,In_4959,In_4960,In_4961,In_4962,In_4963,In_4964,In_4965,In_4966,In_4967,In_4968,In_4969,In_4970,In_4971,In_4972,In_4973,In_4974,In_4975,In_4976,In_4977,In_4978,In_4979,In_4980,In_4981,In_4982,In_4983,In_4984,In_4985,In_4986,In_4987,In_4988,In_4989,In_4990,In_4991,In_4992,In_4993,In_4994,In_4995,In_4996,In_4997,In_4998,In_4999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499,O_3500,O_3501,O_3502,O_3503,O_3504,O_3505,O_3506,O_3507,O_3508,O_3509,O_3510,O_3511,O_3512,O_3513,O_3514,O_3515,O_3516,O_3517,O_3518,O_3519,O_3520,O_3521,O_3522,O_3523,O_3524,O_3525,O_3526,O_3527,O_3528,O_3529,O_3530,O_3531,O_3532,O_3533,O_3534,O_3535,O_3536,O_3537,O_3538,O_3539,O_3540,O_3541,O_3542,O_3543,O_3544,O_3545,O_3546,O_3547,O_3548,O_3549,O_3550,O_3551,O_3552,O_3553,O_3554,O_3555,O_3556,O_3557,O_3558,O_3559,O_3560,O_3561,O_3562,O_3563,O_3564,O_3565,O_3566,O_3567,O_3568,O_3569,O_3570,O_3571,O_3572,O_3573,O_3574,O_3575,O_3576,O_3577,O_3578,O_3579,O_3580,O_3581,O_3582,O_3583,O_3584,O_3585,O_3586,O_3587,O_3588,O_3589,O_3590,O_3591,O_3592,O_3593,O_3594,O_3595,O_3596,O_3597,O_3598,O_3599,O_3600,O_3601,O_3602,O_3603,O_3604,O_3605,O_3606,O_3607,O_3608,O_3609,O_3610,O_3611,O_3612,O_3613,O_3614,O_3615,O_3616,O_3617,O_3618,O_3619,O_3620,O_3621,O_3622,O_3623,O_3624,O_3625,O_3626,O_3627,O_3628,O_3629,O_3630,O_3631,O_3632,O_3633,O_3634,O_3635,O_3636,O_3637,O_3638,O_3639,O_3640,O_3641,O_3642,O_3643,O_3644,O_3645,O_3646,O_3647,O_3648,O_3649,O_3650,O_3651,O_3652,O_3653,O_3654,O_3655,O_3656,O_3657,O_3658,O_3659,O_3660,O_3661,O_3662,O_3663,O_3664,O_3665,O_3666,O_3667,O_3668,O_3669,O_3670,O_3671,O_3672,O_3673,O_3674,O_3675,O_3676,O_3677,O_3678,O_3679,O_3680,O_3681,O_3682,O_3683,O_3684,O_3685,O_3686,O_3687,O_3688,O_3689,O_3690,O_3691,O_3692,O_3693,O_3694,O_3695,O_3696,O_3697,O_3698,O_3699,O_3700,O_3701,O_3702,O_3703,O_3704,O_3705,O_3706,O_3707,O_3708,O_3709,O_3710,O_3711,O_3712,O_3713,O_3714,O_3715,O_3716,O_3717,O_3718,O_3719,O_3720,O_3721,O_3722,O_3723,O_3724,O_3725,O_3726,O_3727,O_3728,O_3729,O_3730,O_3731,O_3732,O_3733,O_3734,O_3735,O_3736,O_3737,O_3738,O_3739,O_3740,O_3741,O_3742,O_3743,O_3744,O_3745,O_3746,O_3747,O_3748,O_3749,O_3750,O_3751,O_3752,O_3753,O_3754,O_3755,O_3756,O_3757,O_3758,O_3759,O_3760,O_3761,O_3762,O_3763,O_3764,O_3765,O_3766,O_3767,O_3768,O_3769,O_3770,O_3771,O_3772,O_3773,O_3774,O_3775,O_3776,O_3777,O_3778,O_3779,O_3780,O_3781,O_3782,O_3783,O_3784,O_3785,O_3786,O_3787,O_3788,O_3789,O_3790,O_3791,O_3792,O_3793,O_3794,O_3795,O_3796,O_3797,O_3798,O_3799,O_3800,O_3801,O_3802,O_3803,O_3804,O_3805,O_3806,O_3807,O_3808,O_3809,O_3810,O_3811,O_3812,O_3813,O_3814,O_3815,O_3816,O_3817,O_3818,O_3819,O_3820,O_3821,O_3822,O_3823,O_3824,O_3825,O_3826,O_3827,O_3828,O_3829,O_3830,O_3831,O_3832,O_3833,O_3834,O_3835,O_3836,O_3837,O_3838,O_3839,O_3840,O_3841,O_3842,O_3843,O_3844,O_3845,O_3846,O_3847,O_3848,O_3849,O_3850,O_3851,O_3852,O_3853,O_3854,O_3855,O_3856,O_3857,O_3858,O_3859,O_3860,O_3861,O_3862,O_3863,O_3864,O_3865,O_3866,O_3867,O_3868,O_3869,O_3870,O_3871,O_3872,O_3873,O_3874,O_3875,O_3876,O_3877,O_3878,O_3879,O_3880,O_3881,O_3882,O_3883,O_3884,O_3885,O_3886,O_3887,O_3888,O_3889,O_3890,O_3891,O_3892,O_3893,O_3894,O_3895,O_3896,O_3897,O_3898,O_3899,O_3900,O_3901,O_3902,O_3903,O_3904,O_3905,O_3906,O_3907,O_3908,O_3909,O_3910,O_3911,O_3912,O_3913,O_3914,O_3915,O_3916,O_3917,O_3918,O_3919,O_3920,O_3921,O_3922,O_3923,O_3924,O_3925,O_3926,O_3927,O_3928,O_3929,O_3930,O_3931,O_3932,O_3933,O_3934,O_3935,O_3936,O_3937,O_3938,O_3939,O_3940,O_3941,O_3942,O_3943,O_3944,O_3945,O_3946,O_3947,O_3948,O_3949,O_3950,O_3951,O_3952,O_3953,O_3954,O_3955,O_3956,O_3957,O_3958,O_3959,O_3960,O_3961,O_3962,O_3963,O_3964,O_3965,O_3966,O_3967,O_3968,O_3969,O_3970,O_3971,O_3972,O_3973,O_3974,O_3975,O_3976,O_3977,O_3978,O_3979,O_3980,O_3981,O_3982,O_3983,O_3984,O_3985,O_3986,O_3987,O_3988,O_3989,O_3990,O_3991,O_3992,O_3993,O_3994,O_3995,O_3996,O_3997,O_3998,O_3999,O_4000,O_4001,O_4002,O_4003,O_4004,O_4005,O_4006,O_4007,O_4008,O_4009,O_4010,O_4011,O_4012,O_4013,O_4014,O_4015,O_4016,O_4017,O_4018,O_4019,O_4020,O_4021,O_4022,O_4023,O_4024,O_4025,O_4026,O_4027,O_4028,O_4029,O_4030,O_4031,O_4032,O_4033,O_4034,O_4035,O_4036,O_4037,O_4038,O_4039,O_4040,O_4041,O_4042,O_4043,O_4044,O_4045,O_4046,O_4047,O_4048,O_4049,O_4050,O_4051,O_4052,O_4053,O_4054,O_4055,O_4056,O_4057,O_4058,O_4059,O_4060,O_4061,O_4062,O_4063,O_4064,O_4065,O_4066,O_4067,O_4068,O_4069,O_4070,O_4071,O_4072,O_4073,O_4074,O_4075,O_4076,O_4077,O_4078,O_4079,O_4080,O_4081,O_4082,O_4083,O_4084,O_4085,O_4086,O_4087,O_4088,O_4089,O_4090,O_4091,O_4092,O_4093,O_4094,O_4095,O_4096,O_4097,O_4098,O_4099,O_4100,O_4101,O_4102,O_4103,O_4104,O_4105,O_4106,O_4107,O_4108,O_4109,O_4110,O_4111,O_4112,O_4113,O_4114,O_4115,O_4116,O_4117,O_4118,O_4119,O_4120,O_4121,O_4122,O_4123,O_4124,O_4125,O_4126,O_4127,O_4128,O_4129,O_4130,O_4131,O_4132,O_4133,O_4134,O_4135,O_4136,O_4137,O_4138,O_4139,O_4140,O_4141,O_4142,O_4143,O_4144,O_4145,O_4146,O_4147,O_4148,O_4149,O_4150,O_4151,O_4152,O_4153,O_4154,O_4155,O_4156,O_4157,O_4158,O_4159,O_4160,O_4161,O_4162,O_4163,O_4164,O_4165,O_4166,O_4167,O_4168,O_4169,O_4170,O_4171,O_4172,O_4173,O_4174,O_4175,O_4176,O_4177,O_4178,O_4179,O_4180,O_4181,O_4182,O_4183,O_4184,O_4185,O_4186,O_4187,O_4188,O_4189,O_4190,O_4191,O_4192,O_4193,O_4194,O_4195,O_4196,O_4197,O_4198,O_4199,O_4200,O_4201,O_4202,O_4203,O_4204,O_4205,O_4206,O_4207,O_4208,O_4209,O_4210,O_4211,O_4212,O_4213,O_4214,O_4215,O_4216,O_4217,O_4218,O_4219,O_4220,O_4221,O_4222,O_4223,O_4224,O_4225,O_4226,O_4227,O_4228,O_4229,O_4230,O_4231,O_4232,O_4233,O_4234,O_4235,O_4236,O_4237,O_4238,O_4239,O_4240,O_4241,O_4242,O_4243,O_4244,O_4245,O_4246,O_4247,O_4248,O_4249,O_4250,O_4251,O_4252,O_4253,O_4254,O_4255,O_4256,O_4257,O_4258,O_4259,O_4260,O_4261,O_4262,O_4263,O_4264,O_4265,O_4266,O_4267,O_4268,O_4269,O_4270,O_4271,O_4272,O_4273,O_4274,O_4275,O_4276,O_4277,O_4278,O_4279,O_4280,O_4281,O_4282,O_4283,O_4284,O_4285,O_4286,O_4287,O_4288,O_4289,O_4290,O_4291,O_4292,O_4293,O_4294,O_4295,O_4296,O_4297,O_4298,O_4299,O_4300,O_4301,O_4302,O_4303,O_4304,O_4305,O_4306,O_4307,O_4308,O_4309,O_4310,O_4311,O_4312,O_4313,O_4314,O_4315,O_4316,O_4317,O_4318,O_4319,O_4320,O_4321,O_4322,O_4323,O_4324,O_4325,O_4326,O_4327,O_4328,O_4329,O_4330,O_4331,O_4332,O_4333,O_4334,O_4335,O_4336,O_4337,O_4338,O_4339,O_4340,O_4341,O_4342,O_4343,O_4344,O_4345,O_4346,O_4347,O_4348,O_4349,O_4350,O_4351,O_4352,O_4353,O_4354,O_4355,O_4356,O_4357,O_4358,O_4359,O_4360,O_4361,O_4362,O_4363,O_4364,O_4365,O_4366,O_4367,O_4368,O_4369,O_4370,O_4371,O_4372,O_4373,O_4374,O_4375,O_4376,O_4377,O_4378,O_4379,O_4380,O_4381,O_4382,O_4383,O_4384,O_4385,O_4386,O_4387,O_4388,O_4389,O_4390,O_4391,O_4392,O_4393,O_4394,O_4395,O_4396,O_4397,O_4398,O_4399,O_4400,O_4401,O_4402,O_4403,O_4404,O_4405,O_4406,O_4407,O_4408,O_4409,O_4410,O_4411,O_4412,O_4413,O_4414,O_4415,O_4416,O_4417,O_4418,O_4419,O_4420,O_4421,O_4422,O_4423,O_4424,O_4425,O_4426,O_4427,O_4428,O_4429,O_4430,O_4431,O_4432,O_4433,O_4434,O_4435,O_4436,O_4437,O_4438,O_4439,O_4440,O_4441,O_4442,O_4443,O_4444,O_4445,O_4446,O_4447,O_4448,O_4449,O_4450,O_4451,O_4452,O_4453,O_4454,O_4455,O_4456,O_4457,O_4458,O_4459,O_4460,O_4461,O_4462,O_4463,O_4464,O_4465,O_4466,O_4467,O_4468,O_4469,O_4470,O_4471,O_4472,O_4473,O_4474,O_4475,O_4476,O_4477,O_4478,O_4479,O_4480,O_4481,O_4482,O_4483,O_4484,O_4485,O_4486,O_4487,O_4488,O_4489,O_4490,O_4491,O_4492,O_4493,O_4494,O_4495,O_4496,O_4497,O_4498,O_4499,O_4500,O_4501,O_4502,O_4503,O_4504,O_4505,O_4506,O_4507,O_4508,O_4509,O_4510,O_4511,O_4512,O_4513,O_4514,O_4515,O_4516,O_4517,O_4518,O_4519,O_4520,O_4521,O_4522,O_4523,O_4524,O_4525,O_4526,O_4527,O_4528,O_4529,O_4530,O_4531,O_4532,O_4533,O_4534,O_4535,O_4536,O_4537,O_4538,O_4539,O_4540,O_4541,O_4542,O_4543,O_4544,O_4545,O_4546,O_4547,O_4548,O_4549,O_4550,O_4551,O_4552,O_4553,O_4554,O_4555,O_4556,O_4557,O_4558,O_4559,O_4560,O_4561,O_4562,O_4563,O_4564,O_4565,O_4566,O_4567,O_4568,O_4569,O_4570,O_4571,O_4572,O_4573,O_4574,O_4575,O_4576,O_4577,O_4578,O_4579,O_4580,O_4581,O_4582,O_4583,O_4584,O_4585,O_4586,O_4587,O_4588,O_4589,O_4590,O_4591,O_4592,O_4593,O_4594,O_4595,O_4596,O_4597,O_4598,O_4599,O_4600,O_4601,O_4602,O_4603,O_4604,O_4605,O_4606,O_4607,O_4608,O_4609,O_4610,O_4611,O_4612,O_4613,O_4614,O_4615,O_4616,O_4617,O_4618,O_4619,O_4620,O_4621,O_4622,O_4623,O_4624,O_4625,O_4626,O_4627,O_4628,O_4629,O_4630,O_4631,O_4632,O_4633,O_4634,O_4635,O_4636,O_4637,O_4638,O_4639,O_4640,O_4641,O_4642,O_4643,O_4644,O_4645,O_4646,O_4647,O_4648,O_4649,O_4650,O_4651,O_4652,O_4653,O_4654,O_4655,O_4656,O_4657,O_4658,O_4659,O_4660,O_4661,O_4662,O_4663,O_4664,O_4665,O_4666,O_4667,O_4668,O_4669,O_4670,O_4671,O_4672,O_4673,O_4674,O_4675,O_4676,O_4677,O_4678,O_4679,O_4680,O_4681,O_4682,O_4683,O_4684,O_4685,O_4686,O_4687,O_4688,O_4689,O_4690,O_4691,O_4692,O_4693,O_4694,O_4695,O_4696,O_4697,O_4698,O_4699,O_4700,O_4701,O_4702,O_4703,O_4704,O_4705,O_4706,O_4707,O_4708,O_4709,O_4710,O_4711,O_4712,O_4713,O_4714,O_4715,O_4716,O_4717,O_4718,O_4719,O_4720,O_4721,O_4722,O_4723,O_4724,O_4725,O_4726,O_4727,O_4728,O_4729,O_4730,O_4731,O_4732,O_4733,O_4734,O_4735,O_4736,O_4737,O_4738,O_4739,O_4740,O_4741,O_4742,O_4743,O_4744,O_4745,O_4746,O_4747,O_4748,O_4749,O_4750,O_4751,O_4752,O_4753,O_4754,O_4755,O_4756,O_4757,O_4758,O_4759,O_4760,O_4761,O_4762,O_4763,O_4764,O_4765,O_4766,O_4767,O_4768,O_4769,O_4770,O_4771,O_4772,O_4773,O_4774,O_4775,O_4776,O_4777,O_4778,O_4779,O_4780,O_4781,O_4782,O_4783,O_4784,O_4785,O_4786,O_4787,O_4788,O_4789,O_4790,O_4791,O_4792,O_4793,O_4794,O_4795,O_4796,O_4797,O_4798,O_4799,O_4800,O_4801,O_4802,O_4803,O_4804,O_4805,O_4806,O_4807,O_4808,O_4809,O_4810,O_4811,O_4812,O_4813,O_4814,O_4815,O_4816,O_4817,O_4818,O_4819,O_4820,O_4821,O_4822,O_4823,O_4824,O_4825,O_4826,O_4827,O_4828,O_4829,O_4830,O_4831,O_4832,O_4833,O_4834,O_4835,O_4836,O_4837,O_4838,O_4839,O_4840,O_4841,O_4842,O_4843,O_4844,O_4845,O_4846,O_4847,O_4848,O_4849,O_4850,O_4851,O_4852,O_4853,O_4854,O_4855,O_4856,O_4857,O_4858,O_4859,O_4860,O_4861,O_4862,O_4863,O_4864,O_4865,O_4866,O_4867,O_4868,O_4869,O_4870,O_4871,O_4872,O_4873,O_4874,O_4875,O_4876,O_4877,O_4878,O_4879,O_4880,O_4881,O_4882,O_4883,O_4884,O_4885,O_4886,O_4887,O_4888,O_4889,O_4890,O_4891,O_4892,O_4893,O_4894,O_4895,O_4896,O_4897,O_4898,O_4899,O_4900,O_4901,O_4902,O_4903,O_4904,O_4905,O_4906,O_4907,O_4908,O_4909,O_4910,O_4911,O_4912,O_4913,O_4914,O_4915,O_4916,O_4917,O_4918,O_4919,O_4920,O_4921,O_4922,O_4923,O_4924,O_4925,O_4926,O_4927,O_4928,O_4929,O_4930,O_4931,O_4932,O_4933,O_4934,O_4935,O_4936,O_4937,O_4938,O_4939,O_4940,O_4941,O_4942,O_4943,O_4944,O_4945,O_4946,O_4947,O_4948,O_4949,O_4950,O_4951,O_4952,O_4953,O_4954,O_4955,O_4956,O_4957,O_4958,O_4959,O_4960,O_4961,O_4962,O_4963,O_4964,O_4965,O_4966,O_4967,O_4968,O_4969,O_4970,O_4971,O_4972,O_4973,O_4974,O_4975,O_4976,O_4977,O_4978,O_4979,O_4980,O_4981,O_4982,O_4983,O_4984,O_4985,O_4986,O_4987,O_4988,O_4989,O_4990,O_4991,O_4992,O_4993,O_4994,O_4995,O_4996,O_4997,O_4998,O_4999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999,N_30000,N_30001,N_30002,N_30003,N_30004,N_30005,N_30006,N_30007,N_30008,N_30009,N_30010,N_30011,N_30012,N_30013,N_30014,N_30015,N_30016,N_30017,N_30018,N_30019,N_30020,N_30021,N_30022,N_30023,N_30024,N_30025,N_30026,N_30027,N_30028,N_30029,N_30030,N_30031,N_30032,N_30033,N_30034,N_30035,N_30036,N_30037,N_30038,N_30039,N_30040,N_30041,N_30042,N_30043,N_30044,N_30045,N_30046,N_30047,N_30048,N_30049,N_30050,N_30051,N_30052,N_30053,N_30054,N_30055,N_30056,N_30057,N_30058,N_30059,N_30060,N_30061,N_30062,N_30063,N_30064,N_30065,N_30066,N_30067,N_30068,N_30069,N_30070,N_30071,N_30072,N_30073,N_30074,N_30075,N_30076,N_30077,N_30078,N_30079,N_30080,N_30081,N_30082,N_30083,N_30084,N_30085,N_30086,N_30087,N_30088,N_30089,N_30090,N_30091,N_30092,N_30093,N_30094,N_30095,N_30096,N_30097,N_30098,N_30099,N_30100,N_30101,N_30102,N_30103,N_30104,N_30105,N_30106,N_30107,N_30108,N_30109,N_30110,N_30111,N_30112,N_30113,N_30114,N_30115,N_30116,N_30117,N_30118,N_30119,N_30120,N_30121,N_30122,N_30123,N_30124,N_30125,N_30126,N_30127,N_30128,N_30129,N_30130,N_30131,N_30132,N_30133,N_30134,N_30135,N_30136,N_30137,N_30138,N_30139,N_30140,N_30141,N_30142,N_30143,N_30144,N_30145,N_30146,N_30147,N_30148,N_30149,N_30150,N_30151,N_30152,N_30153,N_30154,N_30155,N_30156,N_30157,N_30158,N_30159,N_30160,N_30161,N_30162,N_30163,N_30164,N_30165,N_30166,N_30167,N_30168,N_30169,N_30170,N_30171,N_30172,N_30173,N_30174,N_30175,N_30176,N_30177,N_30178,N_30179,N_30180,N_30181,N_30182,N_30183,N_30184,N_30185,N_30186,N_30187,N_30188,N_30189,N_30190,N_30191,N_30192,N_30193,N_30194,N_30195,N_30196,N_30197,N_30198,N_30199,N_30200,N_30201,N_30202,N_30203,N_30204,N_30205,N_30206,N_30207,N_30208,N_30209,N_30210,N_30211,N_30212,N_30213,N_30214,N_30215,N_30216,N_30217,N_30218,N_30219,N_30220,N_30221,N_30222,N_30223,N_30224,N_30225,N_30226,N_30227,N_30228,N_30229,N_30230,N_30231,N_30232,N_30233,N_30234,N_30235,N_30236,N_30237,N_30238,N_30239,N_30240,N_30241,N_30242,N_30243,N_30244,N_30245,N_30246,N_30247,N_30248,N_30249,N_30250,N_30251,N_30252,N_30253,N_30254,N_30255,N_30256,N_30257,N_30258,N_30259,N_30260,N_30261,N_30262,N_30263,N_30264,N_30265,N_30266,N_30267,N_30268,N_30269,N_30270,N_30271,N_30272,N_30273,N_30274,N_30275,N_30276,N_30277,N_30278,N_30279,N_30280,N_30281,N_30282,N_30283,N_30284,N_30285,N_30286,N_30287,N_30288,N_30289,N_30290,N_30291,N_30292,N_30293,N_30294,N_30295,N_30296,N_30297,N_30298,N_30299,N_30300,N_30301,N_30302,N_30303,N_30304,N_30305,N_30306,N_30307,N_30308,N_30309,N_30310,N_30311,N_30312,N_30313,N_30314,N_30315,N_30316,N_30317,N_30318,N_30319,N_30320,N_30321,N_30322,N_30323,N_30324,N_30325,N_30326,N_30327,N_30328,N_30329,N_30330,N_30331,N_30332,N_30333,N_30334,N_30335,N_30336,N_30337,N_30338,N_30339,N_30340,N_30341,N_30342,N_30343,N_30344,N_30345,N_30346,N_30347,N_30348,N_30349,N_30350,N_30351,N_30352,N_30353,N_30354,N_30355,N_30356,N_30357,N_30358,N_30359,N_30360,N_30361,N_30362,N_30363,N_30364,N_30365,N_30366,N_30367,N_30368,N_30369,N_30370,N_30371,N_30372,N_30373,N_30374,N_30375,N_30376,N_30377,N_30378,N_30379,N_30380,N_30381,N_30382,N_30383,N_30384,N_30385,N_30386,N_30387,N_30388,N_30389,N_30390,N_30391,N_30392,N_30393,N_30394,N_30395,N_30396,N_30397,N_30398,N_30399,N_30400,N_30401,N_30402,N_30403,N_30404,N_30405,N_30406,N_30407,N_30408,N_30409,N_30410,N_30411,N_30412,N_30413,N_30414,N_30415,N_30416,N_30417,N_30418,N_30419,N_30420,N_30421,N_30422,N_30423,N_30424,N_30425,N_30426,N_30427,N_30428,N_30429,N_30430,N_30431,N_30432,N_30433,N_30434,N_30435,N_30436,N_30437,N_30438,N_30439,N_30440,N_30441,N_30442,N_30443,N_30444,N_30445,N_30446,N_30447,N_30448,N_30449,N_30450,N_30451,N_30452,N_30453,N_30454,N_30455,N_30456,N_30457,N_30458,N_30459,N_30460,N_30461,N_30462,N_30463,N_30464,N_30465,N_30466,N_30467,N_30468,N_30469,N_30470,N_30471,N_30472,N_30473,N_30474,N_30475,N_30476,N_30477,N_30478,N_30479,N_30480,N_30481,N_30482,N_30483,N_30484,N_30485,N_30486,N_30487,N_30488,N_30489,N_30490,N_30491,N_30492,N_30493,N_30494,N_30495,N_30496,N_30497,N_30498,N_30499,N_30500,N_30501,N_30502,N_30503,N_30504,N_30505,N_30506,N_30507,N_30508,N_30509,N_30510,N_30511,N_30512,N_30513,N_30514,N_30515,N_30516,N_30517,N_30518,N_30519,N_30520,N_30521,N_30522,N_30523,N_30524,N_30525,N_30526,N_30527,N_30528,N_30529,N_30530,N_30531,N_30532,N_30533,N_30534,N_30535,N_30536,N_30537,N_30538,N_30539,N_30540,N_30541,N_30542,N_30543,N_30544,N_30545,N_30546,N_30547,N_30548,N_30549,N_30550,N_30551,N_30552,N_30553,N_30554,N_30555,N_30556,N_30557,N_30558,N_30559,N_30560,N_30561,N_30562,N_30563,N_30564,N_30565,N_30566,N_30567,N_30568,N_30569,N_30570,N_30571,N_30572,N_30573,N_30574,N_30575,N_30576,N_30577,N_30578,N_30579,N_30580,N_30581,N_30582,N_30583,N_30584,N_30585,N_30586,N_30587,N_30588,N_30589,N_30590,N_30591,N_30592,N_30593,N_30594,N_30595,N_30596,N_30597,N_30598,N_30599,N_30600,N_30601,N_30602,N_30603,N_30604,N_30605,N_30606,N_30607,N_30608,N_30609,N_30610,N_30611,N_30612,N_30613,N_30614,N_30615,N_30616,N_30617,N_30618,N_30619,N_30620,N_30621,N_30622,N_30623,N_30624,N_30625,N_30626,N_30627,N_30628,N_30629,N_30630,N_30631,N_30632,N_30633,N_30634,N_30635,N_30636,N_30637,N_30638,N_30639,N_30640,N_30641,N_30642,N_30643,N_30644,N_30645,N_30646,N_30647,N_30648,N_30649,N_30650,N_30651,N_30652,N_30653,N_30654,N_30655,N_30656,N_30657,N_30658,N_30659,N_30660,N_30661,N_30662,N_30663,N_30664,N_30665,N_30666,N_30667,N_30668,N_30669,N_30670,N_30671,N_30672,N_30673,N_30674,N_30675,N_30676,N_30677,N_30678,N_30679,N_30680,N_30681,N_30682,N_30683,N_30684,N_30685,N_30686,N_30687,N_30688,N_30689,N_30690,N_30691,N_30692,N_30693,N_30694,N_30695,N_30696,N_30697,N_30698,N_30699,N_30700,N_30701,N_30702,N_30703,N_30704,N_30705,N_30706,N_30707,N_30708,N_30709,N_30710,N_30711,N_30712,N_30713,N_30714,N_30715,N_30716,N_30717,N_30718,N_30719,N_30720,N_30721,N_30722,N_30723,N_30724,N_30725,N_30726,N_30727,N_30728,N_30729,N_30730,N_30731,N_30732,N_30733,N_30734,N_30735,N_30736,N_30737,N_30738,N_30739,N_30740,N_30741,N_30742,N_30743,N_30744,N_30745,N_30746,N_30747,N_30748,N_30749,N_30750,N_30751,N_30752,N_30753,N_30754,N_30755,N_30756,N_30757,N_30758,N_30759,N_30760,N_30761,N_30762,N_30763,N_30764,N_30765,N_30766,N_30767,N_30768,N_30769,N_30770,N_30771,N_30772,N_30773,N_30774,N_30775,N_30776,N_30777,N_30778,N_30779,N_30780,N_30781,N_30782,N_30783,N_30784,N_30785,N_30786,N_30787,N_30788,N_30789,N_30790,N_30791,N_30792,N_30793,N_30794,N_30795,N_30796,N_30797,N_30798,N_30799,N_30800,N_30801,N_30802,N_30803,N_30804,N_30805,N_30806,N_30807,N_30808,N_30809,N_30810,N_30811,N_30812,N_30813,N_30814,N_30815,N_30816,N_30817,N_30818,N_30819,N_30820,N_30821,N_30822,N_30823,N_30824,N_30825,N_30826,N_30827,N_30828,N_30829,N_30830,N_30831,N_30832,N_30833,N_30834,N_30835,N_30836,N_30837,N_30838,N_30839,N_30840,N_30841,N_30842,N_30843,N_30844,N_30845,N_30846,N_30847,N_30848,N_30849,N_30850,N_30851,N_30852,N_30853,N_30854,N_30855,N_30856,N_30857,N_30858,N_30859,N_30860,N_30861,N_30862,N_30863,N_30864,N_30865,N_30866,N_30867,N_30868,N_30869,N_30870,N_30871,N_30872,N_30873,N_30874,N_30875,N_30876,N_30877,N_30878,N_30879,N_30880,N_30881,N_30882,N_30883,N_30884,N_30885,N_30886,N_30887,N_30888,N_30889,N_30890,N_30891,N_30892,N_30893,N_30894,N_30895,N_30896,N_30897,N_30898,N_30899,N_30900,N_30901,N_30902,N_30903,N_30904,N_30905,N_30906,N_30907,N_30908,N_30909,N_30910,N_30911,N_30912,N_30913,N_30914,N_30915,N_30916,N_30917,N_30918,N_30919,N_30920,N_30921,N_30922,N_30923,N_30924,N_30925,N_30926,N_30927,N_30928,N_30929,N_30930,N_30931,N_30932,N_30933,N_30934,N_30935,N_30936,N_30937,N_30938,N_30939,N_30940,N_30941,N_30942,N_30943,N_30944,N_30945,N_30946,N_30947,N_30948,N_30949,N_30950,N_30951,N_30952,N_30953,N_30954,N_30955,N_30956,N_30957,N_30958,N_30959,N_30960,N_30961,N_30962,N_30963,N_30964,N_30965,N_30966,N_30967,N_30968,N_30969,N_30970,N_30971,N_30972,N_30973,N_30974,N_30975,N_30976,N_30977,N_30978,N_30979,N_30980,N_30981,N_30982,N_30983,N_30984,N_30985,N_30986,N_30987,N_30988,N_30989,N_30990,N_30991,N_30992,N_30993,N_30994,N_30995,N_30996,N_30997,N_30998,N_30999,N_31000,N_31001,N_31002,N_31003,N_31004,N_31005,N_31006,N_31007,N_31008,N_31009,N_31010,N_31011,N_31012,N_31013,N_31014,N_31015,N_31016,N_31017,N_31018,N_31019,N_31020,N_31021,N_31022,N_31023,N_31024,N_31025,N_31026,N_31027,N_31028,N_31029,N_31030,N_31031,N_31032,N_31033,N_31034,N_31035,N_31036,N_31037,N_31038,N_31039,N_31040,N_31041,N_31042,N_31043,N_31044,N_31045,N_31046,N_31047,N_31048,N_31049,N_31050,N_31051,N_31052,N_31053,N_31054,N_31055,N_31056,N_31057,N_31058,N_31059,N_31060,N_31061,N_31062,N_31063,N_31064,N_31065,N_31066,N_31067,N_31068,N_31069,N_31070,N_31071,N_31072,N_31073,N_31074,N_31075,N_31076,N_31077,N_31078,N_31079,N_31080,N_31081,N_31082,N_31083,N_31084,N_31085,N_31086,N_31087,N_31088,N_31089,N_31090,N_31091,N_31092,N_31093,N_31094,N_31095,N_31096,N_31097,N_31098,N_31099,N_31100,N_31101,N_31102,N_31103,N_31104,N_31105,N_31106,N_31107,N_31108,N_31109,N_31110,N_31111,N_31112,N_31113,N_31114,N_31115,N_31116,N_31117,N_31118,N_31119,N_31120,N_31121,N_31122,N_31123,N_31124,N_31125,N_31126,N_31127,N_31128,N_31129,N_31130,N_31131,N_31132,N_31133,N_31134,N_31135,N_31136,N_31137,N_31138,N_31139,N_31140,N_31141,N_31142,N_31143,N_31144,N_31145,N_31146,N_31147,N_31148,N_31149,N_31150,N_31151,N_31152,N_31153,N_31154,N_31155,N_31156,N_31157,N_31158,N_31159,N_31160,N_31161,N_31162,N_31163,N_31164,N_31165,N_31166,N_31167,N_31168,N_31169,N_31170,N_31171,N_31172,N_31173,N_31174,N_31175,N_31176,N_31177,N_31178,N_31179,N_31180,N_31181,N_31182,N_31183,N_31184,N_31185,N_31186,N_31187,N_31188,N_31189,N_31190,N_31191,N_31192,N_31193,N_31194,N_31195,N_31196,N_31197,N_31198,N_31199,N_31200,N_31201,N_31202,N_31203,N_31204,N_31205,N_31206,N_31207,N_31208,N_31209,N_31210,N_31211,N_31212,N_31213,N_31214,N_31215,N_31216,N_31217,N_31218,N_31219,N_31220,N_31221,N_31222,N_31223,N_31224,N_31225,N_31226,N_31227,N_31228,N_31229,N_31230,N_31231,N_31232,N_31233,N_31234,N_31235,N_31236,N_31237,N_31238,N_31239,N_31240,N_31241,N_31242,N_31243,N_31244,N_31245,N_31246,N_31247,N_31248,N_31249,N_31250,N_31251,N_31252,N_31253,N_31254,N_31255,N_31256,N_31257,N_31258,N_31259,N_31260,N_31261,N_31262,N_31263,N_31264,N_31265,N_31266,N_31267,N_31268,N_31269,N_31270,N_31271,N_31272,N_31273,N_31274,N_31275,N_31276,N_31277,N_31278,N_31279,N_31280,N_31281,N_31282,N_31283,N_31284,N_31285,N_31286,N_31287,N_31288,N_31289,N_31290,N_31291,N_31292,N_31293,N_31294,N_31295,N_31296,N_31297,N_31298,N_31299,N_31300,N_31301,N_31302,N_31303,N_31304,N_31305,N_31306,N_31307,N_31308,N_31309,N_31310,N_31311,N_31312,N_31313,N_31314,N_31315,N_31316,N_31317,N_31318,N_31319,N_31320,N_31321,N_31322,N_31323,N_31324,N_31325,N_31326,N_31327,N_31328,N_31329,N_31330,N_31331,N_31332,N_31333,N_31334,N_31335,N_31336,N_31337,N_31338,N_31339,N_31340,N_31341,N_31342,N_31343,N_31344,N_31345,N_31346,N_31347,N_31348,N_31349,N_31350,N_31351,N_31352,N_31353,N_31354,N_31355,N_31356,N_31357,N_31358,N_31359,N_31360,N_31361,N_31362,N_31363,N_31364,N_31365,N_31366,N_31367,N_31368,N_31369,N_31370,N_31371,N_31372,N_31373,N_31374,N_31375,N_31376,N_31377,N_31378,N_31379,N_31380,N_31381,N_31382,N_31383,N_31384,N_31385,N_31386,N_31387,N_31388,N_31389,N_31390,N_31391,N_31392,N_31393,N_31394,N_31395,N_31396,N_31397,N_31398,N_31399,N_31400,N_31401,N_31402,N_31403,N_31404,N_31405,N_31406,N_31407,N_31408,N_31409,N_31410,N_31411,N_31412,N_31413,N_31414,N_31415,N_31416,N_31417,N_31418,N_31419,N_31420,N_31421,N_31422,N_31423,N_31424,N_31425,N_31426,N_31427,N_31428,N_31429,N_31430,N_31431,N_31432,N_31433,N_31434,N_31435,N_31436,N_31437,N_31438,N_31439,N_31440,N_31441,N_31442,N_31443,N_31444,N_31445,N_31446,N_31447,N_31448,N_31449,N_31450,N_31451,N_31452,N_31453,N_31454,N_31455,N_31456,N_31457,N_31458,N_31459,N_31460,N_31461,N_31462,N_31463,N_31464,N_31465,N_31466,N_31467,N_31468,N_31469,N_31470,N_31471,N_31472,N_31473,N_31474,N_31475,N_31476,N_31477,N_31478,N_31479,N_31480,N_31481,N_31482,N_31483,N_31484,N_31485,N_31486,N_31487,N_31488,N_31489,N_31490,N_31491,N_31492,N_31493,N_31494,N_31495,N_31496,N_31497,N_31498,N_31499,N_31500,N_31501,N_31502,N_31503,N_31504,N_31505,N_31506,N_31507,N_31508,N_31509,N_31510,N_31511,N_31512,N_31513,N_31514,N_31515,N_31516,N_31517,N_31518,N_31519,N_31520,N_31521,N_31522,N_31523,N_31524,N_31525,N_31526,N_31527,N_31528,N_31529,N_31530,N_31531,N_31532,N_31533,N_31534,N_31535,N_31536,N_31537,N_31538,N_31539,N_31540,N_31541,N_31542,N_31543,N_31544,N_31545,N_31546,N_31547,N_31548,N_31549,N_31550,N_31551,N_31552,N_31553,N_31554,N_31555,N_31556,N_31557,N_31558,N_31559,N_31560,N_31561,N_31562,N_31563,N_31564,N_31565,N_31566,N_31567,N_31568,N_31569,N_31570,N_31571,N_31572,N_31573,N_31574,N_31575,N_31576,N_31577,N_31578,N_31579,N_31580,N_31581,N_31582,N_31583,N_31584,N_31585,N_31586,N_31587,N_31588,N_31589,N_31590,N_31591,N_31592,N_31593,N_31594,N_31595,N_31596,N_31597,N_31598,N_31599,N_31600,N_31601,N_31602,N_31603,N_31604,N_31605,N_31606,N_31607,N_31608,N_31609,N_31610,N_31611,N_31612,N_31613,N_31614,N_31615,N_31616,N_31617,N_31618,N_31619,N_31620,N_31621,N_31622,N_31623,N_31624,N_31625,N_31626,N_31627,N_31628,N_31629,N_31630,N_31631,N_31632,N_31633,N_31634,N_31635,N_31636,N_31637,N_31638,N_31639,N_31640,N_31641,N_31642,N_31643,N_31644,N_31645,N_31646,N_31647,N_31648,N_31649,N_31650,N_31651,N_31652,N_31653,N_31654,N_31655,N_31656,N_31657,N_31658,N_31659,N_31660,N_31661,N_31662,N_31663,N_31664,N_31665,N_31666,N_31667,N_31668,N_31669,N_31670,N_31671,N_31672,N_31673,N_31674,N_31675,N_31676,N_31677,N_31678,N_31679,N_31680,N_31681,N_31682,N_31683,N_31684,N_31685,N_31686,N_31687,N_31688,N_31689,N_31690,N_31691,N_31692,N_31693,N_31694,N_31695,N_31696,N_31697,N_31698,N_31699,N_31700,N_31701,N_31702,N_31703,N_31704,N_31705,N_31706,N_31707,N_31708,N_31709,N_31710,N_31711,N_31712,N_31713,N_31714,N_31715,N_31716,N_31717,N_31718,N_31719,N_31720,N_31721,N_31722,N_31723,N_31724,N_31725,N_31726,N_31727,N_31728,N_31729,N_31730,N_31731,N_31732,N_31733,N_31734,N_31735,N_31736,N_31737,N_31738,N_31739,N_31740,N_31741,N_31742,N_31743,N_31744,N_31745,N_31746,N_31747,N_31748,N_31749,N_31750,N_31751,N_31752,N_31753,N_31754,N_31755,N_31756,N_31757,N_31758,N_31759,N_31760,N_31761,N_31762,N_31763,N_31764,N_31765,N_31766,N_31767,N_31768,N_31769,N_31770,N_31771,N_31772,N_31773,N_31774,N_31775,N_31776,N_31777,N_31778,N_31779,N_31780,N_31781,N_31782,N_31783,N_31784,N_31785,N_31786,N_31787,N_31788,N_31789,N_31790,N_31791,N_31792,N_31793,N_31794,N_31795,N_31796,N_31797,N_31798,N_31799,N_31800,N_31801,N_31802,N_31803,N_31804,N_31805,N_31806,N_31807,N_31808,N_31809,N_31810,N_31811,N_31812,N_31813,N_31814,N_31815,N_31816,N_31817,N_31818,N_31819,N_31820,N_31821,N_31822,N_31823,N_31824,N_31825,N_31826,N_31827,N_31828,N_31829,N_31830,N_31831,N_31832,N_31833,N_31834,N_31835,N_31836,N_31837,N_31838,N_31839,N_31840,N_31841,N_31842,N_31843,N_31844,N_31845,N_31846,N_31847,N_31848,N_31849,N_31850,N_31851,N_31852,N_31853,N_31854,N_31855,N_31856,N_31857,N_31858,N_31859,N_31860,N_31861,N_31862,N_31863,N_31864,N_31865,N_31866,N_31867,N_31868,N_31869,N_31870,N_31871,N_31872,N_31873,N_31874,N_31875,N_31876,N_31877,N_31878,N_31879,N_31880,N_31881,N_31882,N_31883,N_31884,N_31885,N_31886,N_31887,N_31888,N_31889,N_31890,N_31891,N_31892,N_31893,N_31894,N_31895,N_31896,N_31897,N_31898,N_31899,N_31900,N_31901,N_31902,N_31903,N_31904,N_31905,N_31906,N_31907,N_31908,N_31909,N_31910,N_31911,N_31912,N_31913,N_31914,N_31915,N_31916,N_31917,N_31918,N_31919,N_31920,N_31921,N_31922,N_31923,N_31924,N_31925,N_31926,N_31927,N_31928,N_31929,N_31930,N_31931,N_31932,N_31933,N_31934,N_31935,N_31936,N_31937,N_31938,N_31939,N_31940,N_31941,N_31942,N_31943,N_31944,N_31945,N_31946,N_31947,N_31948,N_31949,N_31950,N_31951,N_31952,N_31953,N_31954,N_31955,N_31956,N_31957,N_31958,N_31959,N_31960,N_31961,N_31962,N_31963,N_31964,N_31965,N_31966,N_31967,N_31968,N_31969,N_31970,N_31971,N_31972,N_31973,N_31974,N_31975,N_31976,N_31977,N_31978,N_31979,N_31980,N_31981,N_31982,N_31983,N_31984,N_31985,N_31986,N_31987,N_31988,N_31989,N_31990,N_31991,N_31992,N_31993,N_31994,N_31995,N_31996,N_31997,N_31998,N_31999,N_32000,N_32001,N_32002,N_32003,N_32004,N_32005,N_32006,N_32007,N_32008,N_32009,N_32010,N_32011,N_32012,N_32013,N_32014,N_32015,N_32016,N_32017,N_32018,N_32019,N_32020,N_32021,N_32022,N_32023,N_32024,N_32025,N_32026,N_32027,N_32028,N_32029,N_32030,N_32031,N_32032,N_32033,N_32034,N_32035,N_32036,N_32037,N_32038,N_32039,N_32040,N_32041,N_32042,N_32043,N_32044,N_32045,N_32046,N_32047,N_32048,N_32049,N_32050,N_32051,N_32052,N_32053,N_32054,N_32055,N_32056,N_32057,N_32058,N_32059,N_32060,N_32061,N_32062,N_32063,N_32064,N_32065,N_32066,N_32067,N_32068,N_32069,N_32070,N_32071,N_32072,N_32073,N_32074,N_32075,N_32076,N_32077,N_32078,N_32079,N_32080,N_32081,N_32082,N_32083,N_32084,N_32085,N_32086,N_32087,N_32088,N_32089,N_32090,N_32091,N_32092,N_32093,N_32094,N_32095,N_32096,N_32097,N_32098,N_32099,N_32100,N_32101,N_32102,N_32103,N_32104,N_32105,N_32106,N_32107,N_32108,N_32109,N_32110,N_32111,N_32112,N_32113,N_32114,N_32115,N_32116,N_32117,N_32118,N_32119,N_32120,N_32121,N_32122,N_32123,N_32124,N_32125,N_32126,N_32127,N_32128,N_32129,N_32130,N_32131,N_32132,N_32133,N_32134,N_32135,N_32136,N_32137,N_32138,N_32139,N_32140,N_32141,N_32142,N_32143,N_32144,N_32145,N_32146,N_32147,N_32148,N_32149,N_32150,N_32151,N_32152,N_32153,N_32154,N_32155,N_32156,N_32157,N_32158,N_32159,N_32160,N_32161,N_32162,N_32163,N_32164,N_32165,N_32166,N_32167,N_32168,N_32169,N_32170,N_32171,N_32172,N_32173,N_32174,N_32175,N_32176,N_32177,N_32178,N_32179,N_32180,N_32181,N_32182,N_32183,N_32184,N_32185,N_32186,N_32187,N_32188,N_32189,N_32190,N_32191,N_32192,N_32193,N_32194,N_32195,N_32196,N_32197,N_32198,N_32199,N_32200,N_32201,N_32202,N_32203,N_32204,N_32205,N_32206,N_32207,N_32208,N_32209,N_32210,N_32211,N_32212,N_32213,N_32214,N_32215,N_32216,N_32217,N_32218,N_32219,N_32220,N_32221,N_32222,N_32223,N_32224,N_32225,N_32226,N_32227,N_32228,N_32229,N_32230,N_32231,N_32232,N_32233,N_32234,N_32235,N_32236,N_32237,N_32238,N_32239,N_32240,N_32241,N_32242,N_32243,N_32244,N_32245,N_32246,N_32247,N_32248,N_32249,N_32250,N_32251,N_32252,N_32253,N_32254,N_32255,N_32256,N_32257,N_32258,N_32259,N_32260,N_32261,N_32262,N_32263,N_32264,N_32265,N_32266,N_32267,N_32268,N_32269,N_32270,N_32271,N_32272,N_32273,N_32274,N_32275,N_32276,N_32277,N_32278,N_32279,N_32280,N_32281,N_32282,N_32283,N_32284,N_32285,N_32286,N_32287,N_32288,N_32289,N_32290,N_32291,N_32292,N_32293,N_32294,N_32295,N_32296,N_32297,N_32298,N_32299,N_32300,N_32301,N_32302,N_32303,N_32304,N_32305,N_32306,N_32307,N_32308,N_32309,N_32310,N_32311,N_32312,N_32313,N_32314,N_32315,N_32316,N_32317,N_32318,N_32319,N_32320,N_32321,N_32322,N_32323,N_32324,N_32325,N_32326,N_32327,N_32328,N_32329,N_32330,N_32331,N_32332,N_32333,N_32334,N_32335,N_32336,N_32337,N_32338,N_32339,N_32340,N_32341,N_32342,N_32343,N_32344,N_32345,N_32346,N_32347,N_32348,N_32349,N_32350,N_32351,N_32352,N_32353,N_32354,N_32355,N_32356,N_32357,N_32358,N_32359,N_32360,N_32361,N_32362,N_32363,N_32364,N_32365,N_32366,N_32367,N_32368,N_32369,N_32370,N_32371,N_32372,N_32373,N_32374,N_32375,N_32376,N_32377,N_32378,N_32379,N_32380,N_32381,N_32382,N_32383,N_32384,N_32385,N_32386,N_32387,N_32388,N_32389,N_32390,N_32391,N_32392,N_32393,N_32394,N_32395,N_32396,N_32397,N_32398,N_32399,N_32400,N_32401,N_32402,N_32403,N_32404,N_32405,N_32406,N_32407,N_32408,N_32409,N_32410,N_32411,N_32412,N_32413,N_32414,N_32415,N_32416,N_32417,N_32418,N_32419,N_32420,N_32421,N_32422,N_32423,N_32424,N_32425,N_32426,N_32427,N_32428,N_32429,N_32430,N_32431,N_32432,N_32433,N_32434,N_32435,N_32436,N_32437,N_32438,N_32439,N_32440,N_32441,N_32442,N_32443,N_32444,N_32445,N_32446,N_32447,N_32448,N_32449,N_32450,N_32451,N_32452,N_32453,N_32454,N_32455,N_32456,N_32457,N_32458,N_32459,N_32460,N_32461,N_32462,N_32463,N_32464,N_32465,N_32466,N_32467,N_32468,N_32469,N_32470,N_32471,N_32472,N_32473,N_32474,N_32475,N_32476,N_32477,N_32478,N_32479,N_32480,N_32481,N_32482,N_32483,N_32484,N_32485,N_32486,N_32487,N_32488,N_32489,N_32490,N_32491,N_32492,N_32493,N_32494,N_32495,N_32496,N_32497,N_32498,N_32499,N_32500,N_32501,N_32502,N_32503,N_32504,N_32505,N_32506,N_32507,N_32508,N_32509,N_32510,N_32511,N_32512,N_32513,N_32514,N_32515,N_32516,N_32517,N_32518,N_32519,N_32520,N_32521,N_32522,N_32523,N_32524,N_32525,N_32526,N_32527,N_32528,N_32529,N_32530,N_32531,N_32532,N_32533,N_32534,N_32535,N_32536,N_32537,N_32538,N_32539,N_32540,N_32541,N_32542,N_32543,N_32544,N_32545,N_32546,N_32547,N_32548,N_32549,N_32550,N_32551,N_32552,N_32553,N_32554,N_32555,N_32556,N_32557,N_32558,N_32559,N_32560,N_32561,N_32562,N_32563,N_32564,N_32565,N_32566,N_32567,N_32568,N_32569,N_32570,N_32571,N_32572,N_32573,N_32574,N_32575,N_32576,N_32577,N_32578,N_32579,N_32580,N_32581,N_32582,N_32583,N_32584,N_32585,N_32586,N_32587,N_32588,N_32589,N_32590,N_32591,N_32592,N_32593,N_32594,N_32595,N_32596,N_32597,N_32598,N_32599,N_32600,N_32601,N_32602,N_32603,N_32604,N_32605,N_32606,N_32607,N_32608,N_32609,N_32610,N_32611,N_32612,N_32613,N_32614,N_32615,N_32616,N_32617,N_32618,N_32619,N_32620,N_32621,N_32622,N_32623,N_32624,N_32625,N_32626,N_32627,N_32628,N_32629,N_32630,N_32631,N_32632,N_32633,N_32634,N_32635,N_32636,N_32637,N_32638,N_32639,N_32640,N_32641,N_32642,N_32643,N_32644,N_32645,N_32646,N_32647,N_32648,N_32649,N_32650,N_32651,N_32652,N_32653,N_32654,N_32655,N_32656,N_32657,N_32658,N_32659,N_32660,N_32661,N_32662,N_32663,N_32664,N_32665,N_32666,N_32667,N_32668,N_32669,N_32670,N_32671,N_32672,N_32673,N_32674,N_32675,N_32676,N_32677,N_32678,N_32679,N_32680,N_32681,N_32682,N_32683,N_32684,N_32685,N_32686,N_32687,N_32688,N_32689,N_32690,N_32691,N_32692,N_32693,N_32694,N_32695,N_32696,N_32697,N_32698,N_32699,N_32700,N_32701,N_32702,N_32703,N_32704,N_32705,N_32706,N_32707,N_32708,N_32709,N_32710,N_32711,N_32712,N_32713,N_32714,N_32715,N_32716,N_32717,N_32718,N_32719,N_32720,N_32721,N_32722,N_32723,N_32724,N_32725,N_32726,N_32727,N_32728,N_32729,N_32730,N_32731,N_32732,N_32733,N_32734,N_32735,N_32736,N_32737,N_32738,N_32739,N_32740,N_32741,N_32742,N_32743,N_32744,N_32745,N_32746,N_32747,N_32748,N_32749,N_32750,N_32751,N_32752,N_32753,N_32754,N_32755,N_32756,N_32757,N_32758,N_32759,N_32760,N_32761,N_32762,N_32763,N_32764,N_32765,N_32766,N_32767,N_32768,N_32769,N_32770,N_32771,N_32772,N_32773,N_32774,N_32775,N_32776,N_32777,N_32778,N_32779,N_32780,N_32781,N_32782,N_32783,N_32784,N_32785,N_32786,N_32787,N_32788,N_32789,N_32790,N_32791,N_32792,N_32793,N_32794,N_32795,N_32796,N_32797,N_32798,N_32799,N_32800,N_32801,N_32802,N_32803,N_32804,N_32805,N_32806,N_32807,N_32808,N_32809,N_32810,N_32811,N_32812,N_32813,N_32814,N_32815,N_32816,N_32817,N_32818,N_32819,N_32820,N_32821,N_32822,N_32823,N_32824,N_32825,N_32826,N_32827,N_32828,N_32829,N_32830,N_32831,N_32832,N_32833,N_32834,N_32835,N_32836,N_32837,N_32838,N_32839,N_32840,N_32841,N_32842,N_32843,N_32844,N_32845,N_32846,N_32847,N_32848,N_32849,N_32850,N_32851,N_32852,N_32853,N_32854,N_32855,N_32856,N_32857,N_32858,N_32859,N_32860,N_32861,N_32862,N_32863,N_32864,N_32865,N_32866,N_32867,N_32868,N_32869,N_32870,N_32871,N_32872,N_32873,N_32874,N_32875,N_32876,N_32877,N_32878,N_32879,N_32880,N_32881,N_32882,N_32883,N_32884,N_32885,N_32886,N_32887,N_32888,N_32889,N_32890,N_32891,N_32892,N_32893,N_32894,N_32895,N_32896,N_32897,N_32898,N_32899,N_32900,N_32901,N_32902,N_32903,N_32904,N_32905,N_32906,N_32907,N_32908,N_32909,N_32910,N_32911,N_32912,N_32913,N_32914,N_32915,N_32916,N_32917,N_32918,N_32919,N_32920,N_32921,N_32922,N_32923,N_32924,N_32925,N_32926,N_32927,N_32928,N_32929,N_32930,N_32931,N_32932,N_32933,N_32934,N_32935,N_32936,N_32937,N_32938,N_32939,N_32940,N_32941,N_32942,N_32943,N_32944,N_32945,N_32946,N_32947,N_32948,N_32949,N_32950,N_32951,N_32952,N_32953,N_32954,N_32955,N_32956,N_32957,N_32958,N_32959,N_32960,N_32961,N_32962,N_32963,N_32964,N_32965,N_32966,N_32967,N_32968,N_32969,N_32970,N_32971,N_32972,N_32973,N_32974,N_32975,N_32976,N_32977,N_32978,N_32979,N_32980,N_32981,N_32982,N_32983,N_32984,N_32985,N_32986,N_32987,N_32988,N_32989,N_32990,N_32991,N_32992,N_32993,N_32994,N_32995,N_32996,N_32997,N_32998,N_32999,N_33000,N_33001,N_33002,N_33003,N_33004,N_33005,N_33006,N_33007,N_33008,N_33009,N_33010,N_33011,N_33012,N_33013,N_33014,N_33015,N_33016,N_33017,N_33018,N_33019,N_33020,N_33021,N_33022,N_33023,N_33024,N_33025,N_33026,N_33027,N_33028,N_33029,N_33030,N_33031,N_33032,N_33033,N_33034,N_33035,N_33036,N_33037,N_33038,N_33039,N_33040,N_33041,N_33042,N_33043,N_33044,N_33045,N_33046,N_33047,N_33048,N_33049,N_33050,N_33051,N_33052,N_33053,N_33054,N_33055,N_33056,N_33057,N_33058,N_33059,N_33060,N_33061,N_33062,N_33063,N_33064,N_33065,N_33066,N_33067,N_33068,N_33069,N_33070,N_33071,N_33072,N_33073,N_33074,N_33075,N_33076,N_33077,N_33078,N_33079,N_33080,N_33081,N_33082,N_33083,N_33084,N_33085,N_33086,N_33087,N_33088,N_33089,N_33090,N_33091,N_33092,N_33093,N_33094,N_33095,N_33096,N_33097,N_33098,N_33099,N_33100,N_33101,N_33102,N_33103,N_33104,N_33105,N_33106,N_33107,N_33108,N_33109,N_33110,N_33111,N_33112,N_33113,N_33114,N_33115,N_33116,N_33117,N_33118,N_33119,N_33120,N_33121,N_33122,N_33123,N_33124,N_33125,N_33126,N_33127,N_33128,N_33129,N_33130,N_33131,N_33132,N_33133,N_33134,N_33135,N_33136,N_33137,N_33138,N_33139,N_33140,N_33141,N_33142,N_33143,N_33144,N_33145,N_33146,N_33147,N_33148,N_33149,N_33150,N_33151,N_33152,N_33153,N_33154,N_33155,N_33156,N_33157,N_33158,N_33159,N_33160,N_33161,N_33162,N_33163,N_33164,N_33165,N_33166,N_33167,N_33168,N_33169,N_33170,N_33171,N_33172,N_33173,N_33174,N_33175,N_33176,N_33177,N_33178,N_33179,N_33180,N_33181,N_33182,N_33183,N_33184,N_33185,N_33186,N_33187,N_33188,N_33189,N_33190,N_33191,N_33192,N_33193,N_33194,N_33195,N_33196,N_33197,N_33198,N_33199,N_33200,N_33201,N_33202,N_33203,N_33204,N_33205,N_33206,N_33207,N_33208,N_33209,N_33210,N_33211,N_33212,N_33213,N_33214,N_33215,N_33216,N_33217,N_33218,N_33219,N_33220,N_33221,N_33222,N_33223,N_33224,N_33225,N_33226,N_33227,N_33228,N_33229,N_33230,N_33231,N_33232,N_33233,N_33234,N_33235,N_33236,N_33237,N_33238,N_33239,N_33240,N_33241,N_33242,N_33243,N_33244,N_33245,N_33246,N_33247,N_33248,N_33249,N_33250,N_33251,N_33252,N_33253,N_33254,N_33255,N_33256,N_33257,N_33258,N_33259,N_33260,N_33261,N_33262,N_33263,N_33264,N_33265,N_33266,N_33267,N_33268,N_33269,N_33270,N_33271,N_33272,N_33273,N_33274,N_33275,N_33276,N_33277,N_33278,N_33279,N_33280,N_33281,N_33282,N_33283,N_33284,N_33285,N_33286,N_33287,N_33288,N_33289,N_33290,N_33291,N_33292,N_33293,N_33294,N_33295,N_33296,N_33297,N_33298,N_33299,N_33300,N_33301,N_33302,N_33303,N_33304,N_33305,N_33306,N_33307,N_33308,N_33309,N_33310,N_33311,N_33312,N_33313,N_33314,N_33315,N_33316,N_33317,N_33318,N_33319,N_33320,N_33321,N_33322,N_33323,N_33324,N_33325,N_33326,N_33327,N_33328,N_33329,N_33330,N_33331,N_33332,N_33333,N_33334,N_33335,N_33336,N_33337,N_33338,N_33339,N_33340,N_33341,N_33342,N_33343,N_33344,N_33345,N_33346,N_33347,N_33348,N_33349,N_33350,N_33351,N_33352,N_33353,N_33354,N_33355,N_33356,N_33357,N_33358,N_33359,N_33360,N_33361,N_33362,N_33363,N_33364,N_33365,N_33366,N_33367,N_33368,N_33369,N_33370,N_33371,N_33372,N_33373,N_33374,N_33375,N_33376,N_33377,N_33378,N_33379,N_33380,N_33381,N_33382,N_33383,N_33384,N_33385,N_33386,N_33387,N_33388,N_33389,N_33390,N_33391,N_33392,N_33393,N_33394,N_33395,N_33396,N_33397,N_33398,N_33399,N_33400,N_33401,N_33402,N_33403,N_33404,N_33405,N_33406,N_33407,N_33408,N_33409,N_33410,N_33411,N_33412,N_33413,N_33414,N_33415,N_33416,N_33417,N_33418,N_33419,N_33420,N_33421,N_33422,N_33423,N_33424,N_33425,N_33426,N_33427,N_33428,N_33429,N_33430,N_33431,N_33432,N_33433,N_33434,N_33435,N_33436,N_33437,N_33438,N_33439,N_33440,N_33441,N_33442,N_33443,N_33444,N_33445,N_33446,N_33447,N_33448,N_33449,N_33450,N_33451,N_33452,N_33453,N_33454,N_33455,N_33456,N_33457,N_33458,N_33459,N_33460,N_33461,N_33462,N_33463,N_33464,N_33465,N_33466,N_33467,N_33468,N_33469,N_33470,N_33471,N_33472,N_33473,N_33474,N_33475,N_33476,N_33477,N_33478,N_33479,N_33480,N_33481,N_33482,N_33483,N_33484,N_33485,N_33486,N_33487,N_33488,N_33489,N_33490,N_33491,N_33492,N_33493,N_33494,N_33495,N_33496,N_33497,N_33498,N_33499,N_33500,N_33501,N_33502,N_33503,N_33504,N_33505,N_33506,N_33507,N_33508,N_33509,N_33510,N_33511,N_33512,N_33513,N_33514,N_33515,N_33516,N_33517,N_33518,N_33519,N_33520,N_33521,N_33522,N_33523,N_33524,N_33525,N_33526,N_33527,N_33528,N_33529,N_33530,N_33531,N_33532,N_33533,N_33534,N_33535,N_33536,N_33537,N_33538,N_33539,N_33540,N_33541,N_33542,N_33543,N_33544,N_33545,N_33546,N_33547,N_33548,N_33549,N_33550,N_33551,N_33552,N_33553,N_33554,N_33555,N_33556,N_33557,N_33558,N_33559,N_33560,N_33561,N_33562,N_33563,N_33564,N_33565,N_33566,N_33567,N_33568,N_33569,N_33570,N_33571,N_33572,N_33573,N_33574,N_33575,N_33576,N_33577,N_33578,N_33579,N_33580,N_33581,N_33582,N_33583,N_33584,N_33585,N_33586,N_33587,N_33588,N_33589,N_33590,N_33591,N_33592,N_33593,N_33594,N_33595,N_33596,N_33597,N_33598,N_33599,N_33600,N_33601,N_33602,N_33603,N_33604,N_33605,N_33606,N_33607,N_33608,N_33609,N_33610,N_33611,N_33612,N_33613,N_33614,N_33615,N_33616,N_33617,N_33618,N_33619,N_33620,N_33621,N_33622,N_33623,N_33624,N_33625,N_33626,N_33627,N_33628,N_33629,N_33630,N_33631,N_33632,N_33633,N_33634,N_33635,N_33636,N_33637,N_33638,N_33639,N_33640,N_33641,N_33642,N_33643,N_33644,N_33645,N_33646,N_33647,N_33648,N_33649,N_33650,N_33651,N_33652,N_33653,N_33654,N_33655,N_33656,N_33657,N_33658,N_33659,N_33660,N_33661,N_33662,N_33663,N_33664,N_33665,N_33666,N_33667,N_33668,N_33669,N_33670,N_33671,N_33672,N_33673,N_33674,N_33675,N_33676,N_33677,N_33678,N_33679,N_33680,N_33681,N_33682,N_33683,N_33684,N_33685,N_33686,N_33687,N_33688,N_33689,N_33690,N_33691,N_33692,N_33693,N_33694,N_33695,N_33696,N_33697,N_33698,N_33699,N_33700,N_33701,N_33702,N_33703,N_33704,N_33705,N_33706,N_33707,N_33708,N_33709,N_33710,N_33711,N_33712,N_33713,N_33714,N_33715,N_33716,N_33717,N_33718,N_33719,N_33720,N_33721,N_33722,N_33723,N_33724,N_33725,N_33726,N_33727,N_33728,N_33729,N_33730,N_33731,N_33732,N_33733,N_33734,N_33735,N_33736,N_33737,N_33738,N_33739,N_33740,N_33741,N_33742,N_33743,N_33744,N_33745,N_33746,N_33747,N_33748,N_33749,N_33750,N_33751,N_33752,N_33753,N_33754,N_33755,N_33756,N_33757,N_33758,N_33759,N_33760,N_33761,N_33762,N_33763,N_33764,N_33765,N_33766,N_33767,N_33768,N_33769,N_33770,N_33771,N_33772,N_33773,N_33774,N_33775,N_33776,N_33777,N_33778,N_33779,N_33780,N_33781,N_33782,N_33783,N_33784,N_33785,N_33786,N_33787,N_33788,N_33789,N_33790,N_33791,N_33792,N_33793,N_33794,N_33795,N_33796,N_33797,N_33798,N_33799,N_33800,N_33801,N_33802,N_33803,N_33804,N_33805,N_33806,N_33807,N_33808,N_33809,N_33810,N_33811,N_33812,N_33813,N_33814,N_33815,N_33816,N_33817,N_33818,N_33819,N_33820,N_33821,N_33822,N_33823,N_33824,N_33825,N_33826,N_33827,N_33828,N_33829,N_33830,N_33831,N_33832,N_33833,N_33834,N_33835,N_33836,N_33837,N_33838,N_33839,N_33840,N_33841,N_33842,N_33843,N_33844,N_33845,N_33846,N_33847,N_33848,N_33849,N_33850,N_33851,N_33852,N_33853,N_33854,N_33855,N_33856,N_33857,N_33858,N_33859,N_33860,N_33861,N_33862,N_33863,N_33864,N_33865,N_33866,N_33867,N_33868,N_33869,N_33870,N_33871,N_33872,N_33873,N_33874,N_33875,N_33876,N_33877,N_33878,N_33879,N_33880,N_33881,N_33882,N_33883,N_33884,N_33885,N_33886,N_33887,N_33888,N_33889,N_33890,N_33891,N_33892,N_33893,N_33894,N_33895,N_33896,N_33897,N_33898,N_33899,N_33900,N_33901,N_33902,N_33903,N_33904,N_33905,N_33906,N_33907,N_33908,N_33909,N_33910,N_33911,N_33912,N_33913,N_33914,N_33915,N_33916,N_33917,N_33918,N_33919,N_33920,N_33921,N_33922,N_33923,N_33924,N_33925,N_33926,N_33927,N_33928,N_33929,N_33930,N_33931,N_33932,N_33933,N_33934,N_33935,N_33936,N_33937,N_33938,N_33939,N_33940,N_33941,N_33942,N_33943,N_33944,N_33945,N_33946,N_33947,N_33948,N_33949,N_33950,N_33951,N_33952,N_33953,N_33954,N_33955,N_33956,N_33957,N_33958,N_33959,N_33960,N_33961,N_33962,N_33963,N_33964,N_33965,N_33966,N_33967,N_33968,N_33969,N_33970,N_33971,N_33972,N_33973,N_33974,N_33975,N_33976,N_33977,N_33978,N_33979,N_33980,N_33981,N_33982,N_33983,N_33984,N_33985,N_33986,N_33987,N_33988,N_33989,N_33990,N_33991,N_33992,N_33993,N_33994,N_33995,N_33996,N_33997,N_33998,N_33999,N_34000,N_34001,N_34002,N_34003,N_34004,N_34005,N_34006,N_34007,N_34008,N_34009,N_34010,N_34011,N_34012,N_34013,N_34014,N_34015,N_34016,N_34017,N_34018,N_34019,N_34020,N_34021,N_34022,N_34023,N_34024,N_34025,N_34026,N_34027,N_34028,N_34029,N_34030,N_34031,N_34032,N_34033,N_34034,N_34035,N_34036,N_34037,N_34038,N_34039,N_34040,N_34041,N_34042,N_34043,N_34044,N_34045,N_34046,N_34047,N_34048,N_34049,N_34050,N_34051,N_34052,N_34053,N_34054,N_34055,N_34056,N_34057,N_34058,N_34059,N_34060,N_34061,N_34062,N_34063,N_34064,N_34065,N_34066,N_34067,N_34068,N_34069,N_34070,N_34071,N_34072,N_34073,N_34074,N_34075,N_34076,N_34077,N_34078,N_34079,N_34080,N_34081,N_34082,N_34083,N_34084,N_34085,N_34086,N_34087,N_34088,N_34089,N_34090,N_34091,N_34092,N_34093,N_34094,N_34095,N_34096,N_34097,N_34098,N_34099,N_34100,N_34101,N_34102,N_34103,N_34104,N_34105,N_34106,N_34107,N_34108,N_34109,N_34110,N_34111,N_34112,N_34113,N_34114,N_34115,N_34116,N_34117,N_34118,N_34119,N_34120,N_34121,N_34122,N_34123,N_34124,N_34125,N_34126,N_34127,N_34128,N_34129,N_34130,N_34131,N_34132,N_34133,N_34134,N_34135,N_34136,N_34137,N_34138,N_34139,N_34140,N_34141,N_34142,N_34143,N_34144,N_34145,N_34146,N_34147,N_34148,N_34149,N_34150,N_34151,N_34152,N_34153,N_34154,N_34155,N_34156,N_34157,N_34158,N_34159,N_34160,N_34161,N_34162,N_34163,N_34164,N_34165,N_34166,N_34167,N_34168,N_34169,N_34170,N_34171,N_34172,N_34173,N_34174,N_34175,N_34176,N_34177,N_34178,N_34179,N_34180,N_34181,N_34182,N_34183,N_34184,N_34185,N_34186,N_34187,N_34188,N_34189,N_34190,N_34191,N_34192,N_34193,N_34194,N_34195,N_34196,N_34197,N_34198,N_34199,N_34200,N_34201,N_34202,N_34203,N_34204,N_34205,N_34206,N_34207,N_34208,N_34209,N_34210,N_34211,N_34212,N_34213,N_34214,N_34215,N_34216,N_34217,N_34218,N_34219,N_34220,N_34221,N_34222,N_34223,N_34224,N_34225,N_34226,N_34227,N_34228,N_34229,N_34230,N_34231,N_34232,N_34233,N_34234,N_34235,N_34236,N_34237,N_34238,N_34239,N_34240,N_34241,N_34242,N_34243,N_34244,N_34245,N_34246,N_34247,N_34248,N_34249,N_34250,N_34251,N_34252,N_34253,N_34254,N_34255,N_34256,N_34257,N_34258,N_34259,N_34260,N_34261,N_34262,N_34263,N_34264,N_34265,N_34266,N_34267,N_34268,N_34269,N_34270,N_34271,N_34272,N_34273,N_34274,N_34275,N_34276,N_34277,N_34278,N_34279,N_34280,N_34281,N_34282,N_34283,N_34284,N_34285,N_34286,N_34287,N_34288,N_34289,N_34290,N_34291,N_34292,N_34293,N_34294,N_34295,N_34296,N_34297,N_34298,N_34299,N_34300,N_34301,N_34302,N_34303,N_34304,N_34305,N_34306,N_34307,N_34308,N_34309,N_34310,N_34311,N_34312,N_34313,N_34314,N_34315,N_34316,N_34317,N_34318,N_34319,N_34320,N_34321,N_34322,N_34323,N_34324,N_34325,N_34326,N_34327,N_34328,N_34329,N_34330,N_34331,N_34332,N_34333,N_34334,N_34335,N_34336,N_34337,N_34338,N_34339,N_34340,N_34341,N_34342,N_34343,N_34344,N_34345,N_34346,N_34347,N_34348,N_34349,N_34350,N_34351,N_34352,N_34353,N_34354,N_34355,N_34356,N_34357,N_34358,N_34359,N_34360,N_34361,N_34362,N_34363,N_34364,N_34365,N_34366,N_34367,N_34368,N_34369,N_34370,N_34371,N_34372,N_34373,N_34374,N_34375,N_34376,N_34377,N_34378,N_34379,N_34380,N_34381,N_34382,N_34383,N_34384,N_34385,N_34386,N_34387,N_34388,N_34389,N_34390,N_34391,N_34392,N_34393,N_34394,N_34395,N_34396,N_34397,N_34398,N_34399,N_34400,N_34401,N_34402,N_34403,N_34404,N_34405,N_34406,N_34407,N_34408,N_34409,N_34410,N_34411,N_34412,N_34413,N_34414,N_34415,N_34416,N_34417,N_34418,N_34419,N_34420,N_34421,N_34422,N_34423,N_34424,N_34425,N_34426,N_34427,N_34428,N_34429,N_34430,N_34431,N_34432,N_34433,N_34434,N_34435,N_34436,N_34437,N_34438,N_34439,N_34440,N_34441,N_34442,N_34443,N_34444,N_34445,N_34446,N_34447,N_34448,N_34449,N_34450,N_34451,N_34452,N_34453,N_34454,N_34455,N_34456,N_34457,N_34458,N_34459,N_34460,N_34461,N_34462,N_34463,N_34464,N_34465,N_34466,N_34467,N_34468,N_34469,N_34470,N_34471,N_34472,N_34473,N_34474,N_34475,N_34476,N_34477,N_34478,N_34479,N_34480,N_34481,N_34482,N_34483,N_34484,N_34485,N_34486,N_34487,N_34488,N_34489,N_34490,N_34491,N_34492,N_34493,N_34494,N_34495,N_34496,N_34497,N_34498,N_34499,N_34500,N_34501,N_34502,N_34503,N_34504,N_34505,N_34506,N_34507,N_34508,N_34509,N_34510,N_34511,N_34512,N_34513,N_34514,N_34515,N_34516,N_34517,N_34518,N_34519,N_34520,N_34521,N_34522,N_34523,N_34524,N_34525,N_34526,N_34527,N_34528,N_34529,N_34530,N_34531,N_34532,N_34533,N_34534,N_34535,N_34536,N_34537,N_34538,N_34539,N_34540,N_34541,N_34542,N_34543,N_34544,N_34545,N_34546,N_34547,N_34548,N_34549,N_34550,N_34551,N_34552,N_34553,N_34554,N_34555,N_34556,N_34557,N_34558,N_34559,N_34560,N_34561,N_34562,N_34563,N_34564,N_34565,N_34566,N_34567,N_34568,N_34569,N_34570,N_34571,N_34572,N_34573,N_34574,N_34575,N_34576,N_34577,N_34578,N_34579,N_34580,N_34581,N_34582,N_34583,N_34584,N_34585,N_34586,N_34587,N_34588,N_34589,N_34590,N_34591,N_34592,N_34593,N_34594,N_34595,N_34596,N_34597,N_34598,N_34599,N_34600,N_34601,N_34602,N_34603,N_34604,N_34605,N_34606,N_34607,N_34608,N_34609,N_34610,N_34611,N_34612,N_34613,N_34614,N_34615,N_34616,N_34617,N_34618,N_34619,N_34620,N_34621,N_34622,N_34623,N_34624,N_34625,N_34626,N_34627,N_34628,N_34629,N_34630,N_34631,N_34632,N_34633,N_34634,N_34635,N_34636,N_34637,N_34638,N_34639,N_34640,N_34641,N_34642,N_34643,N_34644,N_34645,N_34646,N_34647,N_34648,N_34649,N_34650,N_34651,N_34652,N_34653,N_34654,N_34655,N_34656,N_34657,N_34658,N_34659,N_34660,N_34661,N_34662,N_34663,N_34664,N_34665,N_34666,N_34667,N_34668,N_34669,N_34670,N_34671,N_34672,N_34673,N_34674,N_34675,N_34676,N_34677,N_34678,N_34679,N_34680,N_34681,N_34682,N_34683,N_34684,N_34685,N_34686,N_34687,N_34688,N_34689,N_34690,N_34691,N_34692,N_34693,N_34694,N_34695,N_34696,N_34697,N_34698,N_34699,N_34700,N_34701,N_34702,N_34703,N_34704,N_34705,N_34706,N_34707,N_34708,N_34709,N_34710,N_34711,N_34712,N_34713,N_34714,N_34715,N_34716,N_34717,N_34718,N_34719,N_34720,N_34721,N_34722,N_34723,N_34724,N_34725,N_34726,N_34727,N_34728,N_34729,N_34730,N_34731,N_34732,N_34733,N_34734,N_34735,N_34736,N_34737,N_34738,N_34739,N_34740,N_34741,N_34742,N_34743,N_34744,N_34745,N_34746,N_34747,N_34748,N_34749,N_34750,N_34751,N_34752,N_34753,N_34754,N_34755,N_34756,N_34757,N_34758,N_34759,N_34760,N_34761,N_34762,N_34763,N_34764,N_34765,N_34766,N_34767,N_34768,N_34769,N_34770,N_34771,N_34772,N_34773,N_34774,N_34775,N_34776,N_34777,N_34778,N_34779,N_34780,N_34781,N_34782,N_34783,N_34784,N_34785,N_34786,N_34787,N_34788,N_34789,N_34790,N_34791,N_34792,N_34793,N_34794,N_34795,N_34796,N_34797,N_34798,N_34799,N_34800,N_34801,N_34802,N_34803,N_34804,N_34805,N_34806,N_34807,N_34808,N_34809,N_34810,N_34811,N_34812,N_34813,N_34814,N_34815,N_34816,N_34817,N_34818,N_34819,N_34820,N_34821,N_34822,N_34823,N_34824,N_34825,N_34826,N_34827,N_34828,N_34829,N_34830,N_34831,N_34832,N_34833,N_34834,N_34835,N_34836,N_34837,N_34838,N_34839,N_34840,N_34841,N_34842,N_34843,N_34844,N_34845,N_34846,N_34847,N_34848,N_34849,N_34850,N_34851,N_34852,N_34853,N_34854,N_34855,N_34856,N_34857,N_34858,N_34859,N_34860,N_34861,N_34862,N_34863,N_34864,N_34865,N_34866,N_34867,N_34868,N_34869,N_34870,N_34871,N_34872,N_34873,N_34874,N_34875,N_34876,N_34877,N_34878,N_34879,N_34880,N_34881,N_34882,N_34883,N_34884,N_34885,N_34886,N_34887,N_34888,N_34889,N_34890,N_34891,N_34892,N_34893,N_34894,N_34895,N_34896,N_34897,N_34898,N_34899,N_34900,N_34901,N_34902,N_34903,N_34904,N_34905,N_34906,N_34907,N_34908,N_34909,N_34910,N_34911,N_34912,N_34913,N_34914,N_34915,N_34916,N_34917,N_34918,N_34919,N_34920,N_34921,N_34922,N_34923,N_34924,N_34925,N_34926,N_34927,N_34928,N_34929,N_34930,N_34931,N_34932,N_34933,N_34934,N_34935,N_34936,N_34937,N_34938,N_34939,N_34940,N_34941,N_34942,N_34943,N_34944,N_34945,N_34946,N_34947,N_34948,N_34949,N_34950,N_34951,N_34952,N_34953,N_34954,N_34955,N_34956,N_34957,N_34958,N_34959,N_34960,N_34961,N_34962,N_34963,N_34964,N_34965,N_34966,N_34967,N_34968,N_34969,N_34970,N_34971,N_34972,N_34973,N_34974,N_34975,N_34976,N_34977,N_34978,N_34979,N_34980,N_34981,N_34982,N_34983,N_34984,N_34985,N_34986,N_34987,N_34988,N_34989,N_34990,N_34991,N_34992,N_34993,N_34994,N_34995,N_34996,N_34997,N_34998,N_34999,N_35000,N_35001,N_35002,N_35003,N_35004,N_35005,N_35006,N_35007,N_35008,N_35009,N_35010,N_35011,N_35012,N_35013,N_35014,N_35015,N_35016,N_35017,N_35018,N_35019,N_35020,N_35021,N_35022,N_35023,N_35024,N_35025,N_35026,N_35027,N_35028,N_35029,N_35030,N_35031,N_35032,N_35033,N_35034,N_35035,N_35036,N_35037,N_35038,N_35039,N_35040,N_35041,N_35042,N_35043,N_35044,N_35045,N_35046,N_35047,N_35048,N_35049,N_35050,N_35051,N_35052,N_35053,N_35054,N_35055,N_35056,N_35057,N_35058,N_35059,N_35060,N_35061,N_35062,N_35063,N_35064,N_35065,N_35066,N_35067,N_35068,N_35069,N_35070,N_35071,N_35072,N_35073,N_35074,N_35075,N_35076,N_35077,N_35078,N_35079,N_35080,N_35081,N_35082,N_35083,N_35084,N_35085,N_35086,N_35087,N_35088,N_35089,N_35090,N_35091,N_35092,N_35093,N_35094,N_35095,N_35096,N_35097,N_35098,N_35099,N_35100,N_35101,N_35102,N_35103,N_35104,N_35105,N_35106,N_35107,N_35108,N_35109,N_35110,N_35111,N_35112,N_35113,N_35114,N_35115,N_35116,N_35117,N_35118,N_35119,N_35120,N_35121,N_35122,N_35123,N_35124,N_35125,N_35126,N_35127,N_35128,N_35129,N_35130,N_35131,N_35132,N_35133,N_35134,N_35135,N_35136,N_35137,N_35138,N_35139,N_35140,N_35141,N_35142,N_35143,N_35144,N_35145,N_35146,N_35147,N_35148,N_35149,N_35150,N_35151,N_35152,N_35153,N_35154,N_35155,N_35156,N_35157,N_35158,N_35159,N_35160,N_35161,N_35162,N_35163,N_35164,N_35165,N_35166,N_35167,N_35168,N_35169,N_35170,N_35171,N_35172,N_35173,N_35174,N_35175,N_35176,N_35177,N_35178,N_35179,N_35180,N_35181,N_35182,N_35183,N_35184,N_35185,N_35186,N_35187,N_35188,N_35189,N_35190,N_35191,N_35192,N_35193,N_35194,N_35195,N_35196,N_35197,N_35198,N_35199,N_35200,N_35201,N_35202,N_35203,N_35204,N_35205,N_35206,N_35207,N_35208,N_35209,N_35210,N_35211,N_35212,N_35213,N_35214,N_35215,N_35216,N_35217,N_35218,N_35219,N_35220,N_35221,N_35222,N_35223,N_35224,N_35225,N_35226,N_35227,N_35228,N_35229,N_35230,N_35231,N_35232,N_35233,N_35234,N_35235,N_35236,N_35237,N_35238,N_35239,N_35240,N_35241,N_35242,N_35243,N_35244,N_35245,N_35246,N_35247,N_35248,N_35249,N_35250,N_35251,N_35252,N_35253,N_35254,N_35255,N_35256,N_35257,N_35258,N_35259,N_35260,N_35261,N_35262,N_35263,N_35264,N_35265,N_35266,N_35267,N_35268,N_35269,N_35270,N_35271,N_35272,N_35273,N_35274,N_35275,N_35276,N_35277,N_35278,N_35279,N_35280,N_35281,N_35282,N_35283,N_35284,N_35285,N_35286,N_35287,N_35288,N_35289,N_35290,N_35291,N_35292,N_35293,N_35294,N_35295,N_35296,N_35297,N_35298,N_35299,N_35300,N_35301,N_35302,N_35303,N_35304,N_35305,N_35306,N_35307,N_35308,N_35309,N_35310,N_35311,N_35312,N_35313,N_35314,N_35315,N_35316,N_35317,N_35318,N_35319,N_35320,N_35321,N_35322,N_35323,N_35324,N_35325,N_35326,N_35327,N_35328,N_35329,N_35330,N_35331,N_35332,N_35333,N_35334,N_35335,N_35336,N_35337,N_35338,N_35339,N_35340,N_35341,N_35342,N_35343,N_35344,N_35345,N_35346,N_35347,N_35348,N_35349,N_35350,N_35351,N_35352,N_35353,N_35354,N_35355,N_35356,N_35357,N_35358,N_35359,N_35360,N_35361,N_35362,N_35363,N_35364,N_35365,N_35366,N_35367,N_35368,N_35369,N_35370,N_35371,N_35372,N_35373,N_35374,N_35375,N_35376,N_35377,N_35378,N_35379,N_35380,N_35381,N_35382,N_35383,N_35384,N_35385,N_35386,N_35387,N_35388,N_35389,N_35390,N_35391,N_35392,N_35393,N_35394,N_35395,N_35396,N_35397,N_35398,N_35399,N_35400,N_35401,N_35402,N_35403,N_35404,N_35405,N_35406,N_35407,N_35408,N_35409,N_35410,N_35411,N_35412,N_35413,N_35414,N_35415,N_35416,N_35417,N_35418,N_35419,N_35420,N_35421,N_35422,N_35423,N_35424,N_35425,N_35426,N_35427,N_35428,N_35429,N_35430,N_35431,N_35432,N_35433,N_35434,N_35435,N_35436,N_35437,N_35438,N_35439,N_35440,N_35441,N_35442,N_35443,N_35444,N_35445,N_35446,N_35447,N_35448,N_35449,N_35450,N_35451,N_35452,N_35453,N_35454,N_35455,N_35456,N_35457,N_35458,N_35459,N_35460,N_35461,N_35462,N_35463,N_35464,N_35465,N_35466,N_35467,N_35468,N_35469,N_35470,N_35471,N_35472,N_35473,N_35474,N_35475,N_35476,N_35477,N_35478,N_35479,N_35480,N_35481,N_35482,N_35483,N_35484,N_35485,N_35486,N_35487,N_35488,N_35489,N_35490,N_35491,N_35492,N_35493,N_35494,N_35495,N_35496,N_35497,N_35498,N_35499,N_35500,N_35501,N_35502,N_35503,N_35504,N_35505,N_35506,N_35507,N_35508,N_35509,N_35510,N_35511,N_35512,N_35513,N_35514,N_35515,N_35516,N_35517,N_35518,N_35519,N_35520,N_35521,N_35522,N_35523,N_35524,N_35525,N_35526,N_35527,N_35528,N_35529,N_35530,N_35531,N_35532,N_35533,N_35534,N_35535,N_35536,N_35537,N_35538,N_35539,N_35540,N_35541,N_35542,N_35543,N_35544,N_35545,N_35546,N_35547,N_35548,N_35549,N_35550,N_35551,N_35552,N_35553,N_35554,N_35555,N_35556,N_35557,N_35558,N_35559,N_35560,N_35561,N_35562,N_35563,N_35564,N_35565,N_35566,N_35567,N_35568,N_35569,N_35570,N_35571,N_35572,N_35573,N_35574,N_35575,N_35576,N_35577,N_35578,N_35579,N_35580,N_35581,N_35582,N_35583,N_35584,N_35585,N_35586,N_35587,N_35588,N_35589,N_35590,N_35591,N_35592,N_35593,N_35594,N_35595,N_35596,N_35597,N_35598,N_35599,N_35600,N_35601,N_35602,N_35603,N_35604,N_35605,N_35606,N_35607,N_35608,N_35609,N_35610,N_35611,N_35612,N_35613,N_35614,N_35615,N_35616,N_35617,N_35618,N_35619,N_35620,N_35621,N_35622,N_35623,N_35624,N_35625,N_35626,N_35627,N_35628,N_35629,N_35630,N_35631,N_35632,N_35633,N_35634,N_35635,N_35636,N_35637,N_35638,N_35639,N_35640,N_35641,N_35642,N_35643,N_35644,N_35645,N_35646,N_35647,N_35648,N_35649,N_35650,N_35651,N_35652,N_35653,N_35654,N_35655,N_35656,N_35657,N_35658,N_35659,N_35660,N_35661,N_35662,N_35663,N_35664,N_35665,N_35666,N_35667,N_35668,N_35669,N_35670,N_35671,N_35672,N_35673,N_35674,N_35675,N_35676,N_35677,N_35678,N_35679,N_35680,N_35681,N_35682,N_35683,N_35684,N_35685,N_35686,N_35687,N_35688,N_35689,N_35690,N_35691,N_35692,N_35693,N_35694,N_35695,N_35696,N_35697,N_35698,N_35699,N_35700,N_35701,N_35702,N_35703,N_35704,N_35705,N_35706,N_35707,N_35708,N_35709,N_35710,N_35711,N_35712,N_35713,N_35714,N_35715,N_35716,N_35717,N_35718,N_35719,N_35720,N_35721,N_35722,N_35723,N_35724,N_35725,N_35726,N_35727,N_35728,N_35729,N_35730,N_35731,N_35732,N_35733,N_35734,N_35735,N_35736,N_35737,N_35738,N_35739,N_35740,N_35741,N_35742,N_35743,N_35744,N_35745,N_35746,N_35747,N_35748,N_35749,N_35750,N_35751,N_35752,N_35753,N_35754,N_35755,N_35756,N_35757,N_35758,N_35759,N_35760,N_35761,N_35762,N_35763,N_35764,N_35765,N_35766,N_35767,N_35768,N_35769,N_35770,N_35771,N_35772,N_35773,N_35774,N_35775,N_35776,N_35777,N_35778,N_35779,N_35780,N_35781,N_35782,N_35783,N_35784,N_35785,N_35786,N_35787,N_35788,N_35789,N_35790,N_35791,N_35792,N_35793,N_35794,N_35795,N_35796,N_35797,N_35798,N_35799,N_35800,N_35801,N_35802,N_35803,N_35804,N_35805,N_35806,N_35807,N_35808,N_35809,N_35810,N_35811,N_35812,N_35813,N_35814,N_35815,N_35816,N_35817,N_35818,N_35819,N_35820,N_35821,N_35822,N_35823,N_35824,N_35825,N_35826,N_35827,N_35828,N_35829,N_35830,N_35831,N_35832,N_35833,N_35834,N_35835,N_35836,N_35837,N_35838,N_35839,N_35840,N_35841,N_35842,N_35843,N_35844,N_35845,N_35846,N_35847,N_35848,N_35849,N_35850,N_35851,N_35852,N_35853,N_35854,N_35855,N_35856,N_35857,N_35858,N_35859,N_35860,N_35861,N_35862,N_35863,N_35864,N_35865,N_35866,N_35867,N_35868,N_35869,N_35870,N_35871,N_35872,N_35873,N_35874,N_35875,N_35876,N_35877,N_35878,N_35879,N_35880,N_35881,N_35882,N_35883,N_35884,N_35885,N_35886,N_35887,N_35888,N_35889,N_35890,N_35891,N_35892,N_35893,N_35894,N_35895,N_35896,N_35897,N_35898,N_35899,N_35900,N_35901,N_35902,N_35903,N_35904,N_35905,N_35906,N_35907,N_35908,N_35909,N_35910,N_35911,N_35912,N_35913,N_35914,N_35915,N_35916,N_35917,N_35918,N_35919,N_35920,N_35921,N_35922,N_35923,N_35924,N_35925,N_35926,N_35927,N_35928,N_35929,N_35930,N_35931,N_35932,N_35933,N_35934,N_35935,N_35936,N_35937,N_35938,N_35939,N_35940,N_35941,N_35942,N_35943,N_35944,N_35945,N_35946,N_35947,N_35948,N_35949,N_35950,N_35951,N_35952,N_35953,N_35954,N_35955,N_35956,N_35957,N_35958,N_35959,N_35960,N_35961,N_35962,N_35963,N_35964,N_35965,N_35966,N_35967,N_35968,N_35969,N_35970,N_35971,N_35972,N_35973,N_35974,N_35975,N_35976,N_35977,N_35978,N_35979,N_35980,N_35981,N_35982,N_35983,N_35984,N_35985,N_35986,N_35987,N_35988,N_35989,N_35990,N_35991,N_35992,N_35993,N_35994,N_35995,N_35996,N_35997,N_35998,N_35999,N_36000,N_36001,N_36002,N_36003,N_36004,N_36005,N_36006,N_36007,N_36008,N_36009,N_36010,N_36011,N_36012,N_36013,N_36014,N_36015,N_36016,N_36017,N_36018,N_36019,N_36020,N_36021,N_36022,N_36023,N_36024,N_36025,N_36026,N_36027,N_36028,N_36029,N_36030,N_36031,N_36032,N_36033,N_36034,N_36035,N_36036,N_36037,N_36038,N_36039,N_36040,N_36041,N_36042,N_36043,N_36044,N_36045,N_36046,N_36047,N_36048,N_36049,N_36050,N_36051,N_36052,N_36053,N_36054,N_36055,N_36056,N_36057,N_36058,N_36059,N_36060,N_36061,N_36062,N_36063,N_36064,N_36065,N_36066,N_36067,N_36068,N_36069,N_36070,N_36071,N_36072,N_36073,N_36074,N_36075,N_36076,N_36077,N_36078,N_36079,N_36080,N_36081,N_36082,N_36083,N_36084,N_36085,N_36086,N_36087,N_36088,N_36089,N_36090,N_36091,N_36092,N_36093,N_36094,N_36095,N_36096,N_36097,N_36098,N_36099,N_36100,N_36101,N_36102,N_36103,N_36104,N_36105,N_36106,N_36107,N_36108,N_36109,N_36110,N_36111,N_36112,N_36113,N_36114,N_36115,N_36116,N_36117,N_36118,N_36119,N_36120,N_36121,N_36122,N_36123,N_36124,N_36125,N_36126,N_36127,N_36128,N_36129,N_36130,N_36131,N_36132,N_36133,N_36134,N_36135,N_36136,N_36137,N_36138,N_36139,N_36140,N_36141,N_36142,N_36143,N_36144,N_36145,N_36146,N_36147,N_36148,N_36149,N_36150,N_36151,N_36152,N_36153,N_36154,N_36155,N_36156,N_36157,N_36158,N_36159,N_36160,N_36161,N_36162,N_36163,N_36164,N_36165,N_36166,N_36167,N_36168,N_36169,N_36170,N_36171,N_36172,N_36173,N_36174,N_36175,N_36176,N_36177,N_36178,N_36179,N_36180,N_36181,N_36182,N_36183,N_36184,N_36185,N_36186,N_36187,N_36188,N_36189,N_36190,N_36191,N_36192,N_36193,N_36194,N_36195,N_36196,N_36197,N_36198,N_36199,N_36200,N_36201,N_36202,N_36203,N_36204,N_36205,N_36206,N_36207,N_36208,N_36209,N_36210,N_36211,N_36212,N_36213,N_36214,N_36215,N_36216,N_36217,N_36218,N_36219,N_36220,N_36221,N_36222,N_36223,N_36224,N_36225,N_36226,N_36227,N_36228,N_36229,N_36230,N_36231,N_36232,N_36233,N_36234,N_36235,N_36236,N_36237,N_36238,N_36239,N_36240,N_36241,N_36242,N_36243,N_36244,N_36245,N_36246,N_36247,N_36248,N_36249,N_36250,N_36251,N_36252,N_36253,N_36254,N_36255,N_36256,N_36257,N_36258,N_36259,N_36260,N_36261,N_36262,N_36263,N_36264,N_36265,N_36266,N_36267,N_36268,N_36269,N_36270,N_36271,N_36272,N_36273,N_36274,N_36275,N_36276,N_36277,N_36278,N_36279,N_36280,N_36281,N_36282,N_36283,N_36284,N_36285,N_36286,N_36287,N_36288,N_36289,N_36290,N_36291,N_36292,N_36293,N_36294,N_36295,N_36296,N_36297,N_36298,N_36299,N_36300,N_36301,N_36302,N_36303,N_36304,N_36305,N_36306,N_36307,N_36308,N_36309,N_36310,N_36311,N_36312,N_36313,N_36314,N_36315,N_36316,N_36317,N_36318,N_36319,N_36320,N_36321,N_36322,N_36323,N_36324,N_36325,N_36326,N_36327,N_36328,N_36329,N_36330,N_36331,N_36332,N_36333,N_36334,N_36335,N_36336,N_36337,N_36338,N_36339,N_36340,N_36341,N_36342,N_36343,N_36344,N_36345,N_36346,N_36347,N_36348,N_36349,N_36350,N_36351,N_36352,N_36353,N_36354,N_36355,N_36356,N_36357,N_36358,N_36359,N_36360,N_36361,N_36362,N_36363,N_36364,N_36365,N_36366,N_36367,N_36368,N_36369,N_36370,N_36371,N_36372,N_36373,N_36374,N_36375,N_36376,N_36377,N_36378,N_36379,N_36380,N_36381,N_36382,N_36383,N_36384,N_36385,N_36386,N_36387,N_36388,N_36389,N_36390,N_36391,N_36392,N_36393,N_36394,N_36395,N_36396,N_36397,N_36398,N_36399,N_36400,N_36401,N_36402,N_36403,N_36404,N_36405,N_36406,N_36407,N_36408,N_36409,N_36410,N_36411,N_36412,N_36413,N_36414,N_36415,N_36416,N_36417,N_36418,N_36419,N_36420,N_36421,N_36422,N_36423,N_36424,N_36425,N_36426,N_36427,N_36428,N_36429,N_36430,N_36431,N_36432,N_36433,N_36434,N_36435,N_36436,N_36437,N_36438,N_36439,N_36440,N_36441,N_36442,N_36443,N_36444,N_36445,N_36446,N_36447,N_36448,N_36449,N_36450,N_36451,N_36452,N_36453,N_36454,N_36455,N_36456,N_36457,N_36458,N_36459,N_36460,N_36461,N_36462,N_36463,N_36464,N_36465,N_36466,N_36467,N_36468,N_36469,N_36470,N_36471,N_36472,N_36473,N_36474,N_36475,N_36476,N_36477,N_36478,N_36479,N_36480,N_36481,N_36482,N_36483,N_36484,N_36485,N_36486,N_36487,N_36488,N_36489,N_36490,N_36491,N_36492,N_36493,N_36494,N_36495,N_36496,N_36497,N_36498,N_36499,N_36500,N_36501,N_36502,N_36503,N_36504,N_36505,N_36506,N_36507,N_36508,N_36509,N_36510,N_36511,N_36512,N_36513,N_36514,N_36515,N_36516,N_36517,N_36518,N_36519,N_36520,N_36521,N_36522,N_36523,N_36524,N_36525,N_36526,N_36527,N_36528,N_36529,N_36530,N_36531,N_36532,N_36533,N_36534,N_36535,N_36536,N_36537,N_36538,N_36539,N_36540,N_36541,N_36542,N_36543,N_36544,N_36545,N_36546,N_36547,N_36548,N_36549,N_36550,N_36551,N_36552,N_36553,N_36554,N_36555,N_36556,N_36557,N_36558,N_36559,N_36560,N_36561,N_36562,N_36563,N_36564,N_36565,N_36566,N_36567,N_36568,N_36569,N_36570,N_36571,N_36572,N_36573,N_36574,N_36575,N_36576,N_36577,N_36578,N_36579,N_36580,N_36581,N_36582,N_36583,N_36584,N_36585,N_36586,N_36587,N_36588,N_36589,N_36590,N_36591,N_36592,N_36593,N_36594,N_36595,N_36596,N_36597,N_36598,N_36599,N_36600,N_36601,N_36602,N_36603,N_36604,N_36605,N_36606,N_36607,N_36608,N_36609,N_36610,N_36611,N_36612,N_36613,N_36614,N_36615,N_36616,N_36617,N_36618,N_36619,N_36620,N_36621,N_36622,N_36623,N_36624,N_36625,N_36626,N_36627,N_36628,N_36629,N_36630,N_36631,N_36632,N_36633,N_36634,N_36635,N_36636,N_36637,N_36638,N_36639,N_36640,N_36641,N_36642,N_36643,N_36644,N_36645,N_36646,N_36647,N_36648,N_36649,N_36650,N_36651,N_36652,N_36653,N_36654,N_36655,N_36656,N_36657,N_36658,N_36659,N_36660,N_36661,N_36662,N_36663,N_36664,N_36665,N_36666,N_36667,N_36668,N_36669,N_36670,N_36671,N_36672,N_36673,N_36674,N_36675,N_36676,N_36677,N_36678,N_36679,N_36680,N_36681,N_36682,N_36683,N_36684,N_36685,N_36686,N_36687,N_36688,N_36689,N_36690,N_36691,N_36692,N_36693,N_36694,N_36695,N_36696,N_36697,N_36698,N_36699,N_36700,N_36701,N_36702,N_36703,N_36704,N_36705,N_36706,N_36707,N_36708,N_36709,N_36710,N_36711,N_36712,N_36713,N_36714,N_36715,N_36716,N_36717,N_36718,N_36719,N_36720,N_36721,N_36722,N_36723,N_36724,N_36725,N_36726,N_36727,N_36728,N_36729,N_36730,N_36731,N_36732,N_36733,N_36734,N_36735,N_36736,N_36737,N_36738,N_36739,N_36740,N_36741,N_36742,N_36743,N_36744,N_36745,N_36746,N_36747,N_36748,N_36749,N_36750,N_36751,N_36752,N_36753,N_36754,N_36755,N_36756,N_36757,N_36758,N_36759,N_36760,N_36761,N_36762,N_36763,N_36764,N_36765,N_36766,N_36767,N_36768,N_36769,N_36770,N_36771,N_36772,N_36773,N_36774,N_36775,N_36776,N_36777,N_36778,N_36779,N_36780,N_36781,N_36782,N_36783,N_36784,N_36785,N_36786,N_36787,N_36788,N_36789,N_36790,N_36791,N_36792,N_36793,N_36794,N_36795,N_36796,N_36797,N_36798,N_36799,N_36800,N_36801,N_36802,N_36803,N_36804,N_36805,N_36806,N_36807,N_36808,N_36809,N_36810,N_36811,N_36812,N_36813,N_36814,N_36815,N_36816,N_36817,N_36818,N_36819,N_36820,N_36821,N_36822,N_36823,N_36824,N_36825,N_36826,N_36827,N_36828,N_36829,N_36830,N_36831,N_36832,N_36833,N_36834,N_36835,N_36836,N_36837,N_36838,N_36839,N_36840,N_36841,N_36842,N_36843,N_36844,N_36845,N_36846,N_36847,N_36848,N_36849,N_36850,N_36851,N_36852,N_36853,N_36854,N_36855,N_36856,N_36857,N_36858,N_36859,N_36860,N_36861,N_36862,N_36863,N_36864,N_36865,N_36866,N_36867,N_36868,N_36869,N_36870,N_36871,N_36872,N_36873,N_36874,N_36875,N_36876,N_36877,N_36878,N_36879,N_36880,N_36881,N_36882,N_36883,N_36884,N_36885,N_36886,N_36887,N_36888,N_36889,N_36890,N_36891,N_36892,N_36893,N_36894,N_36895,N_36896,N_36897,N_36898,N_36899,N_36900,N_36901,N_36902,N_36903,N_36904,N_36905,N_36906,N_36907,N_36908,N_36909,N_36910,N_36911,N_36912,N_36913,N_36914,N_36915,N_36916,N_36917,N_36918,N_36919,N_36920,N_36921,N_36922,N_36923,N_36924,N_36925,N_36926,N_36927,N_36928,N_36929,N_36930,N_36931,N_36932,N_36933,N_36934,N_36935,N_36936,N_36937,N_36938,N_36939,N_36940,N_36941,N_36942,N_36943,N_36944,N_36945,N_36946,N_36947,N_36948,N_36949,N_36950,N_36951,N_36952,N_36953,N_36954,N_36955,N_36956,N_36957,N_36958,N_36959,N_36960,N_36961,N_36962,N_36963,N_36964,N_36965,N_36966,N_36967,N_36968,N_36969,N_36970,N_36971,N_36972,N_36973,N_36974,N_36975,N_36976,N_36977,N_36978,N_36979,N_36980,N_36981,N_36982,N_36983,N_36984,N_36985,N_36986,N_36987,N_36988,N_36989,N_36990,N_36991,N_36992,N_36993,N_36994,N_36995,N_36996,N_36997,N_36998,N_36999,N_37000,N_37001,N_37002,N_37003,N_37004,N_37005,N_37006,N_37007,N_37008,N_37009,N_37010,N_37011,N_37012,N_37013,N_37014,N_37015,N_37016,N_37017,N_37018,N_37019,N_37020,N_37021,N_37022,N_37023,N_37024,N_37025,N_37026,N_37027,N_37028,N_37029,N_37030,N_37031,N_37032,N_37033,N_37034,N_37035,N_37036,N_37037,N_37038,N_37039,N_37040,N_37041,N_37042,N_37043,N_37044,N_37045,N_37046,N_37047,N_37048,N_37049,N_37050,N_37051,N_37052,N_37053,N_37054,N_37055,N_37056,N_37057,N_37058,N_37059,N_37060,N_37061,N_37062,N_37063,N_37064,N_37065,N_37066,N_37067,N_37068,N_37069,N_37070,N_37071,N_37072,N_37073,N_37074,N_37075,N_37076,N_37077,N_37078,N_37079,N_37080,N_37081,N_37082,N_37083,N_37084,N_37085,N_37086,N_37087,N_37088,N_37089,N_37090,N_37091,N_37092,N_37093,N_37094,N_37095,N_37096,N_37097,N_37098,N_37099,N_37100,N_37101,N_37102,N_37103,N_37104,N_37105,N_37106,N_37107,N_37108,N_37109,N_37110,N_37111,N_37112,N_37113,N_37114,N_37115,N_37116,N_37117,N_37118,N_37119,N_37120,N_37121,N_37122,N_37123,N_37124,N_37125,N_37126,N_37127,N_37128,N_37129,N_37130,N_37131,N_37132,N_37133,N_37134,N_37135,N_37136,N_37137,N_37138,N_37139,N_37140,N_37141,N_37142,N_37143,N_37144,N_37145,N_37146,N_37147,N_37148,N_37149,N_37150,N_37151,N_37152,N_37153,N_37154,N_37155,N_37156,N_37157,N_37158,N_37159,N_37160,N_37161,N_37162,N_37163,N_37164,N_37165,N_37166,N_37167,N_37168,N_37169,N_37170,N_37171,N_37172,N_37173,N_37174,N_37175,N_37176,N_37177,N_37178,N_37179,N_37180,N_37181,N_37182,N_37183,N_37184,N_37185,N_37186,N_37187,N_37188,N_37189,N_37190,N_37191,N_37192,N_37193,N_37194,N_37195,N_37196,N_37197,N_37198,N_37199,N_37200,N_37201,N_37202,N_37203,N_37204,N_37205,N_37206,N_37207,N_37208,N_37209,N_37210,N_37211,N_37212,N_37213,N_37214,N_37215,N_37216,N_37217,N_37218,N_37219,N_37220,N_37221,N_37222,N_37223,N_37224,N_37225,N_37226,N_37227,N_37228,N_37229,N_37230,N_37231,N_37232,N_37233,N_37234,N_37235,N_37236,N_37237,N_37238,N_37239,N_37240,N_37241,N_37242,N_37243,N_37244,N_37245,N_37246,N_37247,N_37248,N_37249,N_37250,N_37251,N_37252,N_37253,N_37254,N_37255,N_37256,N_37257,N_37258,N_37259,N_37260,N_37261,N_37262,N_37263,N_37264,N_37265,N_37266,N_37267,N_37268,N_37269,N_37270,N_37271,N_37272,N_37273,N_37274,N_37275,N_37276,N_37277,N_37278,N_37279,N_37280,N_37281,N_37282,N_37283,N_37284,N_37285,N_37286,N_37287,N_37288,N_37289,N_37290,N_37291,N_37292,N_37293,N_37294,N_37295,N_37296,N_37297,N_37298,N_37299,N_37300,N_37301,N_37302,N_37303,N_37304,N_37305,N_37306,N_37307,N_37308,N_37309,N_37310,N_37311,N_37312,N_37313,N_37314,N_37315,N_37316,N_37317,N_37318,N_37319,N_37320,N_37321,N_37322,N_37323,N_37324,N_37325,N_37326,N_37327,N_37328,N_37329,N_37330,N_37331,N_37332,N_37333,N_37334,N_37335,N_37336,N_37337,N_37338,N_37339,N_37340,N_37341,N_37342,N_37343,N_37344,N_37345,N_37346,N_37347,N_37348,N_37349,N_37350,N_37351,N_37352,N_37353,N_37354,N_37355,N_37356,N_37357,N_37358,N_37359,N_37360,N_37361,N_37362,N_37363,N_37364,N_37365,N_37366,N_37367,N_37368,N_37369,N_37370,N_37371,N_37372,N_37373,N_37374,N_37375,N_37376,N_37377,N_37378,N_37379,N_37380,N_37381,N_37382,N_37383,N_37384,N_37385,N_37386,N_37387,N_37388,N_37389,N_37390,N_37391,N_37392,N_37393,N_37394,N_37395,N_37396,N_37397,N_37398,N_37399,N_37400,N_37401,N_37402,N_37403,N_37404,N_37405,N_37406,N_37407,N_37408,N_37409,N_37410,N_37411,N_37412,N_37413,N_37414,N_37415,N_37416,N_37417,N_37418,N_37419,N_37420,N_37421,N_37422,N_37423,N_37424,N_37425,N_37426,N_37427,N_37428,N_37429,N_37430,N_37431,N_37432,N_37433,N_37434,N_37435,N_37436,N_37437,N_37438,N_37439,N_37440,N_37441,N_37442,N_37443,N_37444,N_37445,N_37446,N_37447,N_37448,N_37449,N_37450,N_37451,N_37452,N_37453,N_37454,N_37455,N_37456,N_37457,N_37458,N_37459,N_37460,N_37461,N_37462,N_37463,N_37464,N_37465,N_37466,N_37467,N_37468,N_37469,N_37470,N_37471,N_37472,N_37473,N_37474,N_37475,N_37476,N_37477,N_37478,N_37479,N_37480,N_37481,N_37482,N_37483,N_37484,N_37485,N_37486,N_37487,N_37488,N_37489,N_37490,N_37491,N_37492,N_37493,N_37494,N_37495,N_37496,N_37497,N_37498,N_37499,N_37500,N_37501,N_37502,N_37503,N_37504,N_37505,N_37506,N_37507,N_37508,N_37509,N_37510,N_37511,N_37512,N_37513,N_37514,N_37515,N_37516,N_37517,N_37518,N_37519,N_37520,N_37521,N_37522,N_37523,N_37524,N_37525,N_37526,N_37527,N_37528,N_37529,N_37530,N_37531,N_37532,N_37533,N_37534,N_37535,N_37536,N_37537,N_37538,N_37539,N_37540,N_37541,N_37542,N_37543,N_37544,N_37545,N_37546,N_37547,N_37548,N_37549,N_37550,N_37551,N_37552,N_37553,N_37554,N_37555,N_37556,N_37557,N_37558,N_37559,N_37560,N_37561,N_37562,N_37563,N_37564,N_37565,N_37566,N_37567,N_37568,N_37569,N_37570,N_37571,N_37572,N_37573,N_37574,N_37575,N_37576,N_37577,N_37578,N_37579,N_37580,N_37581,N_37582,N_37583,N_37584,N_37585,N_37586,N_37587,N_37588,N_37589,N_37590,N_37591,N_37592,N_37593,N_37594,N_37595,N_37596,N_37597,N_37598,N_37599,N_37600,N_37601,N_37602,N_37603,N_37604,N_37605,N_37606,N_37607,N_37608,N_37609,N_37610,N_37611,N_37612,N_37613,N_37614,N_37615,N_37616,N_37617,N_37618,N_37619,N_37620,N_37621,N_37622,N_37623,N_37624,N_37625,N_37626,N_37627,N_37628,N_37629,N_37630,N_37631,N_37632,N_37633,N_37634,N_37635,N_37636,N_37637,N_37638,N_37639,N_37640,N_37641,N_37642,N_37643,N_37644,N_37645,N_37646,N_37647,N_37648,N_37649,N_37650,N_37651,N_37652,N_37653,N_37654,N_37655,N_37656,N_37657,N_37658,N_37659,N_37660,N_37661,N_37662,N_37663,N_37664,N_37665,N_37666,N_37667,N_37668,N_37669,N_37670,N_37671,N_37672,N_37673,N_37674,N_37675,N_37676,N_37677,N_37678,N_37679,N_37680,N_37681,N_37682,N_37683,N_37684,N_37685,N_37686,N_37687,N_37688,N_37689,N_37690,N_37691,N_37692,N_37693,N_37694,N_37695,N_37696,N_37697,N_37698,N_37699,N_37700,N_37701,N_37702,N_37703,N_37704,N_37705,N_37706,N_37707,N_37708,N_37709,N_37710,N_37711,N_37712,N_37713,N_37714,N_37715,N_37716,N_37717,N_37718,N_37719,N_37720,N_37721,N_37722,N_37723,N_37724,N_37725,N_37726,N_37727,N_37728,N_37729,N_37730,N_37731,N_37732,N_37733,N_37734,N_37735,N_37736,N_37737,N_37738,N_37739,N_37740,N_37741,N_37742,N_37743,N_37744,N_37745,N_37746,N_37747,N_37748,N_37749,N_37750,N_37751,N_37752,N_37753,N_37754,N_37755,N_37756,N_37757,N_37758,N_37759,N_37760,N_37761,N_37762,N_37763,N_37764,N_37765,N_37766,N_37767,N_37768,N_37769,N_37770,N_37771,N_37772,N_37773,N_37774,N_37775,N_37776,N_37777,N_37778,N_37779,N_37780,N_37781,N_37782,N_37783,N_37784,N_37785,N_37786,N_37787,N_37788,N_37789,N_37790,N_37791,N_37792,N_37793,N_37794,N_37795,N_37796,N_37797,N_37798,N_37799,N_37800,N_37801,N_37802,N_37803,N_37804,N_37805,N_37806,N_37807,N_37808,N_37809,N_37810,N_37811,N_37812,N_37813,N_37814,N_37815,N_37816,N_37817,N_37818,N_37819,N_37820,N_37821,N_37822,N_37823,N_37824,N_37825,N_37826,N_37827,N_37828,N_37829,N_37830,N_37831,N_37832,N_37833,N_37834,N_37835,N_37836,N_37837,N_37838,N_37839,N_37840,N_37841,N_37842,N_37843,N_37844,N_37845,N_37846,N_37847,N_37848,N_37849,N_37850,N_37851,N_37852,N_37853,N_37854,N_37855,N_37856,N_37857,N_37858,N_37859,N_37860,N_37861,N_37862,N_37863,N_37864,N_37865,N_37866,N_37867,N_37868,N_37869,N_37870,N_37871,N_37872,N_37873,N_37874,N_37875,N_37876,N_37877,N_37878,N_37879,N_37880,N_37881,N_37882,N_37883,N_37884,N_37885,N_37886,N_37887,N_37888,N_37889,N_37890,N_37891,N_37892,N_37893,N_37894,N_37895,N_37896,N_37897,N_37898,N_37899,N_37900,N_37901,N_37902,N_37903,N_37904,N_37905,N_37906,N_37907,N_37908,N_37909,N_37910,N_37911,N_37912,N_37913,N_37914,N_37915,N_37916,N_37917,N_37918,N_37919,N_37920,N_37921,N_37922,N_37923,N_37924,N_37925,N_37926,N_37927,N_37928,N_37929,N_37930,N_37931,N_37932,N_37933,N_37934,N_37935,N_37936,N_37937,N_37938,N_37939,N_37940,N_37941,N_37942,N_37943,N_37944,N_37945,N_37946,N_37947,N_37948,N_37949,N_37950,N_37951,N_37952,N_37953,N_37954,N_37955,N_37956,N_37957,N_37958,N_37959,N_37960,N_37961,N_37962,N_37963,N_37964,N_37965,N_37966,N_37967,N_37968,N_37969,N_37970,N_37971,N_37972,N_37973,N_37974,N_37975,N_37976,N_37977,N_37978,N_37979,N_37980,N_37981,N_37982,N_37983,N_37984,N_37985,N_37986,N_37987,N_37988,N_37989,N_37990,N_37991,N_37992,N_37993,N_37994,N_37995,N_37996,N_37997,N_37998,N_37999,N_38000,N_38001,N_38002,N_38003,N_38004,N_38005,N_38006,N_38007,N_38008,N_38009,N_38010,N_38011,N_38012,N_38013,N_38014,N_38015,N_38016,N_38017,N_38018,N_38019,N_38020,N_38021,N_38022,N_38023,N_38024,N_38025,N_38026,N_38027,N_38028,N_38029,N_38030,N_38031,N_38032,N_38033,N_38034,N_38035,N_38036,N_38037,N_38038,N_38039,N_38040,N_38041,N_38042,N_38043,N_38044,N_38045,N_38046,N_38047,N_38048,N_38049,N_38050,N_38051,N_38052,N_38053,N_38054,N_38055,N_38056,N_38057,N_38058,N_38059,N_38060,N_38061,N_38062,N_38063,N_38064,N_38065,N_38066,N_38067,N_38068,N_38069,N_38070,N_38071,N_38072,N_38073,N_38074,N_38075,N_38076,N_38077,N_38078,N_38079,N_38080,N_38081,N_38082,N_38083,N_38084,N_38085,N_38086,N_38087,N_38088,N_38089,N_38090,N_38091,N_38092,N_38093,N_38094,N_38095,N_38096,N_38097,N_38098,N_38099,N_38100,N_38101,N_38102,N_38103,N_38104,N_38105,N_38106,N_38107,N_38108,N_38109,N_38110,N_38111,N_38112,N_38113,N_38114,N_38115,N_38116,N_38117,N_38118,N_38119,N_38120,N_38121,N_38122,N_38123,N_38124,N_38125,N_38126,N_38127,N_38128,N_38129,N_38130,N_38131,N_38132,N_38133,N_38134,N_38135,N_38136,N_38137,N_38138,N_38139,N_38140,N_38141,N_38142,N_38143,N_38144,N_38145,N_38146,N_38147,N_38148,N_38149,N_38150,N_38151,N_38152,N_38153,N_38154,N_38155,N_38156,N_38157,N_38158,N_38159,N_38160,N_38161,N_38162,N_38163,N_38164,N_38165,N_38166,N_38167,N_38168,N_38169,N_38170,N_38171,N_38172,N_38173,N_38174,N_38175,N_38176,N_38177,N_38178,N_38179,N_38180,N_38181,N_38182,N_38183,N_38184,N_38185,N_38186,N_38187,N_38188,N_38189,N_38190,N_38191,N_38192,N_38193,N_38194,N_38195,N_38196,N_38197,N_38198,N_38199,N_38200,N_38201,N_38202,N_38203,N_38204,N_38205,N_38206,N_38207,N_38208,N_38209,N_38210,N_38211,N_38212,N_38213,N_38214,N_38215,N_38216,N_38217,N_38218,N_38219,N_38220,N_38221,N_38222,N_38223,N_38224,N_38225,N_38226,N_38227,N_38228,N_38229,N_38230,N_38231,N_38232,N_38233,N_38234,N_38235,N_38236,N_38237,N_38238,N_38239,N_38240,N_38241,N_38242,N_38243,N_38244,N_38245,N_38246,N_38247,N_38248,N_38249,N_38250,N_38251,N_38252,N_38253,N_38254,N_38255,N_38256,N_38257,N_38258,N_38259,N_38260,N_38261,N_38262,N_38263,N_38264,N_38265,N_38266,N_38267,N_38268,N_38269,N_38270,N_38271,N_38272,N_38273,N_38274,N_38275,N_38276,N_38277,N_38278,N_38279,N_38280,N_38281,N_38282,N_38283,N_38284,N_38285,N_38286,N_38287,N_38288,N_38289,N_38290,N_38291,N_38292,N_38293,N_38294,N_38295,N_38296,N_38297,N_38298,N_38299,N_38300,N_38301,N_38302,N_38303,N_38304,N_38305,N_38306,N_38307,N_38308,N_38309,N_38310,N_38311,N_38312,N_38313,N_38314,N_38315,N_38316,N_38317,N_38318,N_38319,N_38320,N_38321,N_38322,N_38323,N_38324,N_38325,N_38326,N_38327,N_38328,N_38329,N_38330,N_38331,N_38332,N_38333,N_38334,N_38335,N_38336,N_38337,N_38338,N_38339,N_38340,N_38341,N_38342,N_38343,N_38344,N_38345,N_38346,N_38347,N_38348,N_38349,N_38350,N_38351,N_38352,N_38353,N_38354,N_38355,N_38356,N_38357,N_38358,N_38359,N_38360,N_38361,N_38362,N_38363,N_38364,N_38365,N_38366,N_38367,N_38368,N_38369,N_38370,N_38371,N_38372,N_38373,N_38374,N_38375,N_38376,N_38377,N_38378,N_38379,N_38380,N_38381,N_38382,N_38383,N_38384,N_38385,N_38386,N_38387,N_38388,N_38389,N_38390,N_38391,N_38392,N_38393,N_38394,N_38395,N_38396,N_38397,N_38398,N_38399,N_38400,N_38401,N_38402,N_38403,N_38404,N_38405,N_38406,N_38407,N_38408,N_38409,N_38410,N_38411,N_38412,N_38413,N_38414,N_38415,N_38416,N_38417,N_38418,N_38419,N_38420,N_38421,N_38422,N_38423,N_38424,N_38425,N_38426,N_38427,N_38428,N_38429,N_38430,N_38431,N_38432,N_38433,N_38434,N_38435,N_38436,N_38437,N_38438,N_38439,N_38440,N_38441,N_38442,N_38443,N_38444,N_38445,N_38446,N_38447,N_38448,N_38449,N_38450,N_38451,N_38452,N_38453,N_38454,N_38455,N_38456,N_38457,N_38458,N_38459,N_38460,N_38461,N_38462,N_38463,N_38464,N_38465,N_38466,N_38467,N_38468,N_38469,N_38470,N_38471,N_38472,N_38473,N_38474,N_38475,N_38476,N_38477,N_38478,N_38479,N_38480,N_38481,N_38482,N_38483,N_38484,N_38485,N_38486,N_38487,N_38488,N_38489,N_38490,N_38491,N_38492,N_38493,N_38494,N_38495,N_38496,N_38497,N_38498,N_38499,N_38500,N_38501,N_38502,N_38503,N_38504,N_38505,N_38506,N_38507,N_38508,N_38509,N_38510,N_38511,N_38512,N_38513,N_38514,N_38515,N_38516,N_38517,N_38518,N_38519,N_38520,N_38521,N_38522,N_38523,N_38524,N_38525,N_38526,N_38527,N_38528,N_38529,N_38530,N_38531,N_38532,N_38533,N_38534,N_38535,N_38536,N_38537,N_38538,N_38539,N_38540,N_38541,N_38542,N_38543,N_38544,N_38545,N_38546,N_38547,N_38548,N_38549,N_38550,N_38551,N_38552,N_38553,N_38554,N_38555,N_38556,N_38557,N_38558,N_38559,N_38560,N_38561,N_38562,N_38563,N_38564,N_38565,N_38566,N_38567,N_38568,N_38569,N_38570,N_38571,N_38572,N_38573,N_38574,N_38575,N_38576,N_38577,N_38578,N_38579,N_38580,N_38581,N_38582,N_38583,N_38584,N_38585,N_38586,N_38587,N_38588,N_38589,N_38590,N_38591,N_38592,N_38593,N_38594,N_38595,N_38596,N_38597,N_38598,N_38599,N_38600,N_38601,N_38602,N_38603,N_38604,N_38605,N_38606,N_38607,N_38608,N_38609,N_38610,N_38611,N_38612,N_38613,N_38614,N_38615,N_38616,N_38617,N_38618,N_38619,N_38620,N_38621,N_38622,N_38623,N_38624,N_38625,N_38626,N_38627,N_38628,N_38629,N_38630,N_38631,N_38632,N_38633,N_38634,N_38635,N_38636,N_38637,N_38638,N_38639,N_38640,N_38641,N_38642,N_38643,N_38644,N_38645,N_38646,N_38647,N_38648,N_38649,N_38650,N_38651,N_38652,N_38653,N_38654,N_38655,N_38656,N_38657,N_38658,N_38659,N_38660,N_38661,N_38662,N_38663,N_38664,N_38665,N_38666,N_38667,N_38668,N_38669,N_38670,N_38671,N_38672,N_38673,N_38674,N_38675,N_38676,N_38677,N_38678,N_38679,N_38680,N_38681,N_38682,N_38683,N_38684,N_38685,N_38686,N_38687,N_38688,N_38689,N_38690,N_38691,N_38692,N_38693,N_38694,N_38695,N_38696,N_38697,N_38698,N_38699,N_38700,N_38701,N_38702,N_38703,N_38704,N_38705,N_38706,N_38707,N_38708,N_38709,N_38710,N_38711,N_38712,N_38713,N_38714,N_38715,N_38716,N_38717,N_38718,N_38719,N_38720,N_38721,N_38722,N_38723,N_38724,N_38725,N_38726,N_38727,N_38728,N_38729,N_38730,N_38731,N_38732,N_38733,N_38734,N_38735,N_38736,N_38737,N_38738,N_38739,N_38740,N_38741,N_38742,N_38743,N_38744,N_38745,N_38746,N_38747,N_38748,N_38749,N_38750,N_38751,N_38752,N_38753,N_38754,N_38755,N_38756,N_38757,N_38758,N_38759,N_38760,N_38761,N_38762,N_38763,N_38764,N_38765,N_38766,N_38767,N_38768,N_38769,N_38770,N_38771,N_38772,N_38773,N_38774,N_38775,N_38776,N_38777,N_38778,N_38779,N_38780,N_38781,N_38782,N_38783,N_38784,N_38785,N_38786,N_38787,N_38788,N_38789,N_38790,N_38791,N_38792,N_38793,N_38794,N_38795,N_38796,N_38797,N_38798,N_38799,N_38800,N_38801,N_38802,N_38803,N_38804,N_38805,N_38806,N_38807,N_38808,N_38809,N_38810,N_38811,N_38812,N_38813,N_38814,N_38815,N_38816,N_38817,N_38818,N_38819,N_38820,N_38821,N_38822,N_38823,N_38824,N_38825,N_38826,N_38827,N_38828,N_38829,N_38830,N_38831,N_38832,N_38833,N_38834,N_38835,N_38836,N_38837,N_38838,N_38839,N_38840,N_38841,N_38842,N_38843,N_38844,N_38845,N_38846,N_38847,N_38848,N_38849,N_38850,N_38851,N_38852,N_38853,N_38854,N_38855,N_38856,N_38857,N_38858,N_38859,N_38860,N_38861,N_38862,N_38863,N_38864,N_38865,N_38866,N_38867,N_38868,N_38869,N_38870,N_38871,N_38872,N_38873,N_38874,N_38875,N_38876,N_38877,N_38878,N_38879,N_38880,N_38881,N_38882,N_38883,N_38884,N_38885,N_38886,N_38887,N_38888,N_38889,N_38890,N_38891,N_38892,N_38893,N_38894,N_38895,N_38896,N_38897,N_38898,N_38899,N_38900,N_38901,N_38902,N_38903,N_38904,N_38905,N_38906,N_38907,N_38908,N_38909,N_38910,N_38911,N_38912,N_38913,N_38914,N_38915,N_38916,N_38917,N_38918,N_38919,N_38920,N_38921,N_38922,N_38923,N_38924,N_38925,N_38926,N_38927,N_38928,N_38929,N_38930,N_38931,N_38932,N_38933,N_38934,N_38935,N_38936,N_38937,N_38938,N_38939,N_38940,N_38941,N_38942,N_38943,N_38944,N_38945,N_38946,N_38947,N_38948,N_38949,N_38950,N_38951,N_38952,N_38953,N_38954,N_38955,N_38956,N_38957,N_38958,N_38959,N_38960,N_38961,N_38962,N_38963,N_38964,N_38965,N_38966,N_38967,N_38968,N_38969,N_38970,N_38971,N_38972,N_38973,N_38974,N_38975,N_38976,N_38977,N_38978,N_38979,N_38980,N_38981,N_38982,N_38983,N_38984,N_38985,N_38986,N_38987,N_38988,N_38989,N_38990,N_38991,N_38992,N_38993,N_38994,N_38995,N_38996,N_38997,N_38998,N_38999,N_39000,N_39001,N_39002,N_39003,N_39004,N_39005,N_39006,N_39007,N_39008,N_39009,N_39010,N_39011,N_39012,N_39013,N_39014,N_39015,N_39016,N_39017,N_39018,N_39019,N_39020,N_39021,N_39022,N_39023,N_39024,N_39025,N_39026,N_39027,N_39028,N_39029,N_39030,N_39031,N_39032,N_39033,N_39034,N_39035,N_39036,N_39037,N_39038,N_39039,N_39040,N_39041,N_39042,N_39043,N_39044,N_39045,N_39046,N_39047,N_39048,N_39049,N_39050,N_39051,N_39052,N_39053,N_39054,N_39055,N_39056,N_39057,N_39058,N_39059,N_39060,N_39061,N_39062,N_39063,N_39064,N_39065,N_39066,N_39067,N_39068,N_39069,N_39070,N_39071,N_39072,N_39073,N_39074,N_39075,N_39076,N_39077,N_39078,N_39079,N_39080,N_39081,N_39082,N_39083,N_39084,N_39085,N_39086,N_39087,N_39088,N_39089,N_39090,N_39091,N_39092,N_39093,N_39094,N_39095,N_39096,N_39097,N_39098,N_39099,N_39100,N_39101,N_39102,N_39103,N_39104,N_39105,N_39106,N_39107,N_39108,N_39109,N_39110,N_39111,N_39112,N_39113,N_39114,N_39115,N_39116,N_39117,N_39118,N_39119,N_39120,N_39121,N_39122,N_39123,N_39124,N_39125,N_39126,N_39127,N_39128,N_39129,N_39130,N_39131,N_39132,N_39133,N_39134,N_39135,N_39136,N_39137,N_39138,N_39139,N_39140,N_39141,N_39142,N_39143,N_39144,N_39145,N_39146,N_39147,N_39148,N_39149,N_39150,N_39151,N_39152,N_39153,N_39154,N_39155,N_39156,N_39157,N_39158,N_39159,N_39160,N_39161,N_39162,N_39163,N_39164,N_39165,N_39166,N_39167,N_39168,N_39169,N_39170,N_39171,N_39172,N_39173,N_39174,N_39175,N_39176,N_39177,N_39178,N_39179,N_39180,N_39181,N_39182,N_39183,N_39184,N_39185,N_39186,N_39187,N_39188,N_39189,N_39190,N_39191,N_39192,N_39193,N_39194,N_39195,N_39196,N_39197,N_39198,N_39199,N_39200,N_39201,N_39202,N_39203,N_39204,N_39205,N_39206,N_39207,N_39208,N_39209,N_39210,N_39211,N_39212,N_39213,N_39214,N_39215,N_39216,N_39217,N_39218,N_39219,N_39220,N_39221,N_39222,N_39223,N_39224,N_39225,N_39226,N_39227,N_39228,N_39229,N_39230,N_39231,N_39232,N_39233,N_39234,N_39235,N_39236,N_39237,N_39238,N_39239,N_39240,N_39241,N_39242,N_39243,N_39244,N_39245,N_39246,N_39247,N_39248,N_39249,N_39250,N_39251,N_39252,N_39253,N_39254,N_39255,N_39256,N_39257,N_39258,N_39259,N_39260,N_39261,N_39262,N_39263,N_39264,N_39265,N_39266,N_39267,N_39268,N_39269,N_39270,N_39271,N_39272,N_39273,N_39274,N_39275,N_39276,N_39277,N_39278,N_39279,N_39280,N_39281,N_39282,N_39283,N_39284,N_39285,N_39286,N_39287,N_39288,N_39289,N_39290,N_39291,N_39292,N_39293,N_39294,N_39295,N_39296,N_39297,N_39298,N_39299,N_39300,N_39301,N_39302,N_39303,N_39304,N_39305,N_39306,N_39307,N_39308,N_39309,N_39310,N_39311,N_39312,N_39313,N_39314,N_39315,N_39316,N_39317,N_39318,N_39319,N_39320,N_39321,N_39322,N_39323,N_39324,N_39325,N_39326,N_39327,N_39328,N_39329,N_39330,N_39331,N_39332,N_39333,N_39334,N_39335,N_39336,N_39337,N_39338,N_39339,N_39340,N_39341,N_39342,N_39343,N_39344,N_39345,N_39346,N_39347,N_39348,N_39349,N_39350,N_39351,N_39352,N_39353,N_39354,N_39355,N_39356,N_39357,N_39358,N_39359,N_39360,N_39361,N_39362,N_39363,N_39364,N_39365,N_39366,N_39367,N_39368,N_39369,N_39370,N_39371,N_39372,N_39373,N_39374,N_39375,N_39376,N_39377,N_39378,N_39379,N_39380,N_39381,N_39382,N_39383,N_39384,N_39385,N_39386,N_39387,N_39388,N_39389,N_39390,N_39391,N_39392,N_39393,N_39394,N_39395,N_39396,N_39397,N_39398,N_39399,N_39400,N_39401,N_39402,N_39403,N_39404,N_39405,N_39406,N_39407,N_39408,N_39409,N_39410,N_39411,N_39412,N_39413,N_39414,N_39415,N_39416,N_39417,N_39418,N_39419,N_39420,N_39421,N_39422,N_39423,N_39424,N_39425,N_39426,N_39427,N_39428,N_39429,N_39430,N_39431,N_39432,N_39433,N_39434,N_39435,N_39436,N_39437,N_39438,N_39439,N_39440,N_39441,N_39442,N_39443,N_39444,N_39445,N_39446,N_39447,N_39448,N_39449,N_39450,N_39451,N_39452,N_39453,N_39454,N_39455,N_39456,N_39457,N_39458,N_39459,N_39460,N_39461,N_39462,N_39463,N_39464,N_39465,N_39466,N_39467,N_39468,N_39469,N_39470,N_39471,N_39472,N_39473,N_39474,N_39475,N_39476,N_39477,N_39478,N_39479,N_39480,N_39481,N_39482,N_39483,N_39484,N_39485,N_39486,N_39487,N_39488,N_39489,N_39490,N_39491,N_39492,N_39493,N_39494,N_39495,N_39496,N_39497,N_39498,N_39499,N_39500,N_39501,N_39502,N_39503,N_39504,N_39505,N_39506,N_39507,N_39508,N_39509,N_39510,N_39511,N_39512,N_39513,N_39514,N_39515,N_39516,N_39517,N_39518,N_39519,N_39520,N_39521,N_39522,N_39523,N_39524,N_39525,N_39526,N_39527,N_39528,N_39529,N_39530,N_39531,N_39532,N_39533,N_39534,N_39535,N_39536,N_39537,N_39538,N_39539,N_39540,N_39541,N_39542,N_39543,N_39544,N_39545,N_39546,N_39547,N_39548,N_39549,N_39550,N_39551,N_39552,N_39553,N_39554,N_39555,N_39556,N_39557,N_39558,N_39559,N_39560,N_39561,N_39562,N_39563,N_39564,N_39565,N_39566,N_39567,N_39568,N_39569,N_39570,N_39571,N_39572,N_39573,N_39574,N_39575,N_39576,N_39577,N_39578,N_39579,N_39580,N_39581,N_39582,N_39583,N_39584,N_39585,N_39586,N_39587,N_39588,N_39589,N_39590,N_39591,N_39592,N_39593,N_39594,N_39595,N_39596,N_39597,N_39598,N_39599,N_39600,N_39601,N_39602,N_39603,N_39604,N_39605,N_39606,N_39607,N_39608,N_39609,N_39610,N_39611,N_39612,N_39613,N_39614,N_39615,N_39616,N_39617,N_39618,N_39619,N_39620,N_39621,N_39622,N_39623,N_39624,N_39625,N_39626,N_39627,N_39628,N_39629,N_39630,N_39631,N_39632,N_39633,N_39634,N_39635,N_39636,N_39637,N_39638,N_39639,N_39640,N_39641,N_39642,N_39643,N_39644,N_39645,N_39646,N_39647,N_39648,N_39649,N_39650,N_39651,N_39652,N_39653,N_39654,N_39655,N_39656,N_39657,N_39658,N_39659,N_39660,N_39661,N_39662,N_39663,N_39664,N_39665,N_39666,N_39667,N_39668,N_39669,N_39670,N_39671,N_39672,N_39673,N_39674,N_39675,N_39676,N_39677,N_39678,N_39679,N_39680,N_39681,N_39682,N_39683,N_39684,N_39685,N_39686,N_39687,N_39688,N_39689,N_39690,N_39691,N_39692,N_39693,N_39694,N_39695,N_39696,N_39697,N_39698,N_39699,N_39700,N_39701,N_39702,N_39703,N_39704,N_39705,N_39706,N_39707,N_39708,N_39709,N_39710,N_39711,N_39712,N_39713,N_39714,N_39715,N_39716,N_39717,N_39718,N_39719,N_39720,N_39721,N_39722,N_39723,N_39724,N_39725,N_39726,N_39727,N_39728,N_39729,N_39730,N_39731,N_39732,N_39733,N_39734,N_39735,N_39736,N_39737,N_39738,N_39739,N_39740,N_39741,N_39742,N_39743,N_39744,N_39745,N_39746,N_39747,N_39748,N_39749,N_39750,N_39751,N_39752,N_39753,N_39754,N_39755,N_39756,N_39757,N_39758,N_39759,N_39760,N_39761,N_39762,N_39763,N_39764,N_39765,N_39766,N_39767,N_39768,N_39769,N_39770,N_39771,N_39772,N_39773,N_39774,N_39775,N_39776,N_39777,N_39778,N_39779,N_39780,N_39781,N_39782,N_39783,N_39784,N_39785,N_39786,N_39787,N_39788,N_39789,N_39790,N_39791,N_39792,N_39793,N_39794,N_39795,N_39796,N_39797,N_39798,N_39799,N_39800,N_39801,N_39802,N_39803,N_39804,N_39805,N_39806,N_39807,N_39808,N_39809,N_39810,N_39811,N_39812,N_39813,N_39814,N_39815,N_39816,N_39817,N_39818,N_39819,N_39820,N_39821,N_39822,N_39823,N_39824,N_39825,N_39826,N_39827,N_39828,N_39829,N_39830,N_39831,N_39832,N_39833,N_39834,N_39835,N_39836,N_39837,N_39838,N_39839,N_39840,N_39841,N_39842,N_39843,N_39844,N_39845,N_39846,N_39847,N_39848,N_39849,N_39850,N_39851,N_39852,N_39853,N_39854,N_39855,N_39856,N_39857,N_39858,N_39859,N_39860,N_39861,N_39862,N_39863,N_39864,N_39865,N_39866,N_39867,N_39868,N_39869,N_39870,N_39871,N_39872,N_39873,N_39874,N_39875,N_39876,N_39877,N_39878,N_39879,N_39880,N_39881,N_39882,N_39883,N_39884,N_39885,N_39886,N_39887,N_39888,N_39889,N_39890,N_39891,N_39892,N_39893,N_39894,N_39895,N_39896,N_39897,N_39898,N_39899,N_39900,N_39901,N_39902,N_39903,N_39904,N_39905,N_39906,N_39907,N_39908,N_39909,N_39910,N_39911,N_39912,N_39913,N_39914,N_39915,N_39916,N_39917,N_39918,N_39919,N_39920,N_39921,N_39922,N_39923,N_39924,N_39925,N_39926,N_39927,N_39928,N_39929,N_39930,N_39931,N_39932,N_39933,N_39934,N_39935,N_39936,N_39937,N_39938,N_39939,N_39940,N_39941,N_39942,N_39943,N_39944,N_39945,N_39946,N_39947,N_39948,N_39949,N_39950,N_39951,N_39952,N_39953,N_39954,N_39955,N_39956,N_39957,N_39958,N_39959,N_39960,N_39961,N_39962,N_39963,N_39964,N_39965,N_39966,N_39967,N_39968,N_39969,N_39970,N_39971,N_39972,N_39973,N_39974,N_39975,N_39976,N_39977,N_39978,N_39979,N_39980,N_39981,N_39982,N_39983,N_39984,N_39985,N_39986,N_39987,N_39988,N_39989,N_39990,N_39991,N_39992,N_39993,N_39994,N_39995,N_39996,N_39997,N_39998,N_39999,N_40000,N_40001,N_40002,N_40003,N_40004,N_40005,N_40006,N_40007,N_40008,N_40009,N_40010,N_40011,N_40012,N_40013,N_40014,N_40015,N_40016,N_40017,N_40018,N_40019,N_40020,N_40021,N_40022,N_40023,N_40024,N_40025,N_40026,N_40027,N_40028,N_40029,N_40030,N_40031,N_40032,N_40033,N_40034,N_40035,N_40036,N_40037,N_40038,N_40039,N_40040,N_40041,N_40042,N_40043,N_40044,N_40045,N_40046,N_40047,N_40048,N_40049,N_40050,N_40051,N_40052,N_40053,N_40054,N_40055,N_40056,N_40057,N_40058,N_40059,N_40060,N_40061,N_40062,N_40063,N_40064,N_40065,N_40066,N_40067,N_40068,N_40069,N_40070,N_40071,N_40072,N_40073,N_40074,N_40075,N_40076,N_40077,N_40078,N_40079,N_40080,N_40081,N_40082,N_40083,N_40084,N_40085,N_40086,N_40087,N_40088,N_40089,N_40090,N_40091,N_40092,N_40093,N_40094,N_40095,N_40096,N_40097,N_40098,N_40099,N_40100,N_40101,N_40102,N_40103,N_40104,N_40105,N_40106,N_40107,N_40108,N_40109,N_40110,N_40111,N_40112,N_40113,N_40114,N_40115,N_40116,N_40117,N_40118,N_40119,N_40120,N_40121,N_40122,N_40123,N_40124,N_40125,N_40126,N_40127,N_40128,N_40129,N_40130,N_40131,N_40132,N_40133,N_40134,N_40135,N_40136,N_40137,N_40138,N_40139,N_40140,N_40141,N_40142,N_40143,N_40144,N_40145,N_40146,N_40147,N_40148,N_40149,N_40150,N_40151,N_40152,N_40153,N_40154,N_40155,N_40156,N_40157,N_40158,N_40159,N_40160,N_40161,N_40162,N_40163,N_40164,N_40165,N_40166,N_40167,N_40168,N_40169,N_40170,N_40171,N_40172,N_40173,N_40174,N_40175,N_40176,N_40177,N_40178,N_40179,N_40180,N_40181,N_40182,N_40183,N_40184,N_40185,N_40186,N_40187,N_40188,N_40189,N_40190,N_40191,N_40192,N_40193,N_40194,N_40195,N_40196,N_40197,N_40198,N_40199,N_40200,N_40201,N_40202,N_40203,N_40204,N_40205,N_40206,N_40207,N_40208,N_40209,N_40210,N_40211,N_40212,N_40213,N_40214,N_40215,N_40216,N_40217,N_40218,N_40219,N_40220,N_40221,N_40222,N_40223,N_40224,N_40225,N_40226,N_40227,N_40228,N_40229,N_40230,N_40231,N_40232,N_40233,N_40234,N_40235,N_40236,N_40237,N_40238,N_40239,N_40240,N_40241,N_40242,N_40243,N_40244,N_40245,N_40246,N_40247,N_40248,N_40249,N_40250,N_40251,N_40252,N_40253,N_40254,N_40255,N_40256,N_40257,N_40258,N_40259,N_40260,N_40261,N_40262,N_40263,N_40264,N_40265,N_40266,N_40267,N_40268,N_40269,N_40270,N_40271,N_40272,N_40273,N_40274,N_40275,N_40276,N_40277,N_40278,N_40279,N_40280,N_40281,N_40282,N_40283,N_40284,N_40285,N_40286,N_40287,N_40288,N_40289,N_40290,N_40291,N_40292,N_40293,N_40294,N_40295,N_40296,N_40297,N_40298,N_40299,N_40300,N_40301,N_40302,N_40303,N_40304,N_40305,N_40306,N_40307,N_40308,N_40309,N_40310,N_40311,N_40312,N_40313,N_40314,N_40315,N_40316,N_40317,N_40318,N_40319,N_40320,N_40321,N_40322,N_40323,N_40324,N_40325,N_40326,N_40327,N_40328,N_40329,N_40330,N_40331,N_40332,N_40333,N_40334,N_40335,N_40336,N_40337,N_40338,N_40339,N_40340,N_40341,N_40342,N_40343,N_40344,N_40345,N_40346,N_40347,N_40348,N_40349,N_40350,N_40351,N_40352,N_40353,N_40354,N_40355,N_40356,N_40357,N_40358,N_40359,N_40360,N_40361,N_40362,N_40363,N_40364,N_40365,N_40366,N_40367,N_40368,N_40369,N_40370,N_40371,N_40372,N_40373,N_40374,N_40375,N_40376,N_40377,N_40378,N_40379,N_40380,N_40381,N_40382,N_40383,N_40384,N_40385,N_40386,N_40387,N_40388,N_40389,N_40390,N_40391,N_40392,N_40393,N_40394,N_40395,N_40396,N_40397,N_40398,N_40399,N_40400,N_40401,N_40402,N_40403,N_40404,N_40405,N_40406,N_40407,N_40408,N_40409,N_40410,N_40411,N_40412,N_40413,N_40414,N_40415,N_40416,N_40417,N_40418,N_40419,N_40420,N_40421,N_40422,N_40423,N_40424,N_40425,N_40426,N_40427,N_40428,N_40429,N_40430,N_40431,N_40432,N_40433,N_40434,N_40435,N_40436,N_40437,N_40438,N_40439,N_40440,N_40441,N_40442,N_40443,N_40444,N_40445,N_40446,N_40447,N_40448,N_40449,N_40450,N_40451,N_40452,N_40453,N_40454,N_40455,N_40456,N_40457,N_40458,N_40459,N_40460,N_40461,N_40462,N_40463,N_40464,N_40465,N_40466,N_40467,N_40468,N_40469,N_40470,N_40471,N_40472,N_40473,N_40474,N_40475,N_40476,N_40477,N_40478,N_40479,N_40480,N_40481,N_40482,N_40483,N_40484,N_40485,N_40486,N_40487,N_40488,N_40489,N_40490,N_40491,N_40492,N_40493,N_40494,N_40495,N_40496,N_40497,N_40498,N_40499,N_40500,N_40501,N_40502,N_40503,N_40504,N_40505,N_40506,N_40507,N_40508,N_40509,N_40510,N_40511,N_40512,N_40513,N_40514,N_40515,N_40516,N_40517,N_40518,N_40519,N_40520,N_40521,N_40522,N_40523,N_40524,N_40525,N_40526,N_40527,N_40528,N_40529,N_40530,N_40531,N_40532,N_40533,N_40534,N_40535,N_40536,N_40537,N_40538,N_40539,N_40540,N_40541,N_40542,N_40543,N_40544,N_40545,N_40546,N_40547,N_40548,N_40549,N_40550,N_40551,N_40552,N_40553,N_40554,N_40555,N_40556,N_40557,N_40558,N_40559,N_40560,N_40561,N_40562,N_40563,N_40564,N_40565,N_40566,N_40567,N_40568,N_40569,N_40570,N_40571,N_40572,N_40573,N_40574,N_40575,N_40576,N_40577,N_40578,N_40579,N_40580,N_40581,N_40582,N_40583,N_40584,N_40585,N_40586,N_40587,N_40588,N_40589,N_40590,N_40591,N_40592,N_40593,N_40594,N_40595,N_40596,N_40597,N_40598,N_40599,N_40600,N_40601,N_40602,N_40603,N_40604,N_40605,N_40606,N_40607,N_40608,N_40609,N_40610,N_40611,N_40612,N_40613,N_40614,N_40615,N_40616,N_40617,N_40618,N_40619,N_40620,N_40621,N_40622,N_40623,N_40624,N_40625,N_40626,N_40627,N_40628,N_40629,N_40630,N_40631,N_40632,N_40633,N_40634,N_40635,N_40636,N_40637,N_40638,N_40639,N_40640,N_40641,N_40642,N_40643,N_40644,N_40645,N_40646,N_40647,N_40648,N_40649,N_40650,N_40651,N_40652,N_40653,N_40654,N_40655,N_40656,N_40657,N_40658,N_40659,N_40660,N_40661,N_40662,N_40663,N_40664,N_40665,N_40666,N_40667,N_40668,N_40669,N_40670,N_40671,N_40672,N_40673,N_40674,N_40675,N_40676,N_40677,N_40678,N_40679,N_40680,N_40681,N_40682,N_40683,N_40684,N_40685,N_40686,N_40687,N_40688,N_40689,N_40690,N_40691,N_40692,N_40693,N_40694,N_40695,N_40696,N_40697,N_40698,N_40699,N_40700,N_40701,N_40702,N_40703,N_40704,N_40705,N_40706,N_40707,N_40708,N_40709,N_40710,N_40711,N_40712,N_40713,N_40714,N_40715,N_40716,N_40717,N_40718,N_40719,N_40720,N_40721,N_40722,N_40723,N_40724,N_40725,N_40726,N_40727,N_40728,N_40729,N_40730,N_40731,N_40732,N_40733,N_40734,N_40735,N_40736,N_40737,N_40738,N_40739,N_40740,N_40741,N_40742,N_40743,N_40744,N_40745,N_40746,N_40747,N_40748,N_40749,N_40750,N_40751,N_40752,N_40753,N_40754,N_40755,N_40756,N_40757,N_40758,N_40759,N_40760,N_40761,N_40762,N_40763,N_40764,N_40765,N_40766,N_40767,N_40768,N_40769,N_40770,N_40771,N_40772,N_40773,N_40774,N_40775,N_40776,N_40777,N_40778,N_40779,N_40780,N_40781,N_40782,N_40783,N_40784,N_40785,N_40786,N_40787,N_40788,N_40789,N_40790,N_40791,N_40792,N_40793,N_40794,N_40795,N_40796,N_40797,N_40798,N_40799,N_40800,N_40801,N_40802,N_40803,N_40804,N_40805,N_40806,N_40807,N_40808,N_40809,N_40810,N_40811,N_40812,N_40813,N_40814,N_40815,N_40816,N_40817,N_40818,N_40819,N_40820,N_40821,N_40822,N_40823,N_40824,N_40825,N_40826,N_40827,N_40828,N_40829,N_40830,N_40831,N_40832,N_40833,N_40834,N_40835,N_40836,N_40837,N_40838,N_40839,N_40840,N_40841,N_40842,N_40843,N_40844,N_40845,N_40846,N_40847,N_40848,N_40849,N_40850,N_40851,N_40852,N_40853,N_40854,N_40855,N_40856,N_40857,N_40858,N_40859,N_40860,N_40861,N_40862,N_40863,N_40864,N_40865,N_40866,N_40867,N_40868,N_40869,N_40870,N_40871,N_40872,N_40873,N_40874,N_40875,N_40876,N_40877,N_40878,N_40879,N_40880,N_40881,N_40882,N_40883,N_40884,N_40885,N_40886,N_40887,N_40888,N_40889,N_40890,N_40891,N_40892,N_40893,N_40894,N_40895,N_40896,N_40897,N_40898,N_40899,N_40900,N_40901,N_40902,N_40903,N_40904,N_40905,N_40906,N_40907,N_40908,N_40909,N_40910,N_40911,N_40912,N_40913,N_40914,N_40915,N_40916,N_40917,N_40918,N_40919,N_40920,N_40921,N_40922,N_40923,N_40924,N_40925,N_40926,N_40927,N_40928,N_40929,N_40930,N_40931,N_40932,N_40933,N_40934,N_40935,N_40936,N_40937,N_40938,N_40939,N_40940,N_40941,N_40942,N_40943,N_40944,N_40945,N_40946,N_40947,N_40948,N_40949,N_40950,N_40951,N_40952,N_40953,N_40954,N_40955,N_40956,N_40957,N_40958,N_40959,N_40960,N_40961,N_40962,N_40963,N_40964,N_40965,N_40966,N_40967,N_40968,N_40969,N_40970,N_40971,N_40972,N_40973,N_40974,N_40975,N_40976,N_40977,N_40978,N_40979,N_40980,N_40981,N_40982,N_40983,N_40984,N_40985,N_40986,N_40987,N_40988,N_40989,N_40990,N_40991,N_40992,N_40993,N_40994,N_40995,N_40996,N_40997,N_40998,N_40999,N_41000,N_41001,N_41002,N_41003,N_41004,N_41005,N_41006,N_41007,N_41008,N_41009,N_41010,N_41011,N_41012,N_41013,N_41014,N_41015,N_41016,N_41017,N_41018,N_41019,N_41020,N_41021,N_41022,N_41023,N_41024,N_41025,N_41026,N_41027,N_41028,N_41029,N_41030,N_41031,N_41032,N_41033,N_41034,N_41035,N_41036,N_41037,N_41038,N_41039,N_41040,N_41041,N_41042,N_41043,N_41044,N_41045,N_41046,N_41047,N_41048,N_41049,N_41050,N_41051,N_41052,N_41053,N_41054,N_41055,N_41056,N_41057,N_41058,N_41059,N_41060,N_41061,N_41062,N_41063,N_41064,N_41065,N_41066,N_41067,N_41068,N_41069,N_41070,N_41071,N_41072,N_41073,N_41074,N_41075,N_41076,N_41077,N_41078,N_41079,N_41080,N_41081,N_41082,N_41083,N_41084,N_41085,N_41086,N_41087,N_41088,N_41089,N_41090,N_41091,N_41092,N_41093,N_41094,N_41095,N_41096,N_41097,N_41098,N_41099,N_41100,N_41101,N_41102,N_41103,N_41104,N_41105,N_41106,N_41107,N_41108,N_41109,N_41110,N_41111,N_41112,N_41113,N_41114,N_41115,N_41116,N_41117,N_41118,N_41119,N_41120,N_41121,N_41122,N_41123,N_41124,N_41125,N_41126,N_41127,N_41128,N_41129,N_41130,N_41131,N_41132,N_41133,N_41134,N_41135,N_41136,N_41137,N_41138,N_41139,N_41140,N_41141,N_41142,N_41143,N_41144,N_41145,N_41146,N_41147,N_41148,N_41149,N_41150,N_41151,N_41152,N_41153,N_41154,N_41155,N_41156,N_41157,N_41158,N_41159,N_41160,N_41161,N_41162,N_41163,N_41164,N_41165,N_41166,N_41167,N_41168,N_41169,N_41170,N_41171,N_41172,N_41173,N_41174,N_41175,N_41176,N_41177,N_41178,N_41179,N_41180,N_41181,N_41182,N_41183,N_41184,N_41185,N_41186,N_41187,N_41188,N_41189,N_41190,N_41191,N_41192,N_41193,N_41194,N_41195,N_41196,N_41197,N_41198,N_41199,N_41200,N_41201,N_41202,N_41203,N_41204,N_41205,N_41206,N_41207,N_41208,N_41209,N_41210,N_41211,N_41212,N_41213,N_41214,N_41215,N_41216,N_41217,N_41218,N_41219,N_41220,N_41221,N_41222,N_41223,N_41224,N_41225,N_41226,N_41227,N_41228,N_41229,N_41230,N_41231,N_41232,N_41233,N_41234,N_41235,N_41236,N_41237,N_41238,N_41239,N_41240,N_41241,N_41242,N_41243,N_41244,N_41245,N_41246,N_41247,N_41248,N_41249,N_41250,N_41251,N_41252,N_41253,N_41254,N_41255,N_41256,N_41257,N_41258,N_41259,N_41260,N_41261,N_41262,N_41263,N_41264,N_41265,N_41266,N_41267,N_41268,N_41269,N_41270,N_41271,N_41272,N_41273,N_41274,N_41275,N_41276,N_41277,N_41278,N_41279,N_41280,N_41281,N_41282,N_41283,N_41284,N_41285,N_41286,N_41287,N_41288,N_41289,N_41290,N_41291,N_41292,N_41293,N_41294,N_41295,N_41296,N_41297,N_41298,N_41299,N_41300,N_41301,N_41302,N_41303,N_41304,N_41305,N_41306,N_41307,N_41308,N_41309,N_41310,N_41311,N_41312,N_41313,N_41314,N_41315,N_41316,N_41317,N_41318,N_41319,N_41320,N_41321,N_41322,N_41323,N_41324,N_41325,N_41326,N_41327,N_41328,N_41329,N_41330,N_41331,N_41332,N_41333,N_41334,N_41335,N_41336,N_41337,N_41338,N_41339,N_41340,N_41341,N_41342,N_41343,N_41344,N_41345,N_41346,N_41347,N_41348,N_41349,N_41350,N_41351,N_41352,N_41353,N_41354,N_41355,N_41356,N_41357,N_41358,N_41359,N_41360,N_41361,N_41362,N_41363,N_41364,N_41365,N_41366,N_41367,N_41368,N_41369,N_41370,N_41371,N_41372,N_41373,N_41374,N_41375,N_41376,N_41377,N_41378,N_41379,N_41380,N_41381,N_41382,N_41383,N_41384,N_41385,N_41386,N_41387,N_41388,N_41389,N_41390,N_41391,N_41392,N_41393,N_41394,N_41395,N_41396,N_41397,N_41398,N_41399,N_41400,N_41401,N_41402,N_41403,N_41404,N_41405,N_41406,N_41407,N_41408,N_41409,N_41410,N_41411,N_41412,N_41413,N_41414,N_41415,N_41416,N_41417,N_41418,N_41419,N_41420,N_41421,N_41422,N_41423,N_41424,N_41425,N_41426,N_41427,N_41428,N_41429,N_41430,N_41431,N_41432,N_41433,N_41434,N_41435,N_41436,N_41437,N_41438,N_41439,N_41440,N_41441,N_41442,N_41443,N_41444,N_41445,N_41446,N_41447,N_41448,N_41449,N_41450,N_41451,N_41452,N_41453,N_41454,N_41455,N_41456,N_41457,N_41458,N_41459,N_41460,N_41461,N_41462,N_41463,N_41464,N_41465,N_41466,N_41467,N_41468,N_41469,N_41470,N_41471,N_41472,N_41473,N_41474,N_41475,N_41476,N_41477,N_41478,N_41479,N_41480,N_41481,N_41482,N_41483,N_41484,N_41485,N_41486,N_41487,N_41488,N_41489,N_41490,N_41491,N_41492,N_41493,N_41494,N_41495,N_41496,N_41497,N_41498,N_41499,N_41500,N_41501,N_41502,N_41503,N_41504,N_41505,N_41506,N_41507,N_41508,N_41509,N_41510,N_41511,N_41512,N_41513,N_41514,N_41515,N_41516,N_41517,N_41518,N_41519,N_41520,N_41521,N_41522,N_41523,N_41524,N_41525,N_41526,N_41527,N_41528,N_41529,N_41530,N_41531,N_41532,N_41533,N_41534,N_41535,N_41536,N_41537,N_41538,N_41539,N_41540,N_41541,N_41542,N_41543,N_41544,N_41545,N_41546,N_41547,N_41548,N_41549,N_41550,N_41551,N_41552,N_41553,N_41554,N_41555,N_41556,N_41557,N_41558,N_41559,N_41560,N_41561,N_41562,N_41563,N_41564,N_41565,N_41566,N_41567,N_41568,N_41569,N_41570,N_41571,N_41572,N_41573,N_41574,N_41575,N_41576,N_41577,N_41578,N_41579,N_41580,N_41581,N_41582,N_41583,N_41584,N_41585,N_41586,N_41587,N_41588,N_41589,N_41590,N_41591,N_41592,N_41593,N_41594,N_41595,N_41596,N_41597,N_41598,N_41599,N_41600,N_41601,N_41602,N_41603,N_41604,N_41605,N_41606,N_41607,N_41608,N_41609,N_41610,N_41611,N_41612,N_41613,N_41614,N_41615,N_41616,N_41617,N_41618,N_41619,N_41620,N_41621,N_41622,N_41623,N_41624,N_41625,N_41626,N_41627,N_41628,N_41629,N_41630,N_41631,N_41632,N_41633,N_41634,N_41635,N_41636,N_41637,N_41638,N_41639,N_41640,N_41641,N_41642,N_41643,N_41644,N_41645,N_41646,N_41647,N_41648,N_41649,N_41650,N_41651,N_41652,N_41653,N_41654,N_41655,N_41656,N_41657,N_41658,N_41659,N_41660,N_41661,N_41662,N_41663,N_41664,N_41665,N_41666,N_41667,N_41668,N_41669,N_41670,N_41671,N_41672,N_41673,N_41674,N_41675,N_41676,N_41677,N_41678,N_41679,N_41680,N_41681,N_41682,N_41683,N_41684,N_41685,N_41686,N_41687,N_41688,N_41689,N_41690,N_41691,N_41692,N_41693,N_41694,N_41695,N_41696,N_41697,N_41698,N_41699,N_41700,N_41701,N_41702,N_41703,N_41704,N_41705,N_41706,N_41707,N_41708,N_41709,N_41710,N_41711,N_41712,N_41713,N_41714,N_41715,N_41716,N_41717,N_41718,N_41719,N_41720,N_41721,N_41722,N_41723,N_41724,N_41725,N_41726,N_41727,N_41728,N_41729,N_41730,N_41731,N_41732,N_41733,N_41734,N_41735,N_41736,N_41737,N_41738,N_41739,N_41740,N_41741,N_41742,N_41743,N_41744,N_41745,N_41746,N_41747,N_41748,N_41749,N_41750,N_41751,N_41752,N_41753,N_41754,N_41755,N_41756,N_41757,N_41758,N_41759,N_41760,N_41761,N_41762,N_41763,N_41764,N_41765,N_41766,N_41767,N_41768,N_41769,N_41770,N_41771,N_41772,N_41773,N_41774,N_41775,N_41776,N_41777,N_41778,N_41779,N_41780,N_41781,N_41782,N_41783,N_41784,N_41785,N_41786,N_41787,N_41788,N_41789,N_41790,N_41791,N_41792,N_41793,N_41794,N_41795,N_41796,N_41797,N_41798,N_41799,N_41800,N_41801,N_41802,N_41803,N_41804,N_41805,N_41806,N_41807,N_41808,N_41809,N_41810,N_41811,N_41812,N_41813,N_41814,N_41815,N_41816,N_41817,N_41818,N_41819,N_41820,N_41821,N_41822,N_41823,N_41824,N_41825,N_41826,N_41827,N_41828,N_41829,N_41830,N_41831,N_41832,N_41833,N_41834,N_41835,N_41836,N_41837,N_41838,N_41839,N_41840,N_41841,N_41842,N_41843,N_41844,N_41845,N_41846,N_41847,N_41848,N_41849,N_41850,N_41851,N_41852,N_41853,N_41854,N_41855,N_41856,N_41857,N_41858,N_41859,N_41860,N_41861,N_41862,N_41863,N_41864,N_41865,N_41866,N_41867,N_41868,N_41869,N_41870,N_41871,N_41872,N_41873,N_41874,N_41875,N_41876,N_41877,N_41878,N_41879,N_41880,N_41881,N_41882,N_41883,N_41884,N_41885,N_41886,N_41887,N_41888,N_41889,N_41890,N_41891,N_41892,N_41893,N_41894,N_41895,N_41896,N_41897,N_41898,N_41899,N_41900,N_41901,N_41902,N_41903,N_41904,N_41905,N_41906,N_41907,N_41908,N_41909,N_41910,N_41911,N_41912,N_41913,N_41914,N_41915,N_41916,N_41917,N_41918,N_41919,N_41920,N_41921,N_41922,N_41923,N_41924,N_41925,N_41926,N_41927,N_41928,N_41929,N_41930,N_41931,N_41932,N_41933,N_41934,N_41935,N_41936,N_41937,N_41938,N_41939,N_41940,N_41941,N_41942,N_41943,N_41944,N_41945,N_41946,N_41947,N_41948,N_41949,N_41950,N_41951,N_41952,N_41953,N_41954,N_41955,N_41956,N_41957,N_41958,N_41959,N_41960,N_41961,N_41962,N_41963,N_41964,N_41965,N_41966,N_41967,N_41968,N_41969,N_41970,N_41971,N_41972,N_41973,N_41974,N_41975,N_41976,N_41977,N_41978,N_41979,N_41980,N_41981,N_41982,N_41983,N_41984,N_41985,N_41986,N_41987,N_41988,N_41989,N_41990,N_41991,N_41992,N_41993,N_41994,N_41995,N_41996,N_41997,N_41998,N_41999,N_42000,N_42001,N_42002,N_42003,N_42004,N_42005,N_42006,N_42007,N_42008,N_42009,N_42010,N_42011,N_42012,N_42013,N_42014,N_42015,N_42016,N_42017,N_42018,N_42019,N_42020,N_42021,N_42022,N_42023,N_42024,N_42025,N_42026,N_42027,N_42028,N_42029,N_42030,N_42031,N_42032,N_42033,N_42034,N_42035,N_42036,N_42037,N_42038,N_42039,N_42040,N_42041,N_42042,N_42043,N_42044,N_42045,N_42046,N_42047,N_42048,N_42049,N_42050,N_42051,N_42052,N_42053,N_42054,N_42055,N_42056,N_42057,N_42058,N_42059,N_42060,N_42061,N_42062,N_42063,N_42064,N_42065,N_42066,N_42067,N_42068,N_42069,N_42070,N_42071,N_42072,N_42073,N_42074,N_42075,N_42076,N_42077,N_42078,N_42079,N_42080,N_42081,N_42082,N_42083,N_42084,N_42085,N_42086,N_42087,N_42088,N_42089,N_42090,N_42091,N_42092,N_42093,N_42094,N_42095,N_42096,N_42097,N_42098,N_42099,N_42100,N_42101,N_42102,N_42103,N_42104,N_42105,N_42106,N_42107,N_42108,N_42109,N_42110,N_42111,N_42112,N_42113,N_42114,N_42115,N_42116,N_42117,N_42118,N_42119,N_42120,N_42121,N_42122,N_42123,N_42124,N_42125,N_42126,N_42127,N_42128,N_42129,N_42130,N_42131,N_42132,N_42133,N_42134,N_42135,N_42136,N_42137,N_42138,N_42139,N_42140,N_42141,N_42142,N_42143,N_42144,N_42145,N_42146,N_42147,N_42148,N_42149,N_42150,N_42151,N_42152,N_42153,N_42154,N_42155,N_42156,N_42157,N_42158,N_42159,N_42160,N_42161,N_42162,N_42163,N_42164,N_42165,N_42166,N_42167,N_42168,N_42169,N_42170,N_42171,N_42172,N_42173,N_42174,N_42175,N_42176,N_42177,N_42178,N_42179,N_42180,N_42181,N_42182,N_42183,N_42184,N_42185,N_42186,N_42187,N_42188,N_42189,N_42190,N_42191,N_42192,N_42193,N_42194,N_42195,N_42196,N_42197,N_42198,N_42199,N_42200,N_42201,N_42202,N_42203,N_42204,N_42205,N_42206,N_42207,N_42208,N_42209,N_42210,N_42211,N_42212,N_42213,N_42214,N_42215,N_42216,N_42217,N_42218,N_42219,N_42220,N_42221,N_42222,N_42223,N_42224,N_42225,N_42226,N_42227,N_42228,N_42229,N_42230,N_42231,N_42232,N_42233,N_42234,N_42235,N_42236,N_42237,N_42238,N_42239,N_42240,N_42241,N_42242,N_42243,N_42244,N_42245,N_42246,N_42247,N_42248,N_42249,N_42250,N_42251,N_42252,N_42253,N_42254,N_42255,N_42256,N_42257,N_42258,N_42259,N_42260,N_42261,N_42262,N_42263,N_42264,N_42265,N_42266,N_42267,N_42268,N_42269,N_42270,N_42271,N_42272,N_42273,N_42274,N_42275,N_42276,N_42277,N_42278,N_42279,N_42280,N_42281,N_42282,N_42283,N_42284,N_42285,N_42286,N_42287,N_42288,N_42289,N_42290,N_42291,N_42292,N_42293,N_42294,N_42295,N_42296,N_42297,N_42298,N_42299,N_42300,N_42301,N_42302,N_42303,N_42304,N_42305,N_42306,N_42307,N_42308,N_42309,N_42310,N_42311,N_42312,N_42313,N_42314,N_42315,N_42316,N_42317,N_42318,N_42319,N_42320,N_42321,N_42322,N_42323,N_42324,N_42325,N_42326,N_42327,N_42328,N_42329,N_42330,N_42331,N_42332,N_42333,N_42334,N_42335,N_42336,N_42337,N_42338,N_42339,N_42340,N_42341,N_42342,N_42343,N_42344,N_42345,N_42346,N_42347,N_42348,N_42349,N_42350,N_42351,N_42352,N_42353,N_42354,N_42355,N_42356,N_42357,N_42358,N_42359,N_42360,N_42361,N_42362,N_42363,N_42364,N_42365,N_42366,N_42367,N_42368,N_42369,N_42370,N_42371,N_42372,N_42373,N_42374,N_42375,N_42376,N_42377,N_42378,N_42379,N_42380,N_42381,N_42382,N_42383,N_42384,N_42385,N_42386,N_42387,N_42388,N_42389,N_42390,N_42391,N_42392,N_42393,N_42394,N_42395,N_42396,N_42397,N_42398,N_42399,N_42400,N_42401,N_42402,N_42403,N_42404,N_42405,N_42406,N_42407,N_42408,N_42409,N_42410,N_42411,N_42412,N_42413,N_42414,N_42415,N_42416,N_42417,N_42418,N_42419,N_42420,N_42421,N_42422,N_42423,N_42424,N_42425,N_42426,N_42427,N_42428,N_42429,N_42430,N_42431,N_42432,N_42433,N_42434,N_42435,N_42436,N_42437,N_42438,N_42439,N_42440,N_42441,N_42442,N_42443,N_42444,N_42445,N_42446,N_42447,N_42448,N_42449,N_42450,N_42451,N_42452,N_42453,N_42454,N_42455,N_42456,N_42457,N_42458,N_42459,N_42460,N_42461,N_42462,N_42463,N_42464,N_42465,N_42466,N_42467,N_42468,N_42469,N_42470,N_42471,N_42472,N_42473,N_42474,N_42475,N_42476,N_42477,N_42478,N_42479,N_42480,N_42481,N_42482,N_42483,N_42484,N_42485,N_42486,N_42487,N_42488,N_42489,N_42490,N_42491,N_42492,N_42493,N_42494,N_42495,N_42496,N_42497,N_42498,N_42499,N_42500,N_42501,N_42502,N_42503,N_42504,N_42505,N_42506,N_42507,N_42508,N_42509,N_42510,N_42511,N_42512,N_42513,N_42514,N_42515,N_42516,N_42517,N_42518,N_42519,N_42520,N_42521,N_42522,N_42523,N_42524,N_42525,N_42526,N_42527,N_42528,N_42529,N_42530,N_42531,N_42532,N_42533,N_42534,N_42535,N_42536,N_42537,N_42538,N_42539,N_42540,N_42541,N_42542,N_42543,N_42544,N_42545,N_42546,N_42547,N_42548,N_42549,N_42550,N_42551,N_42552,N_42553,N_42554,N_42555,N_42556,N_42557,N_42558,N_42559,N_42560,N_42561,N_42562,N_42563,N_42564,N_42565,N_42566,N_42567,N_42568,N_42569,N_42570,N_42571,N_42572,N_42573,N_42574,N_42575,N_42576,N_42577,N_42578,N_42579,N_42580,N_42581,N_42582,N_42583,N_42584,N_42585,N_42586,N_42587,N_42588,N_42589,N_42590,N_42591,N_42592,N_42593,N_42594,N_42595,N_42596,N_42597,N_42598,N_42599,N_42600,N_42601,N_42602,N_42603,N_42604,N_42605,N_42606,N_42607,N_42608,N_42609,N_42610,N_42611,N_42612,N_42613,N_42614,N_42615,N_42616,N_42617,N_42618,N_42619,N_42620,N_42621,N_42622,N_42623,N_42624,N_42625,N_42626,N_42627,N_42628,N_42629,N_42630,N_42631,N_42632,N_42633,N_42634,N_42635,N_42636,N_42637,N_42638,N_42639,N_42640,N_42641,N_42642,N_42643,N_42644,N_42645,N_42646,N_42647,N_42648,N_42649,N_42650,N_42651,N_42652,N_42653,N_42654,N_42655,N_42656,N_42657,N_42658,N_42659,N_42660,N_42661,N_42662,N_42663,N_42664,N_42665,N_42666,N_42667,N_42668,N_42669,N_42670,N_42671,N_42672,N_42673,N_42674,N_42675,N_42676,N_42677,N_42678,N_42679,N_42680,N_42681,N_42682,N_42683,N_42684,N_42685,N_42686,N_42687,N_42688,N_42689,N_42690,N_42691,N_42692,N_42693,N_42694,N_42695,N_42696,N_42697,N_42698,N_42699,N_42700,N_42701,N_42702,N_42703,N_42704,N_42705,N_42706,N_42707,N_42708,N_42709,N_42710,N_42711,N_42712,N_42713,N_42714,N_42715,N_42716,N_42717,N_42718,N_42719,N_42720,N_42721,N_42722,N_42723,N_42724,N_42725,N_42726,N_42727,N_42728,N_42729,N_42730,N_42731,N_42732,N_42733,N_42734,N_42735,N_42736,N_42737,N_42738,N_42739,N_42740,N_42741,N_42742,N_42743,N_42744,N_42745,N_42746,N_42747,N_42748,N_42749,N_42750,N_42751,N_42752,N_42753,N_42754,N_42755,N_42756,N_42757,N_42758,N_42759,N_42760,N_42761,N_42762,N_42763,N_42764,N_42765,N_42766,N_42767,N_42768,N_42769,N_42770,N_42771,N_42772,N_42773,N_42774,N_42775,N_42776,N_42777,N_42778,N_42779,N_42780,N_42781,N_42782,N_42783,N_42784,N_42785,N_42786,N_42787,N_42788,N_42789,N_42790,N_42791,N_42792,N_42793,N_42794,N_42795,N_42796,N_42797,N_42798,N_42799,N_42800,N_42801,N_42802,N_42803,N_42804,N_42805,N_42806,N_42807,N_42808,N_42809,N_42810,N_42811,N_42812,N_42813,N_42814,N_42815,N_42816,N_42817,N_42818,N_42819,N_42820,N_42821,N_42822,N_42823,N_42824,N_42825,N_42826,N_42827,N_42828,N_42829,N_42830,N_42831,N_42832,N_42833,N_42834,N_42835,N_42836,N_42837,N_42838,N_42839,N_42840,N_42841,N_42842,N_42843,N_42844,N_42845,N_42846,N_42847,N_42848,N_42849,N_42850,N_42851,N_42852,N_42853,N_42854,N_42855,N_42856,N_42857,N_42858,N_42859,N_42860,N_42861,N_42862,N_42863,N_42864,N_42865,N_42866,N_42867,N_42868,N_42869,N_42870,N_42871,N_42872,N_42873,N_42874,N_42875,N_42876,N_42877,N_42878,N_42879,N_42880,N_42881,N_42882,N_42883,N_42884,N_42885,N_42886,N_42887,N_42888,N_42889,N_42890,N_42891,N_42892,N_42893,N_42894,N_42895,N_42896,N_42897,N_42898,N_42899,N_42900,N_42901,N_42902,N_42903,N_42904,N_42905,N_42906,N_42907,N_42908,N_42909,N_42910,N_42911,N_42912,N_42913,N_42914,N_42915,N_42916,N_42917,N_42918,N_42919,N_42920,N_42921,N_42922,N_42923,N_42924,N_42925,N_42926,N_42927,N_42928,N_42929,N_42930,N_42931,N_42932,N_42933,N_42934,N_42935,N_42936,N_42937,N_42938,N_42939,N_42940,N_42941,N_42942,N_42943,N_42944,N_42945,N_42946,N_42947,N_42948,N_42949,N_42950,N_42951,N_42952,N_42953,N_42954,N_42955,N_42956,N_42957,N_42958,N_42959,N_42960,N_42961,N_42962,N_42963,N_42964,N_42965,N_42966,N_42967,N_42968,N_42969,N_42970,N_42971,N_42972,N_42973,N_42974,N_42975,N_42976,N_42977,N_42978,N_42979,N_42980,N_42981,N_42982,N_42983,N_42984,N_42985,N_42986,N_42987,N_42988,N_42989,N_42990,N_42991,N_42992,N_42993,N_42994,N_42995,N_42996,N_42997,N_42998,N_42999,N_43000,N_43001,N_43002,N_43003,N_43004,N_43005,N_43006,N_43007,N_43008,N_43009,N_43010,N_43011,N_43012,N_43013,N_43014,N_43015,N_43016,N_43017,N_43018,N_43019,N_43020,N_43021,N_43022,N_43023,N_43024,N_43025,N_43026,N_43027,N_43028,N_43029,N_43030,N_43031,N_43032,N_43033,N_43034,N_43035,N_43036,N_43037,N_43038,N_43039,N_43040,N_43041,N_43042,N_43043,N_43044,N_43045,N_43046,N_43047,N_43048,N_43049,N_43050,N_43051,N_43052,N_43053,N_43054,N_43055,N_43056,N_43057,N_43058,N_43059,N_43060,N_43061,N_43062,N_43063,N_43064,N_43065,N_43066,N_43067,N_43068,N_43069,N_43070,N_43071,N_43072,N_43073,N_43074,N_43075,N_43076,N_43077,N_43078,N_43079,N_43080,N_43081,N_43082,N_43083,N_43084,N_43085,N_43086,N_43087,N_43088,N_43089,N_43090,N_43091,N_43092,N_43093,N_43094,N_43095,N_43096,N_43097,N_43098,N_43099,N_43100,N_43101,N_43102,N_43103,N_43104,N_43105,N_43106,N_43107,N_43108,N_43109,N_43110,N_43111,N_43112,N_43113,N_43114,N_43115,N_43116,N_43117,N_43118,N_43119,N_43120,N_43121,N_43122,N_43123,N_43124,N_43125,N_43126,N_43127,N_43128,N_43129,N_43130,N_43131,N_43132,N_43133,N_43134,N_43135,N_43136,N_43137,N_43138,N_43139,N_43140,N_43141,N_43142,N_43143,N_43144,N_43145,N_43146,N_43147,N_43148,N_43149,N_43150,N_43151,N_43152,N_43153,N_43154,N_43155,N_43156,N_43157,N_43158,N_43159,N_43160,N_43161,N_43162,N_43163,N_43164,N_43165,N_43166,N_43167,N_43168,N_43169,N_43170,N_43171,N_43172,N_43173,N_43174,N_43175,N_43176,N_43177,N_43178,N_43179,N_43180,N_43181,N_43182,N_43183,N_43184,N_43185,N_43186,N_43187,N_43188,N_43189,N_43190,N_43191,N_43192,N_43193,N_43194,N_43195,N_43196,N_43197,N_43198,N_43199,N_43200,N_43201,N_43202,N_43203,N_43204,N_43205,N_43206,N_43207,N_43208,N_43209,N_43210,N_43211,N_43212,N_43213,N_43214,N_43215,N_43216,N_43217,N_43218,N_43219,N_43220,N_43221,N_43222,N_43223,N_43224,N_43225,N_43226,N_43227,N_43228,N_43229,N_43230,N_43231,N_43232,N_43233,N_43234,N_43235,N_43236,N_43237,N_43238,N_43239,N_43240,N_43241,N_43242,N_43243,N_43244,N_43245,N_43246,N_43247,N_43248,N_43249,N_43250,N_43251,N_43252,N_43253,N_43254,N_43255,N_43256,N_43257,N_43258,N_43259,N_43260,N_43261,N_43262,N_43263,N_43264,N_43265,N_43266,N_43267,N_43268,N_43269,N_43270,N_43271,N_43272,N_43273,N_43274,N_43275,N_43276,N_43277,N_43278,N_43279,N_43280,N_43281,N_43282,N_43283,N_43284,N_43285,N_43286,N_43287,N_43288,N_43289,N_43290,N_43291,N_43292,N_43293,N_43294,N_43295,N_43296,N_43297,N_43298,N_43299,N_43300,N_43301,N_43302,N_43303,N_43304,N_43305,N_43306,N_43307,N_43308,N_43309,N_43310,N_43311,N_43312,N_43313,N_43314,N_43315,N_43316,N_43317,N_43318,N_43319,N_43320,N_43321,N_43322,N_43323,N_43324,N_43325,N_43326,N_43327,N_43328,N_43329,N_43330,N_43331,N_43332,N_43333,N_43334,N_43335,N_43336,N_43337,N_43338,N_43339,N_43340,N_43341,N_43342,N_43343,N_43344,N_43345,N_43346,N_43347,N_43348,N_43349,N_43350,N_43351,N_43352,N_43353,N_43354,N_43355,N_43356,N_43357,N_43358,N_43359,N_43360,N_43361,N_43362,N_43363,N_43364,N_43365,N_43366,N_43367,N_43368,N_43369,N_43370,N_43371,N_43372,N_43373,N_43374,N_43375,N_43376,N_43377,N_43378,N_43379,N_43380,N_43381,N_43382,N_43383,N_43384,N_43385,N_43386,N_43387,N_43388,N_43389,N_43390,N_43391,N_43392,N_43393,N_43394,N_43395,N_43396,N_43397,N_43398,N_43399,N_43400,N_43401,N_43402,N_43403,N_43404,N_43405,N_43406,N_43407,N_43408,N_43409,N_43410,N_43411,N_43412,N_43413,N_43414,N_43415,N_43416,N_43417,N_43418,N_43419,N_43420,N_43421,N_43422,N_43423,N_43424,N_43425,N_43426,N_43427,N_43428,N_43429,N_43430,N_43431,N_43432,N_43433,N_43434,N_43435,N_43436,N_43437,N_43438,N_43439,N_43440,N_43441,N_43442,N_43443,N_43444,N_43445,N_43446,N_43447,N_43448,N_43449,N_43450,N_43451,N_43452,N_43453,N_43454,N_43455,N_43456,N_43457,N_43458,N_43459,N_43460,N_43461,N_43462,N_43463,N_43464,N_43465,N_43466,N_43467,N_43468,N_43469,N_43470,N_43471,N_43472,N_43473,N_43474,N_43475,N_43476,N_43477,N_43478,N_43479,N_43480,N_43481,N_43482,N_43483,N_43484,N_43485,N_43486,N_43487,N_43488,N_43489,N_43490,N_43491,N_43492,N_43493,N_43494,N_43495,N_43496,N_43497,N_43498,N_43499,N_43500,N_43501,N_43502,N_43503,N_43504,N_43505,N_43506,N_43507,N_43508,N_43509,N_43510,N_43511,N_43512,N_43513,N_43514,N_43515,N_43516,N_43517,N_43518,N_43519,N_43520,N_43521,N_43522,N_43523,N_43524,N_43525,N_43526,N_43527,N_43528,N_43529,N_43530,N_43531,N_43532,N_43533,N_43534,N_43535,N_43536,N_43537,N_43538,N_43539,N_43540,N_43541,N_43542,N_43543,N_43544,N_43545,N_43546,N_43547,N_43548,N_43549,N_43550,N_43551,N_43552,N_43553,N_43554,N_43555,N_43556,N_43557,N_43558,N_43559,N_43560,N_43561,N_43562,N_43563,N_43564,N_43565,N_43566,N_43567,N_43568,N_43569,N_43570,N_43571,N_43572,N_43573,N_43574,N_43575,N_43576,N_43577,N_43578,N_43579,N_43580,N_43581,N_43582,N_43583,N_43584,N_43585,N_43586,N_43587,N_43588,N_43589,N_43590,N_43591,N_43592,N_43593,N_43594,N_43595,N_43596,N_43597,N_43598,N_43599,N_43600,N_43601,N_43602,N_43603,N_43604,N_43605,N_43606,N_43607,N_43608,N_43609,N_43610,N_43611,N_43612,N_43613,N_43614,N_43615,N_43616,N_43617,N_43618,N_43619,N_43620,N_43621,N_43622,N_43623,N_43624,N_43625,N_43626,N_43627,N_43628,N_43629,N_43630,N_43631,N_43632,N_43633,N_43634,N_43635,N_43636,N_43637,N_43638,N_43639,N_43640,N_43641,N_43642,N_43643,N_43644,N_43645,N_43646,N_43647,N_43648,N_43649,N_43650,N_43651,N_43652,N_43653,N_43654,N_43655,N_43656,N_43657,N_43658,N_43659,N_43660,N_43661,N_43662,N_43663,N_43664,N_43665,N_43666,N_43667,N_43668,N_43669,N_43670,N_43671,N_43672,N_43673,N_43674,N_43675,N_43676,N_43677,N_43678,N_43679,N_43680,N_43681,N_43682,N_43683,N_43684,N_43685,N_43686,N_43687,N_43688,N_43689,N_43690,N_43691,N_43692,N_43693,N_43694,N_43695,N_43696,N_43697,N_43698,N_43699,N_43700,N_43701,N_43702,N_43703,N_43704,N_43705,N_43706,N_43707,N_43708,N_43709,N_43710,N_43711,N_43712,N_43713,N_43714,N_43715,N_43716,N_43717,N_43718,N_43719,N_43720,N_43721,N_43722,N_43723,N_43724,N_43725,N_43726,N_43727,N_43728,N_43729,N_43730,N_43731,N_43732,N_43733,N_43734,N_43735,N_43736,N_43737,N_43738,N_43739,N_43740,N_43741,N_43742,N_43743,N_43744,N_43745,N_43746,N_43747,N_43748,N_43749,N_43750,N_43751,N_43752,N_43753,N_43754,N_43755,N_43756,N_43757,N_43758,N_43759,N_43760,N_43761,N_43762,N_43763,N_43764,N_43765,N_43766,N_43767,N_43768,N_43769,N_43770,N_43771,N_43772,N_43773,N_43774,N_43775,N_43776,N_43777,N_43778,N_43779,N_43780,N_43781,N_43782,N_43783,N_43784,N_43785,N_43786,N_43787,N_43788,N_43789,N_43790,N_43791,N_43792,N_43793,N_43794,N_43795,N_43796,N_43797,N_43798,N_43799,N_43800,N_43801,N_43802,N_43803,N_43804,N_43805,N_43806,N_43807,N_43808,N_43809,N_43810,N_43811,N_43812,N_43813,N_43814,N_43815,N_43816,N_43817,N_43818,N_43819,N_43820,N_43821,N_43822,N_43823,N_43824,N_43825,N_43826,N_43827,N_43828,N_43829,N_43830,N_43831,N_43832,N_43833,N_43834,N_43835,N_43836,N_43837,N_43838,N_43839,N_43840,N_43841,N_43842,N_43843,N_43844,N_43845,N_43846,N_43847,N_43848,N_43849,N_43850,N_43851,N_43852,N_43853,N_43854,N_43855,N_43856,N_43857,N_43858,N_43859,N_43860,N_43861,N_43862,N_43863,N_43864,N_43865,N_43866,N_43867,N_43868,N_43869,N_43870,N_43871,N_43872,N_43873,N_43874,N_43875,N_43876,N_43877,N_43878,N_43879,N_43880,N_43881,N_43882,N_43883,N_43884,N_43885,N_43886,N_43887,N_43888,N_43889,N_43890,N_43891,N_43892,N_43893,N_43894,N_43895,N_43896,N_43897,N_43898,N_43899,N_43900,N_43901,N_43902,N_43903,N_43904,N_43905,N_43906,N_43907,N_43908,N_43909,N_43910,N_43911,N_43912,N_43913,N_43914,N_43915,N_43916,N_43917,N_43918,N_43919,N_43920,N_43921,N_43922,N_43923,N_43924,N_43925,N_43926,N_43927,N_43928,N_43929,N_43930,N_43931,N_43932,N_43933,N_43934,N_43935,N_43936,N_43937,N_43938,N_43939,N_43940,N_43941,N_43942,N_43943,N_43944,N_43945,N_43946,N_43947,N_43948,N_43949,N_43950,N_43951,N_43952,N_43953,N_43954,N_43955,N_43956,N_43957,N_43958,N_43959,N_43960,N_43961,N_43962,N_43963,N_43964,N_43965,N_43966,N_43967,N_43968,N_43969,N_43970,N_43971,N_43972,N_43973,N_43974,N_43975,N_43976,N_43977,N_43978,N_43979,N_43980,N_43981,N_43982,N_43983,N_43984,N_43985,N_43986,N_43987,N_43988,N_43989,N_43990,N_43991,N_43992,N_43993,N_43994,N_43995,N_43996,N_43997,N_43998,N_43999,N_44000,N_44001,N_44002,N_44003,N_44004,N_44005,N_44006,N_44007,N_44008,N_44009,N_44010,N_44011,N_44012,N_44013,N_44014,N_44015,N_44016,N_44017,N_44018,N_44019,N_44020,N_44021,N_44022,N_44023,N_44024,N_44025,N_44026,N_44027,N_44028,N_44029,N_44030,N_44031,N_44032,N_44033,N_44034,N_44035,N_44036,N_44037,N_44038,N_44039,N_44040,N_44041,N_44042,N_44043,N_44044,N_44045,N_44046,N_44047,N_44048,N_44049,N_44050,N_44051,N_44052,N_44053,N_44054,N_44055,N_44056,N_44057,N_44058,N_44059,N_44060,N_44061,N_44062,N_44063,N_44064,N_44065,N_44066,N_44067,N_44068,N_44069,N_44070,N_44071,N_44072,N_44073,N_44074,N_44075,N_44076,N_44077,N_44078,N_44079,N_44080,N_44081,N_44082,N_44083,N_44084,N_44085,N_44086,N_44087,N_44088,N_44089,N_44090,N_44091,N_44092,N_44093,N_44094,N_44095,N_44096,N_44097,N_44098,N_44099,N_44100,N_44101,N_44102,N_44103,N_44104,N_44105,N_44106,N_44107,N_44108,N_44109,N_44110,N_44111,N_44112,N_44113,N_44114,N_44115,N_44116,N_44117,N_44118,N_44119,N_44120,N_44121,N_44122,N_44123,N_44124,N_44125,N_44126,N_44127,N_44128,N_44129,N_44130,N_44131,N_44132,N_44133,N_44134,N_44135,N_44136,N_44137,N_44138,N_44139,N_44140,N_44141,N_44142,N_44143,N_44144,N_44145,N_44146,N_44147,N_44148,N_44149,N_44150,N_44151,N_44152,N_44153,N_44154,N_44155,N_44156,N_44157,N_44158,N_44159,N_44160,N_44161,N_44162,N_44163,N_44164,N_44165,N_44166,N_44167,N_44168,N_44169,N_44170,N_44171,N_44172,N_44173,N_44174,N_44175,N_44176,N_44177,N_44178,N_44179,N_44180,N_44181,N_44182,N_44183,N_44184,N_44185,N_44186,N_44187,N_44188,N_44189,N_44190,N_44191,N_44192,N_44193,N_44194,N_44195,N_44196,N_44197,N_44198,N_44199,N_44200,N_44201,N_44202,N_44203,N_44204,N_44205,N_44206,N_44207,N_44208,N_44209,N_44210,N_44211,N_44212,N_44213,N_44214,N_44215,N_44216,N_44217,N_44218,N_44219,N_44220,N_44221,N_44222,N_44223,N_44224,N_44225,N_44226,N_44227,N_44228,N_44229,N_44230,N_44231,N_44232,N_44233,N_44234,N_44235,N_44236,N_44237,N_44238,N_44239,N_44240,N_44241,N_44242,N_44243,N_44244,N_44245,N_44246,N_44247,N_44248,N_44249,N_44250,N_44251,N_44252,N_44253,N_44254,N_44255,N_44256,N_44257,N_44258,N_44259,N_44260,N_44261,N_44262,N_44263,N_44264,N_44265,N_44266,N_44267,N_44268,N_44269,N_44270,N_44271,N_44272,N_44273,N_44274,N_44275,N_44276,N_44277,N_44278,N_44279,N_44280,N_44281,N_44282,N_44283,N_44284,N_44285,N_44286,N_44287,N_44288,N_44289,N_44290,N_44291,N_44292,N_44293,N_44294,N_44295,N_44296,N_44297,N_44298,N_44299,N_44300,N_44301,N_44302,N_44303,N_44304,N_44305,N_44306,N_44307,N_44308,N_44309,N_44310,N_44311,N_44312,N_44313,N_44314,N_44315,N_44316,N_44317,N_44318,N_44319,N_44320,N_44321,N_44322,N_44323,N_44324,N_44325,N_44326,N_44327,N_44328,N_44329,N_44330,N_44331,N_44332,N_44333,N_44334,N_44335,N_44336,N_44337,N_44338,N_44339,N_44340,N_44341,N_44342,N_44343,N_44344,N_44345,N_44346,N_44347,N_44348,N_44349,N_44350,N_44351,N_44352,N_44353,N_44354,N_44355,N_44356,N_44357,N_44358,N_44359,N_44360,N_44361,N_44362,N_44363,N_44364,N_44365,N_44366,N_44367,N_44368,N_44369,N_44370,N_44371,N_44372,N_44373,N_44374,N_44375,N_44376,N_44377,N_44378,N_44379,N_44380,N_44381,N_44382,N_44383,N_44384,N_44385,N_44386,N_44387,N_44388,N_44389,N_44390,N_44391,N_44392,N_44393,N_44394,N_44395,N_44396,N_44397,N_44398,N_44399,N_44400,N_44401,N_44402,N_44403,N_44404,N_44405,N_44406,N_44407,N_44408,N_44409,N_44410,N_44411,N_44412,N_44413,N_44414,N_44415,N_44416,N_44417,N_44418,N_44419,N_44420,N_44421,N_44422,N_44423,N_44424,N_44425,N_44426,N_44427,N_44428,N_44429,N_44430,N_44431,N_44432,N_44433,N_44434,N_44435,N_44436,N_44437,N_44438,N_44439,N_44440,N_44441,N_44442,N_44443,N_44444,N_44445,N_44446,N_44447,N_44448,N_44449,N_44450,N_44451,N_44452,N_44453,N_44454,N_44455,N_44456,N_44457,N_44458,N_44459,N_44460,N_44461,N_44462,N_44463,N_44464,N_44465,N_44466,N_44467,N_44468,N_44469,N_44470,N_44471,N_44472,N_44473,N_44474,N_44475,N_44476,N_44477,N_44478,N_44479,N_44480,N_44481,N_44482,N_44483,N_44484,N_44485,N_44486,N_44487,N_44488,N_44489,N_44490,N_44491,N_44492,N_44493,N_44494,N_44495,N_44496,N_44497,N_44498,N_44499,N_44500,N_44501,N_44502,N_44503,N_44504,N_44505,N_44506,N_44507,N_44508,N_44509,N_44510,N_44511,N_44512,N_44513,N_44514,N_44515,N_44516,N_44517,N_44518,N_44519,N_44520,N_44521,N_44522,N_44523,N_44524,N_44525,N_44526,N_44527,N_44528,N_44529,N_44530,N_44531,N_44532,N_44533,N_44534,N_44535,N_44536,N_44537,N_44538,N_44539,N_44540,N_44541,N_44542,N_44543,N_44544,N_44545,N_44546,N_44547,N_44548,N_44549,N_44550,N_44551,N_44552,N_44553,N_44554,N_44555,N_44556,N_44557,N_44558,N_44559,N_44560,N_44561,N_44562,N_44563,N_44564,N_44565,N_44566,N_44567,N_44568,N_44569,N_44570,N_44571,N_44572,N_44573,N_44574,N_44575,N_44576,N_44577,N_44578,N_44579,N_44580,N_44581,N_44582,N_44583,N_44584,N_44585,N_44586,N_44587,N_44588,N_44589,N_44590,N_44591,N_44592,N_44593,N_44594,N_44595,N_44596,N_44597,N_44598,N_44599,N_44600,N_44601,N_44602,N_44603,N_44604,N_44605,N_44606,N_44607,N_44608,N_44609,N_44610,N_44611,N_44612,N_44613,N_44614,N_44615,N_44616,N_44617,N_44618,N_44619,N_44620,N_44621,N_44622,N_44623,N_44624,N_44625,N_44626,N_44627,N_44628,N_44629,N_44630,N_44631,N_44632,N_44633,N_44634,N_44635,N_44636,N_44637,N_44638,N_44639,N_44640,N_44641,N_44642,N_44643,N_44644,N_44645,N_44646,N_44647,N_44648,N_44649,N_44650,N_44651,N_44652,N_44653,N_44654,N_44655,N_44656,N_44657,N_44658,N_44659,N_44660,N_44661,N_44662,N_44663,N_44664,N_44665,N_44666,N_44667,N_44668,N_44669,N_44670,N_44671,N_44672,N_44673,N_44674,N_44675,N_44676,N_44677,N_44678,N_44679,N_44680,N_44681,N_44682,N_44683,N_44684,N_44685,N_44686,N_44687,N_44688,N_44689,N_44690,N_44691,N_44692,N_44693,N_44694,N_44695,N_44696,N_44697,N_44698,N_44699,N_44700,N_44701,N_44702,N_44703,N_44704,N_44705,N_44706,N_44707,N_44708,N_44709,N_44710,N_44711,N_44712,N_44713,N_44714,N_44715,N_44716,N_44717,N_44718,N_44719,N_44720,N_44721,N_44722,N_44723,N_44724,N_44725,N_44726,N_44727,N_44728,N_44729,N_44730,N_44731,N_44732,N_44733,N_44734,N_44735,N_44736,N_44737,N_44738,N_44739,N_44740,N_44741,N_44742,N_44743,N_44744,N_44745,N_44746,N_44747,N_44748,N_44749,N_44750,N_44751,N_44752,N_44753,N_44754,N_44755,N_44756,N_44757,N_44758,N_44759,N_44760,N_44761,N_44762,N_44763,N_44764,N_44765,N_44766,N_44767,N_44768,N_44769,N_44770,N_44771,N_44772,N_44773,N_44774,N_44775,N_44776,N_44777,N_44778,N_44779,N_44780,N_44781,N_44782,N_44783,N_44784,N_44785,N_44786,N_44787,N_44788,N_44789,N_44790,N_44791,N_44792,N_44793,N_44794,N_44795,N_44796,N_44797,N_44798,N_44799,N_44800,N_44801,N_44802,N_44803,N_44804,N_44805,N_44806,N_44807,N_44808,N_44809,N_44810,N_44811,N_44812,N_44813,N_44814,N_44815,N_44816,N_44817,N_44818,N_44819,N_44820,N_44821,N_44822,N_44823,N_44824,N_44825,N_44826,N_44827,N_44828,N_44829,N_44830,N_44831,N_44832,N_44833,N_44834,N_44835,N_44836,N_44837,N_44838,N_44839,N_44840,N_44841,N_44842,N_44843,N_44844,N_44845,N_44846,N_44847,N_44848,N_44849,N_44850,N_44851,N_44852,N_44853,N_44854,N_44855,N_44856,N_44857,N_44858,N_44859,N_44860,N_44861,N_44862,N_44863,N_44864,N_44865,N_44866,N_44867,N_44868,N_44869,N_44870,N_44871,N_44872,N_44873,N_44874,N_44875,N_44876,N_44877,N_44878,N_44879,N_44880,N_44881,N_44882,N_44883,N_44884,N_44885,N_44886,N_44887,N_44888,N_44889,N_44890,N_44891,N_44892,N_44893,N_44894,N_44895,N_44896,N_44897,N_44898,N_44899,N_44900,N_44901,N_44902,N_44903,N_44904,N_44905,N_44906,N_44907,N_44908,N_44909,N_44910,N_44911,N_44912,N_44913,N_44914,N_44915,N_44916,N_44917,N_44918,N_44919,N_44920,N_44921,N_44922,N_44923,N_44924,N_44925,N_44926,N_44927,N_44928,N_44929,N_44930,N_44931,N_44932,N_44933,N_44934,N_44935,N_44936,N_44937,N_44938,N_44939,N_44940,N_44941,N_44942,N_44943,N_44944,N_44945,N_44946,N_44947,N_44948,N_44949,N_44950,N_44951,N_44952,N_44953,N_44954,N_44955,N_44956,N_44957,N_44958,N_44959,N_44960,N_44961,N_44962,N_44963,N_44964,N_44965,N_44966,N_44967,N_44968,N_44969,N_44970,N_44971,N_44972,N_44973,N_44974,N_44975,N_44976,N_44977,N_44978,N_44979,N_44980,N_44981,N_44982,N_44983,N_44984,N_44985,N_44986,N_44987,N_44988,N_44989,N_44990,N_44991,N_44992,N_44993,N_44994,N_44995,N_44996,N_44997,N_44998,N_44999,N_45000,N_45001,N_45002,N_45003,N_45004,N_45005,N_45006,N_45007,N_45008,N_45009,N_45010,N_45011,N_45012,N_45013,N_45014,N_45015,N_45016,N_45017,N_45018,N_45019,N_45020,N_45021,N_45022,N_45023,N_45024,N_45025,N_45026,N_45027,N_45028,N_45029,N_45030,N_45031,N_45032,N_45033,N_45034,N_45035,N_45036,N_45037,N_45038,N_45039,N_45040,N_45041,N_45042,N_45043,N_45044,N_45045,N_45046,N_45047,N_45048,N_45049,N_45050,N_45051,N_45052,N_45053,N_45054,N_45055,N_45056,N_45057,N_45058,N_45059,N_45060,N_45061,N_45062,N_45063,N_45064,N_45065,N_45066,N_45067,N_45068,N_45069,N_45070,N_45071,N_45072,N_45073,N_45074,N_45075,N_45076,N_45077,N_45078,N_45079,N_45080,N_45081,N_45082,N_45083,N_45084,N_45085,N_45086,N_45087,N_45088,N_45089,N_45090,N_45091,N_45092,N_45093,N_45094,N_45095,N_45096,N_45097,N_45098,N_45099,N_45100,N_45101,N_45102,N_45103,N_45104,N_45105,N_45106,N_45107,N_45108,N_45109,N_45110,N_45111,N_45112,N_45113,N_45114,N_45115,N_45116,N_45117,N_45118,N_45119,N_45120,N_45121,N_45122,N_45123,N_45124,N_45125,N_45126,N_45127,N_45128,N_45129,N_45130,N_45131,N_45132,N_45133,N_45134,N_45135,N_45136,N_45137,N_45138,N_45139,N_45140,N_45141,N_45142,N_45143,N_45144,N_45145,N_45146,N_45147,N_45148,N_45149,N_45150,N_45151,N_45152,N_45153,N_45154,N_45155,N_45156,N_45157,N_45158,N_45159,N_45160,N_45161,N_45162,N_45163,N_45164,N_45165,N_45166,N_45167,N_45168,N_45169,N_45170,N_45171,N_45172,N_45173,N_45174,N_45175,N_45176,N_45177,N_45178,N_45179,N_45180,N_45181,N_45182,N_45183,N_45184,N_45185,N_45186,N_45187,N_45188,N_45189,N_45190,N_45191,N_45192,N_45193,N_45194,N_45195,N_45196,N_45197,N_45198,N_45199,N_45200,N_45201,N_45202,N_45203,N_45204,N_45205,N_45206,N_45207,N_45208,N_45209,N_45210,N_45211,N_45212,N_45213,N_45214,N_45215,N_45216,N_45217,N_45218,N_45219,N_45220,N_45221,N_45222,N_45223,N_45224,N_45225,N_45226,N_45227,N_45228,N_45229,N_45230,N_45231,N_45232,N_45233,N_45234,N_45235,N_45236,N_45237,N_45238,N_45239,N_45240,N_45241,N_45242,N_45243,N_45244,N_45245,N_45246,N_45247,N_45248,N_45249,N_45250,N_45251,N_45252,N_45253,N_45254,N_45255,N_45256,N_45257,N_45258,N_45259,N_45260,N_45261,N_45262,N_45263,N_45264,N_45265,N_45266,N_45267,N_45268,N_45269,N_45270,N_45271,N_45272,N_45273,N_45274,N_45275,N_45276,N_45277,N_45278,N_45279,N_45280,N_45281,N_45282,N_45283,N_45284,N_45285,N_45286,N_45287,N_45288,N_45289,N_45290,N_45291,N_45292,N_45293,N_45294,N_45295,N_45296,N_45297,N_45298,N_45299,N_45300,N_45301,N_45302,N_45303,N_45304,N_45305,N_45306,N_45307,N_45308,N_45309,N_45310,N_45311,N_45312,N_45313,N_45314,N_45315,N_45316,N_45317,N_45318,N_45319,N_45320,N_45321,N_45322,N_45323,N_45324,N_45325,N_45326,N_45327,N_45328,N_45329,N_45330,N_45331,N_45332,N_45333,N_45334,N_45335,N_45336,N_45337,N_45338,N_45339,N_45340,N_45341,N_45342,N_45343,N_45344,N_45345,N_45346,N_45347,N_45348,N_45349,N_45350,N_45351,N_45352,N_45353,N_45354,N_45355,N_45356,N_45357,N_45358,N_45359,N_45360,N_45361,N_45362,N_45363,N_45364,N_45365,N_45366,N_45367,N_45368,N_45369,N_45370,N_45371,N_45372,N_45373,N_45374,N_45375,N_45376,N_45377,N_45378,N_45379,N_45380,N_45381,N_45382,N_45383,N_45384,N_45385,N_45386,N_45387,N_45388,N_45389,N_45390,N_45391,N_45392,N_45393,N_45394,N_45395,N_45396,N_45397,N_45398,N_45399,N_45400,N_45401,N_45402,N_45403,N_45404,N_45405,N_45406,N_45407,N_45408,N_45409,N_45410,N_45411,N_45412,N_45413,N_45414,N_45415,N_45416,N_45417,N_45418,N_45419,N_45420,N_45421,N_45422,N_45423,N_45424,N_45425,N_45426,N_45427,N_45428,N_45429,N_45430,N_45431,N_45432,N_45433,N_45434,N_45435,N_45436,N_45437,N_45438,N_45439,N_45440,N_45441,N_45442,N_45443,N_45444,N_45445,N_45446,N_45447,N_45448,N_45449,N_45450,N_45451,N_45452,N_45453,N_45454,N_45455,N_45456,N_45457,N_45458,N_45459,N_45460,N_45461,N_45462,N_45463,N_45464,N_45465,N_45466,N_45467,N_45468,N_45469,N_45470,N_45471,N_45472,N_45473,N_45474,N_45475,N_45476,N_45477,N_45478,N_45479,N_45480,N_45481,N_45482,N_45483,N_45484,N_45485,N_45486,N_45487,N_45488,N_45489,N_45490,N_45491,N_45492,N_45493,N_45494,N_45495,N_45496,N_45497,N_45498,N_45499,N_45500,N_45501,N_45502,N_45503,N_45504,N_45505,N_45506,N_45507,N_45508,N_45509,N_45510,N_45511,N_45512,N_45513,N_45514,N_45515,N_45516,N_45517,N_45518,N_45519,N_45520,N_45521,N_45522,N_45523,N_45524,N_45525,N_45526,N_45527,N_45528,N_45529,N_45530,N_45531,N_45532,N_45533,N_45534,N_45535,N_45536,N_45537,N_45538,N_45539,N_45540,N_45541,N_45542,N_45543,N_45544,N_45545,N_45546,N_45547,N_45548,N_45549,N_45550,N_45551,N_45552,N_45553,N_45554,N_45555,N_45556,N_45557,N_45558,N_45559,N_45560,N_45561,N_45562,N_45563,N_45564,N_45565,N_45566,N_45567,N_45568,N_45569,N_45570,N_45571,N_45572,N_45573,N_45574,N_45575,N_45576,N_45577,N_45578,N_45579,N_45580,N_45581,N_45582,N_45583,N_45584,N_45585,N_45586,N_45587,N_45588,N_45589,N_45590,N_45591,N_45592,N_45593,N_45594,N_45595,N_45596,N_45597,N_45598,N_45599,N_45600,N_45601,N_45602,N_45603,N_45604,N_45605,N_45606,N_45607,N_45608,N_45609,N_45610,N_45611,N_45612,N_45613,N_45614,N_45615,N_45616,N_45617,N_45618,N_45619,N_45620,N_45621,N_45622,N_45623,N_45624,N_45625,N_45626,N_45627,N_45628,N_45629,N_45630,N_45631,N_45632,N_45633,N_45634,N_45635,N_45636,N_45637,N_45638,N_45639,N_45640,N_45641,N_45642,N_45643,N_45644,N_45645,N_45646,N_45647,N_45648,N_45649,N_45650,N_45651,N_45652,N_45653,N_45654,N_45655,N_45656,N_45657,N_45658,N_45659,N_45660,N_45661,N_45662,N_45663,N_45664,N_45665,N_45666,N_45667,N_45668,N_45669,N_45670,N_45671,N_45672,N_45673,N_45674,N_45675,N_45676,N_45677,N_45678,N_45679,N_45680,N_45681,N_45682,N_45683,N_45684,N_45685,N_45686,N_45687,N_45688,N_45689,N_45690,N_45691,N_45692,N_45693,N_45694,N_45695,N_45696,N_45697,N_45698,N_45699,N_45700,N_45701,N_45702,N_45703,N_45704,N_45705,N_45706,N_45707,N_45708,N_45709,N_45710,N_45711,N_45712,N_45713,N_45714,N_45715,N_45716,N_45717,N_45718,N_45719,N_45720,N_45721,N_45722,N_45723,N_45724,N_45725,N_45726,N_45727,N_45728,N_45729,N_45730,N_45731,N_45732,N_45733,N_45734,N_45735,N_45736,N_45737,N_45738,N_45739,N_45740,N_45741,N_45742,N_45743,N_45744,N_45745,N_45746,N_45747,N_45748,N_45749,N_45750,N_45751,N_45752,N_45753,N_45754,N_45755,N_45756,N_45757,N_45758,N_45759,N_45760,N_45761,N_45762,N_45763,N_45764,N_45765,N_45766,N_45767,N_45768,N_45769,N_45770,N_45771,N_45772,N_45773,N_45774,N_45775,N_45776,N_45777,N_45778,N_45779,N_45780,N_45781,N_45782,N_45783,N_45784,N_45785,N_45786,N_45787,N_45788,N_45789,N_45790,N_45791,N_45792,N_45793,N_45794,N_45795,N_45796,N_45797,N_45798,N_45799,N_45800,N_45801,N_45802,N_45803,N_45804,N_45805,N_45806,N_45807,N_45808,N_45809,N_45810,N_45811,N_45812,N_45813,N_45814,N_45815,N_45816,N_45817,N_45818,N_45819,N_45820,N_45821,N_45822,N_45823,N_45824,N_45825,N_45826,N_45827,N_45828,N_45829,N_45830,N_45831,N_45832,N_45833,N_45834,N_45835,N_45836,N_45837,N_45838,N_45839,N_45840,N_45841,N_45842,N_45843,N_45844,N_45845,N_45846,N_45847,N_45848,N_45849,N_45850,N_45851,N_45852,N_45853,N_45854,N_45855,N_45856,N_45857,N_45858,N_45859,N_45860,N_45861,N_45862,N_45863,N_45864,N_45865,N_45866,N_45867,N_45868,N_45869,N_45870,N_45871,N_45872,N_45873,N_45874,N_45875,N_45876,N_45877,N_45878,N_45879,N_45880,N_45881,N_45882,N_45883,N_45884,N_45885,N_45886,N_45887,N_45888,N_45889,N_45890,N_45891,N_45892,N_45893,N_45894,N_45895,N_45896,N_45897,N_45898,N_45899,N_45900,N_45901,N_45902,N_45903,N_45904,N_45905,N_45906,N_45907,N_45908,N_45909,N_45910,N_45911,N_45912,N_45913,N_45914,N_45915,N_45916,N_45917,N_45918,N_45919,N_45920,N_45921,N_45922,N_45923,N_45924,N_45925,N_45926,N_45927,N_45928,N_45929,N_45930,N_45931,N_45932,N_45933,N_45934,N_45935,N_45936,N_45937,N_45938,N_45939,N_45940,N_45941,N_45942,N_45943,N_45944,N_45945,N_45946,N_45947,N_45948,N_45949,N_45950,N_45951,N_45952,N_45953,N_45954,N_45955,N_45956,N_45957,N_45958,N_45959,N_45960,N_45961,N_45962,N_45963,N_45964,N_45965,N_45966,N_45967,N_45968,N_45969,N_45970,N_45971,N_45972,N_45973,N_45974,N_45975,N_45976,N_45977,N_45978,N_45979,N_45980,N_45981,N_45982,N_45983,N_45984,N_45985,N_45986,N_45987,N_45988,N_45989,N_45990,N_45991,N_45992,N_45993,N_45994,N_45995,N_45996,N_45997,N_45998,N_45999,N_46000,N_46001,N_46002,N_46003,N_46004,N_46005,N_46006,N_46007,N_46008,N_46009,N_46010,N_46011,N_46012,N_46013,N_46014,N_46015,N_46016,N_46017,N_46018,N_46019,N_46020,N_46021,N_46022,N_46023,N_46024,N_46025,N_46026,N_46027,N_46028,N_46029,N_46030,N_46031,N_46032,N_46033,N_46034,N_46035,N_46036,N_46037,N_46038,N_46039,N_46040,N_46041,N_46042,N_46043,N_46044,N_46045,N_46046,N_46047,N_46048,N_46049,N_46050,N_46051,N_46052,N_46053,N_46054,N_46055,N_46056,N_46057,N_46058,N_46059,N_46060,N_46061,N_46062,N_46063,N_46064,N_46065,N_46066,N_46067,N_46068,N_46069,N_46070,N_46071,N_46072,N_46073,N_46074,N_46075,N_46076,N_46077,N_46078,N_46079,N_46080,N_46081,N_46082,N_46083,N_46084,N_46085,N_46086,N_46087,N_46088,N_46089,N_46090,N_46091,N_46092,N_46093,N_46094,N_46095,N_46096,N_46097,N_46098,N_46099,N_46100,N_46101,N_46102,N_46103,N_46104,N_46105,N_46106,N_46107,N_46108,N_46109,N_46110,N_46111,N_46112,N_46113,N_46114,N_46115,N_46116,N_46117,N_46118,N_46119,N_46120,N_46121,N_46122,N_46123,N_46124,N_46125,N_46126,N_46127,N_46128,N_46129,N_46130,N_46131,N_46132,N_46133,N_46134,N_46135,N_46136,N_46137,N_46138,N_46139,N_46140,N_46141,N_46142,N_46143,N_46144,N_46145,N_46146,N_46147,N_46148,N_46149,N_46150,N_46151,N_46152,N_46153,N_46154,N_46155,N_46156,N_46157,N_46158,N_46159,N_46160,N_46161,N_46162,N_46163,N_46164,N_46165,N_46166,N_46167,N_46168,N_46169,N_46170,N_46171,N_46172,N_46173,N_46174,N_46175,N_46176,N_46177,N_46178,N_46179,N_46180,N_46181,N_46182,N_46183,N_46184,N_46185,N_46186,N_46187,N_46188,N_46189,N_46190,N_46191,N_46192,N_46193,N_46194,N_46195,N_46196,N_46197,N_46198,N_46199,N_46200,N_46201,N_46202,N_46203,N_46204,N_46205,N_46206,N_46207,N_46208,N_46209,N_46210,N_46211,N_46212,N_46213,N_46214,N_46215,N_46216,N_46217,N_46218,N_46219,N_46220,N_46221,N_46222,N_46223,N_46224,N_46225,N_46226,N_46227,N_46228,N_46229,N_46230,N_46231,N_46232,N_46233,N_46234,N_46235,N_46236,N_46237,N_46238,N_46239,N_46240,N_46241,N_46242,N_46243,N_46244,N_46245,N_46246,N_46247,N_46248,N_46249,N_46250,N_46251,N_46252,N_46253,N_46254,N_46255,N_46256,N_46257,N_46258,N_46259,N_46260,N_46261,N_46262,N_46263,N_46264,N_46265,N_46266,N_46267,N_46268,N_46269,N_46270,N_46271,N_46272,N_46273,N_46274,N_46275,N_46276,N_46277,N_46278,N_46279,N_46280,N_46281,N_46282,N_46283,N_46284,N_46285,N_46286,N_46287,N_46288,N_46289,N_46290,N_46291,N_46292,N_46293,N_46294,N_46295,N_46296,N_46297,N_46298,N_46299,N_46300,N_46301,N_46302,N_46303,N_46304,N_46305,N_46306,N_46307,N_46308,N_46309,N_46310,N_46311,N_46312,N_46313,N_46314,N_46315,N_46316,N_46317,N_46318,N_46319,N_46320,N_46321,N_46322,N_46323,N_46324,N_46325,N_46326,N_46327,N_46328,N_46329,N_46330,N_46331,N_46332,N_46333,N_46334,N_46335,N_46336,N_46337,N_46338,N_46339,N_46340,N_46341,N_46342,N_46343,N_46344,N_46345,N_46346,N_46347,N_46348,N_46349,N_46350,N_46351,N_46352,N_46353,N_46354,N_46355,N_46356,N_46357,N_46358,N_46359,N_46360,N_46361,N_46362,N_46363,N_46364,N_46365,N_46366,N_46367,N_46368,N_46369,N_46370,N_46371,N_46372,N_46373,N_46374,N_46375,N_46376,N_46377,N_46378,N_46379,N_46380,N_46381,N_46382,N_46383,N_46384,N_46385,N_46386,N_46387,N_46388,N_46389,N_46390,N_46391,N_46392,N_46393,N_46394,N_46395,N_46396,N_46397,N_46398,N_46399,N_46400,N_46401,N_46402,N_46403,N_46404,N_46405,N_46406,N_46407,N_46408,N_46409,N_46410,N_46411,N_46412,N_46413,N_46414,N_46415,N_46416,N_46417,N_46418,N_46419,N_46420,N_46421,N_46422,N_46423,N_46424,N_46425,N_46426,N_46427,N_46428,N_46429,N_46430,N_46431,N_46432,N_46433,N_46434,N_46435,N_46436,N_46437,N_46438,N_46439,N_46440,N_46441,N_46442,N_46443,N_46444,N_46445,N_46446,N_46447,N_46448,N_46449,N_46450,N_46451,N_46452,N_46453,N_46454,N_46455,N_46456,N_46457,N_46458,N_46459,N_46460,N_46461,N_46462,N_46463,N_46464,N_46465,N_46466,N_46467,N_46468,N_46469,N_46470,N_46471,N_46472,N_46473,N_46474,N_46475,N_46476,N_46477,N_46478,N_46479,N_46480,N_46481,N_46482,N_46483,N_46484,N_46485,N_46486,N_46487,N_46488,N_46489,N_46490,N_46491,N_46492,N_46493,N_46494,N_46495,N_46496,N_46497,N_46498,N_46499,N_46500,N_46501,N_46502,N_46503,N_46504,N_46505,N_46506,N_46507,N_46508,N_46509,N_46510,N_46511,N_46512,N_46513,N_46514,N_46515,N_46516,N_46517,N_46518,N_46519,N_46520,N_46521,N_46522,N_46523,N_46524,N_46525,N_46526,N_46527,N_46528,N_46529,N_46530,N_46531,N_46532,N_46533,N_46534,N_46535,N_46536,N_46537,N_46538,N_46539,N_46540,N_46541,N_46542,N_46543,N_46544,N_46545,N_46546,N_46547,N_46548,N_46549,N_46550,N_46551,N_46552,N_46553,N_46554,N_46555,N_46556,N_46557,N_46558,N_46559,N_46560,N_46561,N_46562,N_46563,N_46564,N_46565,N_46566,N_46567,N_46568,N_46569,N_46570,N_46571,N_46572,N_46573,N_46574,N_46575,N_46576,N_46577,N_46578,N_46579,N_46580,N_46581,N_46582,N_46583,N_46584,N_46585,N_46586,N_46587,N_46588,N_46589,N_46590,N_46591,N_46592,N_46593,N_46594,N_46595,N_46596,N_46597,N_46598,N_46599,N_46600,N_46601,N_46602,N_46603,N_46604,N_46605,N_46606,N_46607,N_46608,N_46609,N_46610,N_46611,N_46612,N_46613,N_46614,N_46615,N_46616,N_46617,N_46618,N_46619,N_46620,N_46621,N_46622,N_46623,N_46624,N_46625,N_46626,N_46627,N_46628,N_46629,N_46630,N_46631,N_46632,N_46633,N_46634,N_46635,N_46636,N_46637,N_46638,N_46639,N_46640,N_46641,N_46642,N_46643,N_46644,N_46645,N_46646,N_46647,N_46648,N_46649,N_46650,N_46651,N_46652,N_46653,N_46654,N_46655,N_46656,N_46657,N_46658,N_46659,N_46660,N_46661,N_46662,N_46663,N_46664,N_46665,N_46666,N_46667,N_46668,N_46669,N_46670,N_46671,N_46672,N_46673,N_46674,N_46675,N_46676,N_46677,N_46678,N_46679,N_46680,N_46681,N_46682,N_46683,N_46684,N_46685,N_46686,N_46687,N_46688,N_46689,N_46690,N_46691,N_46692,N_46693,N_46694,N_46695,N_46696,N_46697,N_46698,N_46699,N_46700,N_46701,N_46702,N_46703,N_46704,N_46705,N_46706,N_46707,N_46708,N_46709,N_46710,N_46711,N_46712,N_46713,N_46714,N_46715,N_46716,N_46717,N_46718,N_46719,N_46720,N_46721,N_46722,N_46723,N_46724,N_46725,N_46726,N_46727,N_46728,N_46729,N_46730,N_46731,N_46732,N_46733,N_46734,N_46735,N_46736,N_46737,N_46738,N_46739,N_46740,N_46741,N_46742,N_46743,N_46744,N_46745,N_46746,N_46747,N_46748,N_46749,N_46750,N_46751,N_46752,N_46753,N_46754,N_46755,N_46756,N_46757,N_46758,N_46759,N_46760,N_46761,N_46762,N_46763,N_46764,N_46765,N_46766,N_46767,N_46768,N_46769,N_46770,N_46771,N_46772,N_46773,N_46774,N_46775,N_46776,N_46777,N_46778,N_46779,N_46780,N_46781,N_46782,N_46783,N_46784,N_46785,N_46786,N_46787,N_46788,N_46789,N_46790,N_46791,N_46792,N_46793,N_46794,N_46795,N_46796,N_46797,N_46798,N_46799,N_46800,N_46801,N_46802,N_46803,N_46804,N_46805,N_46806,N_46807,N_46808,N_46809,N_46810,N_46811,N_46812,N_46813,N_46814,N_46815,N_46816,N_46817,N_46818,N_46819,N_46820,N_46821,N_46822,N_46823,N_46824,N_46825,N_46826,N_46827,N_46828,N_46829,N_46830,N_46831,N_46832,N_46833,N_46834,N_46835,N_46836,N_46837,N_46838,N_46839,N_46840,N_46841,N_46842,N_46843,N_46844,N_46845,N_46846,N_46847,N_46848,N_46849,N_46850,N_46851,N_46852,N_46853,N_46854,N_46855,N_46856,N_46857,N_46858,N_46859,N_46860,N_46861,N_46862,N_46863,N_46864,N_46865,N_46866,N_46867,N_46868,N_46869,N_46870,N_46871,N_46872,N_46873,N_46874,N_46875,N_46876,N_46877,N_46878,N_46879,N_46880,N_46881,N_46882,N_46883,N_46884,N_46885,N_46886,N_46887,N_46888,N_46889,N_46890,N_46891,N_46892,N_46893,N_46894,N_46895,N_46896,N_46897,N_46898,N_46899,N_46900,N_46901,N_46902,N_46903,N_46904,N_46905,N_46906,N_46907,N_46908,N_46909,N_46910,N_46911,N_46912,N_46913,N_46914,N_46915,N_46916,N_46917,N_46918,N_46919,N_46920,N_46921,N_46922,N_46923,N_46924,N_46925,N_46926,N_46927,N_46928,N_46929,N_46930,N_46931,N_46932,N_46933,N_46934,N_46935,N_46936,N_46937,N_46938,N_46939,N_46940,N_46941,N_46942,N_46943,N_46944,N_46945,N_46946,N_46947,N_46948,N_46949,N_46950,N_46951,N_46952,N_46953,N_46954,N_46955,N_46956,N_46957,N_46958,N_46959,N_46960,N_46961,N_46962,N_46963,N_46964,N_46965,N_46966,N_46967,N_46968,N_46969,N_46970,N_46971,N_46972,N_46973,N_46974,N_46975,N_46976,N_46977,N_46978,N_46979,N_46980,N_46981,N_46982,N_46983,N_46984,N_46985,N_46986,N_46987,N_46988,N_46989,N_46990,N_46991,N_46992,N_46993,N_46994,N_46995,N_46996,N_46997,N_46998,N_46999,N_47000,N_47001,N_47002,N_47003,N_47004,N_47005,N_47006,N_47007,N_47008,N_47009,N_47010,N_47011,N_47012,N_47013,N_47014,N_47015,N_47016,N_47017,N_47018,N_47019,N_47020,N_47021,N_47022,N_47023,N_47024,N_47025,N_47026,N_47027,N_47028,N_47029,N_47030,N_47031,N_47032,N_47033,N_47034,N_47035,N_47036,N_47037,N_47038,N_47039,N_47040,N_47041,N_47042,N_47043,N_47044,N_47045,N_47046,N_47047,N_47048,N_47049,N_47050,N_47051,N_47052,N_47053,N_47054,N_47055,N_47056,N_47057,N_47058,N_47059,N_47060,N_47061,N_47062,N_47063,N_47064,N_47065,N_47066,N_47067,N_47068,N_47069,N_47070,N_47071,N_47072,N_47073,N_47074,N_47075,N_47076,N_47077,N_47078,N_47079,N_47080,N_47081,N_47082,N_47083,N_47084,N_47085,N_47086,N_47087,N_47088,N_47089,N_47090,N_47091,N_47092,N_47093,N_47094,N_47095,N_47096,N_47097,N_47098,N_47099,N_47100,N_47101,N_47102,N_47103,N_47104,N_47105,N_47106,N_47107,N_47108,N_47109,N_47110,N_47111,N_47112,N_47113,N_47114,N_47115,N_47116,N_47117,N_47118,N_47119,N_47120,N_47121,N_47122,N_47123,N_47124,N_47125,N_47126,N_47127,N_47128,N_47129,N_47130,N_47131,N_47132,N_47133,N_47134,N_47135,N_47136,N_47137,N_47138,N_47139,N_47140,N_47141,N_47142,N_47143,N_47144,N_47145,N_47146,N_47147,N_47148,N_47149,N_47150,N_47151,N_47152,N_47153,N_47154,N_47155,N_47156,N_47157,N_47158,N_47159,N_47160,N_47161,N_47162,N_47163,N_47164,N_47165,N_47166,N_47167,N_47168,N_47169,N_47170,N_47171,N_47172,N_47173,N_47174,N_47175,N_47176,N_47177,N_47178,N_47179,N_47180,N_47181,N_47182,N_47183,N_47184,N_47185,N_47186,N_47187,N_47188,N_47189,N_47190,N_47191,N_47192,N_47193,N_47194,N_47195,N_47196,N_47197,N_47198,N_47199,N_47200,N_47201,N_47202,N_47203,N_47204,N_47205,N_47206,N_47207,N_47208,N_47209,N_47210,N_47211,N_47212,N_47213,N_47214,N_47215,N_47216,N_47217,N_47218,N_47219,N_47220,N_47221,N_47222,N_47223,N_47224,N_47225,N_47226,N_47227,N_47228,N_47229,N_47230,N_47231,N_47232,N_47233,N_47234,N_47235,N_47236,N_47237,N_47238,N_47239,N_47240,N_47241,N_47242,N_47243,N_47244,N_47245,N_47246,N_47247,N_47248,N_47249,N_47250,N_47251,N_47252,N_47253,N_47254,N_47255,N_47256,N_47257,N_47258,N_47259,N_47260,N_47261,N_47262,N_47263,N_47264,N_47265,N_47266,N_47267,N_47268,N_47269,N_47270,N_47271,N_47272,N_47273,N_47274,N_47275,N_47276,N_47277,N_47278,N_47279,N_47280,N_47281,N_47282,N_47283,N_47284,N_47285,N_47286,N_47287,N_47288,N_47289,N_47290,N_47291,N_47292,N_47293,N_47294,N_47295,N_47296,N_47297,N_47298,N_47299,N_47300,N_47301,N_47302,N_47303,N_47304,N_47305,N_47306,N_47307,N_47308,N_47309,N_47310,N_47311,N_47312,N_47313,N_47314,N_47315,N_47316,N_47317,N_47318,N_47319,N_47320,N_47321,N_47322,N_47323,N_47324,N_47325,N_47326,N_47327,N_47328,N_47329,N_47330,N_47331,N_47332,N_47333,N_47334,N_47335,N_47336,N_47337,N_47338,N_47339,N_47340,N_47341,N_47342,N_47343,N_47344,N_47345,N_47346,N_47347,N_47348,N_47349,N_47350,N_47351,N_47352,N_47353,N_47354,N_47355,N_47356,N_47357,N_47358,N_47359,N_47360,N_47361,N_47362,N_47363,N_47364,N_47365,N_47366,N_47367,N_47368,N_47369,N_47370,N_47371,N_47372,N_47373,N_47374,N_47375,N_47376,N_47377,N_47378,N_47379,N_47380,N_47381,N_47382,N_47383,N_47384,N_47385,N_47386,N_47387,N_47388,N_47389,N_47390,N_47391,N_47392,N_47393,N_47394,N_47395,N_47396,N_47397,N_47398,N_47399,N_47400,N_47401,N_47402,N_47403,N_47404,N_47405,N_47406,N_47407,N_47408,N_47409,N_47410,N_47411,N_47412,N_47413,N_47414,N_47415,N_47416,N_47417,N_47418,N_47419,N_47420,N_47421,N_47422,N_47423,N_47424,N_47425,N_47426,N_47427,N_47428,N_47429,N_47430,N_47431,N_47432,N_47433,N_47434,N_47435,N_47436,N_47437,N_47438,N_47439,N_47440,N_47441,N_47442,N_47443,N_47444,N_47445,N_47446,N_47447,N_47448,N_47449,N_47450,N_47451,N_47452,N_47453,N_47454,N_47455,N_47456,N_47457,N_47458,N_47459,N_47460,N_47461,N_47462,N_47463,N_47464,N_47465,N_47466,N_47467,N_47468,N_47469,N_47470,N_47471,N_47472,N_47473,N_47474,N_47475,N_47476,N_47477,N_47478,N_47479,N_47480,N_47481,N_47482,N_47483,N_47484,N_47485,N_47486,N_47487,N_47488,N_47489,N_47490,N_47491,N_47492,N_47493,N_47494,N_47495,N_47496,N_47497,N_47498,N_47499,N_47500,N_47501,N_47502,N_47503,N_47504,N_47505,N_47506,N_47507,N_47508,N_47509,N_47510,N_47511,N_47512,N_47513,N_47514,N_47515,N_47516,N_47517,N_47518,N_47519,N_47520,N_47521,N_47522,N_47523,N_47524,N_47525,N_47526,N_47527,N_47528,N_47529,N_47530,N_47531,N_47532,N_47533,N_47534,N_47535,N_47536,N_47537,N_47538,N_47539,N_47540,N_47541,N_47542,N_47543,N_47544,N_47545,N_47546,N_47547,N_47548,N_47549,N_47550,N_47551,N_47552,N_47553,N_47554,N_47555,N_47556,N_47557,N_47558,N_47559,N_47560,N_47561,N_47562,N_47563,N_47564,N_47565,N_47566,N_47567,N_47568,N_47569,N_47570,N_47571,N_47572,N_47573,N_47574,N_47575,N_47576,N_47577,N_47578,N_47579,N_47580,N_47581,N_47582,N_47583,N_47584,N_47585,N_47586,N_47587,N_47588,N_47589,N_47590,N_47591,N_47592,N_47593,N_47594,N_47595,N_47596,N_47597,N_47598,N_47599,N_47600,N_47601,N_47602,N_47603,N_47604,N_47605,N_47606,N_47607,N_47608,N_47609,N_47610,N_47611,N_47612,N_47613,N_47614,N_47615,N_47616,N_47617,N_47618,N_47619,N_47620,N_47621,N_47622,N_47623,N_47624,N_47625,N_47626,N_47627,N_47628,N_47629,N_47630,N_47631,N_47632,N_47633,N_47634,N_47635,N_47636,N_47637,N_47638,N_47639,N_47640,N_47641,N_47642,N_47643,N_47644,N_47645,N_47646,N_47647,N_47648,N_47649,N_47650,N_47651,N_47652,N_47653,N_47654,N_47655,N_47656,N_47657,N_47658,N_47659,N_47660,N_47661,N_47662,N_47663,N_47664,N_47665,N_47666,N_47667,N_47668,N_47669,N_47670,N_47671,N_47672,N_47673,N_47674,N_47675,N_47676,N_47677,N_47678,N_47679,N_47680,N_47681,N_47682,N_47683,N_47684,N_47685,N_47686,N_47687,N_47688,N_47689,N_47690,N_47691,N_47692,N_47693,N_47694,N_47695,N_47696,N_47697,N_47698,N_47699,N_47700,N_47701,N_47702,N_47703,N_47704,N_47705,N_47706,N_47707,N_47708,N_47709,N_47710,N_47711,N_47712,N_47713,N_47714,N_47715,N_47716,N_47717,N_47718,N_47719,N_47720,N_47721,N_47722,N_47723,N_47724,N_47725,N_47726,N_47727,N_47728,N_47729,N_47730,N_47731,N_47732,N_47733,N_47734,N_47735,N_47736,N_47737,N_47738,N_47739,N_47740,N_47741,N_47742,N_47743,N_47744,N_47745,N_47746,N_47747,N_47748,N_47749,N_47750,N_47751,N_47752,N_47753,N_47754,N_47755,N_47756,N_47757,N_47758,N_47759,N_47760,N_47761,N_47762,N_47763,N_47764,N_47765,N_47766,N_47767,N_47768,N_47769,N_47770,N_47771,N_47772,N_47773,N_47774,N_47775,N_47776,N_47777,N_47778,N_47779,N_47780,N_47781,N_47782,N_47783,N_47784,N_47785,N_47786,N_47787,N_47788,N_47789,N_47790,N_47791,N_47792,N_47793,N_47794,N_47795,N_47796,N_47797,N_47798,N_47799,N_47800,N_47801,N_47802,N_47803,N_47804,N_47805,N_47806,N_47807,N_47808,N_47809,N_47810,N_47811,N_47812,N_47813,N_47814,N_47815,N_47816,N_47817,N_47818,N_47819,N_47820,N_47821,N_47822,N_47823,N_47824,N_47825,N_47826,N_47827,N_47828,N_47829,N_47830,N_47831,N_47832,N_47833,N_47834,N_47835,N_47836,N_47837,N_47838,N_47839,N_47840,N_47841,N_47842,N_47843,N_47844,N_47845,N_47846,N_47847,N_47848,N_47849,N_47850,N_47851,N_47852,N_47853,N_47854,N_47855,N_47856,N_47857,N_47858,N_47859,N_47860,N_47861,N_47862,N_47863,N_47864,N_47865,N_47866,N_47867,N_47868,N_47869,N_47870,N_47871,N_47872,N_47873,N_47874,N_47875,N_47876,N_47877,N_47878,N_47879,N_47880,N_47881,N_47882,N_47883,N_47884,N_47885,N_47886,N_47887,N_47888,N_47889,N_47890,N_47891,N_47892,N_47893,N_47894,N_47895,N_47896,N_47897,N_47898,N_47899,N_47900,N_47901,N_47902,N_47903,N_47904,N_47905,N_47906,N_47907,N_47908,N_47909,N_47910,N_47911,N_47912,N_47913,N_47914,N_47915,N_47916,N_47917,N_47918,N_47919,N_47920,N_47921,N_47922,N_47923,N_47924,N_47925,N_47926,N_47927,N_47928,N_47929,N_47930,N_47931,N_47932,N_47933,N_47934,N_47935,N_47936,N_47937,N_47938,N_47939,N_47940,N_47941,N_47942,N_47943,N_47944,N_47945,N_47946,N_47947,N_47948,N_47949,N_47950,N_47951,N_47952,N_47953,N_47954,N_47955,N_47956,N_47957,N_47958,N_47959,N_47960,N_47961,N_47962,N_47963,N_47964,N_47965,N_47966,N_47967,N_47968,N_47969,N_47970,N_47971,N_47972,N_47973,N_47974,N_47975,N_47976,N_47977,N_47978,N_47979,N_47980,N_47981,N_47982,N_47983,N_47984,N_47985,N_47986,N_47987,N_47988,N_47989,N_47990,N_47991,N_47992,N_47993,N_47994,N_47995,N_47996,N_47997,N_47998,N_47999,N_48000,N_48001,N_48002,N_48003,N_48004,N_48005,N_48006,N_48007,N_48008,N_48009,N_48010,N_48011,N_48012,N_48013,N_48014,N_48015,N_48016,N_48017,N_48018,N_48019,N_48020,N_48021,N_48022,N_48023,N_48024,N_48025,N_48026,N_48027,N_48028,N_48029,N_48030,N_48031,N_48032,N_48033,N_48034,N_48035,N_48036,N_48037,N_48038,N_48039,N_48040,N_48041,N_48042,N_48043,N_48044,N_48045,N_48046,N_48047,N_48048,N_48049,N_48050,N_48051,N_48052,N_48053,N_48054,N_48055,N_48056,N_48057,N_48058,N_48059,N_48060,N_48061,N_48062,N_48063,N_48064,N_48065,N_48066,N_48067,N_48068,N_48069,N_48070,N_48071,N_48072,N_48073,N_48074,N_48075,N_48076,N_48077,N_48078,N_48079,N_48080,N_48081,N_48082,N_48083,N_48084,N_48085,N_48086,N_48087,N_48088,N_48089,N_48090,N_48091,N_48092,N_48093,N_48094,N_48095,N_48096,N_48097,N_48098,N_48099,N_48100,N_48101,N_48102,N_48103,N_48104,N_48105,N_48106,N_48107,N_48108,N_48109,N_48110,N_48111,N_48112,N_48113,N_48114,N_48115,N_48116,N_48117,N_48118,N_48119,N_48120,N_48121,N_48122,N_48123,N_48124,N_48125,N_48126,N_48127,N_48128,N_48129,N_48130,N_48131,N_48132,N_48133,N_48134,N_48135,N_48136,N_48137,N_48138,N_48139,N_48140,N_48141,N_48142,N_48143,N_48144,N_48145,N_48146,N_48147,N_48148,N_48149,N_48150,N_48151,N_48152,N_48153,N_48154,N_48155,N_48156,N_48157,N_48158,N_48159,N_48160,N_48161,N_48162,N_48163,N_48164,N_48165,N_48166,N_48167,N_48168,N_48169,N_48170,N_48171,N_48172,N_48173,N_48174,N_48175,N_48176,N_48177,N_48178,N_48179,N_48180,N_48181,N_48182,N_48183,N_48184,N_48185,N_48186,N_48187,N_48188,N_48189,N_48190,N_48191,N_48192,N_48193,N_48194,N_48195,N_48196,N_48197,N_48198,N_48199,N_48200,N_48201,N_48202,N_48203,N_48204,N_48205,N_48206,N_48207,N_48208,N_48209,N_48210,N_48211,N_48212,N_48213,N_48214,N_48215,N_48216,N_48217,N_48218,N_48219,N_48220,N_48221,N_48222,N_48223,N_48224,N_48225,N_48226,N_48227,N_48228,N_48229,N_48230,N_48231,N_48232,N_48233,N_48234,N_48235,N_48236,N_48237,N_48238,N_48239,N_48240,N_48241,N_48242,N_48243,N_48244,N_48245,N_48246,N_48247,N_48248,N_48249,N_48250,N_48251,N_48252,N_48253,N_48254,N_48255,N_48256,N_48257,N_48258,N_48259,N_48260,N_48261,N_48262,N_48263,N_48264,N_48265,N_48266,N_48267,N_48268,N_48269,N_48270,N_48271,N_48272,N_48273,N_48274,N_48275,N_48276,N_48277,N_48278,N_48279,N_48280,N_48281,N_48282,N_48283,N_48284,N_48285,N_48286,N_48287,N_48288,N_48289,N_48290,N_48291,N_48292,N_48293,N_48294,N_48295,N_48296,N_48297,N_48298,N_48299,N_48300,N_48301,N_48302,N_48303,N_48304,N_48305,N_48306,N_48307,N_48308,N_48309,N_48310,N_48311,N_48312,N_48313,N_48314,N_48315,N_48316,N_48317,N_48318,N_48319,N_48320,N_48321,N_48322,N_48323,N_48324,N_48325,N_48326,N_48327,N_48328,N_48329,N_48330,N_48331,N_48332,N_48333,N_48334,N_48335,N_48336,N_48337,N_48338,N_48339,N_48340,N_48341,N_48342,N_48343,N_48344,N_48345,N_48346,N_48347,N_48348,N_48349,N_48350,N_48351,N_48352,N_48353,N_48354,N_48355,N_48356,N_48357,N_48358,N_48359,N_48360,N_48361,N_48362,N_48363,N_48364,N_48365,N_48366,N_48367,N_48368,N_48369,N_48370,N_48371,N_48372,N_48373,N_48374,N_48375,N_48376,N_48377,N_48378,N_48379,N_48380,N_48381,N_48382,N_48383,N_48384,N_48385,N_48386,N_48387,N_48388,N_48389,N_48390,N_48391,N_48392,N_48393,N_48394,N_48395,N_48396,N_48397,N_48398,N_48399,N_48400,N_48401,N_48402,N_48403,N_48404,N_48405,N_48406,N_48407,N_48408,N_48409,N_48410,N_48411,N_48412,N_48413,N_48414,N_48415,N_48416,N_48417,N_48418,N_48419,N_48420,N_48421,N_48422,N_48423,N_48424,N_48425,N_48426,N_48427,N_48428,N_48429,N_48430,N_48431,N_48432,N_48433,N_48434,N_48435,N_48436,N_48437,N_48438,N_48439,N_48440,N_48441,N_48442,N_48443,N_48444,N_48445,N_48446,N_48447,N_48448,N_48449,N_48450,N_48451,N_48452,N_48453,N_48454,N_48455,N_48456,N_48457,N_48458,N_48459,N_48460,N_48461,N_48462,N_48463,N_48464,N_48465,N_48466,N_48467,N_48468,N_48469,N_48470,N_48471,N_48472,N_48473,N_48474,N_48475,N_48476,N_48477,N_48478,N_48479,N_48480,N_48481,N_48482,N_48483,N_48484,N_48485,N_48486,N_48487,N_48488,N_48489,N_48490,N_48491,N_48492,N_48493,N_48494,N_48495,N_48496,N_48497,N_48498,N_48499,N_48500,N_48501,N_48502,N_48503,N_48504,N_48505,N_48506,N_48507,N_48508,N_48509,N_48510,N_48511,N_48512,N_48513,N_48514,N_48515,N_48516,N_48517,N_48518,N_48519,N_48520,N_48521,N_48522,N_48523,N_48524,N_48525,N_48526,N_48527,N_48528,N_48529,N_48530,N_48531,N_48532,N_48533,N_48534,N_48535,N_48536,N_48537,N_48538,N_48539,N_48540,N_48541,N_48542,N_48543,N_48544,N_48545,N_48546,N_48547,N_48548,N_48549,N_48550,N_48551,N_48552,N_48553,N_48554,N_48555,N_48556,N_48557,N_48558,N_48559,N_48560,N_48561,N_48562,N_48563,N_48564,N_48565,N_48566,N_48567,N_48568,N_48569,N_48570,N_48571,N_48572,N_48573,N_48574,N_48575,N_48576,N_48577,N_48578,N_48579,N_48580,N_48581,N_48582,N_48583,N_48584,N_48585,N_48586,N_48587,N_48588,N_48589,N_48590,N_48591,N_48592,N_48593,N_48594,N_48595,N_48596,N_48597,N_48598,N_48599,N_48600,N_48601,N_48602,N_48603,N_48604,N_48605,N_48606,N_48607,N_48608,N_48609,N_48610,N_48611,N_48612,N_48613,N_48614,N_48615,N_48616,N_48617,N_48618,N_48619,N_48620,N_48621,N_48622,N_48623,N_48624,N_48625,N_48626,N_48627,N_48628,N_48629,N_48630,N_48631,N_48632,N_48633,N_48634,N_48635,N_48636,N_48637,N_48638,N_48639,N_48640,N_48641,N_48642,N_48643,N_48644,N_48645,N_48646,N_48647,N_48648,N_48649,N_48650,N_48651,N_48652,N_48653,N_48654,N_48655,N_48656,N_48657,N_48658,N_48659,N_48660,N_48661,N_48662,N_48663,N_48664,N_48665,N_48666,N_48667,N_48668,N_48669,N_48670,N_48671,N_48672,N_48673,N_48674,N_48675,N_48676,N_48677,N_48678,N_48679,N_48680,N_48681,N_48682,N_48683,N_48684,N_48685,N_48686,N_48687,N_48688,N_48689,N_48690,N_48691,N_48692,N_48693,N_48694,N_48695,N_48696,N_48697,N_48698,N_48699,N_48700,N_48701,N_48702,N_48703,N_48704,N_48705,N_48706,N_48707,N_48708,N_48709,N_48710,N_48711,N_48712,N_48713,N_48714,N_48715,N_48716,N_48717,N_48718,N_48719,N_48720,N_48721,N_48722,N_48723,N_48724,N_48725,N_48726,N_48727,N_48728,N_48729,N_48730,N_48731,N_48732,N_48733,N_48734,N_48735,N_48736,N_48737,N_48738,N_48739,N_48740,N_48741,N_48742,N_48743,N_48744,N_48745,N_48746,N_48747,N_48748,N_48749,N_48750,N_48751,N_48752,N_48753,N_48754,N_48755,N_48756,N_48757,N_48758,N_48759,N_48760,N_48761,N_48762,N_48763,N_48764,N_48765,N_48766,N_48767,N_48768,N_48769,N_48770,N_48771,N_48772,N_48773,N_48774,N_48775,N_48776,N_48777,N_48778,N_48779,N_48780,N_48781,N_48782,N_48783,N_48784,N_48785,N_48786,N_48787,N_48788,N_48789,N_48790,N_48791,N_48792,N_48793,N_48794,N_48795,N_48796,N_48797,N_48798,N_48799,N_48800,N_48801,N_48802,N_48803,N_48804,N_48805,N_48806,N_48807,N_48808,N_48809,N_48810,N_48811,N_48812,N_48813,N_48814,N_48815,N_48816,N_48817,N_48818,N_48819,N_48820,N_48821,N_48822,N_48823,N_48824,N_48825,N_48826,N_48827,N_48828,N_48829,N_48830,N_48831,N_48832,N_48833,N_48834,N_48835,N_48836,N_48837,N_48838,N_48839,N_48840,N_48841,N_48842,N_48843,N_48844,N_48845,N_48846,N_48847,N_48848,N_48849,N_48850,N_48851,N_48852,N_48853,N_48854,N_48855,N_48856,N_48857,N_48858,N_48859,N_48860,N_48861,N_48862,N_48863,N_48864,N_48865,N_48866,N_48867,N_48868,N_48869,N_48870,N_48871,N_48872,N_48873,N_48874,N_48875,N_48876,N_48877,N_48878,N_48879,N_48880,N_48881,N_48882,N_48883,N_48884,N_48885,N_48886,N_48887,N_48888,N_48889,N_48890,N_48891,N_48892,N_48893,N_48894,N_48895,N_48896,N_48897,N_48898,N_48899,N_48900,N_48901,N_48902,N_48903,N_48904,N_48905,N_48906,N_48907,N_48908,N_48909,N_48910,N_48911,N_48912,N_48913,N_48914,N_48915,N_48916,N_48917,N_48918,N_48919,N_48920,N_48921,N_48922,N_48923,N_48924,N_48925,N_48926,N_48927,N_48928,N_48929,N_48930,N_48931,N_48932,N_48933,N_48934,N_48935,N_48936,N_48937,N_48938,N_48939,N_48940,N_48941,N_48942,N_48943,N_48944,N_48945,N_48946,N_48947,N_48948,N_48949,N_48950,N_48951,N_48952,N_48953,N_48954,N_48955,N_48956,N_48957,N_48958,N_48959,N_48960,N_48961,N_48962,N_48963,N_48964,N_48965,N_48966,N_48967,N_48968,N_48969,N_48970,N_48971,N_48972,N_48973,N_48974,N_48975,N_48976,N_48977,N_48978,N_48979,N_48980,N_48981,N_48982,N_48983,N_48984,N_48985,N_48986,N_48987,N_48988,N_48989,N_48990,N_48991,N_48992,N_48993,N_48994,N_48995,N_48996,N_48997,N_48998,N_48999,N_49000,N_49001,N_49002,N_49003,N_49004,N_49005,N_49006,N_49007,N_49008,N_49009,N_49010,N_49011,N_49012,N_49013,N_49014,N_49015,N_49016,N_49017,N_49018,N_49019,N_49020,N_49021,N_49022,N_49023,N_49024,N_49025,N_49026,N_49027,N_49028,N_49029,N_49030,N_49031,N_49032,N_49033,N_49034,N_49035,N_49036,N_49037,N_49038,N_49039,N_49040,N_49041,N_49042,N_49043,N_49044,N_49045,N_49046,N_49047,N_49048,N_49049,N_49050,N_49051,N_49052,N_49053,N_49054,N_49055,N_49056,N_49057,N_49058,N_49059,N_49060,N_49061,N_49062,N_49063,N_49064,N_49065,N_49066,N_49067,N_49068,N_49069,N_49070,N_49071,N_49072,N_49073,N_49074,N_49075,N_49076,N_49077,N_49078,N_49079,N_49080,N_49081,N_49082,N_49083,N_49084,N_49085,N_49086,N_49087,N_49088,N_49089,N_49090,N_49091,N_49092,N_49093,N_49094,N_49095,N_49096,N_49097,N_49098,N_49099,N_49100,N_49101,N_49102,N_49103,N_49104,N_49105,N_49106,N_49107,N_49108,N_49109,N_49110,N_49111,N_49112,N_49113,N_49114,N_49115,N_49116,N_49117,N_49118,N_49119,N_49120,N_49121,N_49122,N_49123,N_49124,N_49125,N_49126,N_49127,N_49128,N_49129,N_49130,N_49131,N_49132,N_49133,N_49134,N_49135,N_49136,N_49137,N_49138,N_49139,N_49140,N_49141,N_49142,N_49143,N_49144,N_49145,N_49146,N_49147,N_49148,N_49149,N_49150,N_49151,N_49152,N_49153,N_49154,N_49155,N_49156,N_49157,N_49158,N_49159,N_49160,N_49161,N_49162,N_49163,N_49164,N_49165,N_49166,N_49167,N_49168,N_49169,N_49170,N_49171,N_49172,N_49173,N_49174,N_49175,N_49176,N_49177,N_49178,N_49179,N_49180,N_49181,N_49182,N_49183,N_49184,N_49185,N_49186,N_49187,N_49188,N_49189,N_49190,N_49191,N_49192,N_49193,N_49194,N_49195,N_49196,N_49197,N_49198,N_49199,N_49200,N_49201,N_49202,N_49203,N_49204,N_49205,N_49206,N_49207,N_49208,N_49209,N_49210,N_49211,N_49212,N_49213,N_49214,N_49215,N_49216,N_49217,N_49218,N_49219,N_49220,N_49221,N_49222,N_49223,N_49224,N_49225,N_49226,N_49227,N_49228,N_49229,N_49230,N_49231,N_49232,N_49233,N_49234,N_49235,N_49236,N_49237,N_49238,N_49239,N_49240,N_49241,N_49242,N_49243,N_49244,N_49245,N_49246,N_49247,N_49248,N_49249,N_49250,N_49251,N_49252,N_49253,N_49254,N_49255,N_49256,N_49257,N_49258,N_49259,N_49260,N_49261,N_49262,N_49263,N_49264,N_49265,N_49266,N_49267,N_49268,N_49269,N_49270,N_49271,N_49272,N_49273,N_49274,N_49275,N_49276,N_49277,N_49278,N_49279,N_49280,N_49281,N_49282,N_49283,N_49284,N_49285,N_49286,N_49287,N_49288,N_49289,N_49290,N_49291,N_49292,N_49293,N_49294,N_49295,N_49296,N_49297,N_49298,N_49299,N_49300,N_49301,N_49302,N_49303,N_49304,N_49305,N_49306,N_49307,N_49308,N_49309,N_49310,N_49311,N_49312,N_49313,N_49314,N_49315,N_49316,N_49317,N_49318,N_49319,N_49320,N_49321,N_49322,N_49323,N_49324,N_49325,N_49326,N_49327,N_49328,N_49329,N_49330,N_49331,N_49332,N_49333,N_49334,N_49335,N_49336,N_49337,N_49338,N_49339,N_49340,N_49341,N_49342,N_49343,N_49344,N_49345,N_49346,N_49347,N_49348,N_49349,N_49350,N_49351,N_49352,N_49353,N_49354,N_49355,N_49356,N_49357,N_49358,N_49359,N_49360,N_49361,N_49362,N_49363,N_49364,N_49365,N_49366,N_49367,N_49368,N_49369,N_49370,N_49371,N_49372,N_49373,N_49374,N_49375,N_49376,N_49377,N_49378,N_49379,N_49380,N_49381,N_49382,N_49383,N_49384,N_49385,N_49386,N_49387,N_49388,N_49389,N_49390,N_49391,N_49392,N_49393,N_49394,N_49395,N_49396,N_49397,N_49398,N_49399,N_49400,N_49401,N_49402,N_49403,N_49404,N_49405,N_49406,N_49407,N_49408,N_49409,N_49410,N_49411,N_49412,N_49413,N_49414,N_49415,N_49416,N_49417,N_49418,N_49419,N_49420,N_49421,N_49422,N_49423,N_49424,N_49425,N_49426,N_49427,N_49428,N_49429,N_49430,N_49431,N_49432,N_49433,N_49434,N_49435,N_49436,N_49437,N_49438,N_49439,N_49440,N_49441,N_49442,N_49443,N_49444,N_49445,N_49446,N_49447,N_49448,N_49449,N_49450,N_49451,N_49452,N_49453,N_49454,N_49455,N_49456,N_49457,N_49458,N_49459,N_49460,N_49461,N_49462,N_49463,N_49464,N_49465,N_49466,N_49467,N_49468,N_49469,N_49470,N_49471,N_49472,N_49473,N_49474,N_49475,N_49476,N_49477,N_49478,N_49479,N_49480,N_49481,N_49482,N_49483,N_49484,N_49485,N_49486,N_49487,N_49488,N_49489,N_49490,N_49491,N_49492,N_49493,N_49494,N_49495,N_49496,N_49497,N_49498,N_49499,N_49500,N_49501,N_49502,N_49503,N_49504,N_49505,N_49506,N_49507,N_49508,N_49509,N_49510,N_49511,N_49512,N_49513,N_49514,N_49515,N_49516,N_49517,N_49518,N_49519,N_49520,N_49521,N_49522,N_49523,N_49524,N_49525,N_49526,N_49527,N_49528,N_49529,N_49530,N_49531,N_49532,N_49533,N_49534,N_49535,N_49536,N_49537,N_49538,N_49539,N_49540,N_49541,N_49542,N_49543,N_49544,N_49545,N_49546,N_49547,N_49548,N_49549,N_49550,N_49551,N_49552,N_49553,N_49554,N_49555,N_49556,N_49557,N_49558,N_49559,N_49560,N_49561,N_49562,N_49563,N_49564,N_49565,N_49566,N_49567,N_49568,N_49569,N_49570,N_49571,N_49572,N_49573,N_49574,N_49575,N_49576,N_49577,N_49578,N_49579,N_49580,N_49581,N_49582,N_49583,N_49584,N_49585,N_49586,N_49587,N_49588,N_49589,N_49590,N_49591,N_49592,N_49593,N_49594,N_49595,N_49596,N_49597,N_49598,N_49599,N_49600,N_49601,N_49602,N_49603,N_49604,N_49605,N_49606,N_49607,N_49608,N_49609,N_49610,N_49611,N_49612,N_49613,N_49614,N_49615,N_49616,N_49617,N_49618,N_49619,N_49620,N_49621,N_49622,N_49623,N_49624,N_49625,N_49626,N_49627,N_49628,N_49629,N_49630,N_49631,N_49632,N_49633,N_49634,N_49635,N_49636,N_49637,N_49638,N_49639,N_49640,N_49641,N_49642,N_49643,N_49644,N_49645,N_49646,N_49647,N_49648,N_49649,N_49650,N_49651,N_49652,N_49653,N_49654,N_49655,N_49656,N_49657,N_49658,N_49659,N_49660,N_49661,N_49662,N_49663,N_49664,N_49665,N_49666,N_49667,N_49668,N_49669,N_49670,N_49671,N_49672,N_49673,N_49674,N_49675,N_49676,N_49677,N_49678,N_49679,N_49680,N_49681,N_49682,N_49683,N_49684,N_49685,N_49686,N_49687,N_49688,N_49689,N_49690,N_49691,N_49692,N_49693,N_49694,N_49695,N_49696,N_49697,N_49698,N_49699,N_49700,N_49701,N_49702,N_49703,N_49704,N_49705,N_49706,N_49707,N_49708,N_49709,N_49710,N_49711,N_49712,N_49713,N_49714,N_49715,N_49716,N_49717,N_49718,N_49719,N_49720,N_49721,N_49722,N_49723,N_49724,N_49725,N_49726,N_49727,N_49728,N_49729,N_49730,N_49731,N_49732,N_49733,N_49734,N_49735,N_49736,N_49737,N_49738,N_49739,N_49740,N_49741,N_49742,N_49743,N_49744,N_49745,N_49746,N_49747,N_49748,N_49749,N_49750,N_49751,N_49752,N_49753,N_49754,N_49755,N_49756,N_49757,N_49758,N_49759,N_49760,N_49761,N_49762,N_49763,N_49764,N_49765,N_49766,N_49767,N_49768,N_49769,N_49770,N_49771,N_49772,N_49773,N_49774,N_49775,N_49776,N_49777,N_49778,N_49779,N_49780,N_49781,N_49782,N_49783,N_49784,N_49785,N_49786,N_49787,N_49788,N_49789,N_49790,N_49791,N_49792,N_49793,N_49794,N_49795,N_49796,N_49797,N_49798,N_49799,N_49800,N_49801,N_49802,N_49803,N_49804,N_49805,N_49806,N_49807,N_49808,N_49809,N_49810,N_49811,N_49812,N_49813,N_49814,N_49815,N_49816,N_49817,N_49818,N_49819,N_49820,N_49821,N_49822,N_49823,N_49824,N_49825,N_49826,N_49827,N_49828,N_49829,N_49830,N_49831,N_49832,N_49833,N_49834,N_49835,N_49836,N_49837,N_49838,N_49839,N_49840,N_49841,N_49842,N_49843,N_49844,N_49845,N_49846,N_49847,N_49848,N_49849,N_49850,N_49851,N_49852,N_49853,N_49854,N_49855,N_49856,N_49857,N_49858,N_49859,N_49860,N_49861,N_49862,N_49863,N_49864,N_49865,N_49866,N_49867,N_49868,N_49869,N_49870,N_49871,N_49872,N_49873,N_49874,N_49875,N_49876,N_49877,N_49878,N_49879,N_49880,N_49881,N_49882,N_49883,N_49884,N_49885,N_49886,N_49887,N_49888,N_49889,N_49890,N_49891,N_49892,N_49893,N_49894,N_49895,N_49896,N_49897,N_49898,N_49899,N_49900,N_49901,N_49902,N_49903,N_49904,N_49905,N_49906,N_49907,N_49908,N_49909,N_49910,N_49911,N_49912,N_49913,N_49914,N_49915,N_49916,N_49917,N_49918,N_49919,N_49920,N_49921,N_49922,N_49923,N_49924,N_49925,N_49926,N_49927,N_49928,N_49929,N_49930,N_49931,N_49932,N_49933,N_49934,N_49935,N_49936,N_49937,N_49938,N_49939,N_49940,N_49941,N_49942,N_49943,N_49944,N_49945,N_49946,N_49947,N_49948,N_49949,N_49950,N_49951,N_49952,N_49953,N_49954,N_49955,N_49956,N_49957,N_49958,N_49959,N_49960,N_49961,N_49962,N_49963,N_49964,N_49965,N_49966,N_49967,N_49968,N_49969,N_49970,N_49971,N_49972,N_49973,N_49974,N_49975,N_49976,N_49977,N_49978,N_49979,N_49980,N_49981,N_49982,N_49983,N_49984,N_49985,N_49986,N_49987,N_49988,N_49989,N_49990,N_49991,N_49992,N_49993,N_49994,N_49995,N_49996,N_49997,N_49998,N_49999;
xor U0 (N_0,In_3669,In_314);
nand U1 (N_1,In_895,In_2757);
or U2 (N_2,In_1418,In_4701);
and U3 (N_3,In_3643,In_105);
and U4 (N_4,In_4120,In_2412);
nand U5 (N_5,In_3059,In_3313);
xor U6 (N_6,In_1885,In_3563);
nand U7 (N_7,In_4610,In_2064);
nand U8 (N_8,In_946,In_4257);
and U9 (N_9,In_1486,In_3180);
nand U10 (N_10,In_2114,In_2785);
nand U11 (N_11,In_2448,In_1149);
or U12 (N_12,In_1485,In_682);
nor U13 (N_13,In_4385,In_4739);
or U14 (N_14,In_741,In_776);
and U15 (N_15,In_2328,In_2449);
nor U16 (N_16,In_4083,In_3256);
xnor U17 (N_17,In_3414,In_3510);
nor U18 (N_18,In_4964,In_2823);
nor U19 (N_19,In_399,In_3079);
and U20 (N_20,In_2165,In_4322);
nor U21 (N_21,In_3092,In_3885);
or U22 (N_22,In_3266,In_1631);
xor U23 (N_23,In_2827,In_4266);
or U24 (N_24,In_566,In_2811);
nor U25 (N_25,In_4277,In_952);
xnor U26 (N_26,In_4161,In_2754);
or U27 (N_27,In_4505,In_1771);
nor U28 (N_28,In_4521,In_1323);
nand U29 (N_29,In_1077,In_1652);
nand U30 (N_30,In_3432,In_1571);
and U31 (N_31,In_1180,In_322);
xor U32 (N_32,In_1721,In_4095);
or U33 (N_33,In_3802,In_785);
or U34 (N_34,In_2805,In_4822);
and U35 (N_35,In_2526,In_1752);
or U36 (N_36,In_2461,In_2280);
and U37 (N_37,In_2340,In_902);
nand U38 (N_38,In_1927,In_2696);
and U39 (N_39,In_1737,In_2564);
nand U40 (N_40,In_1881,In_3649);
and U41 (N_41,In_2523,In_466);
and U42 (N_42,In_3868,In_1165);
and U43 (N_43,In_2062,In_2762);
and U44 (N_44,In_860,In_2494);
nand U45 (N_45,In_2671,In_2489);
or U46 (N_46,In_2109,In_4057);
nor U47 (N_47,In_2532,In_1032);
or U48 (N_48,In_1179,In_1932);
nor U49 (N_49,In_2744,In_3975);
or U50 (N_50,In_1171,In_655);
and U51 (N_51,In_3769,In_4354);
or U52 (N_52,In_131,In_4980);
nor U53 (N_53,In_1675,In_1280);
xnor U54 (N_54,In_2535,In_4147);
or U55 (N_55,In_1569,In_1953);
or U56 (N_56,In_2385,In_2045);
nor U57 (N_57,In_1139,In_3762);
and U58 (N_58,In_1957,In_2123);
and U59 (N_59,In_4604,In_667);
and U60 (N_60,In_1519,In_3168);
and U61 (N_61,In_2843,In_3956);
or U62 (N_62,In_1369,In_3612);
nand U63 (N_63,In_1501,In_1582);
or U64 (N_64,In_4539,In_3654);
and U65 (N_65,In_4410,In_4416);
and U66 (N_66,In_751,In_3228);
nand U67 (N_67,In_2253,In_732);
and U68 (N_68,In_2998,In_2760);
and U69 (N_69,In_1005,In_3562);
or U70 (N_70,In_4127,In_2091);
and U71 (N_71,In_1056,In_675);
nand U72 (N_72,In_3992,In_2575);
and U73 (N_73,In_1952,In_443);
and U74 (N_74,In_101,In_2437);
or U75 (N_75,In_893,In_4986);
or U76 (N_76,In_1460,In_4085);
or U77 (N_77,In_109,In_3897);
and U78 (N_78,In_1722,In_3344);
and U79 (N_79,In_4729,In_2089);
nor U80 (N_80,In_1900,In_2358);
nand U81 (N_81,In_330,In_1894);
xor U82 (N_82,In_4152,In_4634);
and U83 (N_83,In_3797,In_118);
nor U84 (N_84,In_1660,In_4495);
or U85 (N_85,In_4482,In_4246);
or U86 (N_86,In_1630,In_4655);
xnor U87 (N_87,In_875,In_4946);
or U88 (N_88,In_4900,In_2577);
and U89 (N_89,In_2189,In_1792);
nor U90 (N_90,In_4567,In_733);
or U91 (N_91,In_520,In_3829);
nand U92 (N_92,In_4696,In_1753);
and U93 (N_93,In_4578,In_1616);
or U94 (N_94,In_2224,In_3295);
nor U95 (N_95,In_1956,In_4299);
or U96 (N_96,In_332,In_4254);
and U97 (N_97,In_1539,In_1201);
and U98 (N_98,In_4538,In_980);
xnor U99 (N_99,In_397,In_4396);
nand U100 (N_100,In_2044,In_2073);
nand U101 (N_101,In_851,In_1639);
and U102 (N_102,In_2383,In_3949);
or U103 (N_103,In_3292,In_3105);
and U104 (N_104,In_1524,In_653);
nor U105 (N_105,In_3358,In_3022);
xor U106 (N_106,In_1839,In_1846);
and U107 (N_107,In_2422,In_1347);
nand U108 (N_108,In_1271,In_1218);
xnor U109 (N_109,In_3318,In_1831);
nand U110 (N_110,In_2630,In_4800);
and U111 (N_111,In_2271,In_1859);
or U112 (N_112,In_1277,In_2341);
or U113 (N_113,In_3923,In_4660);
nor U114 (N_114,In_2215,In_2281);
nand U115 (N_115,In_2239,In_251);
nand U116 (N_116,In_1591,In_344);
and U117 (N_117,In_3666,In_4288);
nand U118 (N_118,In_1686,In_2423);
nand U119 (N_119,In_3693,In_4930);
nand U120 (N_120,In_831,In_4039);
xor U121 (N_121,In_4767,In_4869);
or U122 (N_122,In_4312,In_808);
nor U123 (N_123,In_54,In_759);
and U124 (N_124,In_4341,In_3320);
nor U125 (N_125,In_765,In_2065);
or U126 (N_126,In_3844,In_4422);
nor U127 (N_127,In_3484,In_3623);
nand U128 (N_128,In_222,In_4892);
or U129 (N_129,In_1739,In_1095);
and U130 (N_130,In_3466,In_1961);
nand U131 (N_131,In_1468,In_3127);
xnor U132 (N_132,In_703,In_1573);
and U133 (N_133,In_1680,In_2953);
or U134 (N_134,In_2618,In_3396);
and U135 (N_135,In_4215,In_2395);
nor U136 (N_136,In_4021,In_1597);
or U137 (N_137,In_4185,In_4172);
or U138 (N_138,In_1785,In_658);
and U139 (N_139,In_3103,In_3547);
nor U140 (N_140,In_4731,In_422);
nor U141 (N_141,In_3359,In_3705);
nand U142 (N_142,In_1258,In_3821);
or U143 (N_143,In_3545,In_2158);
and U144 (N_144,In_1210,In_3773);
nand U145 (N_145,In_1405,In_237);
nand U146 (N_146,In_3345,In_689);
nand U147 (N_147,In_3519,In_2324);
nor U148 (N_148,In_429,In_2132);
or U149 (N_149,In_4265,In_1465);
nor U150 (N_150,In_2504,In_4972);
nor U151 (N_151,In_958,In_1995);
nor U152 (N_152,In_2695,In_3459);
and U153 (N_153,In_1029,In_4323);
and U154 (N_154,In_1640,In_1034);
nand U155 (N_155,In_1925,In_3481);
nand U156 (N_156,In_778,In_1615);
nand U157 (N_157,In_3700,In_4174);
nand U158 (N_158,In_1408,In_2600);
or U159 (N_159,In_1584,In_3579);
nand U160 (N_160,In_2162,In_1970);
nor U161 (N_161,In_93,In_925);
nand U162 (N_162,In_1624,In_2539);
xnor U163 (N_163,In_2362,In_218);
nor U164 (N_164,In_3641,In_3187);
nand U165 (N_165,In_1004,In_2635);
or U166 (N_166,In_4712,In_2590);
or U167 (N_167,In_994,In_1420);
or U168 (N_168,In_1434,In_3701);
or U169 (N_169,In_2674,In_3647);
or U170 (N_170,In_4998,In_4674);
nor U171 (N_171,In_3381,In_4641);
xor U172 (N_172,In_3793,In_240);
nand U173 (N_173,In_2741,In_2317);
xnor U174 (N_174,In_4652,In_1607);
nand U175 (N_175,In_4788,In_2105);
and U176 (N_176,In_1883,In_1802);
and U177 (N_177,In_4625,In_691);
nand U178 (N_178,In_4280,In_3073);
and U179 (N_179,In_1200,In_3512);
nand U180 (N_180,In_4398,In_66);
or U181 (N_181,In_1132,In_3915);
nor U182 (N_182,In_3747,In_1195);
nand U183 (N_183,In_511,In_1471);
nor U184 (N_184,In_227,In_320);
nor U185 (N_185,In_3041,In_2899);
and U186 (N_186,In_2425,In_4278);
nand U187 (N_187,In_2081,In_4020);
or U188 (N_188,In_4995,In_1414);
nand U189 (N_189,In_777,In_4596);
nor U190 (N_190,In_2690,In_1107);
and U191 (N_191,In_2483,In_1751);
nand U192 (N_192,In_4591,In_4957);
nor U193 (N_193,In_91,In_4094);
or U194 (N_194,In_3901,In_4823);
or U195 (N_195,In_297,In_4461);
or U196 (N_196,In_56,In_666);
and U197 (N_197,In_628,In_2392);
nor U198 (N_198,In_4633,In_3928);
and U199 (N_199,In_3518,In_1728);
or U200 (N_200,In_4983,In_1151);
and U201 (N_201,In_2058,In_2439);
and U202 (N_202,In_3816,In_53);
nand U203 (N_203,In_3549,In_2351);
nor U204 (N_204,In_990,In_2829);
or U205 (N_205,In_2705,In_362);
or U206 (N_206,In_180,In_413);
nand U207 (N_207,In_1764,In_4353);
nand U208 (N_208,In_2841,In_3446);
nand U209 (N_209,In_4916,In_680);
nand U210 (N_210,In_4044,In_2624);
nand U211 (N_211,In_4409,In_3882);
nand U212 (N_212,In_1554,In_2487);
or U213 (N_213,In_3469,In_4207);
nand U214 (N_214,In_474,In_2180);
xor U215 (N_215,In_2731,In_3158);
or U216 (N_216,In_2751,In_4019);
and U217 (N_217,In_3390,In_458);
xor U218 (N_218,In_571,In_3837);
nor U219 (N_219,In_2502,In_4979);
or U220 (N_220,In_1143,In_3270);
or U221 (N_221,In_700,In_3148);
or U222 (N_222,In_1295,In_1740);
nor U223 (N_223,In_4522,In_3768);
and U224 (N_224,In_1160,In_4588);
xnor U225 (N_225,In_873,In_4009);
nor U226 (N_226,In_727,In_1819);
nor U227 (N_227,In_4038,In_38);
and U228 (N_228,In_683,In_70);
xor U229 (N_229,In_4327,In_992);
and U230 (N_230,In_1581,In_1007);
or U231 (N_231,In_4252,In_4412);
nor U232 (N_232,In_304,In_3688);
or U233 (N_233,In_419,In_4781);
or U234 (N_234,In_418,In_3221);
and U235 (N_235,In_0,In_1701);
nor U236 (N_236,In_1069,In_1497);
or U237 (N_237,In_4001,In_2868);
and U238 (N_238,In_4585,In_3796);
nor U239 (N_239,In_86,In_991);
or U240 (N_240,In_1436,In_2225);
nor U241 (N_241,In_2272,In_2913);
or U242 (N_242,In_1334,In_1243);
nand U243 (N_243,In_4303,In_3465);
nor U244 (N_244,In_2090,In_4846);
or U245 (N_245,In_623,In_1493);
nor U246 (N_246,In_3817,In_200);
nor U247 (N_247,In_3565,In_1134);
nand U248 (N_248,In_145,In_1789);
xor U249 (N_249,In_1480,In_934);
and U250 (N_250,In_4157,In_4561);
nor U251 (N_251,In_4008,In_3633);
or U252 (N_252,In_266,In_1102);
and U253 (N_253,In_3822,In_341);
or U254 (N_254,In_194,In_1801);
and U255 (N_255,In_4201,In_4586);
nand U256 (N_256,In_2071,In_4669);
nor U257 (N_257,In_3902,In_1184);
and U258 (N_258,In_3974,In_2581);
or U259 (N_259,In_4308,In_1767);
nor U260 (N_260,In_46,In_2048);
and U261 (N_261,In_4414,In_4883);
nor U262 (N_262,In_3124,In_3775);
nand U263 (N_263,In_4294,In_3767);
or U264 (N_264,In_2547,In_477);
nand U265 (N_265,In_1230,In_3751);
and U266 (N_266,In_1459,In_2921);
xor U267 (N_267,In_1013,In_4379);
or U268 (N_268,In_868,In_4186);
and U269 (N_269,In_2770,In_837);
or U270 (N_270,In_47,In_253);
or U271 (N_271,In_625,In_2778);
nor U272 (N_272,In_1656,In_4237);
and U273 (N_273,In_4352,In_3514);
or U274 (N_274,In_4090,In_166);
or U275 (N_275,In_4273,In_196);
nor U276 (N_276,In_2792,In_2984);
nand U277 (N_277,In_2236,In_4780);
and U278 (N_278,In_3392,In_4132);
and U279 (N_279,In_3401,In_4702);
or U280 (N_280,In_1805,In_4974);
nor U281 (N_281,In_2981,In_4269);
xnor U282 (N_282,In_4098,In_4305);
and U283 (N_283,In_2597,In_1137);
or U284 (N_284,In_1912,In_258);
nand U285 (N_285,In_192,In_2380);
nand U286 (N_286,In_4238,In_4901);
or U287 (N_287,In_2312,In_3941);
nand U288 (N_288,In_4650,In_165);
nor U289 (N_289,In_1400,In_4545);
nor U290 (N_290,In_4343,In_2306);
and U291 (N_291,In_2148,In_311);
nor U292 (N_292,In_1833,In_3687);
nor U293 (N_293,In_3722,In_871);
nand U294 (N_294,In_168,In_306);
or U295 (N_295,In_242,In_4829);
nand U296 (N_296,In_1193,In_3890);
nand U297 (N_297,In_2691,In_4785);
xor U298 (N_298,In_2398,In_2936);
or U299 (N_299,In_2815,In_1491);
nand U300 (N_300,In_1352,In_4677);
nand U301 (N_301,In_1228,In_4332);
nand U302 (N_302,In_3347,In_3239);
or U303 (N_303,In_4629,In_877);
nor U304 (N_304,In_3752,In_788);
nor U305 (N_305,In_4300,In_4827);
nand U306 (N_306,In_554,In_3717);
and U307 (N_307,In_3606,In_4486);
nand U308 (N_308,In_2254,In_2402);
nand U309 (N_309,In_2401,In_688);
or U310 (N_310,In_1301,In_190);
or U311 (N_311,In_2520,In_1272);
or U312 (N_312,In_2017,In_1240);
nor U313 (N_313,In_4720,In_3896);
or U314 (N_314,In_770,In_2150);
nor U315 (N_315,In_1663,In_1169);
nand U316 (N_316,In_4199,In_1495);
xnor U317 (N_317,In_2801,In_4871);
or U318 (N_318,In_23,In_722);
nor U319 (N_319,In_1550,In_1517);
nor U320 (N_320,In_4915,In_4377);
and U321 (N_321,In_507,In_3942);
and U322 (N_322,In_3792,In_2780);
nor U323 (N_323,In_2349,In_4443);
nor U324 (N_324,In_4760,In_4140);
xnor U325 (N_325,In_4188,In_1067);
nor U326 (N_326,In_2686,In_212);
nor U327 (N_327,In_671,In_1768);
or U328 (N_328,In_512,In_360);
and U329 (N_329,In_2659,In_1489);
and U330 (N_330,In_2846,In_4684);
nand U331 (N_331,In_3405,In_544);
or U332 (N_332,In_1211,In_1838);
and U333 (N_333,In_3900,In_1657);
nor U334 (N_334,In_3978,In_734);
nand U335 (N_335,In_3471,In_3013);
or U336 (N_336,In_3998,In_1628);
nand U337 (N_337,In_3575,In_4584);
or U338 (N_338,In_3778,In_1367);
or U339 (N_339,In_4181,In_2554);
or U340 (N_340,In_880,In_4411);
nor U341 (N_341,In_2376,In_2442);
or U342 (N_342,In_2995,In_3939);
or U343 (N_343,In_1183,In_2693);
xnor U344 (N_344,In_1142,In_3480);
xor U345 (N_345,In_2453,In_1800);
or U346 (N_346,In_3293,In_2146);
or U347 (N_347,In_2452,In_197);
xnor U348 (N_348,In_3936,In_3002);
nor U349 (N_349,In_4158,In_3726);
or U350 (N_350,In_3290,In_4481);
and U351 (N_351,In_2202,In_3452);
nor U352 (N_352,In_1181,In_3611);
or U353 (N_353,In_4600,In_3570);
or U354 (N_354,In_4944,In_2832);
nor U355 (N_355,In_562,In_4046);
nor U356 (N_356,In_3141,In_3819);
nand U357 (N_357,In_21,In_356);
or U358 (N_358,In_2692,In_793);
nand U359 (N_359,In_2491,In_3912);
nor U360 (N_360,In_3801,In_3393);
nor U361 (N_361,In_2923,In_164);
or U362 (N_362,In_3966,In_3404);
and U363 (N_363,In_3468,In_669);
nor U364 (N_364,In_959,In_2192);
xnor U365 (N_365,In_2291,In_4241);
or U366 (N_366,In_420,In_2164);
or U367 (N_367,In_264,In_4786);
xor U368 (N_368,In_715,In_4507);
and U369 (N_369,In_1969,In_87);
and U370 (N_370,In_4648,In_545);
nand U371 (N_371,In_1936,In_2752);
nand U372 (N_372,In_431,In_2725);
nand U373 (N_373,In_2916,In_1076);
nor U374 (N_374,In_2332,In_1563);
or U375 (N_375,In_2381,In_1915);
and U376 (N_376,In_4839,In_521);
or U377 (N_377,In_4123,In_4212);
or U378 (N_378,In_4790,In_2125);
nand U379 (N_379,In_567,In_2416);
nand U380 (N_380,In_4420,In_3587);
nor U381 (N_381,In_2078,In_1156);
nand U382 (N_382,In_866,In_3208);
and U383 (N_383,In_1828,In_2495);
xnor U384 (N_384,In_321,In_430);
nor U385 (N_385,In_2826,In_1733);
nor U386 (N_386,In_2582,In_3232);
or U387 (N_387,In_3810,In_1208);
or U388 (N_388,In_930,In_743);
and U389 (N_389,In_1377,In_4198);
nor U390 (N_390,In_2382,In_2473);
xor U391 (N_391,In_2002,In_1855);
or U392 (N_392,In_2596,In_772);
xnor U393 (N_393,In_1669,In_3494);
xnor U394 (N_394,In_588,In_1246);
or U395 (N_395,In_4755,In_2290);
nor U396 (N_396,In_2963,In_469);
or U397 (N_397,In_4251,In_3996);
nand U398 (N_398,In_1786,In_3489);
nor U399 (N_399,In_681,In_4439);
nand U400 (N_400,In_4320,In_1769);
or U401 (N_401,In_3425,In_3033);
xnor U402 (N_402,In_494,In_2276);
nor U403 (N_403,In_1641,In_1710);
and U404 (N_404,In_2643,In_3248);
nor U405 (N_405,In_1507,In_300);
nand U406 (N_406,In_2768,In_532);
or U407 (N_407,In_2061,In_393);
and U408 (N_408,In_1115,In_490);
or U409 (N_409,In_3388,In_2262);
xnor U410 (N_410,In_1560,In_3615);
nor U411 (N_411,In_117,In_3617);
nor U412 (N_412,In_4518,In_665);
nand U413 (N_413,In_2086,In_695);
nor U414 (N_414,In_2040,In_2032);
nor U415 (N_415,In_207,In_3324);
or U416 (N_416,In_905,In_1646);
and U417 (N_417,In_1928,In_2168);
or U418 (N_418,In_4993,In_3916);
nor U419 (N_419,In_3970,In_2703);
nand U420 (N_420,In_1298,In_4070);
nor U421 (N_421,In_811,In_1820);
and U422 (N_422,In_878,In_88);
nand U423 (N_423,In_523,In_2972);
xor U424 (N_424,In_637,In_3375);
and U425 (N_425,In_1446,In_2756);
and U426 (N_426,In_4465,In_684);
nor U427 (N_427,In_1121,In_1297);
nand U428 (N_428,In_1758,In_3330);
nand U429 (N_429,In_1697,In_4097);
nand U430 (N_430,In_259,In_1252);
nor U431 (N_431,In_854,In_3950);
nor U432 (N_432,In_2458,In_668);
or U433 (N_433,In_2873,In_2052);
xnor U434 (N_434,In_135,In_3235);
xnor U435 (N_435,In_2640,In_3500);
and U436 (N_436,In_4483,In_4870);
and U437 (N_437,In_4,In_1694);
nand U438 (N_438,In_4874,In_2675);
and U439 (N_439,In_1225,In_2068);
nor U440 (N_440,In_3675,In_1985);
or U441 (N_441,In_517,In_2314);
nor U442 (N_442,In_4073,In_172);
nand U443 (N_443,In_1877,In_1330);
and U444 (N_444,In_576,In_3542);
nand U445 (N_445,In_4649,In_4381);
or U446 (N_446,In_4575,In_2279);
or U447 (N_447,In_3094,In_3102);
or U448 (N_448,In_2011,In_1747);
or U449 (N_449,In_1215,In_1515);
or U450 (N_450,In_3543,In_4244);
nand U451 (N_451,In_2796,In_1566);
and U452 (N_452,In_986,In_3648);
or U453 (N_453,In_3082,In_3569);
and U454 (N_454,In_3275,In_204);
and U455 (N_455,In_1110,In_94);
or U456 (N_456,In_3370,In_40);
nor U457 (N_457,In_847,In_3918);
nand U458 (N_458,In_2576,In_3457);
nand U459 (N_459,In_2110,In_1916);
nor U460 (N_460,In_3663,In_1555);
or U461 (N_461,In_2355,In_916);
nand U462 (N_462,In_4137,In_775);
nor U463 (N_463,In_2015,In_3034);
and U464 (N_464,In_2599,In_1627);
nand U465 (N_465,In_2707,In_2560);
and U466 (N_466,In_2233,In_4920);
xnor U467 (N_467,In_2617,In_2014);
and U468 (N_468,In_4214,In_1278);
or U469 (N_469,In_1714,In_4010);
nand U470 (N_470,In_3642,In_2335);
nor U471 (N_471,In_3028,In_4066);
or U472 (N_472,In_1540,In_833);
xnor U473 (N_473,In_4110,In_4961);
nor U474 (N_474,In_1790,In_758);
nand U475 (N_475,In_3558,In_4535);
nand U476 (N_476,In_4654,In_2625);
and U477 (N_477,In_236,In_1306);
or U478 (N_478,In_3965,In_2931);
and U479 (N_479,In_505,In_1466);
or U480 (N_480,In_2793,In_1065);
and U481 (N_481,In_3302,In_1386);
and U482 (N_482,In_2396,In_3618);
and U483 (N_483,In_106,In_1084);
nand U484 (N_484,In_4705,In_1396);
xnor U485 (N_485,In_630,In_896);
and U486 (N_486,In_1175,In_3952);
nand U487 (N_487,In_997,In_1853);
nand U488 (N_488,In_4836,In_823);
nor U489 (N_489,In_3433,In_4223);
or U490 (N_490,In_2639,In_537);
and U491 (N_491,In_453,In_4032);
nand U492 (N_492,In_739,In_2460);
nand U493 (N_493,In_3739,In_1882);
nor U494 (N_494,In_3153,In_646);
nand U495 (N_495,In_714,In_3534);
or U496 (N_496,In_1062,In_2622);
nor U497 (N_497,In_181,In_3220);
and U498 (N_498,In_112,In_2070);
xnor U499 (N_499,In_976,In_4072);
xor U500 (N_500,In_4494,In_2157);
and U501 (N_501,In_801,In_257);
or U502 (N_502,In_2544,In_1073);
and U503 (N_503,In_234,In_4084);
or U504 (N_504,In_2108,In_98);
nor U505 (N_505,In_1217,In_4792);
nand U506 (N_506,In_5,In_1903);
and U507 (N_507,In_4356,In_1270);
or U508 (N_508,In_1637,In_2047);
or U509 (N_509,In_229,In_725);
nand U510 (N_510,In_4509,In_1850);
xor U511 (N_511,In_4463,In_1050);
nand U512 (N_512,In_4844,In_4142);
nand U513 (N_513,In_4177,In_3068);
nor U514 (N_514,In_4745,In_2211);
nor U515 (N_515,In_4382,In_742);
nor U516 (N_516,In_3284,In_4959);
nand U517 (N_517,In_4024,In_4653);
nand U518 (N_518,In_3878,In_4193);
xnor U519 (N_519,In_2568,In_1717);
nor U520 (N_520,In_4275,In_1177);
xnor U521 (N_521,In_3316,In_3682);
and U522 (N_522,In_1033,In_3530);
or U523 (N_523,In_3930,In_2714);
and U524 (N_524,In_2628,In_4096);
and U525 (N_525,In_3496,In_3824);
nor U526 (N_526,In_1579,In_2018);
nor U527 (N_527,In_767,In_699);
nand U528 (N_528,In_3177,In_2912);
or U529 (N_529,In_1196,In_3229);
or U530 (N_530,In_4872,In_3921);
xnor U531 (N_531,In_4344,In_446);
xnor U532 (N_532,In_4963,In_2870);
nor U533 (N_533,In_4782,In_3025);
nor U534 (N_534,In_4063,In_2210);
nor U535 (N_535,In_3639,In_2704);
and U536 (N_536,In_915,In_1542);
nand U537 (N_537,In_1152,In_4852);
nor U538 (N_538,In_3886,In_4805);
and U539 (N_539,In_2585,In_2137);
nor U540 (N_540,In_2948,In_4012);
xnor U541 (N_541,In_272,In_1036);
and U542 (N_542,In_3287,In_403);
and U543 (N_543,In_3438,In_2025);
and U544 (N_544,In_186,In_3668);
and U545 (N_545,In_2144,In_2720);
and U546 (N_546,In_271,In_1212);
or U547 (N_547,In_4552,In_376);
xnor U548 (N_548,In_3352,In_4290);
nor U549 (N_549,In_1242,In_4803);
or U550 (N_550,In_559,In_2806);
xor U551 (N_551,In_1422,In_3760);
or U552 (N_552,In_632,In_3800);
nor U553 (N_553,In_2964,In_2897);
and U554 (N_554,In_4703,In_2173);
nand U555 (N_555,In_3554,In_1692);
nor U556 (N_556,In_4816,In_4687);
or U557 (N_557,In_846,In_2456);
or U558 (N_558,In_3826,In_3353);
or U559 (N_559,In_4878,In_904);
nand U560 (N_560,In_3993,In_648);
and U561 (N_561,In_987,In_2240);
nand U562 (N_562,In_4747,In_3559);
and U563 (N_563,In_4611,In_4408);
nor U564 (N_564,In_1051,In_2463);
and U565 (N_565,In_2862,In_3478);
nand U566 (N_566,In_4889,In_4017);
nand U567 (N_567,In_2263,In_4457);
xor U568 (N_568,In_3211,In_1781);
nand U569 (N_569,In_4962,In_4955);
nand U570 (N_570,In_882,In_629);
or U571 (N_571,In_1285,In_3066);
and U572 (N_572,In_4334,In_301);
nor U573 (N_573,In_1112,In_2493);
nor U574 (N_574,In_964,In_1625);
nand U575 (N_575,In_764,In_4933);
and U576 (N_576,In_2669,In_2571);
nand U577 (N_577,In_14,In_3467);
nand U578 (N_578,In_3131,In_522);
xnor U579 (N_579,In_3012,In_1318);
or U580 (N_580,In_2377,In_2863);
nand U581 (N_581,In_911,In_731);
xnor U582 (N_582,In_4316,In_4401);
or U583 (N_583,In_4319,In_4500);
and U584 (N_584,In_4115,In_4282);
nand U585 (N_585,In_2097,In_4813);
nand U586 (N_586,In_3948,In_3738);
nand U587 (N_587,In_260,In_3458);
nand U588 (N_588,In_3753,In_3014);
nor U589 (N_589,In_2877,In_4884);
nor U590 (N_590,In_1836,In_1376);
or U591 (N_591,In_3605,In_3134);
and U592 (N_592,In_4061,In_3441);
or U593 (N_593,In_1287,In_3185);
or U594 (N_594,In_1930,In_2771);
nand U595 (N_595,In_1002,In_2219);
and U596 (N_596,In_4574,In_1594);
or U597 (N_597,In_2814,In_897);
xnor U598 (N_598,In_1075,In_4715);
and U599 (N_599,In_2131,In_1987);
and U600 (N_600,In_2683,In_2858);
xnor U601 (N_601,In_1707,In_4245);
and U602 (N_602,In_3334,In_3166);
or U603 (N_603,In_932,In_3764);
and U604 (N_604,In_1220,In_2946);
xnor U605 (N_605,In_2440,In_3454);
nand U606 (N_606,In_3529,In_4270);
nand U607 (N_607,In_2417,In_4954);
and U608 (N_608,In_1945,In_221);
nor U609 (N_609,In_4003,In_3280);
and U610 (N_610,In_820,In_3445);
or U611 (N_611,In_163,In_1487);
and U612 (N_612,In_1689,In_2433);
nor U613 (N_613,In_1397,In_921);
or U614 (N_614,In_2153,In_3737);
nand U615 (N_615,In_4202,In_4903);
or U616 (N_616,In_2536,In_1696);
and U617 (N_617,In_3110,In_1437);
or U618 (N_618,In_44,In_4092);
nor U619 (N_619,In_4065,In_295);
nor U620 (N_620,In_1719,In_4514);
and U621 (N_621,In_752,In_3046);
nor U622 (N_622,In_1326,In_488);
or U623 (N_623,In_3790,In_2926);
nor U624 (N_624,In_533,In_4490);
xnor U625 (N_625,In_2094,In_3969);
and U626 (N_626,In_139,In_2035);
xor U627 (N_627,In_2727,In_2346);
nor U628 (N_628,In_886,In_4195);
and U629 (N_629,In_1089,In_2724);
and U630 (N_630,In_3342,In_1104);
nor U631 (N_631,In_557,In_607);
nor U632 (N_632,In_2645,In_2797);
nor U633 (N_633,In_4919,In_3779);
and U634 (N_634,In_2432,In_3413);
and U635 (N_635,In_401,In_906);
xor U636 (N_636,In_67,In_31);
nor U637 (N_637,In_3325,In_2302);
or U638 (N_638,In_1724,In_4796);
and U639 (N_639,In_1066,In_4886);
nor U640 (N_640,In_435,In_4736);
or U641 (N_641,In_122,In_3354);
xnor U642 (N_642,In_392,In_1);
nor U643 (N_643,In_2282,In_1843);
nor U644 (N_644,In_1449,In_1251);
or U645 (N_645,In_713,In_427);
or U646 (N_646,In_1390,In_1118);
nor U647 (N_647,In_2486,In_2359);
or U648 (N_648,In_3204,In_2000);
nor U649 (N_649,In_1671,In_4240);
nand U650 (N_650,In_2134,In_3178);
nor U651 (N_651,In_3323,In_1357);
and U652 (N_652,In_1094,In_1531);
nor U653 (N_653,In_4858,In_1250);
nand U654 (N_654,In_3294,In_1552);
and U655 (N_655,In_4311,In_2026);
nand U656 (N_656,In_2779,In_387);
or U657 (N_657,In_924,In_4221);
nor U658 (N_658,In_4004,In_4607);
nand U659 (N_659,In_1754,In_1070);
and U660 (N_660,In_262,In_706);
nand U661 (N_661,In_4367,In_3661);
or U662 (N_662,In_586,In_1974);
nand U663 (N_663,In_1027,In_4564);
nand U664 (N_664,In_595,In_1947);
nor U665 (N_665,In_1809,In_1138);
and U666 (N_666,In_120,In_4166);
or U667 (N_667,In_3994,In_498);
nand U668 (N_668,In_380,In_497);
nand U669 (N_669,In_216,In_719);
and U670 (N_670,In_1990,In_2885);
or U671 (N_671,In_4885,In_4342);
and U672 (N_672,In_3834,In_836);
nor U673 (N_673,In_2126,In_1880);
and U674 (N_674,In_4173,In_1320);
xor U675 (N_675,In_3659,In_4866);
nand U676 (N_676,In_4664,In_2184);
nand U677 (N_677,In_3249,In_104);
nor U678 (N_678,In_351,In_4899);
nor U679 (N_679,In_797,In_3442);
nand U680 (N_680,In_1477,In_3814);
and U681 (N_681,In_3638,In_3464);
nand U682 (N_682,In_1888,In_2550);
or U683 (N_683,In_3268,In_1923);
and U684 (N_684,In_4007,In_290);
nor U685 (N_685,In_410,In_2649);
nor U686 (N_686,In_3015,In_1950);
nand U687 (N_687,In_3116,In_4330);
nor U688 (N_688,In_2830,In_598);
or U689 (N_689,In_4491,In_3156);
or U690 (N_690,In_838,In_2289);
or U691 (N_691,In_1635,In_2787);
or U692 (N_692,In_4225,In_2517);
and U693 (N_693,In_3664,In_535);
xor U694 (N_694,In_3531,In_3273);
or U695 (N_695,In_3195,In_2364);
or U696 (N_696,In_3734,In_3355);
or U697 (N_697,In_2907,In_4417);
or U698 (N_698,In_3190,In_381);
and U699 (N_699,In_2594,In_1281);
nor U700 (N_700,In_1374,In_888);
or U701 (N_701,In_319,In_1901);
nor U702 (N_702,In_4426,In_128);
nor U703 (N_703,In_1958,In_3272);
nand U704 (N_704,In_2501,In_502);
nor U705 (N_705,In_3237,In_4873);
or U706 (N_706,In_1897,In_2020);
nor U707 (N_707,In_383,In_4267);
nand U708 (N_708,In_395,In_2318);
nand U709 (N_709,In_55,In_4013);
nand U710 (N_710,In_3067,In_184);
or U711 (N_711,In_4848,In_729);
nand U712 (N_712,In_3088,In_2733);
nor U713 (N_713,In_2056,In_4773);
nand U714 (N_714,In_1204,In_2053);
and U715 (N_715,In_3555,In_891);
nand U716 (N_716,In_3036,In_790);
nand U717 (N_717,In_4346,In_1962);
and U718 (N_718,In_3703,In_141);
xnor U719 (N_719,In_687,In_1852);
nand U720 (N_720,In_1353,In_3550);
nand U721 (N_721,In_4691,In_3696);
xor U722 (N_722,In_3716,In_2961);
or U723 (N_723,In_136,In_2859);
and U724 (N_724,In_4051,In_2226);
and U725 (N_725,In_3879,In_966);
nor U726 (N_726,In_4154,In_1576);
or U727 (N_727,In_3870,In_1162);
xor U728 (N_728,In_1650,In_3176);
and U729 (N_729,In_1568,In_3182);
and U730 (N_730,In_3805,In_3622);
or U731 (N_731,In_2589,In_3276);
nand U732 (N_732,In_340,In_3244);
or U733 (N_733,In_4717,In_3260);
nor U734 (N_734,In_1079,In_2135);
and U735 (N_735,In_1858,In_175);
nor U736 (N_736,In_2277,In_2718);
or U737 (N_737,In_2687,In_3803);
nand U738 (N_738,In_1049,In_2369);
and U739 (N_739,In_1834,In_3198);
nand U740 (N_740,In_3096,In_1470);
and U741 (N_741,In_493,In_4402);
and U742 (N_742,In_1934,In_350);
nand U743 (N_743,In_4643,In_4975);
nand U744 (N_744,In_3874,In_2566);
nor U745 (N_745,In_1484,In_4474);
or U746 (N_746,In_4243,In_2869);
nand U747 (N_747,In_4456,In_4080);
and U748 (N_748,In_2974,In_4671);
or U749 (N_749,In_2932,In_841);
and U750 (N_750,In_3597,In_1770);
or U751 (N_751,In_4970,In_4622);
xnor U752 (N_752,In_1265,In_972);
nor U753 (N_753,In_4301,In_1048);
or U754 (N_754,In_3078,In_4479);
xor U755 (N_755,In_1025,In_2915);
nor U756 (N_756,In_3426,In_2084);
nand U757 (N_757,In_451,In_3548);
and U758 (N_758,In_3608,In_4666);
or U759 (N_759,In_773,In_3610);
nand U760 (N_760,In_71,In_3264);
nor U761 (N_761,In_3893,In_4546);
and U762 (N_762,In_2049,In_3508);
nand U763 (N_763,In_4116,In_198);
or U764 (N_764,In_4438,In_132);
or U765 (N_765,In_2304,In_1423);
or U766 (N_766,In_918,In_781);
or U767 (N_767,In_556,In_674);
and U768 (N_768,In_4793,In_4118);
and U769 (N_769,In_1023,In_2530);
or U770 (N_770,In_317,In_2206);
nor U771 (N_771,In_3042,In_2372);
and U772 (N_772,In_426,In_2260);
and U773 (N_773,In_587,In_876);
and U774 (N_774,In_444,In_1508);
nand U775 (N_775,In_4960,In_3856);
or U776 (N_776,In_4102,In_771);
nand U777 (N_777,In_2664,In_1014);
nor U778 (N_778,In_102,In_4645);
and U779 (N_779,In_509,In_1182);
or U780 (N_780,In_578,In_369);
xnor U781 (N_781,In_4138,In_4618);
nor U782 (N_782,In_1268,In_1998);
xnor U783 (N_783,In_296,In_4642);
nand U784 (N_784,In_4397,In_2283);
or U785 (N_785,In_3833,In_1302);
and U786 (N_786,In_1308,In_2824);
nand U787 (N_787,In_3009,In_3707);
and U788 (N_788,In_2270,In_3864);
xor U789 (N_789,In_4328,In_649);
or U790 (N_790,In_2209,In_3130);
or U791 (N_791,In_4317,In_4751);
or U792 (N_792,In_4842,In_2378);
and U793 (N_793,In_1018,In_1989);
and U794 (N_794,In_2481,In_2939);
or U795 (N_795,In_3492,In_2336);
or U796 (N_796,In_1924,In_881);
or U797 (N_797,In_4106,In_2986);
and U798 (N_798,In_4714,In_2941);
nand U799 (N_799,In_4931,In_3212);
xnor U800 (N_800,In_1409,In_2652);
xor U801 (N_801,In_2531,In_4383);
or U802 (N_802,In_2075,In_4124);
nand U803 (N_803,In_4325,In_365);
or U804 (N_804,In_2682,In_819);
nand U805 (N_805,In_2023,In_90);
nor U806 (N_806,In_4089,In_3586);
or U807 (N_807,In_4446,In_1835);
and U808 (N_808,In_276,In_1463);
nand U809 (N_809,In_223,In_2738);
xnor U810 (N_810,In_3343,In_4499);
and U811 (N_811,In_1614,In_4726);
nand U812 (N_812,In_2990,In_64);
and U813 (N_813,In_1725,In_3788);
and U814 (N_814,In_3278,In_3876);
or U815 (N_815,In_4378,In_3098);
or U816 (N_816,In_2565,In_1741);
nor U817 (N_817,In_252,In_2997);
nand U818 (N_818,In_909,In_597);
and U819 (N_819,In_3340,In_2394);
nand U820 (N_820,In_3660,In_4847);
nor U821 (N_821,In_2525,In_3578);
nand U822 (N_822,In_981,In_39);
xor U823 (N_823,In_279,In_3486);
nand U824 (N_824,In_2592,In_3524);
nor U825 (N_825,In_929,In_1166);
and U826 (N_826,In_4700,In_57);
nand U827 (N_827,In_1804,In_756);
nand U828 (N_828,In_2679,In_3947);
and U829 (N_829,In_4526,In_4131);
or U830 (N_830,In_1329,In_1467);
or U831 (N_831,In_4637,In_3511);
nand U832 (N_832,In_4756,In_3372);
or U833 (N_833,In_326,In_263);
nor U834 (N_834,In_470,In_1174);
and U835 (N_835,In_3332,In_4476);
or U836 (N_836,In_4776,In_3924);
nand U837 (N_837,In_1009,In_4468);
nand U838 (N_838,In_2204,In_373);
nor U839 (N_839,In_1873,In_2930);
nor U840 (N_840,In_1481,In_334);
nand U841 (N_841,In_4725,In_347);
xor U842 (N_842,In_2191,In_483);
nand U843 (N_843,In_445,In_2900);
or U844 (N_844,In_1511,In_4197);
or U845 (N_845,In_3999,In_3245);
and U846 (N_846,In_538,In_4860);
or U847 (N_847,In_4554,In_230);
nor U848 (N_848,In_2786,In_581);
or U849 (N_849,In_3713,In_3593);
xnor U850 (N_850,In_254,In_4361);
nor U851 (N_851,In_1441,In_2287);
nand U852 (N_852,In_3851,In_670);
and U853 (N_853,In_1564,In_1403);
xor U854 (N_854,In_3382,In_1321);
nand U855 (N_855,In_89,In_1535);
nor U856 (N_856,In_2667,In_2745);
nand U857 (N_857,In_1083,In_2769);
nand U858 (N_858,In_1577,In_1059);
and U859 (N_859,In_3146,In_696);
and U860 (N_860,In_1824,In_1223);
nor U861 (N_861,In_1911,In_3730);
or U862 (N_862,In_2753,In_4488);
nor U863 (N_863,In_3285,In_2866);
nand U864 (N_864,In_4440,In_1148);
and U865 (N_865,In_2156,In_3410);
and U866 (N_866,In_1345,In_2444);
or U867 (N_867,In_4028,In_1673);
xor U868 (N_868,In_4890,In_150);
nor U869 (N_869,In_1042,In_1920);
nor U870 (N_870,In_3429,In_2430);
or U871 (N_871,In_2472,In_643);
and U872 (N_872,In_324,In_3364);
and U873 (N_873,In_3646,In_3624);
and U874 (N_874,In_162,In_3054);
nand U875 (N_875,In_28,In_4162);
or U876 (N_876,In_920,In_379);
nand U877 (N_877,In_4108,In_3321);
nor U878 (N_878,In_2216,In_3908);
or U879 (N_879,In_478,In_812);
nand U880 (N_880,In_3616,In_2878);
and U881 (N_881,In_558,In_4218);
nor U882 (N_882,In_1186,In_4689);
and U883 (N_883,In_111,In_2772);
or U884 (N_884,In_2400,In_485);
nand U885 (N_885,In_783,In_3818);
xor U886 (N_886,In_182,In_2019);
xor U887 (N_887,In_2098,In_2777);
and U888 (N_888,In_4555,In_539);
nand U889 (N_889,In_4469,In_3919);
and U890 (N_890,In_1862,In_2259);
and U891 (N_891,In_1026,In_4911);
and U892 (N_892,In_3958,In_1865);
nor U893 (N_893,In_4171,In_2464);
nand U894 (N_894,In_2169,In_2527);
xor U895 (N_895,In_1411,In_354);
and U896 (N_896,In_3741,In_1712);
nand U897 (N_897,In_2205,In_489);
or U898 (N_898,In_3378,In_4935);
nand U899 (N_899,In_4496,In_4708);
or U900 (N_900,In_4929,In_1274);
nor U901 (N_901,In_2072,In_763);
nor U902 (N_902,In_813,In_3411);
nand U903 (N_903,In_2194,In_3697);
xnor U904 (N_904,In_3384,In_4504);
or U905 (N_905,In_4798,In_3194);
nand U906 (N_906,In_35,In_1310);
nand U907 (N_907,In_1203,In_3183);
or U908 (N_908,In_3422,In_4524);
nor U909 (N_909,In_3255,In_885);
nand U910 (N_910,In_766,In_2457);
xnor U911 (N_911,In_2166,In_1399);
and U912 (N_912,In_4058,In_3231);
nor U913 (N_913,In_4838,In_4924);
nand U914 (N_914,In_17,In_4807);
nor U915 (N_915,In_482,In_2713);
nor U916 (N_916,In_697,In_4351);
and U917 (N_917,In_414,In_726);
nand U918 (N_918,In_1327,In_3379);
nor U919 (N_919,In_2408,In_1365);
nor U920 (N_920,In_3718,In_1603);
or U921 (N_921,In_3895,In_4403);
or U922 (N_922,In_516,In_1558);
nand U923 (N_923,In_596,In_402);
nand U924 (N_924,In_3683,In_1978);
nand U925 (N_925,In_3759,In_2909);
and U926 (N_926,In_3304,In_2069);
nor U927 (N_927,In_4307,In_386);
and U928 (N_928,In_1780,In_3126);
nor U929 (N_929,In_1890,In_1682);
or U930 (N_930,In_2285,In_3953);
or U931 (N_931,In_2155,In_1889);
xnor U932 (N_932,In_2882,In_1039);
or U933 (N_933,In_1933,In_928);
xor U934 (N_934,In_1071,In_2563);
or U935 (N_935,In_579,In_400);
and U936 (N_936,In_1054,In_3571);
and U937 (N_937,In_4180,In_352);
nor U938 (N_938,In_3546,In_2817);
xor U939 (N_939,In_4027,In_3576);
and U940 (N_940,In_248,In_2776);
nor U941 (N_941,In_2235,In_3163);
or U942 (N_942,In_1127,In_4182);
nor U943 (N_943,In_2584,In_592);
or U944 (N_944,In_3836,In_900);
xnor U945 (N_945,In_33,In_3356);
nand U946 (N_946,In_4272,In_806);
and U947 (N_947,In_1848,In_1942);
nor U948 (N_948,In_2516,In_789);
nor U949 (N_949,In_2199,In_2106);
nand U950 (N_950,In_2513,In_391);
and U951 (N_951,In_2124,In_1774);
nand U952 (N_952,In_3590,In_1807);
nand U953 (N_953,In_720,In_4375);
nor U954 (N_954,In_3673,In_4248);
nor U955 (N_955,In_4321,In_2537);
and U956 (N_956,In_913,In_1311);
nor U957 (N_957,In_2767,In_3725);
nand U958 (N_958,In_2121,In_4867);
nor U959 (N_959,In_2033,In_503);
nor U960 (N_960,In_4734,In_844);
or U961 (N_961,In_2740,In_4897);
and U962 (N_962,In_2413,In_1312);
xor U963 (N_963,In_22,In_4430);
or U964 (N_964,In_4863,In_270);
or U965 (N_965,In_1700,In_4122);
nor U966 (N_966,In_747,In_1305);
or U967 (N_967,In_1621,In_462);
xor U968 (N_968,In_590,In_2092);
or U969 (N_969,In_4676,In_4029);
xnor U970 (N_970,In_3651,In_985);
or U971 (N_971,In_4542,In_4937);
and U972 (N_972,In_892,In_4169);
nand U973 (N_973,In_977,In_705);
nor U974 (N_974,In_4662,In_2013);
or U975 (N_975,In_3035,In_4289);
nor U976 (N_976,In_157,In_3455);
nand U977 (N_977,In_1126,In_3216);
or U978 (N_978,In_3490,In_3932);
and U979 (N_979,In_2354,In_1100);
and U980 (N_980,In_1583,In_563);
or U981 (N_981,In_1991,In_2147);
nor U982 (N_982,In_2934,In_1672);
or U983 (N_983,In_1793,In_2055);
xor U984 (N_984,In_154,In_1022);
and U985 (N_985,In_267,In_529);
or U986 (N_986,In_3997,In_4042);
and U987 (N_987,In_3416,In_3491);
nand U988 (N_988,In_4145,In_1875);
and U989 (N_989,In_1693,In_2203);
or U990 (N_990,In_1666,In_126);
and U991 (N_991,In_4424,In_2804);
nor U992 (N_992,In_2303,In_3064);
nor U993 (N_993,In_4460,In_2141);
or U994 (N_994,In_1735,In_3667);
nand U995 (N_995,In_3219,In_4828);
nor U996 (N_996,In_476,In_1378);
nand U997 (N_997,In_4617,In_3566);
xor U998 (N_998,In_287,In_1325);
and U999 (N_999,In_2099,In_4286);
and U1000 (N_1000,In_2036,In_4784);
nor U1001 (N_1001,In_3487,In_2888);
and U1002 (N_1002,In_4722,In_2737);
nor U1003 (N_1003,In_3614,In_4907);
or U1004 (N_1004,In_548,In_1053);
nor U1005 (N_1005,In_1081,In_1363);
nand U1006 (N_1006,In_3240,In_515);
nand U1007 (N_1007,In_1784,In_4415);
nand U1008 (N_1008,In_3241,In_824);
nor U1009 (N_1009,In_3253,In_2419);
nor U1010 (N_1010,In_2996,In_1668);
nand U1011 (N_1011,In_616,In_4030);
or U1012 (N_1012,In_2208,In_4508);
nor U1013 (N_1013,In_3044,In_2595);
nor U1014 (N_1014,In_3258,In_2128);
nand U1015 (N_1015,In_4967,In_1986);
xor U1016 (N_1016,In_746,In_2746);
nand U1017 (N_1017,In_848,In_2010);
and U1018 (N_1018,In_4769,In_4076);
or U1019 (N_1019,In_686,In_1949);
nor U1020 (N_1020,In_531,In_707);
xnor U1021 (N_1021,In_2305,In_3269);
and U1022 (N_1022,In_4619,In_1057);
nor U1023 (N_1023,In_3644,In_3813);
nor U1024 (N_1024,In_3326,In_3119);
and U1025 (N_1025,In_4927,In_1226);
nand U1026 (N_1026,In_275,In_457);
nand U1027 (N_1027,In_491,In_3809);
nand U1028 (N_1028,In_3881,In_3463);
nor U1029 (N_1029,In_3420,In_2969);
nand U1030 (N_1030,In_834,In_4121);
nor U1031 (N_1031,In_757,In_1574);
nand U1032 (N_1032,In_4940,In_4608);
and U1033 (N_1033,In_3596,In_60);
and U1034 (N_1034,In_4513,In_43);
and U1035 (N_1035,In_3289,In_4117);
nor U1036 (N_1036,In_4568,In_1307);
nor U1037 (N_1037,In_2267,In_936);
or U1038 (N_1038,In_4636,In_4820);
nand U1039 (N_1039,In_2174,In_4431);
or U1040 (N_1040,In_138,In_541);
or U1041 (N_1041,In_3857,In_4388);
and U1042 (N_1042,In_1647,In_461);
nor U1043 (N_1043,In_979,In_375);
and U1044 (N_1044,In_1871,In_2891);
nor U1045 (N_1045,In_95,In_2037);
nand U1046 (N_1046,In_1851,In_4335);
or U1047 (N_1047,In_217,In_1443);
and U1048 (N_1048,In_3815,In_1266);
nor U1049 (N_1049,In_995,In_3907);
nor U1050 (N_1050,In_2701,In_4732);
nand U1051 (N_1051,In_3020,In_2498);
nand U1052 (N_1052,In_1000,In_3503);
nand U1053 (N_1053,In_1941,In_4393);
nor U1054 (N_1054,In_2195,In_3516);
nor U1055 (N_1055,In_336,In_1937);
or U1056 (N_1056,In_2938,In_2492);
xor U1057 (N_1057,In_2298,In_3781);
nor U1058 (N_1058,In_2313,In_3462);
nand U1059 (N_1059,In_4906,In_3552);
and U1060 (N_1060,In_3679,In_2587);
nand U1061 (N_1061,In_3572,In_233);
or U1062 (N_1062,In_4149,In_191);
or U1063 (N_1063,In_574,In_3303);
or U1064 (N_1064,In_1720,In_472);
xor U1065 (N_1065,In_3845,In_4179);
or U1066 (N_1066,In_3858,In_1021);
nor U1067 (N_1067,In_2562,In_908);
xor U1068 (N_1068,In_3595,In_1561);
nand U1069 (N_1069,In_3074,In_4926);
nor U1070 (N_1070,In_4190,In_4040);
or U1071 (N_1071,In_2821,In_1530);
and U1072 (N_1072,In_454,In_1731);
nand U1073 (N_1073,In_2991,In_2356);
or U1074 (N_1074,In_2136,In_2475);
and U1075 (N_1075,In_1490,In_3029);
and U1076 (N_1076,In_2076,In_2238);
or U1077 (N_1077,In_1430,In_609);
and U1078 (N_1078,In_2427,In_1144);
nor U1079 (N_1079,In_1544,In_2251);
or U1080 (N_1080,In_716,In_3132);
and U1081 (N_1081,In_433,In_2258);
or U1082 (N_1082,In_940,In_4875);
nor U1083 (N_1083,In_2895,In_3440);
and U1084 (N_1084,In_829,In_2288);
or U1085 (N_1085,In_1473,In_4592);
xor U1086 (N_1086,In_3327,In_2102);
nor U1087 (N_1087,In_4743,In_2003);
nand U1088 (N_1088,In_2470,In_4104);
nor U1089 (N_1089,In_2231,In_659);
nor U1090 (N_1090,In_202,In_3746);
and U1091 (N_1091,In_1336,In_2955);
nand U1092 (N_1092,In_4298,In_151);
nor U1093 (N_1093,In_2593,In_2605);
or U1094 (N_1094,In_1011,In_4532);
nor U1095 (N_1095,In_4153,In_1759);
nand U1096 (N_1096,In_4812,In_2338);
xor U1097 (N_1097,In_2883,In_4263);
nor U1098 (N_1098,In_3888,In_2989);
nand U1099 (N_1099,In_280,In_65);
nand U1100 (N_1100,In_3210,In_2227);
nand U1101 (N_1101,In_4216,In_3357);
nor U1102 (N_1102,In_4577,In_754);
and U1103 (N_1103,In_1380,In_3374);
nand U1104 (N_1104,In_2672,In_1994);
nor U1105 (N_1105,In_1972,In_4938);
or U1106 (N_1106,In_1370,In_2904);
nor U1107 (N_1107,In_1091,In_782);
nand U1108 (N_1108,In_3338,In_2120);
nor U1109 (N_1109,In_4544,In_3899);
or U1110 (N_1110,In_899,In_2129);
and U1111 (N_1111,In_148,In_2295);
nand U1112 (N_1112,In_4380,In_1111);
or U1113 (N_1113,In_4833,In_2558);
or U1114 (N_1114,In_1314,In_2087);
nand U1115 (N_1115,In_4923,In_1346);
or U1116 (N_1116,In_1529,In_779);
nor U1117 (N_1117,In_998,In_2951);
or U1118 (N_1118,In_4896,In_1438);
and U1119 (N_1119,In_4372,In_3795);
and U1120 (N_1120,In_1261,In_2043);
or U1121 (N_1121,In_1041,In_2774);
nand U1122 (N_1122,In_4768,In_1665);
xnor U1123 (N_1123,In_4052,In_600);
nand U1124 (N_1124,In_499,In_3955);
nand U1125 (N_1125,In_3300,In_1585);
and U1126 (N_1126,In_1812,In_4562);
or U1127 (N_1127,In_4531,In_2570);
and U1128 (N_1128,In_1454,In_3085);
and U1129 (N_1129,In_3867,In_1092);
or U1130 (N_1130,In_2008,In_2755);
and U1131 (N_1131,In_2807,In_1366);
and U1132 (N_1132,In_1727,In_1854);
nand U1133 (N_1133,In_4587,In_4167);
nor U1134 (N_1134,In_3283,In_2249);
nor U1135 (N_1135,In_3140,In_3634);
nand U1136 (N_1136,In_3005,In_3756);
and U1137 (N_1137,In_3509,In_4614);
xor U1138 (N_1138,In_1259,In_2875);
and U1139 (N_1139,In_367,In_2245);
nand U1140 (N_1140,In_411,In_1061);
or U1141 (N_1141,In_800,In_1653);
or U1142 (N_1142,In_2038,In_4754);
or U1143 (N_1143,In_4595,In_2925);
nand U1144 (N_1144,In_4310,In_1757);
nor U1145 (N_1145,In_1500,In_467);
nor U1146 (N_1146,In_1244,In_2538);
and U1147 (N_1147,In_3181,In_147);
nor U1148 (N_1148,In_2663,In_2296);
nand U1149 (N_1149,In_1350,In_3252);
nor U1150 (N_1150,In_103,In_2009);
or U1151 (N_1151,In_1233,In_1249);
or U1152 (N_1152,In_4506,In_2881);
and U1153 (N_1153,In_3225,In_124);
nor U1154 (N_1154,In_1513,In_3672);
and U1155 (N_1155,In_3307,In_2297);
xor U1156 (N_1156,In_2499,In_859);
or U1157 (N_1157,In_361,In_549);
and U1158 (N_1158,In_2161,In_4296);
or U1159 (N_1159,In_3843,In_4125);
and U1160 (N_1160,In_1795,In_2623);
nand U1161 (N_1161,In_4156,In_434);
or U1162 (N_1162,In_2046,In_3058);
nand U1163 (N_1163,In_1860,In_2021);
nand U1164 (N_1164,In_4534,In_3904);
nand U1165 (N_1165,In_2976,In_3472);
nand U1166 (N_1166,In_3935,In_2528);
and U1167 (N_1167,In_999,In_2943);
and U1168 (N_1168,In_4753,In_635);
nand U1169 (N_1169,In_2060,In_4541);
xnor U1170 (N_1170,In_1527,In_2542);
nand U1171 (N_1171,In_1404,In_3349);
or U1172 (N_1172,In_1661,In_3424);
and U1173 (N_1173,In_3341,In_2799);
or U1174 (N_1174,In_4060,In_2889);
nand U1175 (N_1175,In_534,In_4450);
or U1176 (N_1176,In_4437,In_4570);
or U1177 (N_1177,In_3709,In_4247);
nand U1178 (N_1178,In_4170,In_4191);
and U1179 (N_1179,In_1205,In_4859);
and U1180 (N_1180,In_3447,In_3408);
and U1181 (N_1181,In_1736,In_2171);
nor U1182 (N_1182,In_2610,In_1996);
nand U1183 (N_1183,In_4484,In_4394);
nand U1184 (N_1184,In_4413,In_4069);
and U1185 (N_1185,In_4765,In_3564);
or U1186 (N_1186,In_4730,In_4616);
nand U1187 (N_1187,In_3417,In_721);
nand U1188 (N_1188,In_2005,In_1921);
nand U1189 (N_1189,In_3674,In_3206);
and U1190 (N_1190,In_4160,In_4349);
and U1191 (N_1191,In_2145,In_3037);
nor U1192 (N_1192,In_1706,In_36);
xor U1193 (N_1193,In_1221,In_2529);
nor U1194 (N_1194,In_2308,In_3159);
nand U1195 (N_1195,In_408,In_2406);
nor U1196 (N_1196,In_7,In_645);
and U1197 (N_1197,In_4693,In_249);
nor U1198 (N_1198,In_3541,In_1387);
nand U1199 (N_1199,In_1476,In_4996);
nand U1200 (N_1200,In_4037,In_2063);
and U1201 (N_1201,In_4054,In_1821);
nor U1202 (N_1202,In_63,In_1690);
xor U1203 (N_1203,In_817,In_4143);
nor U1204 (N_1204,In_1543,In_3823);
and U1205 (N_1205,In_4268,In_2337);
nand U1206 (N_1206,In_1504,In_1772);
nand U1207 (N_1207,In_1154,In_1440);
and U1208 (N_1208,In_2833,In_3106);
nor U1209 (N_1209,In_970,In_3783);
nor U1210 (N_1210,In_961,In_4621);
and U1211 (N_1211,In_4406,In_724);
xnor U1212 (N_1212,In_1783,In_4520);
xor U1213 (N_1213,In_4824,In_633);
nand U1214 (N_1214,In_4449,In_3113);
nor U1215 (N_1215,In_1289,In_247);
nor U1216 (N_1216,In_805,In_3981);
and U1217 (N_1217,In_2968,In_2506);
nand U1218 (N_1218,In_1602,In_1749);
nor U1219 (N_1219,In_1185,In_4880);
xor U1220 (N_1220,In_496,In_1827);
and U1221 (N_1221,In_75,In_3003);
or U1222 (N_1222,In_97,In_2117);
and U1223 (N_1223,In_372,In_717);
and U1224 (N_1224,In_4752,In_1633);
or U1225 (N_1225,In_4219,In_1045);
nand U1226 (N_1226,In_2415,In_815);
and U1227 (N_1227,In_1632,In_604);
nand U1228 (N_1228,In_2451,In_3265);
or U1229 (N_1229,In_12,In_2782);
and U1230 (N_1230,In_4675,In_1264);
nor U1231 (N_1231,In_2027,In_3883);
or U1232 (N_1232,In_3335,In_328);
xor U1233 (N_1233,In_4908,In_177);
xnor U1234 (N_1234,In_2694,In_2971);
xor U1235 (N_1235,In_255,In_3560);
and U1236 (N_1236,In_1840,In_1384);
xor U1237 (N_1237,In_1514,In_3913);
nand U1238 (N_1238,In_792,In_956);
nor U1239 (N_1239,In_310,In_3125);
and U1240 (N_1240,In_3581,In_2212);
nor U1241 (N_1241,In_2831,In_2041);
xor U1242 (N_1242,In_4639,In_473);
or U1243 (N_1243,In_3267,In_3314);
and U1244 (N_1244,In_3678,In_3620);
xor U1245 (N_1245,In_358,In_1167);
or U1246 (N_1246,In_3430,In_3785);
or U1247 (N_1247,In_2924,In_4744);
nand U1248 (N_1248,In_2001,In_1526);
and U1249 (N_1249,In_780,In_3840);
and U1250 (N_1250,In_1030,In_1609);
and U1251 (N_1251,In_3161,In_1150);
or U1252 (N_1252,In_3386,In_2329);
and U1253 (N_1253,In_3279,In_4235);
xnor U1254 (N_1254,In_2636,In_1322);
and U1255 (N_1255,In_3691,In_4783);
and U1256 (N_1256,In_4336,In_639);
xor U1257 (N_1257,In_2836,In_1518);
and U1258 (N_1258,In_504,In_4306);
and U1259 (N_1259,In_464,In_2431);
xor U1260 (N_1260,In_4795,In_4656);
and U1261 (N_1261,In_4801,In_1649);
xor U1262 (N_1262,In_744,In_405);
or U1263 (N_1263,In_428,In_842);
nand U1264 (N_1264,In_1522,In_1416);
and U1265 (N_1265,In_2838,In_4830);
nand U1266 (N_1266,In_3537,In_787);
and U1267 (N_1267,In_552,In_3766);
or U1268 (N_1268,In_4026,In_61);
and U1269 (N_1269,In_2244,In_3677);
nor U1270 (N_1270,In_1797,In_2662);
nand U1271 (N_1271,In_513,In_2301);
and U1272 (N_1272,In_4467,In_738);
or U1273 (N_1273,In_528,In_2644);
nand U1274 (N_1274,In_4918,In_3117);
nor U1275 (N_1275,In_4492,In_4779);
nor U1276 (N_1276,In_1362,In_3436);
nand U1277 (N_1277,In_2928,In_1525);
or U1278 (N_1278,In_3,In_281);
nor U1279 (N_1279,In_3118,In_4271);
and U1280 (N_1280,In_73,In_385);
nand U1281 (N_1281,In_3377,In_331);
or U1282 (N_1282,In_4549,In_1643);
and U1283 (N_1283,In_3891,In_1168);
nand U1284 (N_1284,In_506,In_3319);
nand U1285 (N_1285,In_4627,In_1164);
or U1286 (N_1286,In_3427,In_2598);
or U1287 (N_1287,In_1176,In_2107);
or U1288 (N_1288,In_606,In_4895);
xor U1289 (N_1289,In_4242,In_2474);
nor U1290 (N_1290,In_1533,In_41);
nand U1291 (N_1291,In_3019,In_4200);
or U1292 (N_1292,In_398,In_3328);
xor U1293 (N_1293,In_855,In_3761);
and U1294 (N_1294,In_436,In_3515);
or U1295 (N_1295,In_3164,In_3719);
and U1296 (N_1296,In_107,In_2246);
or U1297 (N_1297,In_2865,In_3083);
and U1298 (N_1298,In_3582,In_243);
nand U1299 (N_1299,In_1114,In_2330);
and U1300 (N_1300,In_1892,In_1681);
or U1301 (N_1301,In_620,In_4350);
nor U1302 (N_1302,In_1593,In_3039);
xnor U1303 (N_1303,In_4433,In_1335);
nor U1304 (N_1304,In_1761,In_3360);
or U1305 (N_1305,In_4681,In_1427);
or U1306 (N_1306,In_2847,In_1296);
or U1307 (N_1307,In_110,In_611);
nor U1308 (N_1308,In_3706,In_3812);
nand U1309 (N_1309,In_1213,In_4683);
nand U1310 (N_1310,In_2678,In_3142);
nor U1311 (N_1311,In_302,In_939);
and U1312 (N_1312,In_2229,In_1448);
nor U1313 (N_1313,In_525,In_4419);
and U1314 (N_1314,In_4559,In_2761);
nor U1315 (N_1315,In_1537,In_3665);
and U1316 (N_1316,In_342,In_1087);
nor U1317 (N_1317,In_2803,In_1019);
nand U1318 (N_1318,In_4302,In_2299);
nor U1319 (N_1319,In_1068,In_4360);
or U1320 (N_1320,In_3310,In_4074);
nor U1321 (N_1321,In_4997,In_2794);
or U1322 (N_1322,In_864,In_2637);
nand U1323 (N_1323,In_617,In_2348);
or U1324 (N_1324,In_4285,In_3317);
or U1325 (N_1325,In_1239,In_690);
or U1326 (N_1326,In_3087,In_3120);
nand U1327 (N_1327,In_1082,In_907);
nand U1328 (N_1328,In_239,In_4357);
xor U1329 (N_1329,In_51,In_974);
and U1330 (N_1330,In_1699,In_437);
or U1331 (N_1331,In_4602,In_1456);
and U1332 (N_1332,In_736,In_2812);
nor U1333 (N_1333,In_1907,In_1447);
nand U1334 (N_1334,In_4571,In_826);
and U1335 (N_1335,In_4119,In_4711);
nor U1336 (N_1336,In_1123,In_3742);
nor U1337 (N_1337,In_3418,In_2676);
and U1338 (N_1338,In_346,In_2490);
or U1339 (N_1339,In_2384,In_2809);
and U1340 (N_1340,In_18,In_1284);
nand U1341 (N_1341,In_2732,In_4657);
nand U1342 (N_1342,In_2193,In_1975);
xor U1343 (N_1343,In_526,In_1172);
and U1344 (N_1344,In_1283,In_1412);
or U1345 (N_1345,In_4452,In_4857);
nor U1346 (N_1346,In_3169,In_4392);
nand U1347 (N_1347,In_3282,In_1872);
and U1348 (N_1348,In_968,In_2519);
xor U1349 (N_1349,In_2608,In_3789);
nand U1350 (N_1350,In_315,In_3444);
and U1351 (N_1351,In_2478,In_4638);
xor U1352 (N_1352,In_2835,In_3257);
nor U1353 (N_1353,In_3070,In_3782);
and U1354 (N_1354,In_1158,In_1488);
nor U1355 (N_1355,In_4817,In_2388);
or U1356 (N_1356,In_840,In_1870);
nor U1357 (N_1357,In_3892,In_1445);
or U1358 (N_1358,In_4766,In_226);
nand U1359 (N_1359,In_561,In_2552);
nor U1360 (N_1360,In_1662,In_2653);
and U1361 (N_1361,In_540,In_2646);
nand U1362 (N_1362,In_3154,In_4337);
nand U1363 (N_1363,In_3567,In_123);
nor U1364 (N_1364,In_3091,In_1008);
nor U1365 (N_1365,In_4579,In_4719);
and U1366 (N_1366,In_4843,In_3499);
xnor U1367 (N_1367,In_2661,In_2890);
nand U1368 (N_1368,In_2764,In_4359);
nand U1369 (N_1369,In_1299,In_1613);
nor U1370 (N_1370,In_2917,In_487);
or U1371 (N_1371,In_4284,In_2323);
xnor U1372 (N_1372,In_2294,In_1355);
nand U1373 (N_1373,In_2230,In_2633);
and U1374 (N_1374,In_2390,In_1058);
and U1375 (N_1375,In_1197,In_4740);
nand U1376 (N_1376,In_2163,In_1410);
nand U1377 (N_1377,In_2322,In_2665);
nand U1378 (N_1378,In_3847,In_4239);
and U1379 (N_1379,In_2723,In_3584);
and U1380 (N_1380,In_4345,In_1811);
nand U1381 (N_1381,In_1623,In_1676);
or U1382 (N_1382,In_4291,In_1787);
xnor U1383 (N_1383,In_3979,In_1190);
nor U1384 (N_1384,In_1982,In_4876);
nor U1385 (N_1385,In_1893,In_1458);
nand U1386 (N_1386,In_1475,In_4075);
and U1387 (N_1387,In_3841,In_48);
or U1388 (N_1388,In_2556,In_4898);
nand U1389 (N_1389,In_2113,In_2151);
xor U1390 (N_1390,In_3434,In_2657);
and U1391 (N_1391,In_396,In_4853);
xor U1392 (N_1392,In_3702,In_4640);
nand U1393 (N_1393,In_3202,In_4281);
and U1394 (N_1394,In_4888,In_3112);
and U1395 (N_1395,In_2569,In_92);
nand U1396 (N_1396,In_2920,In_799);
xor U1397 (N_1397,In_1159,In_2919);
nand U1398 (N_1398,In_4386,In_4068);
nor U1399 (N_1399,In_957,In_3045);
nand U1400 (N_1400,In_2743,In_74);
or U1401 (N_1401,In_2854,In_1715);
nor U1402 (N_1402,In_2781,In_1955);
xnor U1403 (N_1403,In_4845,In_4209);
or U1404 (N_1404,In_3497,In_4686);
and U1405 (N_1405,In_3875,In_256);
nand U1406 (N_1406,In_3628,In_1263);
and U1407 (N_1407,In_3133,In_2080);
nand U1408 (N_1408,In_4250,In_3306);
or U1409 (N_1409,In_2006,In_2935);
nor U1410 (N_1410,In_1155,In_4949);
xnor U1411 (N_1411,In_4864,In_3007);
nand U1412 (N_1412,In_1826,In_2112);
and U1413 (N_1413,In_3852,In_187);
and U1414 (N_1414,In_3254,In_2994);
nor U1415 (N_1415,In_2748,In_926);
xor U1416 (N_1416,In_3108,In_2952);
nand U1417 (N_1417,In_3808,In_3476);
nor U1418 (N_1418,In_988,In_268);
or U1419 (N_1419,In_455,In_3749);
xor U1420 (N_1420,In_2853,In_285);
nor U1421 (N_1421,In_508,In_3052);
nor U1422 (N_1422,In_3825,In_3711);
nor U1423 (N_1423,In_2315,In_3031);
xor U1424 (N_1424,In_1943,In_2631);
or U1425 (N_1425,In_3456,In_2088);
nand U1426 (N_1426,In_3032,In_3223);
nand U1427 (N_1427,In_2339,In_4647);
and U1428 (N_1428,In_1562,In_292);
nand U1429 (N_1429,In_294,In_887);
nand U1430 (N_1430,In_4502,In_3147);
or U1431 (N_1431,In_2083,In_1256);
and U1432 (N_1432,In_524,In_4550);
and U1433 (N_1433,In_273,In_2668);
and U1434 (N_1434,In_3049,In_3171);
or U1435 (N_1435,In_872,In_1128);
nand U1436 (N_1436,In_3854,In_3076);
or U1437 (N_1437,In_481,In_1521);
and U1438 (N_1438,In_3985,In_4810);
or U1439 (N_1439,In_3488,In_82);
and U1440 (N_1440,In_1502,In_3271);
nor U1441 (N_1441,In_4232,In_2606);
nor U1442 (N_1442,In_3535,In_3371);
nand U1443 (N_1443,In_3188,In_77);
and U1444 (N_1444,In_4688,In_4035);
or U1445 (N_1445,In_4477,In_114);
or U1446 (N_1446,In_231,In_4348);
nor U1447 (N_1447,In_1267,In_4055);
and U1448 (N_1448,In_599,In_4851);
and U1449 (N_1449,In_4749,In_188);
or U1450 (N_1450,In_1743,In_2906);
xor U1451 (N_1451,In_189,In_3604);
or U1452 (N_1452,In_325,In_2200);
nor U1453 (N_1453,In_4309,In_2850);
nor U1454 (N_1454,In_3157,In_1926);
or U1455 (N_1455,In_1479,In_1868);
nand U1456 (N_1456,In_2278,In_2320);
nor U1457 (N_1457,In_3137,In_879);
and U1458 (N_1458,In_3485,In_76);
or U1459 (N_1459,In_3849,In_2480);
or U1460 (N_1460,In_2077,In_1734);
or U1461 (N_1461,In_2232,In_4533);
nand U1462 (N_1462,In_2681,In_816);
nand U1463 (N_1463,In_3362,In_3213);
or U1464 (N_1464,In_4370,In_589);
nand U1465 (N_1465,In_2119,In_4165);
or U1466 (N_1466,In_4144,In_4599);
or U1467 (N_1467,In_839,In_4678);
and U1468 (N_1468,In_4679,In_4988);
and U1469 (N_1469,In_1626,In_4581);
nor U1470 (N_1470,In_3477,In_3754);
nor U1471 (N_1471,In_3602,In_3397);
and U1472 (N_1472,In_1333,In_2405);
and U1473 (N_1473,In_416,In_2221);
nand U1474 (N_1474,In_1688,In_3598);
xnor U1475 (N_1475,In_3128,In_2697);
nor U1476 (N_1476,In_2802,In_1028);
nand U1477 (N_1477,In_3770,In_1291);
nand U1478 (N_1478,In_1017,In_2567);
xnor U1479 (N_1479,In_1702,In_42);
or U1480 (N_1480,In_3681,In_1364);
and U1481 (N_1481,In_2360,In_1234);
nor U1482 (N_1482,In_4391,In_3365);
nand U1483 (N_1483,In_2373,In_3715);
or U1484 (N_1484,In_2546,In_1929);
or U1485 (N_1485,In_156,In_4086);
or U1486 (N_1486,In_2443,In_4045);
and U1487 (N_1487,In_1856,In_4389);
or U1488 (N_1488,In_3361,In_2910);
and U1489 (N_1489,In_3872,In_2503);
nand U1490 (N_1490,In_4213,In_1451);
and U1491 (N_1491,In_2307,In_708);
or U1492 (N_1492,In_4716,In_1309);
and U1493 (N_1493,In_2822,In_2937);
and U1494 (N_1494,In_4624,In_662);
or U1495 (N_1495,In_3060,In_2522);
nand U1496 (N_1496,In_1823,In_4913);
nor U1497 (N_1497,In_3200,In_1756);
nor U1498 (N_1498,In_329,In_2673);
nand U1499 (N_1499,In_10,In_2579);
nor U1500 (N_1500,In_2334,In_4593);
and U1501 (N_1501,In_1260,In_4184);
nor U1502 (N_1502,In_828,In_4260);
or U1503 (N_1503,In_2973,In_4811);
nand U1504 (N_1504,In_2750,In_2139);
nand U1505 (N_1505,In_3493,In_3627);
and U1506 (N_1506,In_4868,In_1038);
nor U1507 (N_1507,In_1191,In_2252);
nor U1508 (N_1508,In_4737,In_2319);
or U1509 (N_1509,In_4082,In_355);
nand U1510 (N_1510,In_969,In_2140);
nand U1511 (N_1511,In_3173,In_3423);
nor U1512 (N_1512,In_3855,In_4748);
xnor U1513 (N_1513,In_701,In_3903);
or U1514 (N_1514,In_2722,In_2309);
nor U1515 (N_1515,In_1241,In_1538);
or U1516 (N_1516,In_3051,In_1973);
or U1517 (N_1517,In_3771,In_3591);
and U1518 (N_1518,In_3238,In_3889);
and U1519 (N_1519,In_4976,In_4135);
nand U1520 (N_1520,In_1896,In_2893);
and U1521 (N_1521,In_2284,In_2445);
or U1522 (N_1522,In_4471,In_2170);
nor U1523 (N_1523,In_949,In_286);
or U1524 (N_1524,In_1977,In_2462);
nor U1525 (N_1525,In_3798,In_3502);
or U1526 (N_1526,In_3391,In_3588);
or U1527 (N_1527,In_4943,In_803);
and U1528 (N_1528,In_3629,In_460);
or U1529 (N_1529,In_641,In_4340);
or U1530 (N_1530,In_363,In_4728);
and U1531 (N_1531,In_1006,In_2059);
xnor U1532 (N_1532,In_1878,In_4673);
or U1533 (N_1533,In_4928,In_768);
and U1534 (N_1534,In_2543,In_3403);
and U1535 (N_1535,In_4551,In_2602);
and U1536 (N_1536,In_2286,In_309);
and U1537 (N_1537,In_3657,In_1664);
and U1538 (N_1538,In_3842,In_170);
and U1539 (N_1539,In_1425,In_1219);
nand U1540 (N_1540,In_1055,In_807);
nand U1541 (N_1541,In_3712,In_3369);
nand U1542 (N_1542,In_3174,In_3757);
and U1543 (N_1543,In_898,In_3050);
and U1544 (N_1544,In_3544,In_377);
or U1545 (N_1545,In_692,In_4510);
xnor U1546 (N_1546,In_312,In_2872);
nand U1547 (N_1547,In_4981,In_2484);
or U1548 (N_1548,In_634,In_210);
and U1549 (N_1549,In_1207,In_3144);
and U1550 (N_1550,In_1382,In_337);
nand U1551 (N_1551,In_4079,In_3526);
nor U1552 (N_1552,In_2982,In_889);
and U1553 (N_1553,In_4576,In_1253);
nand U1554 (N_1554,In_4727,In_4231);
nand U1555 (N_1555,In_4043,In_4187);
nand U1556 (N_1556,In_1394,In_1209);
nand U1557 (N_1557,In_2978,In_265);
nor U1558 (N_1558,In_4470,In_121);
nand U1559 (N_1559,In_3483,In_4047);
nor U1560 (N_1560,In_2085,In_3482);
nor U1561 (N_1561,In_441,In_1906);
nand U1562 (N_1562,In_1866,In_1421);
and U1563 (N_1563,In_3680,In_3162);
nor U1564 (N_1564,In_2051,In_299);
nand U1565 (N_1565,In_185,In_2327);
nor U1566 (N_1566,In_1494,In_2933);
nor U1567 (N_1567,In_2031,In_2188);
and U1568 (N_1568,In_421,In_1031);
nand U1569 (N_1569,In_1360,In_867);
nand U1570 (N_1570,In_3461,In_712);
nor U1571 (N_1571,In_1864,In_4466);
nand U1572 (N_1572,In_1869,In_2466);
and U1573 (N_1573,In_2096,In_463);
or U1574 (N_1574,In_4894,In_2621);
and U1575 (N_1575,In_4680,In_2825);
xor U1576 (N_1576,In_4528,In_1415);
nand U1577 (N_1577,In_174,In_737);
nand U1578 (N_1578,In_1337,In_1385);
nand U1579 (N_1579,In_4229,In_2482);
nand U1580 (N_1580,In_1534,In_3291);
nand U1581 (N_1581,In_447,In_3859);
nor U1582 (N_1582,In_1588,In_4418);
xnor U1583 (N_1583,In_3495,In_1604);
and U1584 (N_1584,In_99,In_1047);
xor U1585 (N_1585,In_3848,In_1999);
or U1586 (N_1586,In_3839,In_2389);
nand U1587 (N_1587,In_2848,In_1122);
nor U1588 (N_1588,In_4318,In_4630);
or U1589 (N_1589,In_1229,In_289);
nand U1590 (N_1590,In_3043,In_450);
and U1591 (N_1591,In_30,In_2615);
nand U1592 (N_1592,In_3201,In_3632);
xnor U1593 (N_1593,In_1984,In_3135);
or U1594 (N_1594,In_3504,In_440);
nand U1595 (N_1595,In_4644,In_3145);
nor U1596 (N_1596,In_2685,In_1744);
or U1597 (N_1597,In_3167,In_1685);
nand U1598 (N_1598,In_173,In_2798);
nand U1599 (N_1599,In_3835,In_4856);
and U1600 (N_1600,In_965,In_3873);
or U1601 (N_1601,In_4462,In_4698);
nand U1602 (N_1602,In_591,In_149);
or U1603 (N_1603,In_4365,In_3869);
or U1604 (N_1604,In_3880,In_1891);
and U1605 (N_1605,In_3121,In_1750);
nor U1606 (N_1606,In_1020,In_2819);
nor U1607 (N_1607,In_550,In_3505);
or U1608 (N_1608,In_3607,In_1553);
xor U1609 (N_1609,In_2735,In_1726);
nand U1610 (N_1610,In_672,In_4071);
nand U1611 (N_1611,In_3090,In_1401);
nor U1612 (N_1612,In_4064,In_1096);
nor U1613 (N_1613,In_4862,In_4697);
or U1614 (N_1614,In_155,In_794);
nor U1615 (N_1615,In_4371,In_3224);
nor U1616 (N_1616,In_1235,In_870);
or U1617 (N_1617,In_2886,In_2255);
or U1618 (N_1618,In_2159,In_2218);
xnor U1619 (N_1619,In_2607,In_2441);
and U1620 (N_1620,In_2524,In_3704);
or U1621 (N_1621,In_4148,In_4806);
xnor U1622 (N_1622,In_3450,In_2220);
nand U1623 (N_1623,In_3728,In_2719);
or U1624 (N_1624,In_514,In_3573);
nand U1625 (N_1625,In_2927,In_4208);
nor U1626 (N_1626,In_3727,In_2959);
or U1627 (N_1627,In_4969,In_4256);
nor U1628 (N_1628,In_2903,In_439);
nor U1629 (N_1629,In_3729,In_4434);
and U1630 (N_1630,In_2766,In_274);
nor U1631 (N_1631,In_4329,In_4373);
or U1632 (N_1632,In_152,In_2729);
nor U1633 (N_1633,In_654,In_3322);
xnor U1634 (N_1634,In_3865,In_2350);
nand U1635 (N_1635,In_2783,In_4458);
nor U1636 (N_1636,In_948,In_1474);
or U1637 (N_1637,In_261,In_2292);
and U1638 (N_1638,In_3943,In_1442);
and U1639 (N_1639,In_1294,In_2842);
xor U1640 (N_1640,In_4146,In_4151);
and U1641 (N_1641,In_2677,In_3056);
and U1642 (N_1642,In_4695,In_3191);
nand U1643 (N_1643,In_1206,In_2880);
nand U1644 (N_1644,In_4620,In_1146);
or U1645 (N_1645,In_3350,In_1703);
or U1646 (N_1646,In_2454,In_2234);
nor U1647 (N_1647,In_853,In_378);
nor U1648 (N_1648,In_910,In_762);
and U1649 (N_1649,In_3387,In_4136);
nand U1650 (N_1650,In_1339,In_1510);
and U1651 (N_1651,In_4718,In_370);
nor U1652 (N_1652,In_753,In_3281);
nand U1653 (N_1653,In_2022,In_4958);
nor U1654 (N_1654,In_1349,In_3296);
or U1655 (N_1655,In_760,In_3399);
or U1656 (N_1656,In_3733,In_3553);
nand U1657 (N_1657,In_3218,In_2426);
nor U1658 (N_1658,In_1136,In_1147);
or U1659 (N_1659,In_3828,In_2716);
nor U1660 (N_1660,In_3250,In_3794);
nand U1661 (N_1661,In_501,In_4668);
or U1662 (N_1662,In_971,In_4690);
xnor U1663 (N_1663,In_3517,In_1822);
nand U1664 (N_1664,In_1575,In_4733);
and U1665 (N_1665,In_1810,In_3297);
or U1666 (N_1666,In_1498,In_3877);
or U1667 (N_1667,In_2717,In_4150);
and U1668 (N_1668,In_50,In_2721);
and U1669 (N_1669,In_4400,In_4774);
or U1670 (N_1670,In_923,In_3217);
nand U1671 (N_1671,In_2837,In_1109);
or U1672 (N_1672,In_2632,In_2616);
or U1673 (N_1673,In_3989,In_3971);
and U1674 (N_1674,In_2908,In_1037);
xnor U1675 (N_1675,In_4432,In_3299);
and U1676 (N_1676,In_3030,In_1254);
nor U1677 (N_1677,In_84,In_1600);
nor U1678 (N_1678,In_2511,In_1844);
and U1679 (N_1679,In_832,In_2851);
or U1680 (N_1680,In_2763,In_456);
nand U1681 (N_1681,In_1315,In_4877);
or U1682 (N_1682,In_4834,In_3038);
nand U1683 (N_1683,In_2711,In_3011);
nand U1684 (N_1684,In_4598,In_1392);
or U1685 (N_1685,In_1044,In_3027);
and U1686 (N_1686,In_1257,In_583);
nor U1687 (N_1687,In_3122,In_2788);
nor U1688 (N_1688,In_2179,In_58);
nand U1689 (N_1689,In_1024,In_245);
nor U1690 (N_1690,In_4442,In_3799);
or U1691 (N_1691,In_3460,In_4480);
nor U1692 (N_1692,In_1644,In_4261);
xnor U1693 (N_1693,In_2104,In_4512);
nand U1694 (N_1694,In_651,In_2580);
nor U1695 (N_1695,In_2471,In_1861);
nand U1696 (N_1696,In_1586,In_2247);
nor U1697 (N_1697,In_1619,In_3175);
and U1698 (N_1698,In_3071,In_1505);
nor U1699 (N_1699,In_3954,In_4126);
xor U1700 (N_1700,In_2118,In_382);
nand U1701 (N_1701,In_4609,In_1194);
and U1702 (N_1702,In_3199,In_3021);
xor U1703 (N_1703,In_3274,In_1131);
xor U1704 (N_1704,In_4453,In_1738);
nor U1705 (N_1705,In_4407,In_1012);
nand U1706 (N_1706,In_2514,In_4605);
or U1707 (N_1707,In_3475,In_3474);
nor U1708 (N_1708,In_3561,In_1914);
nand U1709 (N_1709,In_4659,In_2642);
and U1710 (N_1710,In_4670,In_565);
or U1711 (N_1711,In_1141,In_1424);
or U1712 (N_1712,In_615,In_536);
nand U1713 (N_1713,In_220,In_2515);
or U1714 (N_1714,In_3951,In_246);
or U1715 (N_1715,In_307,In_4128);
and U1716 (N_1716,In_3961,In_179);
and U1717 (N_1717,In_2217,In_4699);
xor U1718 (N_1718,In_761,In_1419);
or U1719 (N_1719,In_318,In_1098);
or U1720 (N_1720,In_133,In_3990);
or U1721 (N_1721,In_3215,In_495);
nor U1722 (N_1722,In_582,In_113);
and U1723 (N_1723,In_4258,In_4831);
or U1724 (N_1724,In_774,In_1773);
nor U1725 (N_1725,In_479,In_1589);
nor U1726 (N_1726,In_3363,In_3538);
or U1727 (N_1727,In_4445,In_1413);
nor U1728 (N_1728,In_919,In_4077);
nor U1729 (N_1729,In_1634,In_917);
nor U1730 (N_1730,In_4893,In_1788);
or U1731 (N_1731,In_2534,In_3479);
or U1732 (N_1732,In_3820,In_2066);
nand U1733 (N_1733,In_2710,In_452);
or U1734 (N_1734,In_83,In_2555);
nor U1735 (N_1735,In_3331,In_1492);
nor U1736 (N_1736,In_201,In_4902);
and U1737 (N_1737,In_3115,In_3850);
and U1738 (N_1738,In_1192,In_1368);
and U1739 (N_1739,In_1407,In_3532);
or U1740 (N_1740,In_4573,In_4107);
nand U1741 (N_1741,In_1035,In_1777);
or U1742 (N_1742,In_967,In_1317);
and U1743 (N_1743,In_3101,In_241);
nor U1744 (N_1744,In_313,In_978);
nor U1745 (N_1745,In_407,In_3205);
and U1746 (N_1746,In_975,In_1622);
nor U1747 (N_1747,In_2726,In_59);
and U1748 (N_1748,In_4556,In_2700);
nor U1749 (N_1749,In_277,In_2300);
or U1750 (N_1750,In_2435,In_4472);
nor U1751 (N_1751,In_4850,In_3653);
or U1752 (N_1752,In_1435,In_4881);
nor U1753 (N_1753,In_4405,In_618);
xor U1754 (N_1754,In_3061,In_3129);
and U1755 (N_1755,In_4374,In_3967);
and U1756 (N_1756,In_3689,In_4548);
or U1757 (N_1757,In_1748,In_2795);
and U1758 (N_1758,In_1601,In_673);
nor U1759 (N_1759,In_4632,In_1718);
and U1760 (N_1760,In_3077,In_4952);
or U1761 (N_1761,In_3827,In_2393);
nor U1762 (N_1762,In_2100,In_1674);
nand U1763 (N_1763,In_4368,In_1599);
xnor U1764 (N_1764,In_1375,In_4770);
nand U1765 (N_1765,In_2947,In_4339);
nor U1766 (N_1766,In_678,In_4631);
nand U1767 (N_1767,In_3138,In_4612);
or U1768 (N_1768,In_2583,In_3395);
or U1769 (N_1769,In_1117,In_1922);
or U1770 (N_1770,In_4059,In_3339);
or U1771 (N_1771,In_1432,In_1959);
and U1772 (N_1772,In_3995,In_1556);
and U1773 (N_1773,In_2201,In_4563);
and U1774 (N_1774,In_3853,In_3062);
and U1775 (N_1775,In_4791,In_857);
and U1776 (N_1776,In_2736,In_1429);
nor U1777 (N_1777,In_2410,In_3906);
nand U1778 (N_1778,In_735,In_1433);
nand U1779 (N_1779,In_3589,In_1439);
xor U1780 (N_1780,In_2404,In_4183);
nor U1781 (N_1781,In_1763,In_4056);
or U1782 (N_1782,In_3631,In_1478);
nand U1783 (N_1783,In_4133,In_232);
nor U1784 (N_1784,In_62,In_4404);
nand U1785 (N_1785,In_2197,In_935);
and U1786 (N_1786,In_4000,In_4672);
or U1787 (N_1787,In_4991,In_1080);
nand U1788 (N_1788,In_4601,In_27);
nor U1789 (N_1789,In_4994,In_2574);
nor U1790 (N_1790,In_2103,In_2680);
nand U1791 (N_1791,In_2698,In_1629);
nor U1792 (N_1792,In_4794,In_2874);
and U1793 (N_1793,In_2945,In_480);
and U1794 (N_1794,In_4435,In_425);
nand U1795 (N_1795,In_1389,In_3048);
nand U1796 (N_1796,In_438,In_1371);
nor U1797 (N_1797,In_4723,In_3086);
nor U1798 (N_1798,In_3964,In_3522);
or U1799 (N_1799,In_2758,In_389);
xnor U1800 (N_1800,In_3763,In_2082);
and U1801 (N_1801,In_627,In_4956);
and U1802 (N_1802,In_1766,In_3619);
and U1803 (N_1803,In_2775,In_3373);
nor U1804 (N_1804,In_68,In_3192);
and U1805 (N_1805,In_4176,In_4454);
nor U1806 (N_1806,In_2370,In_129);
nand U1807 (N_1807,In_1248,In_861);
and U1808 (N_1808,In_4112,In_4459);
nand U1809 (N_1809,In_4194,In_2130);
nand U1810 (N_1810,In_448,In_3645);
or U1811 (N_1811,In_4436,In_2892);
or U1812 (N_1812,In_3246,In_4005);
xor U1813 (N_1813,In_228,In_2321);
xnor U1814 (N_1814,In_3621,In_323);
nand U1815 (N_1815,In_1173,In_3832);
or U1816 (N_1816,In_3972,In_2957);
and U1817 (N_1817,In_2207,In_2950);
and U1818 (N_1818,In_1119,In_4050);
and U1819 (N_1819,In_3209,In_2509);
nand U1820 (N_1820,In_2573,In_4709);
and U1821 (N_1821,In_2654,In_3601);
and U1822 (N_1822,In_4293,In_4455);
or U1823 (N_1823,In_1992,In_3909);
nor U1824 (N_1824,In_3786,In_2342);
and U1825 (N_1825,In_1867,In_2638);
nand U1826 (N_1826,In_3723,In_3008);
or U1827 (N_1827,In_553,In_1342);
nand U1828 (N_1828,In_551,In_945);
and U1829 (N_1829,In_4249,In_890);
xnor U1830 (N_1830,In_3470,In_4011);
nand U1831 (N_1831,In_3635,In_208);
xor U1832 (N_1832,In_2497,In_4236);
nor U1833 (N_1833,In_4665,In_2266);
nor U1834 (N_1834,In_4682,In_1570);
nor U1835 (N_1835,In_3114,In_2979);
nand U1836 (N_1836,In_2316,In_1762);
nand U1837 (N_1837,In_4129,In_2142);
nand U1838 (N_1838,In_614,In_3160);
or U1839 (N_1839,In_4771,In_996);
nand U1840 (N_1840,In_2816,In_3348);
nor U1841 (N_1841,In_2418,In_9);
and U1842 (N_1842,In_4558,In_2940);
or U1843 (N_1843,In_711,In_3520);
xnor U1844 (N_1844,In_4925,In_199);
and U1845 (N_1845,In_3670,In_4205);
or U1846 (N_1846,In_914,In_2067);
xor U1847 (N_1847,In_72,In_3977);
nor U1848 (N_1848,In_843,In_2241);
nand U1849 (N_1849,In_2343,In_612);
or U1850 (N_1850,In_1469,In_327);
or U1851 (N_1851,In_37,In_1395);
nor U1852 (N_1852,In_4832,In_492);
or U1853 (N_1853,In_3298,In_960);
xor U1854 (N_1854,In_3894,In_510);
nand U1855 (N_1855,In_1224,In_3437);
xor U1856 (N_1856,In_2154,In_3884);
nor U1857 (N_1857,In_2447,In_25);
nand U1858 (N_1858,In_4826,In_2310);
nor U1859 (N_1859,In_3603,In_709);
nand U1860 (N_1860,In_3368,In_1464);
and U1861 (N_1861,In_2533,In_4966);
or U1862 (N_1862,In_993,In_3072);
nor U1863 (N_1863,In_2742,In_3431);
xnor U1864 (N_1864,In_2918,In_3721);
nand U1865 (N_1865,In_3329,In_3149);
xor U1866 (N_1866,In_1417,In_4423);
or U1867 (N_1867,In_3150,In_3075);
nor U1868 (N_1868,In_3151,In_4603);
and U1869 (N_1869,In_3172,In_4742);
nand U1870 (N_1870,In_3018,In_4661);
nand U1871 (N_1871,In_4560,In_366);
nor U1872 (N_1872,In_1532,In_8);
nor U1873 (N_1873,In_316,In_4255);
and U1874 (N_1874,In_814,In_384);
nor U1875 (N_1875,In_291,In_3398);
nor U1876 (N_1876,In_2050,In_619);
xor U1877 (N_1877,In_1145,In_4233);
and U1878 (N_1878,In_1120,In_1895);
nand U1879 (N_1879,In_305,In_3861);
nor U1880 (N_1880,In_3613,In_2557);
or U1881 (N_1881,In_631,In_2980);
and U1882 (N_1882,In_2353,In_269);
and U1883 (N_1883,In_4999,In_3247);
or U1884 (N_1884,In_4565,In_3236);
nor U1885 (N_1885,In_1269,In_2999);
and U1886 (N_1886,In_4297,In_937);
and U1887 (N_1887,In_4613,In_3233);
and U1888 (N_1888,In_4557,In_2620);
and U1889 (N_1889,In_2993,In_984);
nand U1890 (N_1890,In_4313,In_1993);
nand U1891 (N_1891,In_1964,In_4685);
or U1892 (N_1892,In_4164,In_4358);
nand U1893 (N_1893,In_3791,In_947);
nor U1894 (N_1894,In_3640,In_621);
and U1895 (N_1895,In_3006,In_2429);
or U1896 (N_1896,In_1106,In_2588);
and U1897 (N_1897,In_4114,In_3731);
nand U1898 (N_1898,In_4220,In_3123);
nor U1899 (N_1899,In_388,In_3111);
nand U1900 (N_1900,In_4932,In_1971);
or U1901 (N_1901,In_4078,In_1238);
or U1902 (N_1902,In_2095,In_1939);
nand U1903 (N_1903,In_4192,In_2739);
xor U1904 (N_1904,In_3600,In_749);
or U1905 (N_1905,In_1548,In_3222);
or U1906 (N_1906,In_4253,In_4002);
xor U1907 (N_1907,In_1536,In_573);
nand U1908 (N_1908,In_1052,In_1090);
or U1909 (N_1909,In_2747,In_2265);
nand U1910 (N_1910,In_2641,In_4489);
or U1911 (N_1911,In_1908,In_193);
nor U1912 (N_1912,In_2791,In_1695);
or U1913 (N_1913,In_4977,In_424);
and U1914 (N_1914,In_78,In_2666);
xnor U1915 (N_1915,In_547,In_4163);
xor U1916 (N_1916,In_755,In_16);
nor U1917 (N_1917,In_160,In_3026);
nor U1918 (N_1918,In_2293,In_656);
nand U1919 (N_1919,In_3968,In_3385);
or U1920 (N_1920,In_3506,In_594);
xor U1921 (N_1921,In_4006,In_796);
nand U1922 (N_1922,In_1976,In_3412);
nand U1923 (N_1923,In_1406,In_3926);
or U1924 (N_1924,In_4626,In_3406);
and U1925 (N_1925,In_3577,In_4724);
and U1926 (N_1926,In_1279,In_1874);
or U1927 (N_1927,In_2004,In_3136);
or U1928 (N_1928,In_1545,In_2627);
nor U1929 (N_1929,In_1450,In_2183);
or U1930 (N_1930,In_3308,In_1483);
or U1931 (N_1931,In_2658,In_3000);
and U1932 (N_1932,In_1981,In_4196);
nor U1933 (N_1933,In_4735,In_555);
or U1934 (N_1934,In_2365,In_4710);
and U1935 (N_1935,In_1997,In_2898);
nor U1936 (N_1936,In_3694,In_1960);
and U1937 (N_1937,In_4713,In_3780);
nor U1938 (N_1938,In_1711,In_213);
nor U1939 (N_1939,In_45,In_1590);
and U1940 (N_1940,In_2548,In_1343);
nor U1941 (N_1941,In_2840,In_2712);
or U1942 (N_1942,In_423,In_1245);
nand U1943 (N_1943,In_1670,In_3234);
nand U1944 (N_1944,In_3920,In_636);
and U1945 (N_1945,In_883,In_1140);
and U1946 (N_1946,In_4789,In_1612);
nand U1947 (N_1947,In_2730,In_1658);
nor U1948 (N_1948,In_575,In_3910);
and U1949 (N_1949,In_1963,In_2790);
or U1950 (N_1950,In_4623,In_3288);
nor U1951 (N_1951,In_1817,In_3991);
nor U1952 (N_1952,In_2864,In_622);
and U1953 (N_1953,In_1935,In_3988);
nor U1954 (N_1954,In_3684,In_4178);
nand U1955 (N_1955,In_2029,In_2905);
nor U1956 (N_1956,In_950,In_1016);
or U1957 (N_1957,In_475,In_484);
and U1958 (N_1958,In_2409,In_664);
and U1959 (N_1959,In_1328,In_963);
and U1960 (N_1960,In_390,In_1202);
and U1961 (N_1961,In_1813,In_4948);
nor U1962 (N_1962,In_4189,In_2228);
and U1963 (N_1963,In_1857,In_1373);
nor U1964 (N_1964,In_3333,In_4615);
nor U1965 (N_1965,In_4746,In_2977);
or U1966 (N_1966,In_608,In_884);
xnor U1967 (N_1967,In_1453,In_4230);
and U1968 (N_1968,In_4304,In_4694);
nor U1969 (N_1969,In_2896,In_183);
nand U1970 (N_1970,In_2181,In_3439);
nor U1971 (N_1971,In_2699,In_4569);
or U1972 (N_1972,In_903,In_3263);
and U1973 (N_1973,In_1222,In_3720);
or U1974 (N_1974,In_4276,In_1559);
or U1975 (N_1975,In_2366,In_2325);
or U1976 (N_1976,In_1904,In_442);
and U1977 (N_1977,In_4175,In_1292);
nand U1978 (N_1978,In_449,In_685);
or U1979 (N_1979,In_3193,In_96);
or U1980 (N_1980,In_4978,In_1572);
xor U1981 (N_1981,In_2512,In_3662);
and U1982 (N_1982,In_2476,In_4292);
xor U1983 (N_1983,In_3055,In_343);
nand U1984 (N_1984,In_4211,In_3227);
xor U1985 (N_1985,In_825,In_750);
nor U1986 (N_1986,In_4101,In_235);
nand U1987 (N_1987,In_2024,In_1129);
and U1988 (N_1988,In_1015,In_158);
nor U1989 (N_1989,In_1462,In_1163);
or U1990 (N_1990,In_944,In_1354);
nand U1991 (N_1991,In_1578,In_1595);
or U1992 (N_1992,In_3428,In_1001);
or U1993 (N_1993,In_3380,In_4497);
nor U1994 (N_1994,In_1549,In_4279);
nand U1995 (N_1995,In_1523,In_955);
nand U1996 (N_1996,In_2242,In_710);
nor U1997 (N_1997,In_1088,In_2860);
nand U1998 (N_1998,In_1520,In_1760);
or U1999 (N_1999,In_1966,In_278);
nand U2000 (N_2000,In_1003,In_1086);
nor U2001 (N_2001,In_4355,In_4750);
nor U2002 (N_2002,In_11,In_584);
and U2003 (N_2003,In_4855,In_1431);
or U2004 (N_2004,In_4295,In_863);
xnor U2005 (N_2005,In_602,In_4228);
xor U2006 (N_2006,In_3830,In_4707);
nor U2007 (N_2007,In_852,In_2914);
or U2008 (N_2008,In_2901,In_2273);
nor U2009 (N_2009,In_2311,In_3259);
or U2010 (N_2010,In_4033,In_308);
or U2011 (N_2011,In_4155,In_2975);
and U2012 (N_2012,In_1940,In_2834);
nand U2013 (N_2013,In_4390,In_2326);
or U2014 (N_2014,In_2728,In_822);
nor U2015 (N_2015,In_1516,In_3305);
and U2016 (N_2016,In_303,In_224);
and U2017 (N_2017,In_568,In_593);
xor U2018 (N_2018,In_1887,In_3367);
nand U2019 (N_2019,In_2521,In_4168);
nor U2020 (N_2020,In_2505,In_2844);
or U2021 (N_2021,In_4464,In_167);
or U2022 (N_2022,In_1755,In_4536);
nand U2023 (N_2023,In_2352,In_1729);
and U2024 (N_2024,In_585,In_2922);
or U2025 (N_2025,In_2911,In_2438);
or U2026 (N_2026,In_1178,In_3525);
and U2027 (N_2027,In_2818,In_2101);
and U2028 (N_2028,In_1902,In_542);
nor U2029 (N_2029,In_4519,In_4553);
xor U2030 (N_2030,In_4210,In_3772);
and U2031 (N_2031,In_1426,In_3922);
nor U2032 (N_2032,In_3710,In_704);
and U2033 (N_2033,In_3451,In_115);
nor U2034 (N_2034,In_1293,In_1288);
nand U2035 (N_2035,In_1348,In_2399);
nand U2036 (N_2036,In_1064,In_1303);
nand U2037 (N_2037,In_4909,In_1286);
xnor U2038 (N_2038,In_4016,In_4134);
nor U2039 (N_2039,In_1608,In_1886);
nor U2040 (N_2040,In_3983,In_2198);
and U2041 (N_2041,In_2572,In_4865);
and U2042 (N_2042,In_3927,In_3337);
nor U2043 (N_2043,In_2626,In_3081);
nor U2044 (N_2044,In_2436,In_2894);
or U2045 (N_2045,In_2,In_3351);
and U2046 (N_2046,In_3453,In_922);
nor U2047 (N_2047,In_4099,In_468);
or U2048 (N_2048,In_2387,In_3080);
xnor U2049 (N_2049,In_3539,In_203);
nor U2050 (N_2050,In_1679,In_4429);
nand U2051 (N_2051,In_4363,In_137);
nand U2052 (N_2052,In_4203,In_2357);
nor U2053 (N_2053,In_4217,In_3556);
or U2054 (N_2054,In_81,In_3758);
or U2055 (N_2055,In_1909,In_1499);
or U2056 (N_2056,In_4376,In_3976);
nand U2057 (N_2057,In_4287,In_2485);
xor U2058 (N_2058,In_3389,In_1393);
and U2059 (N_2059,In_4985,In_1765);
nor U2060 (N_2060,In_640,In_206);
nand U2061 (N_2061,In_2367,In_1944);
nor U2062 (N_2062,In_3743,In_3748);
and U2063 (N_2063,In_108,In_3376);
and U2064 (N_2064,In_1842,In_4721);
xnor U2065 (N_2065,In_4100,In_4226);
nor U2066 (N_2066,In_2016,In_2115);
nor U2067 (N_2067,In_4448,In_2386);
or U2068 (N_2068,In_2450,In_1667);
and U2069 (N_2069,In_1125,In_2257);
nand U2070 (N_2070,In_3714,In_2143);
nand U2071 (N_2071,In_4825,In_3498);
and U2072 (N_2072,In_2264,In_159);
nor U2073 (N_2073,In_4444,In_4333);
nand U2074 (N_2074,In_3905,In_2187);
nand U2075 (N_2075,In_1605,In_2884);
xor U2076 (N_2076,In_4478,In_3690);
nand U2077 (N_2077,In_4580,In_2603);
and U2078 (N_2078,In_1965,In_1452);
and U2079 (N_2079,In_862,In_1557);
and U2080 (N_2080,In_3286,In_2942);
nand U2081 (N_2081,In_1472,In_3887);
nand U2082 (N_2082,In_2275,In_1153);
and U2083 (N_2083,In_698,In_2477);
nor U2084 (N_2084,In_2391,In_3626);
or U2085 (N_2085,In_3179,In_4777);
nand U2086 (N_2086,In_1803,In_1808);
or U2087 (N_2087,In_244,In_4441);
or U2088 (N_2088,In_577,In_3521);
nor U2089 (N_2089,In_3097,In_4447);
or U2090 (N_2090,In_394,In_2956);
and U2091 (N_2091,In_3047,In_2688);
and U2092 (N_2092,In_3592,In_1085);
or U2093 (N_2093,In_2459,In_415);
or U2094 (N_2094,In_2734,In_4583);
and U2095 (N_2095,In_1108,In_644);
nor U2096 (N_2096,In_2655,In_2149);
nor U2097 (N_2097,In_3435,In_3650);
nand U2098 (N_2098,In_4764,In_293);
nor U2099 (N_2099,In_3980,In_1099);
or U2100 (N_2100,In_209,In_2407);
nor U2101 (N_2101,In_3443,In_4036);
xor U2102 (N_2102,In_1078,In_3063);
nor U2103 (N_2103,In_4224,In_3917);
or U2104 (N_2104,In_4761,In_3959);
and U2105 (N_2105,In_3139,In_2379);
nand U2106 (N_2106,In_1905,In_3929);
nor U2107 (N_2107,In_2374,In_1917);
xnor U2108 (N_2108,In_2138,In_4451);
xnor U2109 (N_2109,In_2488,In_3301);
nor U2110 (N_2110,In_2749,In_1074);
nor U2111 (N_2111,In_3084,In_941);
or U2112 (N_2112,In_345,In_161);
and U2113 (N_2113,In_24,In_3963);
and U2114 (N_2114,In_3931,In_938);
and U2115 (N_2115,In_4537,In_3536);
nand U2116 (N_2116,In_2261,In_4917);
nor U2117 (N_2117,In_3656,In_748);
or U2118 (N_2118,In_1698,In_1825);
and U2119 (N_2119,In_2611,In_3774);
nor U2120 (N_2120,In_2820,In_2175);
nand U2121 (N_2121,In_3551,In_2054);
or U2122 (N_2122,In_3040,In_284);
nand U2123 (N_2123,In_3860,In_874);
nor U2124 (N_2124,In_2944,In_32);
nor U2125 (N_2125,In_2962,In_3765);
nor U2126 (N_2126,In_349,In_1816);
or U2127 (N_2127,In_4692,In_1799);
nor U2128 (N_2128,In_2030,In_769);
nand U2129 (N_2129,In_4105,In_2553);
and U2130 (N_2130,In_1198,In_1683);
nand U2131 (N_2131,In_4428,In_1863);
nor U2132 (N_2132,In_1642,In_850);
nor U2133 (N_2133,In_1528,In_1324);
nor U2134 (N_2134,In_3568,In_357);
or U2135 (N_2135,In_3309,In_2274);
nor U2136 (N_2136,In_723,In_2250);
nand U2137 (N_2137,In_3937,In_298);
nand U2138 (N_2138,In_225,In_1189);
nand U2139 (N_2139,In_195,In_1723);
and U2140 (N_2140,In_134,In_1255);
xor U2141 (N_2141,In_4315,In_20);
nand U2142 (N_2142,In_4835,In_1611);
nor U2143 (N_2143,In_143,In_2268);
nand U2144 (N_2144,In_333,In_2966);
or U2145 (N_2145,In_3933,In_2856);
and U2146 (N_2146,In_409,In_1133);
and U2147 (N_2147,In_1237,In_1730);
nand U2148 (N_2148,In_3784,In_3776);
or U2149 (N_2149,In_3155,In_4951);
nand U2150 (N_2150,In_1617,In_2965);
nor U2151 (N_2151,In_4934,In_1592);
nand U2152 (N_2152,In_2813,In_26);
and U2153 (N_2153,In_912,In_1331);
nand U2154 (N_2154,In_1262,In_2839);
or U2155 (N_2155,In_1898,In_1782);
and U2156 (N_2156,In_2248,In_2190);
and U2157 (N_2157,In_3449,In_4968);
nand U2158 (N_2158,In_1113,In_1818);
nand U2159 (N_2159,In_1980,In_1216);
nand U2160 (N_2160,In_1541,In_2420);
nor U2161 (N_2161,In_4530,In_3017);
nand U2162 (N_2162,In_2223,In_2186);
nor U2163 (N_2163,In_2960,In_1655);
or U2164 (N_2164,In_931,In_2604);
nor U2165 (N_2165,In_3069,In_676);
nor U2166 (N_2166,In_4331,In_2510);
xnor U2167 (N_2167,In_1332,In_3196);
xor U2168 (N_2168,In_3962,In_2647);
nor U2169 (N_2169,In_2810,In_2057);
nor U2170 (N_2170,In_4912,In_3676);
and U2171 (N_2171,In_4922,In_4088);
nand U2172 (N_2172,In_1745,In_2465);
xnor U2173 (N_2173,In_1379,In_650);
or U2174 (N_2174,In_4362,In_4762);
nor U2175 (N_2175,In_3745,In_4141);
nor U2176 (N_2176,In_2684,In_1830);
or U2177 (N_2177,In_2609,In_3262);
nor U2178 (N_2178,In_4971,In_3636);
nor U2179 (N_2179,In_2479,In_1276);
xnor U2180 (N_2180,In_642,In_2213);
nand U2181 (N_2181,In_4326,In_2541);
nor U2182 (N_2182,In_3023,In_2709);
nand U2183 (N_2183,In_2876,In_1948);
xor U2184 (N_2184,In_3831,In_1806);
nand U2185 (N_2185,In_3724,In_3750);
and U2186 (N_2186,In_1815,In_176);
xnor U2187 (N_2187,In_4942,In_4887);
and U2188 (N_2188,In_4606,In_4091);
or U2189 (N_2189,In_1988,In_1506);
nor U2190 (N_2190,In_3016,In_4527);
and U2191 (N_2191,In_1954,In_4062);
and U2192 (N_2192,In_4840,In_745);
or U2193 (N_2193,In_2347,In_171);
or U2194 (N_2194,In_2612,In_3940);
nor U2195 (N_2195,In_4347,In_3311);
xnor U2196 (N_2196,In_4992,In_2773);
or U2197 (N_2197,In_1313,In_4936);
nor U2198 (N_2198,In_4819,In_1951);
xor U2199 (N_2199,In_601,In_3419);
nand U2200 (N_2200,In_3109,In_1282);
and U2201 (N_2201,In_3609,In_486);
nand U2202 (N_2202,In_1372,In_951);
nand U2203 (N_2203,In_3065,In_2551);
and U2204 (N_2204,In_679,In_3863);
xor U2205 (N_2205,In_624,In_4759);
or U2206 (N_2206,In_1979,In_4384);
or U2207 (N_2207,In_1444,In_2808);
nor U2208 (N_2208,In_3383,In_4861);
nor U2209 (N_2209,In_4987,In_2879);
nor U2210 (N_2210,In_2012,In_2954);
nor U2211 (N_2211,In_2929,In_4540);
and U2212 (N_2212,In_4525,In_1457);
xnor U2213 (N_2213,In_1841,In_2122);
nor U2214 (N_2214,In_2397,In_954);
or U2215 (N_2215,In_2789,In_4757);
nand U2216 (N_2216,In_2689,In_804);
nand U2217 (N_2217,In_530,In_4799);
nor U2218 (N_2218,In_1105,In_2331);
or U2219 (N_2219,In_4628,In_2656);
or U2220 (N_2220,In_4487,In_1794);
nand U2221 (N_2221,In_2784,In_2702);
and U2222 (N_2222,In_1341,In_364);
xnor U2223 (N_2223,In_2185,In_3170);
or U2224 (N_2224,In_2855,In_1187);
or U2225 (N_2225,In_49,In_953);
or U2226 (N_2226,In_4395,In_4582);
nor U2227 (N_2227,In_564,In_2985);
nor U2228 (N_2228,In_79,In_1188);
or U2229 (N_2229,In_4646,In_2614);
and U2230 (N_2230,In_3807,In_983);
or U2231 (N_2231,In_353,In_2414);
nand U2232 (N_2232,In_942,In_211);
or U2233 (N_2233,In_412,In_973);
and U2234 (N_2234,In_4879,In_2765);
or U2235 (N_2235,In_3944,In_2256);
nor U2236 (N_2236,In_1832,In_4809);
and U2237 (N_2237,In_989,In_3911);
nand U2238 (N_2238,In_3984,In_1130);
xnor U2239 (N_2239,In_3735,In_1796);
nand U2240 (N_2240,In_359,In_2660);
nor U2241 (N_2241,In_1170,In_1319);
nor U2242 (N_2242,In_2345,In_2042);
and U2243 (N_2243,In_2344,In_374);
and U2244 (N_2244,In_1654,In_406);
or U2245 (N_2245,In_140,In_933);
nand U2246 (N_2246,In_4227,In_4093);
and U2247 (N_2247,In_3402,In_4658);
or U2248 (N_2248,In_3104,In_2967);
nand U2249 (N_2249,In_3652,In_2152);
nand U2250 (N_2250,In_4775,In_2455);
and U2251 (N_2251,In_119,In_4808);
nor U2252 (N_2252,In_2034,In_1645);
xnor U2253 (N_2253,In_2496,In_2559);
or U2254 (N_2254,In_613,In_1598);
nor U2255 (N_2255,In_3671,In_1580);
nor U2256 (N_2256,In_85,In_3692);
and U2257 (N_2257,In_2857,In_13);
xnor U2258 (N_2258,In_3594,In_818);
nor U2259 (N_2259,In_1344,In_2411);
or U2260 (N_2260,In_2992,In_1876);
nand U2261 (N_2261,In_3585,In_1097);
nand U2262 (N_2262,In_603,In_927);
nand U2263 (N_2263,In_2549,In_2650);
nor U2264 (N_2264,In_1383,In_2861);
nor U2265 (N_2265,In_1791,In_4031);
or U2266 (N_2266,In_3230,In_250);
nor U2267 (N_2267,In_338,In_4503);
nor U2268 (N_2268,In_3057,In_2601);
or U2269 (N_2269,In_3251,In_2613);
nor U2270 (N_2270,In_2368,In_4882);
nor U2271 (N_2271,In_2428,In_1214);
nand U2272 (N_2272,In_1618,In_1124);
or U2273 (N_2273,In_3846,In_1567);
xor U2274 (N_2274,In_1704,In_2651);
nand U2275 (N_2275,In_3658,In_1010);
and U2276 (N_2276,In_3685,In_2007);
or U2277 (N_2277,In_4081,In_901);
or U2278 (N_2278,In_830,In_2949);
xor U2279 (N_2279,In_404,In_2167);
and U2280 (N_2280,In_1847,In_3583);
nand U2281 (N_2281,In_3001,In_1983);
nand U2282 (N_2282,In_371,In_3336);
nor U2283 (N_2283,In_335,In_4566);
and U2284 (N_2284,In_3277,In_1798);
or U2285 (N_2285,In_2371,In_1636);
or U2286 (N_2286,In_4945,In_2708);
or U2287 (N_2287,In_3973,In_3777);
and U2288 (N_2288,In_1638,In_500);
and U2289 (N_2289,In_2434,In_1040);
nor U2290 (N_2290,In_810,In_2424);
xor U2291 (N_2291,In_2670,In_1648);
nor U2292 (N_2292,In_546,In_580);
nand U2293 (N_2293,In_1967,In_4547);
and U2294 (N_2294,In_3507,In_3261);
xnor U2295 (N_2295,In_1275,In_1247);
nor U2296 (N_2296,In_3186,In_3946);
nor U2297 (N_2297,In_728,In_3698);
and U2298 (N_2298,In_519,In_4025);
or U2299 (N_2299,In_2421,In_2468);
and U2300 (N_2300,In_2222,In_1273);
nand U2301 (N_2301,In_4572,In_4818);
xor U2302 (N_2302,In_3197,In_1509);
nor U2303 (N_2303,In_660,In_3100);
xnor U2304 (N_2304,In_4758,In_2269);
nor U2305 (N_2305,In_3695,In_3736);
or U2306 (N_2306,In_786,In_1551);
and U2307 (N_2307,In_3740,In_2852);
and U2308 (N_2308,In_856,In_2160);
and U2309 (N_2309,In_1678,In_3089);
or U2310 (N_2310,In_3312,In_471);
or U2311 (N_2311,In_827,In_4854);
or U2312 (N_2312,In_3152,In_2500);
nor U2313 (N_2313,In_34,In_1290);
and U2314 (N_2314,In_4990,In_4947);
or U2315 (N_2315,In_4103,In_1606);
nor U2316 (N_2316,In_1884,In_1227);
nor U2317 (N_2317,In_2800,In_4772);
and U2318 (N_2318,In_4049,In_4950);
nor U2319 (N_2319,In_730,In_1361);
nor U2320 (N_2320,In_605,In_2116);
nor U2321 (N_2321,In_1691,In_4274);
and U2322 (N_2322,In_4704,In_652);
and U2323 (N_2323,In_1620,In_2074);
nor U2324 (N_2324,In_3804,In_1199);
xnor U2325 (N_2325,In_3528,In_3243);
or U2326 (N_2326,In_4159,In_626);
and U2327 (N_2327,In_1381,In_1161);
and U2328 (N_2328,In_3226,In_2988);
nor U2329 (N_2329,In_3686,In_2363);
and U2330 (N_2330,In_4022,In_4087);
and U2331 (N_2331,In_1547,In_125);
nand U2332 (N_2332,In_3925,In_3093);
and U2333 (N_2333,In_2648,In_3407);
or U2334 (N_2334,In_1482,In_1359);
or U2335 (N_2335,In_3513,In_4738);
or U2336 (N_2336,In_282,In_1063);
or U2337 (N_2337,In_1659,In_3557);
xnor U2338 (N_2338,In_1687,In_4741);
and U2339 (N_2339,In_3366,In_2127);
or U2340 (N_2340,In_2561,In_4590);
or U2341 (N_2341,In_647,In_3165);
and U2342 (N_2342,In_2333,In_4111);
nor U2343 (N_2343,In_572,In_1391);
or U2344 (N_2344,In_518,In_4849);
and U2345 (N_2345,In_368,In_4663);
and U2346 (N_2346,In_1093,In_1677);
and U2347 (N_2347,In_1351,In_1316);
or U2348 (N_2348,In_791,In_2845);
and U2349 (N_2349,In_1837,In_718);
nand U2350 (N_2350,In_3787,In_3184);
nor U2351 (N_2351,In_3574,In_3938);
or U2352 (N_2352,In_3732,In_2172);
nor U2353 (N_2353,In_1565,In_3580);
xnor U2354 (N_2354,In_215,In_4421);
nor U2355 (N_2355,In_1746,In_849);
nor U2356 (N_2356,In_1946,In_4953);
and U2357 (N_2357,In_693,In_3501);
and U2358 (N_2358,In_740,In_661);
xnor U2359 (N_2359,In_2177,In_4234);
and U2360 (N_2360,In_1103,In_3523);
nand U2361 (N_2361,In_1779,In_153);
and U2362 (N_2362,In_4815,In_663);
nor U2363 (N_2363,In_1778,In_2545);
or U2364 (N_2364,In_4802,In_3099);
nor U2365 (N_2365,In_205,In_1918);
or U2366 (N_2366,In_1919,In_1236);
nand U2367 (N_2367,In_3415,In_3214);
or U2368 (N_2368,In_3189,In_2518);
or U2369 (N_2369,In_1231,In_3838);
nand U2370 (N_2370,In_4706,In_4204);
and U2371 (N_2371,In_1496,In_4015);
xor U2372 (N_2372,In_1968,In_835);
nor U2373 (N_2373,In_1304,In_4139);
xor U2374 (N_2374,In_4841,In_1101);
or U2375 (N_2375,In_1742,In_1116);
and U2376 (N_2376,In_142,In_570);
or U2377 (N_2377,In_3448,In_4517);
nor U2378 (N_2378,In_527,In_2178);
nor U2379 (N_2379,In_1913,In_3755);
or U2380 (N_2380,In_4921,In_2759);
xor U2381 (N_2381,In_1356,In_2375);
nor U2382 (N_2382,In_2469,In_127);
xor U2383 (N_2383,In_4891,In_2403);
nand U2384 (N_2384,In_2111,In_2182);
and U2385 (N_2385,In_3811,In_4014);
and U2386 (N_2386,In_4667,In_982);
nand U2387 (N_2387,In_4023,In_3630);
and U2388 (N_2388,In_3699,In_1732);
and U2389 (N_2389,In_2093,In_4984);
nor U2390 (N_2390,In_1232,In_52);
and U2391 (N_2391,In_4041,In_1060);
and U2392 (N_2392,In_4529,In_3421);
or U2393 (N_2393,In_2887,In_2361);
or U2394 (N_2394,In_1879,In_3708);
nor U2395 (N_2395,In_657,In_4821);
and U2396 (N_2396,In_4523,In_2871);
and U2397 (N_2397,In_1388,In_3957);
nand U2398 (N_2398,In_3540,In_4814);
xor U2399 (N_2399,In_4048,In_238);
and U2400 (N_2400,In_802,In_4053);
or U2401 (N_2401,In_4597,In_809);
and U2402 (N_2402,In_465,In_4283);
and U2403 (N_2403,In_2591,In_3394);
and U2404 (N_2404,In_1135,In_1829);
nand U2405 (N_2405,In_3744,In_4651);
or U2406 (N_2406,In_80,In_116);
nor U2407 (N_2407,In_4475,In_19);
nand U2408 (N_2408,In_2849,In_4589);
xnor U2409 (N_2409,In_2243,In_3625);
nor U2410 (N_2410,In_2508,In_1546);
or U2411 (N_2411,In_3527,In_3934);
nand U2412 (N_2412,In_3315,In_2634);
or U2413 (N_2413,In_4804,In_1157);
and U2414 (N_2414,In_4501,In_4324);
nand U2415 (N_2415,In_2970,In_2619);
nand U2416 (N_2416,In_3095,In_4904);
and U2417 (N_2417,In_1849,In_1775);
nand U2418 (N_2418,In_4787,In_2079);
nor U2419 (N_2419,In_3986,In_4594);
and U2420 (N_2420,In_3655,In_4109);
or U2421 (N_2421,In_69,In_4635);
nor U2422 (N_2422,In_569,In_2446);
or U2423 (N_2423,In_3004,In_144);
nand U2424 (N_2424,In_1899,In_3207);
nor U2425 (N_2425,In_3010,In_4113);
and U2426 (N_2426,In_3107,In_417);
nand U2427 (N_2427,In_2039,In_432);
nor U2428 (N_2428,In_1358,In_2958);
nand U2429 (N_2429,In_894,In_4763);
or U2430 (N_2430,In_2715,In_3473);
and U2431 (N_2431,In_4387,In_4493);
nor U2432 (N_2432,In_1713,In_4338);
nor U2433 (N_2433,In_694,In_3945);
nand U2434 (N_2434,In_283,In_4498);
nand U2435 (N_2435,In_4264,In_4910);
nand U2436 (N_2436,In_1300,In_4130);
nor U2437 (N_2437,In_4018,In_4914);
and U2438 (N_2438,In_1402,In_2828);
or U2439 (N_2439,In_100,In_1512);
nor U2440 (N_2440,In_2586,In_4427);
or U2441 (N_2441,In_2987,In_3914);
nor U2442 (N_2442,In_288,In_2196);
and U2443 (N_2443,In_3806,In_4364);
nand U2444 (N_2444,In_3242,In_560);
or U2445 (N_2445,In_4034,In_4485);
nor U2446 (N_2446,In_1461,In_1043);
and U2447 (N_2447,In_3637,In_1340);
nand U2448 (N_2448,In_865,In_3024);
nand U2449 (N_2449,In_3203,In_130);
nor U2450 (N_2450,In_3898,In_4314);
nand U2451 (N_2451,In_1338,In_677);
nand U2452 (N_2452,In_1708,In_4973);
nand U2453 (N_2453,In_219,In_169);
nand U2454 (N_2454,In_3987,In_2176);
and U2455 (N_2455,In_638,In_3866);
and U2456 (N_2456,In_1845,In_3409);
and U2457 (N_2457,In_2133,In_1072);
nand U2458 (N_2458,In_4067,In_3533);
nand U2459 (N_2459,In_1709,In_214);
and U2460 (N_2460,In_1587,In_543);
xnor U2461 (N_2461,In_3960,In_4222);
nand U2462 (N_2462,In_2629,In_4515);
nand U2463 (N_2463,In_869,In_2706);
xnor U2464 (N_2464,In_2507,In_4965);
or U2465 (N_2465,In_821,In_858);
xor U2466 (N_2466,In_459,In_4543);
or U2467 (N_2467,In_1716,In_1651);
nor U2468 (N_2468,In_2867,In_29);
nor U2469 (N_2469,In_702,In_146);
or U2470 (N_2470,In_1596,In_1684);
or U2471 (N_2471,In_2237,In_1705);
nand U2472 (N_2472,In_348,In_1776);
and U2473 (N_2473,In_2578,In_1610);
or U2474 (N_2474,In_4262,In_339);
nor U2475 (N_2475,In_943,In_798);
nor U2476 (N_2476,In_15,In_4982);
nand U2477 (N_2477,In_4941,In_4989);
nand U2478 (N_2478,In_2028,In_784);
and U2479 (N_2479,In_2214,In_4399);
nor U2480 (N_2480,In_4473,In_3862);
nand U2481 (N_2481,In_1046,In_4259);
nand U2482 (N_2482,In_4905,In_6);
xor U2483 (N_2483,In_2467,In_3982);
nand U2484 (N_2484,In_178,In_2983);
xnor U2485 (N_2485,In_3871,In_4425);
or U2486 (N_2486,In_3346,In_4778);
nor U2487 (N_2487,In_4516,In_795);
or U2488 (N_2488,In_4369,In_4939);
nor U2489 (N_2489,In_1938,In_4206);
nor U2490 (N_2490,In_1428,In_610);
nor U2491 (N_2491,In_1503,In_845);
nor U2492 (N_2492,In_1931,In_4837);
nand U2493 (N_2493,In_4366,In_1455);
nand U2494 (N_2494,In_3143,In_1814);
nor U2495 (N_2495,In_3400,In_1398);
nand U2496 (N_2496,In_2540,In_3599);
or U2497 (N_2497,In_2902,In_962);
or U2498 (N_2498,In_4797,In_3053);
nand U2499 (N_2499,In_1910,In_4511);
and U2500 (N_2500,In_2063,In_2318);
nand U2501 (N_2501,In_1926,In_600);
xnor U2502 (N_2502,In_4155,In_1335);
or U2503 (N_2503,In_1177,In_2886);
nand U2504 (N_2504,In_685,In_949);
xnor U2505 (N_2505,In_4432,In_4954);
and U2506 (N_2506,In_729,In_898);
or U2507 (N_2507,In_2661,In_3774);
xnor U2508 (N_2508,In_3205,In_540);
nor U2509 (N_2509,In_1076,In_2575);
or U2510 (N_2510,In_2239,In_3301);
nand U2511 (N_2511,In_3864,In_1020);
and U2512 (N_2512,In_4384,In_4380);
nand U2513 (N_2513,In_3186,In_1563);
nor U2514 (N_2514,In_680,In_1114);
nor U2515 (N_2515,In_1414,In_1640);
or U2516 (N_2516,In_2217,In_4807);
and U2517 (N_2517,In_55,In_4999);
xor U2518 (N_2518,In_3849,In_1579);
nand U2519 (N_2519,In_4312,In_323);
xnor U2520 (N_2520,In_2953,In_3773);
or U2521 (N_2521,In_3942,In_1755);
nand U2522 (N_2522,In_2965,In_3611);
nor U2523 (N_2523,In_2244,In_2754);
nand U2524 (N_2524,In_1829,In_522);
and U2525 (N_2525,In_3285,In_1959);
and U2526 (N_2526,In_1101,In_1279);
nand U2527 (N_2527,In_2013,In_1743);
or U2528 (N_2528,In_4193,In_2792);
and U2529 (N_2529,In_1103,In_3476);
and U2530 (N_2530,In_1895,In_4723);
nor U2531 (N_2531,In_201,In_612);
nand U2532 (N_2532,In_262,In_3312);
or U2533 (N_2533,In_4540,In_4699);
and U2534 (N_2534,In_1365,In_4965);
or U2535 (N_2535,In_1211,In_2406);
nand U2536 (N_2536,In_4740,In_4481);
and U2537 (N_2537,In_4929,In_1621);
xnor U2538 (N_2538,In_2941,In_4228);
or U2539 (N_2539,In_2643,In_4237);
nor U2540 (N_2540,In_4996,In_3580);
nand U2541 (N_2541,In_369,In_1680);
nor U2542 (N_2542,In_3588,In_184);
nand U2543 (N_2543,In_415,In_1358);
nor U2544 (N_2544,In_2517,In_2362);
xnor U2545 (N_2545,In_1130,In_4564);
or U2546 (N_2546,In_2328,In_125);
or U2547 (N_2547,In_2500,In_3602);
nor U2548 (N_2548,In_3342,In_3625);
nand U2549 (N_2549,In_4381,In_202);
xor U2550 (N_2550,In_3240,In_407);
nand U2551 (N_2551,In_4973,In_1048);
xor U2552 (N_2552,In_1724,In_618);
nand U2553 (N_2553,In_3178,In_809);
nor U2554 (N_2554,In_348,In_2689);
nand U2555 (N_2555,In_3743,In_3252);
nor U2556 (N_2556,In_1797,In_4848);
nand U2557 (N_2557,In_1735,In_2713);
nand U2558 (N_2558,In_1046,In_2574);
nor U2559 (N_2559,In_4650,In_2839);
nor U2560 (N_2560,In_4245,In_3617);
nand U2561 (N_2561,In_2100,In_4050);
and U2562 (N_2562,In_4885,In_2109);
nor U2563 (N_2563,In_307,In_3828);
nand U2564 (N_2564,In_4891,In_3619);
nor U2565 (N_2565,In_2222,In_4809);
or U2566 (N_2566,In_4258,In_4453);
nor U2567 (N_2567,In_3625,In_1620);
nor U2568 (N_2568,In_1166,In_4750);
nor U2569 (N_2569,In_3212,In_4658);
and U2570 (N_2570,In_3490,In_1037);
xor U2571 (N_2571,In_4721,In_2801);
xor U2572 (N_2572,In_4825,In_1465);
and U2573 (N_2573,In_703,In_2658);
nand U2574 (N_2574,In_3120,In_578);
nor U2575 (N_2575,In_3928,In_3997);
nand U2576 (N_2576,In_1586,In_309);
or U2577 (N_2577,In_4499,In_1669);
and U2578 (N_2578,In_880,In_1451);
nand U2579 (N_2579,In_1496,In_280);
nor U2580 (N_2580,In_4248,In_1318);
and U2581 (N_2581,In_1998,In_1437);
and U2582 (N_2582,In_4380,In_4630);
xor U2583 (N_2583,In_24,In_308);
or U2584 (N_2584,In_3911,In_882);
xnor U2585 (N_2585,In_326,In_1083);
or U2586 (N_2586,In_4795,In_1384);
nor U2587 (N_2587,In_828,In_4461);
and U2588 (N_2588,In_141,In_2093);
nand U2589 (N_2589,In_3427,In_4768);
or U2590 (N_2590,In_3525,In_3842);
xor U2591 (N_2591,In_2064,In_2663);
nand U2592 (N_2592,In_1490,In_2153);
nand U2593 (N_2593,In_1267,In_3717);
nand U2594 (N_2594,In_4685,In_3823);
nand U2595 (N_2595,In_2924,In_3228);
or U2596 (N_2596,In_41,In_2307);
xor U2597 (N_2597,In_158,In_3191);
nor U2598 (N_2598,In_957,In_4409);
and U2599 (N_2599,In_220,In_1520);
or U2600 (N_2600,In_3731,In_205);
nand U2601 (N_2601,In_4304,In_3451);
or U2602 (N_2602,In_2574,In_883);
and U2603 (N_2603,In_54,In_1038);
and U2604 (N_2604,In_2753,In_57);
and U2605 (N_2605,In_269,In_1971);
or U2606 (N_2606,In_4326,In_3045);
nor U2607 (N_2607,In_1446,In_3314);
and U2608 (N_2608,In_2168,In_3727);
nand U2609 (N_2609,In_2101,In_3585);
or U2610 (N_2610,In_89,In_3668);
and U2611 (N_2611,In_2481,In_111);
xnor U2612 (N_2612,In_1655,In_2910);
and U2613 (N_2613,In_966,In_3509);
nor U2614 (N_2614,In_2314,In_2750);
and U2615 (N_2615,In_4753,In_4475);
and U2616 (N_2616,In_3518,In_1748);
nor U2617 (N_2617,In_4445,In_4339);
or U2618 (N_2618,In_1163,In_3225);
xnor U2619 (N_2619,In_1211,In_524);
and U2620 (N_2620,In_2895,In_1696);
and U2621 (N_2621,In_946,In_3635);
nor U2622 (N_2622,In_3560,In_4608);
nor U2623 (N_2623,In_4445,In_3791);
or U2624 (N_2624,In_1123,In_2575);
nand U2625 (N_2625,In_4419,In_1161);
and U2626 (N_2626,In_4293,In_3291);
or U2627 (N_2627,In_2645,In_2638);
xnor U2628 (N_2628,In_2709,In_4869);
and U2629 (N_2629,In_921,In_400);
or U2630 (N_2630,In_4254,In_2890);
nor U2631 (N_2631,In_3437,In_1206);
nand U2632 (N_2632,In_3544,In_3453);
and U2633 (N_2633,In_4922,In_149);
or U2634 (N_2634,In_1316,In_4575);
xnor U2635 (N_2635,In_4932,In_1160);
or U2636 (N_2636,In_3310,In_631);
nand U2637 (N_2637,In_3144,In_394);
and U2638 (N_2638,In_294,In_3215);
and U2639 (N_2639,In_972,In_4742);
or U2640 (N_2640,In_3080,In_859);
xnor U2641 (N_2641,In_3342,In_1450);
nor U2642 (N_2642,In_3617,In_3067);
and U2643 (N_2643,In_3837,In_3129);
or U2644 (N_2644,In_3601,In_2556);
xnor U2645 (N_2645,In_2596,In_4421);
and U2646 (N_2646,In_3548,In_4641);
and U2647 (N_2647,In_1732,In_1513);
and U2648 (N_2648,In_711,In_3235);
nor U2649 (N_2649,In_3793,In_1099);
xor U2650 (N_2650,In_4053,In_2018);
nand U2651 (N_2651,In_1952,In_2136);
nand U2652 (N_2652,In_1869,In_2759);
xor U2653 (N_2653,In_3615,In_4770);
xor U2654 (N_2654,In_4880,In_1742);
nand U2655 (N_2655,In_2110,In_2505);
nor U2656 (N_2656,In_2093,In_4564);
nand U2657 (N_2657,In_3464,In_666);
and U2658 (N_2658,In_1011,In_267);
or U2659 (N_2659,In_1131,In_4824);
and U2660 (N_2660,In_2888,In_257);
nor U2661 (N_2661,In_2755,In_4481);
nand U2662 (N_2662,In_2561,In_2300);
or U2663 (N_2663,In_1975,In_814);
nand U2664 (N_2664,In_2214,In_4623);
and U2665 (N_2665,In_788,In_542);
or U2666 (N_2666,In_4972,In_2555);
xnor U2667 (N_2667,In_4477,In_2233);
or U2668 (N_2668,In_4697,In_3973);
nor U2669 (N_2669,In_945,In_3770);
nand U2670 (N_2670,In_3176,In_4443);
nand U2671 (N_2671,In_4315,In_3308);
nand U2672 (N_2672,In_1349,In_560);
nand U2673 (N_2673,In_1949,In_3037);
or U2674 (N_2674,In_3659,In_4795);
nor U2675 (N_2675,In_1561,In_120);
nand U2676 (N_2676,In_1806,In_1347);
and U2677 (N_2677,In_4304,In_2572);
and U2678 (N_2678,In_2715,In_4522);
nand U2679 (N_2679,In_391,In_1714);
and U2680 (N_2680,In_4840,In_515);
or U2681 (N_2681,In_278,In_4221);
and U2682 (N_2682,In_1555,In_4010);
or U2683 (N_2683,In_3216,In_1784);
xor U2684 (N_2684,In_4965,In_4569);
nand U2685 (N_2685,In_3275,In_2838);
xnor U2686 (N_2686,In_2487,In_1766);
or U2687 (N_2687,In_4886,In_587);
or U2688 (N_2688,In_1739,In_4648);
nand U2689 (N_2689,In_1619,In_834);
nor U2690 (N_2690,In_7,In_2629);
and U2691 (N_2691,In_3577,In_260);
nor U2692 (N_2692,In_1485,In_1431);
and U2693 (N_2693,In_4336,In_3323);
nand U2694 (N_2694,In_3986,In_4093);
xor U2695 (N_2695,In_381,In_698);
or U2696 (N_2696,In_3931,In_4815);
and U2697 (N_2697,In_4855,In_3601);
or U2698 (N_2698,In_971,In_2227);
nand U2699 (N_2699,In_424,In_3460);
nor U2700 (N_2700,In_961,In_3888);
xor U2701 (N_2701,In_3935,In_1959);
nand U2702 (N_2702,In_1581,In_3802);
xnor U2703 (N_2703,In_2866,In_3447);
nand U2704 (N_2704,In_4922,In_1926);
and U2705 (N_2705,In_2221,In_1446);
nand U2706 (N_2706,In_1124,In_417);
or U2707 (N_2707,In_4508,In_1618);
xnor U2708 (N_2708,In_3753,In_1574);
and U2709 (N_2709,In_3093,In_2305);
xor U2710 (N_2710,In_976,In_3605);
nand U2711 (N_2711,In_3011,In_571);
and U2712 (N_2712,In_3377,In_1439);
or U2713 (N_2713,In_1078,In_2586);
xnor U2714 (N_2714,In_4566,In_1341);
nor U2715 (N_2715,In_1598,In_1107);
or U2716 (N_2716,In_2862,In_3268);
or U2717 (N_2717,In_4807,In_4975);
or U2718 (N_2718,In_2342,In_4618);
or U2719 (N_2719,In_2538,In_3077);
and U2720 (N_2720,In_848,In_1919);
or U2721 (N_2721,In_1280,In_4521);
and U2722 (N_2722,In_881,In_2348);
xnor U2723 (N_2723,In_4988,In_1247);
and U2724 (N_2724,In_623,In_2647);
or U2725 (N_2725,In_2180,In_4258);
nand U2726 (N_2726,In_3657,In_876);
and U2727 (N_2727,In_3814,In_4772);
or U2728 (N_2728,In_3698,In_771);
nor U2729 (N_2729,In_1175,In_4962);
or U2730 (N_2730,In_4809,In_1956);
nor U2731 (N_2731,In_871,In_1908);
nand U2732 (N_2732,In_1782,In_1552);
or U2733 (N_2733,In_4172,In_4634);
nand U2734 (N_2734,In_3045,In_3268);
nor U2735 (N_2735,In_2182,In_2131);
or U2736 (N_2736,In_4441,In_3076);
and U2737 (N_2737,In_2526,In_698);
and U2738 (N_2738,In_4437,In_4382);
nor U2739 (N_2739,In_877,In_3883);
nor U2740 (N_2740,In_3461,In_1578);
nand U2741 (N_2741,In_1831,In_4312);
nand U2742 (N_2742,In_4964,In_1152);
or U2743 (N_2743,In_3974,In_207);
nand U2744 (N_2744,In_2640,In_4485);
nor U2745 (N_2745,In_1931,In_3270);
xnor U2746 (N_2746,In_104,In_3052);
xor U2747 (N_2747,In_2672,In_2360);
nor U2748 (N_2748,In_4065,In_1037);
nand U2749 (N_2749,In_631,In_909);
or U2750 (N_2750,In_1091,In_4067);
and U2751 (N_2751,In_321,In_4738);
and U2752 (N_2752,In_657,In_1108);
nor U2753 (N_2753,In_1439,In_3717);
nand U2754 (N_2754,In_716,In_3358);
nand U2755 (N_2755,In_3069,In_461);
nand U2756 (N_2756,In_1008,In_4604);
nor U2757 (N_2757,In_982,In_3829);
xnor U2758 (N_2758,In_2662,In_3806);
xnor U2759 (N_2759,In_4853,In_2190);
nand U2760 (N_2760,In_229,In_2111);
nand U2761 (N_2761,In_240,In_121);
xnor U2762 (N_2762,In_1802,In_3814);
nand U2763 (N_2763,In_2570,In_1892);
and U2764 (N_2764,In_1906,In_4691);
or U2765 (N_2765,In_3672,In_1404);
nor U2766 (N_2766,In_2052,In_2783);
and U2767 (N_2767,In_1933,In_4327);
and U2768 (N_2768,In_3373,In_3974);
and U2769 (N_2769,In_2637,In_3551);
xor U2770 (N_2770,In_1218,In_879);
or U2771 (N_2771,In_2662,In_4390);
and U2772 (N_2772,In_1472,In_3441);
nand U2773 (N_2773,In_2959,In_1573);
xnor U2774 (N_2774,In_1456,In_508);
and U2775 (N_2775,In_2124,In_2156);
and U2776 (N_2776,In_2787,In_3628);
nor U2777 (N_2777,In_1864,In_3479);
nand U2778 (N_2778,In_4348,In_4954);
nor U2779 (N_2779,In_110,In_1312);
nor U2780 (N_2780,In_2944,In_1231);
xnor U2781 (N_2781,In_1378,In_2098);
or U2782 (N_2782,In_483,In_2987);
nand U2783 (N_2783,In_1447,In_3751);
nor U2784 (N_2784,In_4949,In_867);
xnor U2785 (N_2785,In_3910,In_4782);
or U2786 (N_2786,In_2012,In_3048);
or U2787 (N_2787,In_4687,In_1337);
xor U2788 (N_2788,In_2375,In_4548);
nand U2789 (N_2789,In_4889,In_1191);
or U2790 (N_2790,In_2895,In_4227);
xnor U2791 (N_2791,In_115,In_84);
nor U2792 (N_2792,In_4504,In_1389);
or U2793 (N_2793,In_1541,In_1035);
nor U2794 (N_2794,In_469,In_1379);
nor U2795 (N_2795,In_1752,In_1551);
xnor U2796 (N_2796,In_1469,In_4885);
nand U2797 (N_2797,In_2915,In_2634);
nand U2798 (N_2798,In_862,In_3974);
nand U2799 (N_2799,In_2529,In_3273);
nor U2800 (N_2800,In_96,In_4038);
and U2801 (N_2801,In_2064,In_116);
and U2802 (N_2802,In_1935,In_1252);
or U2803 (N_2803,In_4211,In_1486);
nor U2804 (N_2804,In_3727,In_1586);
xnor U2805 (N_2805,In_3723,In_3995);
nor U2806 (N_2806,In_2083,In_1089);
nand U2807 (N_2807,In_276,In_16);
and U2808 (N_2808,In_2181,In_2447);
and U2809 (N_2809,In_1712,In_3569);
nor U2810 (N_2810,In_23,In_896);
and U2811 (N_2811,In_1807,In_672);
and U2812 (N_2812,In_2573,In_1379);
and U2813 (N_2813,In_3187,In_4063);
nand U2814 (N_2814,In_874,In_3407);
and U2815 (N_2815,In_4990,In_4252);
nor U2816 (N_2816,In_2491,In_4572);
nand U2817 (N_2817,In_731,In_3844);
nand U2818 (N_2818,In_1993,In_4662);
xnor U2819 (N_2819,In_4000,In_4295);
nand U2820 (N_2820,In_3906,In_4432);
nor U2821 (N_2821,In_1498,In_3902);
and U2822 (N_2822,In_4375,In_2264);
nor U2823 (N_2823,In_1278,In_2416);
or U2824 (N_2824,In_2549,In_4712);
and U2825 (N_2825,In_1766,In_2816);
nor U2826 (N_2826,In_3338,In_4131);
nor U2827 (N_2827,In_257,In_1005);
and U2828 (N_2828,In_4815,In_266);
and U2829 (N_2829,In_995,In_3893);
or U2830 (N_2830,In_1418,In_2800);
and U2831 (N_2831,In_322,In_3758);
or U2832 (N_2832,In_1695,In_2492);
nand U2833 (N_2833,In_808,In_1990);
xnor U2834 (N_2834,In_1662,In_250);
or U2835 (N_2835,In_1801,In_4670);
xnor U2836 (N_2836,In_3401,In_3548);
xnor U2837 (N_2837,In_1154,In_3324);
or U2838 (N_2838,In_185,In_2567);
or U2839 (N_2839,In_2180,In_2667);
nor U2840 (N_2840,In_821,In_4339);
nor U2841 (N_2841,In_3195,In_3409);
nor U2842 (N_2842,In_556,In_671);
and U2843 (N_2843,In_2393,In_2543);
and U2844 (N_2844,In_2781,In_417);
nor U2845 (N_2845,In_1456,In_280);
and U2846 (N_2846,In_4437,In_1276);
or U2847 (N_2847,In_83,In_3794);
xnor U2848 (N_2848,In_2318,In_3230);
nand U2849 (N_2849,In_1539,In_1225);
nand U2850 (N_2850,In_2051,In_4168);
or U2851 (N_2851,In_163,In_2536);
and U2852 (N_2852,In_2900,In_4440);
nand U2853 (N_2853,In_584,In_4791);
and U2854 (N_2854,In_3918,In_541);
or U2855 (N_2855,In_2569,In_3029);
nor U2856 (N_2856,In_750,In_261);
nor U2857 (N_2857,In_1541,In_4688);
nor U2858 (N_2858,In_3096,In_2131);
and U2859 (N_2859,In_2927,In_4172);
or U2860 (N_2860,In_2097,In_2648);
or U2861 (N_2861,In_3021,In_838);
or U2862 (N_2862,In_2758,In_237);
nor U2863 (N_2863,In_1717,In_2793);
and U2864 (N_2864,In_4886,In_1475);
or U2865 (N_2865,In_2550,In_3547);
and U2866 (N_2866,In_1309,In_3154);
and U2867 (N_2867,In_1741,In_4530);
nand U2868 (N_2868,In_2564,In_4720);
nor U2869 (N_2869,In_1095,In_2194);
nand U2870 (N_2870,In_2397,In_29);
or U2871 (N_2871,In_1258,In_4445);
or U2872 (N_2872,In_3274,In_2091);
nand U2873 (N_2873,In_3895,In_3185);
nand U2874 (N_2874,In_3390,In_1699);
or U2875 (N_2875,In_1634,In_4150);
xnor U2876 (N_2876,In_2237,In_4362);
nor U2877 (N_2877,In_30,In_1988);
or U2878 (N_2878,In_1239,In_4519);
or U2879 (N_2879,In_2127,In_3590);
xor U2880 (N_2880,In_2288,In_3777);
or U2881 (N_2881,In_2502,In_3740);
or U2882 (N_2882,In_987,In_2483);
and U2883 (N_2883,In_483,In_3551);
nor U2884 (N_2884,In_2933,In_255);
or U2885 (N_2885,In_1500,In_1444);
nor U2886 (N_2886,In_2573,In_177);
and U2887 (N_2887,In_3991,In_3177);
or U2888 (N_2888,In_1179,In_3604);
nor U2889 (N_2889,In_3886,In_320);
nor U2890 (N_2890,In_1083,In_4327);
nor U2891 (N_2891,In_50,In_1631);
or U2892 (N_2892,In_1126,In_4730);
nand U2893 (N_2893,In_3484,In_1126);
nand U2894 (N_2894,In_4854,In_197);
nand U2895 (N_2895,In_3846,In_2475);
xnor U2896 (N_2896,In_1678,In_783);
or U2897 (N_2897,In_1029,In_519);
nand U2898 (N_2898,In_1156,In_3501);
or U2899 (N_2899,In_4689,In_1915);
and U2900 (N_2900,In_4432,In_978);
nor U2901 (N_2901,In_3002,In_4408);
and U2902 (N_2902,In_4468,In_2399);
nand U2903 (N_2903,In_1301,In_3648);
or U2904 (N_2904,In_3101,In_4501);
or U2905 (N_2905,In_4203,In_4239);
or U2906 (N_2906,In_1104,In_1898);
or U2907 (N_2907,In_657,In_2661);
and U2908 (N_2908,In_1473,In_637);
nor U2909 (N_2909,In_4835,In_3954);
nand U2910 (N_2910,In_4816,In_3435);
or U2911 (N_2911,In_3860,In_4314);
and U2912 (N_2912,In_2367,In_3089);
nand U2913 (N_2913,In_3525,In_561);
or U2914 (N_2914,In_2598,In_2276);
xor U2915 (N_2915,In_3358,In_128);
nand U2916 (N_2916,In_2815,In_4342);
xnor U2917 (N_2917,In_1508,In_3954);
and U2918 (N_2918,In_556,In_2029);
or U2919 (N_2919,In_2933,In_1892);
nand U2920 (N_2920,In_4825,In_2501);
or U2921 (N_2921,In_1907,In_33);
nand U2922 (N_2922,In_2271,In_4423);
or U2923 (N_2923,In_3328,In_1028);
or U2924 (N_2924,In_4305,In_4772);
nor U2925 (N_2925,In_4365,In_3510);
or U2926 (N_2926,In_4209,In_3604);
nand U2927 (N_2927,In_807,In_162);
nor U2928 (N_2928,In_2709,In_2032);
nor U2929 (N_2929,In_2711,In_3538);
nand U2930 (N_2930,In_3436,In_3692);
and U2931 (N_2931,In_2524,In_3698);
xnor U2932 (N_2932,In_167,In_290);
or U2933 (N_2933,In_1232,In_2868);
nand U2934 (N_2934,In_3666,In_4437);
nor U2935 (N_2935,In_929,In_4339);
and U2936 (N_2936,In_4338,In_1561);
nor U2937 (N_2937,In_4716,In_903);
and U2938 (N_2938,In_3139,In_340);
nor U2939 (N_2939,In_1437,In_105);
nor U2940 (N_2940,In_635,In_4415);
nand U2941 (N_2941,In_3913,In_3400);
and U2942 (N_2942,In_59,In_4453);
or U2943 (N_2943,In_367,In_4869);
nor U2944 (N_2944,In_1987,In_3523);
xor U2945 (N_2945,In_3466,In_3510);
xnor U2946 (N_2946,In_3193,In_868);
nor U2947 (N_2947,In_4580,In_3084);
nor U2948 (N_2948,In_2291,In_4303);
nor U2949 (N_2949,In_2794,In_2197);
or U2950 (N_2950,In_4794,In_1338);
and U2951 (N_2951,In_2311,In_2805);
or U2952 (N_2952,In_1758,In_37);
xor U2953 (N_2953,In_3784,In_2117);
nor U2954 (N_2954,In_4887,In_305);
or U2955 (N_2955,In_353,In_4487);
nor U2956 (N_2956,In_176,In_272);
nor U2957 (N_2957,In_1140,In_3903);
and U2958 (N_2958,In_3947,In_2751);
and U2959 (N_2959,In_3491,In_19);
or U2960 (N_2960,In_3238,In_1936);
nor U2961 (N_2961,In_3604,In_514);
nor U2962 (N_2962,In_2244,In_3718);
and U2963 (N_2963,In_420,In_4094);
or U2964 (N_2964,In_16,In_4363);
nand U2965 (N_2965,In_3353,In_794);
nor U2966 (N_2966,In_985,In_759);
nand U2967 (N_2967,In_3232,In_3884);
nor U2968 (N_2968,In_4722,In_3276);
nand U2969 (N_2969,In_4320,In_3805);
xnor U2970 (N_2970,In_967,In_436);
and U2971 (N_2971,In_507,In_3498);
and U2972 (N_2972,In_2955,In_805);
and U2973 (N_2973,In_4420,In_320);
xnor U2974 (N_2974,In_882,In_2373);
nor U2975 (N_2975,In_4276,In_872);
or U2976 (N_2976,In_3055,In_2038);
and U2977 (N_2977,In_4956,In_2730);
nor U2978 (N_2978,In_2615,In_3678);
xnor U2979 (N_2979,In_4246,In_3745);
or U2980 (N_2980,In_3693,In_3564);
and U2981 (N_2981,In_3518,In_3592);
or U2982 (N_2982,In_2724,In_3152);
and U2983 (N_2983,In_2151,In_189);
xnor U2984 (N_2984,In_1408,In_884);
nor U2985 (N_2985,In_3218,In_1798);
nor U2986 (N_2986,In_3970,In_770);
nand U2987 (N_2987,In_3958,In_2040);
nand U2988 (N_2988,In_31,In_3674);
nand U2989 (N_2989,In_3431,In_1120);
nand U2990 (N_2990,In_844,In_2601);
and U2991 (N_2991,In_3965,In_4648);
xnor U2992 (N_2992,In_4183,In_773);
nor U2993 (N_2993,In_2538,In_3961);
or U2994 (N_2994,In_3429,In_4489);
xor U2995 (N_2995,In_2446,In_1458);
nor U2996 (N_2996,In_3474,In_422);
nand U2997 (N_2997,In_662,In_2792);
or U2998 (N_2998,In_1595,In_855);
xor U2999 (N_2999,In_3775,In_4304);
nand U3000 (N_3000,In_2979,In_4909);
xnor U3001 (N_3001,In_3045,In_4600);
or U3002 (N_3002,In_470,In_4565);
and U3003 (N_3003,In_3915,In_4743);
nor U3004 (N_3004,In_2605,In_2846);
xnor U3005 (N_3005,In_4159,In_3288);
and U3006 (N_3006,In_4981,In_4214);
nor U3007 (N_3007,In_1997,In_884);
nand U3008 (N_3008,In_484,In_1815);
and U3009 (N_3009,In_265,In_865);
nand U3010 (N_3010,In_2067,In_1453);
nor U3011 (N_3011,In_3844,In_3898);
nand U3012 (N_3012,In_1234,In_664);
nor U3013 (N_3013,In_1430,In_1468);
nor U3014 (N_3014,In_1093,In_2049);
nor U3015 (N_3015,In_2731,In_1945);
or U3016 (N_3016,In_3583,In_456);
xnor U3017 (N_3017,In_1094,In_2467);
nor U3018 (N_3018,In_57,In_1960);
nand U3019 (N_3019,In_2919,In_3367);
or U3020 (N_3020,In_3810,In_1678);
or U3021 (N_3021,In_4259,In_214);
nor U3022 (N_3022,In_1852,In_1819);
xor U3023 (N_3023,In_464,In_2140);
and U3024 (N_3024,In_2880,In_2740);
and U3025 (N_3025,In_1746,In_1452);
nand U3026 (N_3026,In_779,In_519);
nor U3027 (N_3027,In_1287,In_1025);
and U3028 (N_3028,In_1652,In_4325);
nand U3029 (N_3029,In_3668,In_4094);
nand U3030 (N_3030,In_926,In_3717);
nand U3031 (N_3031,In_1394,In_3900);
and U3032 (N_3032,In_3386,In_2056);
and U3033 (N_3033,In_4644,In_149);
nand U3034 (N_3034,In_565,In_4275);
nand U3035 (N_3035,In_2140,In_1641);
or U3036 (N_3036,In_1540,In_4780);
xor U3037 (N_3037,In_3700,In_2289);
and U3038 (N_3038,In_3951,In_4231);
and U3039 (N_3039,In_2992,In_181);
nor U3040 (N_3040,In_3954,In_1591);
nand U3041 (N_3041,In_2521,In_1116);
and U3042 (N_3042,In_3411,In_191);
xor U3043 (N_3043,In_3362,In_1227);
or U3044 (N_3044,In_4362,In_1135);
nand U3045 (N_3045,In_4689,In_3771);
or U3046 (N_3046,In_3544,In_1598);
nor U3047 (N_3047,In_557,In_2824);
and U3048 (N_3048,In_3903,In_3112);
nand U3049 (N_3049,In_550,In_119);
nand U3050 (N_3050,In_3605,In_4744);
nand U3051 (N_3051,In_1115,In_1174);
nand U3052 (N_3052,In_1028,In_1842);
and U3053 (N_3053,In_4194,In_2134);
and U3054 (N_3054,In_9,In_3913);
and U3055 (N_3055,In_846,In_1845);
and U3056 (N_3056,In_2257,In_2803);
nor U3057 (N_3057,In_2231,In_4864);
xnor U3058 (N_3058,In_4402,In_676);
or U3059 (N_3059,In_1450,In_1734);
nand U3060 (N_3060,In_4475,In_1500);
or U3061 (N_3061,In_662,In_1560);
nand U3062 (N_3062,In_797,In_1995);
nor U3063 (N_3063,In_4135,In_4284);
nand U3064 (N_3064,In_1832,In_2366);
and U3065 (N_3065,In_3814,In_4427);
nor U3066 (N_3066,In_4219,In_4044);
nand U3067 (N_3067,In_2675,In_2776);
and U3068 (N_3068,In_4364,In_92);
nand U3069 (N_3069,In_1070,In_3480);
or U3070 (N_3070,In_498,In_1861);
and U3071 (N_3071,In_1004,In_529);
and U3072 (N_3072,In_4232,In_1921);
nand U3073 (N_3073,In_544,In_4279);
or U3074 (N_3074,In_3285,In_4649);
and U3075 (N_3075,In_4227,In_1285);
or U3076 (N_3076,In_3361,In_4483);
and U3077 (N_3077,In_250,In_428);
nand U3078 (N_3078,In_4493,In_2856);
and U3079 (N_3079,In_274,In_3341);
and U3080 (N_3080,In_2765,In_706);
or U3081 (N_3081,In_2757,In_4754);
nor U3082 (N_3082,In_4578,In_1408);
nand U3083 (N_3083,In_1184,In_4873);
nor U3084 (N_3084,In_2841,In_3210);
xnor U3085 (N_3085,In_4465,In_1471);
nand U3086 (N_3086,In_3211,In_2040);
nor U3087 (N_3087,In_4971,In_1600);
or U3088 (N_3088,In_2794,In_3838);
or U3089 (N_3089,In_475,In_2529);
nor U3090 (N_3090,In_4891,In_2771);
or U3091 (N_3091,In_729,In_2660);
xor U3092 (N_3092,In_2968,In_1141);
and U3093 (N_3093,In_478,In_3220);
and U3094 (N_3094,In_2518,In_2894);
or U3095 (N_3095,In_405,In_2847);
and U3096 (N_3096,In_1494,In_1148);
or U3097 (N_3097,In_2530,In_4900);
or U3098 (N_3098,In_1477,In_3913);
or U3099 (N_3099,In_1869,In_2295);
nor U3100 (N_3100,In_2040,In_1816);
and U3101 (N_3101,In_3921,In_639);
or U3102 (N_3102,In_2620,In_4532);
nor U3103 (N_3103,In_3206,In_2384);
xnor U3104 (N_3104,In_704,In_2185);
or U3105 (N_3105,In_1518,In_2842);
and U3106 (N_3106,In_1691,In_4595);
xor U3107 (N_3107,In_3334,In_3349);
nor U3108 (N_3108,In_4447,In_145);
nand U3109 (N_3109,In_3640,In_2843);
and U3110 (N_3110,In_4773,In_2178);
xnor U3111 (N_3111,In_976,In_769);
and U3112 (N_3112,In_3299,In_169);
or U3113 (N_3113,In_2131,In_2438);
nor U3114 (N_3114,In_1473,In_1667);
and U3115 (N_3115,In_884,In_2518);
and U3116 (N_3116,In_2120,In_2094);
nor U3117 (N_3117,In_4736,In_724);
nand U3118 (N_3118,In_1531,In_4312);
nand U3119 (N_3119,In_773,In_2186);
xor U3120 (N_3120,In_3713,In_1429);
or U3121 (N_3121,In_3436,In_2226);
xor U3122 (N_3122,In_971,In_3293);
nor U3123 (N_3123,In_687,In_839);
xor U3124 (N_3124,In_3485,In_3663);
nand U3125 (N_3125,In_3999,In_2666);
nand U3126 (N_3126,In_3242,In_135);
or U3127 (N_3127,In_3430,In_2900);
nand U3128 (N_3128,In_3880,In_3276);
nor U3129 (N_3129,In_3790,In_354);
nor U3130 (N_3130,In_2524,In_4680);
nor U3131 (N_3131,In_469,In_3517);
nor U3132 (N_3132,In_1664,In_3480);
nand U3133 (N_3133,In_3231,In_3026);
and U3134 (N_3134,In_3952,In_3359);
and U3135 (N_3135,In_1695,In_1999);
and U3136 (N_3136,In_723,In_2258);
xnor U3137 (N_3137,In_4847,In_4451);
or U3138 (N_3138,In_1253,In_1171);
nand U3139 (N_3139,In_2438,In_2771);
nand U3140 (N_3140,In_391,In_2457);
or U3141 (N_3141,In_393,In_1118);
xor U3142 (N_3142,In_3649,In_4313);
or U3143 (N_3143,In_31,In_3769);
nand U3144 (N_3144,In_1283,In_3883);
or U3145 (N_3145,In_1156,In_460);
or U3146 (N_3146,In_276,In_2579);
nor U3147 (N_3147,In_143,In_995);
nand U3148 (N_3148,In_775,In_4708);
nor U3149 (N_3149,In_72,In_3857);
xnor U3150 (N_3150,In_2363,In_3793);
or U3151 (N_3151,In_457,In_1548);
or U3152 (N_3152,In_3711,In_1150);
nand U3153 (N_3153,In_1900,In_863);
or U3154 (N_3154,In_3009,In_3400);
nor U3155 (N_3155,In_3765,In_1002);
and U3156 (N_3156,In_3210,In_3975);
nand U3157 (N_3157,In_4640,In_124);
or U3158 (N_3158,In_639,In_2176);
xnor U3159 (N_3159,In_2702,In_3683);
nor U3160 (N_3160,In_1832,In_3168);
or U3161 (N_3161,In_2171,In_4056);
nor U3162 (N_3162,In_3577,In_3366);
nand U3163 (N_3163,In_2327,In_475);
nand U3164 (N_3164,In_3480,In_1200);
or U3165 (N_3165,In_3436,In_4874);
and U3166 (N_3166,In_1188,In_955);
nand U3167 (N_3167,In_3316,In_271);
nand U3168 (N_3168,In_2372,In_3597);
nor U3169 (N_3169,In_2335,In_1376);
and U3170 (N_3170,In_4604,In_820);
nor U3171 (N_3171,In_3683,In_4990);
or U3172 (N_3172,In_680,In_3668);
or U3173 (N_3173,In_438,In_3874);
or U3174 (N_3174,In_1787,In_588);
nor U3175 (N_3175,In_876,In_2056);
xor U3176 (N_3176,In_4526,In_2570);
nor U3177 (N_3177,In_2778,In_2742);
nor U3178 (N_3178,In_2130,In_1115);
and U3179 (N_3179,In_2967,In_4316);
xnor U3180 (N_3180,In_4107,In_1122);
or U3181 (N_3181,In_2181,In_196);
nand U3182 (N_3182,In_93,In_61);
or U3183 (N_3183,In_1570,In_3502);
xnor U3184 (N_3184,In_4901,In_12);
nand U3185 (N_3185,In_658,In_4420);
or U3186 (N_3186,In_2405,In_3120);
nand U3187 (N_3187,In_1365,In_4665);
nor U3188 (N_3188,In_2865,In_94);
or U3189 (N_3189,In_1751,In_2495);
nor U3190 (N_3190,In_2195,In_207);
and U3191 (N_3191,In_1428,In_4214);
nand U3192 (N_3192,In_3545,In_3040);
nor U3193 (N_3193,In_353,In_2008);
nand U3194 (N_3194,In_1511,In_269);
or U3195 (N_3195,In_3444,In_4166);
and U3196 (N_3196,In_2970,In_2074);
nor U3197 (N_3197,In_1973,In_3550);
nand U3198 (N_3198,In_3104,In_363);
nor U3199 (N_3199,In_2785,In_1761);
nand U3200 (N_3200,In_4836,In_4733);
xnor U3201 (N_3201,In_915,In_4824);
nor U3202 (N_3202,In_4775,In_2412);
or U3203 (N_3203,In_3189,In_2116);
nand U3204 (N_3204,In_3023,In_2220);
xor U3205 (N_3205,In_130,In_1644);
nand U3206 (N_3206,In_4253,In_4245);
xnor U3207 (N_3207,In_1150,In_4767);
or U3208 (N_3208,In_3635,In_115);
or U3209 (N_3209,In_2832,In_432);
or U3210 (N_3210,In_277,In_4429);
nand U3211 (N_3211,In_2835,In_4079);
and U3212 (N_3212,In_3052,In_2725);
nand U3213 (N_3213,In_2446,In_4819);
or U3214 (N_3214,In_3298,In_3796);
nand U3215 (N_3215,In_4411,In_3875);
xnor U3216 (N_3216,In_2837,In_4112);
or U3217 (N_3217,In_3245,In_2146);
nor U3218 (N_3218,In_212,In_4246);
nor U3219 (N_3219,In_3552,In_4748);
nand U3220 (N_3220,In_4110,In_3772);
nor U3221 (N_3221,In_4095,In_4963);
nand U3222 (N_3222,In_2289,In_1285);
nand U3223 (N_3223,In_1376,In_519);
nand U3224 (N_3224,In_683,In_808);
xor U3225 (N_3225,In_3034,In_425);
nand U3226 (N_3226,In_549,In_4886);
nand U3227 (N_3227,In_3551,In_474);
nand U3228 (N_3228,In_2968,In_3259);
and U3229 (N_3229,In_3720,In_1223);
and U3230 (N_3230,In_604,In_1929);
and U3231 (N_3231,In_3129,In_556);
or U3232 (N_3232,In_3598,In_3910);
xor U3233 (N_3233,In_3701,In_1334);
and U3234 (N_3234,In_4082,In_3580);
and U3235 (N_3235,In_1773,In_227);
and U3236 (N_3236,In_3890,In_3604);
nor U3237 (N_3237,In_582,In_430);
nand U3238 (N_3238,In_891,In_3931);
and U3239 (N_3239,In_2232,In_1228);
and U3240 (N_3240,In_3980,In_3150);
nor U3241 (N_3241,In_4330,In_4389);
nand U3242 (N_3242,In_3697,In_2509);
and U3243 (N_3243,In_4971,In_3841);
and U3244 (N_3244,In_4102,In_2690);
and U3245 (N_3245,In_4025,In_4971);
or U3246 (N_3246,In_2220,In_2264);
nor U3247 (N_3247,In_776,In_2229);
and U3248 (N_3248,In_4223,In_1204);
nor U3249 (N_3249,In_691,In_3835);
or U3250 (N_3250,In_907,In_2032);
nand U3251 (N_3251,In_2475,In_2033);
nor U3252 (N_3252,In_2445,In_2212);
nand U3253 (N_3253,In_475,In_3310);
nor U3254 (N_3254,In_4938,In_827);
or U3255 (N_3255,In_3771,In_4242);
and U3256 (N_3256,In_4416,In_2207);
nand U3257 (N_3257,In_4017,In_1886);
and U3258 (N_3258,In_3599,In_2859);
nand U3259 (N_3259,In_3168,In_1822);
nand U3260 (N_3260,In_1397,In_3608);
nor U3261 (N_3261,In_3873,In_822);
and U3262 (N_3262,In_2425,In_189);
nand U3263 (N_3263,In_4907,In_4819);
nand U3264 (N_3264,In_3212,In_808);
nor U3265 (N_3265,In_722,In_4267);
xor U3266 (N_3266,In_2325,In_3317);
and U3267 (N_3267,In_1946,In_709);
or U3268 (N_3268,In_3796,In_4471);
xnor U3269 (N_3269,In_1182,In_2507);
nand U3270 (N_3270,In_728,In_3400);
or U3271 (N_3271,In_485,In_1151);
nor U3272 (N_3272,In_2854,In_2358);
nor U3273 (N_3273,In_2167,In_3274);
nor U3274 (N_3274,In_936,In_4847);
and U3275 (N_3275,In_1554,In_1736);
or U3276 (N_3276,In_2710,In_2772);
nand U3277 (N_3277,In_1928,In_3641);
or U3278 (N_3278,In_312,In_2971);
and U3279 (N_3279,In_2073,In_1662);
and U3280 (N_3280,In_4474,In_4060);
nand U3281 (N_3281,In_3523,In_3301);
xnor U3282 (N_3282,In_3400,In_2723);
nor U3283 (N_3283,In_2054,In_3822);
nor U3284 (N_3284,In_72,In_3111);
or U3285 (N_3285,In_894,In_1223);
xnor U3286 (N_3286,In_2234,In_2440);
nor U3287 (N_3287,In_1672,In_979);
nor U3288 (N_3288,In_811,In_4448);
xor U3289 (N_3289,In_4357,In_4566);
or U3290 (N_3290,In_1730,In_3141);
nor U3291 (N_3291,In_4348,In_2632);
and U3292 (N_3292,In_2329,In_1288);
nand U3293 (N_3293,In_2013,In_1555);
nand U3294 (N_3294,In_528,In_2239);
or U3295 (N_3295,In_1073,In_3101);
xor U3296 (N_3296,In_865,In_3083);
or U3297 (N_3297,In_3688,In_4312);
xnor U3298 (N_3298,In_2247,In_964);
nor U3299 (N_3299,In_2640,In_1696);
or U3300 (N_3300,In_1784,In_4188);
or U3301 (N_3301,In_465,In_2646);
nand U3302 (N_3302,In_4987,In_1185);
or U3303 (N_3303,In_3371,In_3071);
and U3304 (N_3304,In_2418,In_1381);
nand U3305 (N_3305,In_1941,In_639);
nand U3306 (N_3306,In_1775,In_1295);
nand U3307 (N_3307,In_574,In_921);
or U3308 (N_3308,In_820,In_1716);
nor U3309 (N_3309,In_2912,In_1306);
nand U3310 (N_3310,In_3341,In_2281);
nor U3311 (N_3311,In_2625,In_3973);
and U3312 (N_3312,In_1328,In_1098);
and U3313 (N_3313,In_3939,In_4180);
and U3314 (N_3314,In_449,In_236);
or U3315 (N_3315,In_1963,In_2386);
and U3316 (N_3316,In_1692,In_855);
nor U3317 (N_3317,In_3757,In_742);
nor U3318 (N_3318,In_4433,In_3209);
and U3319 (N_3319,In_667,In_840);
nand U3320 (N_3320,In_4447,In_4182);
and U3321 (N_3321,In_1950,In_3321);
and U3322 (N_3322,In_2792,In_70);
nand U3323 (N_3323,In_2606,In_408);
nand U3324 (N_3324,In_2416,In_256);
and U3325 (N_3325,In_760,In_3571);
nor U3326 (N_3326,In_3968,In_2316);
and U3327 (N_3327,In_1945,In_1593);
and U3328 (N_3328,In_2899,In_4372);
and U3329 (N_3329,In_1782,In_3679);
xor U3330 (N_3330,In_2950,In_4160);
nand U3331 (N_3331,In_888,In_3021);
nand U3332 (N_3332,In_1618,In_2549);
nand U3333 (N_3333,In_2608,In_1);
and U3334 (N_3334,In_2233,In_3847);
nand U3335 (N_3335,In_4629,In_153);
and U3336 (N_3336,In_925,In_2374);
nand U3337 (N_3337,In_3356,In_2775);
and U3338 (N_3338,In_4908,In_4688);
nor U3339 (N_3339,In_4772,In_2410);
nor U3340 (N_3340,In_44,In_4227);
or U3341 (N_3341,In_4322,In_546);
xnor U3342 (N_3342,In_2965,In_3335);
nand U3343 (N_3343,In_4881,In_4639);
and U3344 (N_3344,In_1208,In_1283);
nor U3345 (N_3345,In_4710,In_632);
xnor U3346 (N_3346,In_2200,In_4284);
nor U3347 (N_3347,In_3395,In_2661);
nand U3348 (N_3348,In_2716,In_4971);
nor U3349 (N_3349,In_1094,In_4300);
nor U3350 (N_3350,In_2235,In_2250);
and U3351 (N_3351,In_1663,In_3758);
nor U3352 (N_3352,In_3390,In_2132);
nor U3353 (N_3353,In_4706,In_4933);
and U3354 (N_3354,In_2545,In_4279);
or U3355 (N_3355,In_2069,In_1850);
or U3356 (N_3356,In_2393,In_320);
and U3357 (N_3357,In_4262,In_3345);
and U3358 (N_3358,In_1387,In_2076);
nand U3359 (N_3359,In_3041,In_645);
and U3360 (N_3360,In_1645,In_2810);
or U3361 (N_3361,In_90,In_506);
nand U3362 (N_3362,In_2414,In_1395);
and U3363 (N_3363,In_4334,In_4785);
and U3364 (N_3364,In_702,In_802);
xor U3365 (N_3365,In_128,In_3076);
nand U3366 (N_3366,In_4817,In_3398);
xor U3367 (N_3367,In_4987,In_183);
or U3368 (N_3368,In_4525,In_252);
or U3369 (N_3369,In_1849,In_1517);
nand U3370 (N_3370,In_4588,In_3328);
nand U3371 (N_3371,In_1986,In_4119);
and U3372 (N_3372,In_2832,In_4677);
and U3373 (N_3373,In_1462,In_1697);
or U3374 (N_3374,In_2385,In_338);
nor U3375 (N_3375,In_4991,In_4215);
or U3376 (N_3376,In_3706,In_465);
and U3377 (N_3377,In_1245,In_4984);
or U3378 (N_3378,In_175,In_3394);
or U3379 (N_3379,In_2264,In_854);
nor U3380 (N_3380,In_4578,In_4230);
xor U3381 (N_3381,In_1335,In_4972);
or U3382 (N_3382,In_4111,In_4377);
nand U3383 (N_3383,In_1999,In_1904);
or U3384 (N_3384,In_3920,In_3211);
nand U3385 (N_3385,In_2366,In_265);
xnor U3386 (N_3386,In_3103,In_1461);
nor U3387 (N_3387,In_3773,In_3022);
nor U3388 (N_3388,In_599,In_229);
and U3389 (N_3389,In_2843,In_685);
nand U3390 (N_3390,In_4201,In_399);
xnor U3391 (N_3391,In_1440,In_546);
and U3392 (N_3392,In_2421,In_3484);
or U3393 (N_3393,In_1798,In_1173);
nor U3394 (N_3394,In_3085,In_206);
nor U3395 (N_3395,In_317,In_4609);
xor U3396 (N_3396,In_191,In_2473);
xor U3397 (N_3397,In_4891,In_4254);
xnor U3398 (N_3398,In_420,In_239);
xnor U3399 (N_3399,In_4597,In_4318);
nor U3400 (N_3400,In_51,In_2812);
nor U3401 (N_3401,In_2089,In_3149);
or U3402 (N_3402,In_4185,In_1737);
nor U3403 (N_3403,In_187,In_4178);
nand U3404 (N_3404,In_2598,In_2185);
and U3405 (N_3405,In_861,In_2448);
nand U3406 (N_3406,In_3148,In_763);
nand U3407 (N_3407,In_3605,In_3781);
nor U3408 (N_3408,In_1113,In_2443);
nand U3409 (N_3409,In_2805,In_159);
or U3410 (N_3410,In_3706,In_4480);
or U3411 (N_3411,In_1443,In_1190);
or U3412 (N_3412,In_3150,In_2617);
nand U3413 (N_3413,In_1241,In_2831);
nor U3414 (N_3414,In_1879,In_1105);
nand U3415 (N_3415,In_1437,In_1212);
or U3416 (N_3416,In_177,In_2667);
and U3417 (N_3417,In_4114,In_489);
nor U3418 (N_3418,In_2297,In_2423);
nor U3419 (N_3419,In_3346,In_4956);
nor U3420 (N_3420,In_291,In_3378);
and U3421 (N_3421,In_4169,In_3390);
nor U3422 (N_3422,In_3108,In_4404);
or U3423 (N_3423,In_4889,In_777);
nor U3424 (N_3424,In_517,In_885);
nand U3425 (N_3425,In_250,In_1298);
xnor U3426 (N_3426,In_106,In_1782);
or U3427 (N_3427,In_4394,In_1044);
nand U3428 (N_3428,In_3733,In_2416);
nor U3429 (N_3429,In_121,In_4927);
nor U3430 (N_3430,In_4283,In_4196);
nand U3431 (N_3431,In_929,In_2828);
nand U3432 (N_3432,In_1668,In_4285);
nand U3433 (N_3433,In_2920,In_1427);
and U3434 (N_3434,In_3677,In_3097);
nor U3435 (N_3435,In_504,In_881);
and U3436 (N_3436,In_3984,In_652);
or U3437 (N_3437,In_1798,In_3226);
xnor U3438 (N_3438,In_353,In_31);
and U3439 (N_3439,In_1329,In_3787);
nand U3440 (N_3440,In_3639,In_4122);
or U3441 (N_3441,In_2878,In_1596);
or U3442 (N_3442,In_4573,In_3500);
nor U3443 (N_3443,In_3723,In_1633);
or U3444 (N_3444,In_4611,In_1743);
nor U3445 (N_3445,In_4454,In_4953);
and U3446 (N_3446,In_4232,In_125);
and U3447 (N_3447,In_4099,In_4741);
nand U3448 (N_3448,In_3946,In_1150);
nand U3449 (N_3449,In_691,In_4780);
nor U3450 (N_3450,In_1556,In_2188);
xor U3451 (N_3451,In_431,In_2143);
and U3452 (N_3452,In_2110,In_3072);
and U3453 (N_3453,In_528,In_4328);
nand U3454 (N_3454,In_1977,In_464);
or U3455 (N_3455,In_4356,In_136);
and U3456 (N_3456,In_2678,In_1533);
or U3457 (N_3457,In_2417,In_3920);
xnor U3458 (N_3458,In_1843,In_3694);
and U3459 (N_3459,In_1263,In_4817);
nand U3460 (N_3460,In_1002,In_4275);
and U3461 (N_3461,In_4926,In_204);
and U3462 (N_3462,In_4743,In_1788);
and U3463 (N_3463,In_1799,In_4848);
nand U3464 (N_3464,In_2535,In_201);
and U3465 (N_3465,In_3777,In_4577);
and U3466 (N_3466,In_2685,In_4342);
or U3467 (N_3467,In_2537,In_2674);
and U3468 (N_3468,In_625,In_3151);
and U3469 (N_3469,In_2490,In_3069);
nor U3470 (N_3470,In_4723,In_20);
xnor U3471 (N_3471,In_250,In_2511);
nor U3472 (N_3472,In_1050,In_2397);
nand U3473 (N_3473,In_1511,In_766);
xor U3474 (N_3474,In_1189,In_3036);
and U3475 (N_3475,In_3043,In_4556);
or U3476 (N_3476,In_3338,In_2110);
or U3477 (N_3477,In_3136,In_1082);
nand U3478 (N_3478,In_814,In_2432);
and U3479 (N_3479,In_4124,In_3684);
nand U3480 (N_3480,In_2204,In_4176);
or U3481 (N_3481,In_1287,In_4372);
nor U3482 (N_3482,In_1431,In_49);
nand U3483 (N_3483,In_3003,In_4507);
or U3484 (N_3484,In_4222,In_4124);
nor U3485 (N_3485,In_3368,In_1252);
nor U3486 (N_3486,In_168,In_92);
nand U3487 (N_3487,In_1946,In_4250);
nor U3488 (N_3488,In_3936,In_3400);
nor U3489 (N_3489,In_3885,In_4882);
nand U3490 (N_3490,In_3428,In_269);
nand U3491 (N_3491,In_4945,In_4677);
nand U3492 (N_3492,In_2056,In_137);
xor U3493 (N_3493,In_4375,In_3648);
xor U3494 (N_3494,In_4985,In_646);
nand U3495 (N_3495,In_4062,In_2415);
and U3496 (N_3496,In_1374,In_590);
or U3497 (N_3497,In_2529,In_4027);
nand U3498 (N_3498,In_4734,In_2536);
or U3499 (N_3499,In_31,In_3000);
nor U3500 (N_3500,In_2188,In_4796);
and U3501 (N_3501,In_73,In_1667);
nand U3502 (N_3502,In_1263,In_3734);
and U3503 (N_3503,In_4760,In_2641);
or U3504 (N_3504,In_797,In_2746);
nand U3505 (N_3505,In_3574,In_2255);
and U3506 (N_3506,In_2818,In_2619);
or U3507 (N_3507,In_1711,In_3369);
nor U3508 (N_3508,In_4482,In_3854);
or U3509 (N_3509,In_433,In_1384);
and U3510 (N_3510,In_58,In_2696);
nor U3511 (N_3511,In_3528,In_4100);
nand U3512 (N_3512,In_4126,In_2425);
or U3513 (N_3513,In_1142,In_1046);
nand U3514 (N_3514,In_409,In_1608);
and U3515 (N_3515,In_1579,In_2157);
xnor U3516 (N_3516,In_1041,In_4781);
and U3517 (N_3517,In_4842,In_1323);
or U3518 (N_3518,In_791,In_4105);
or U3519 (N_3519,In_865,In_2217);
or U3520 (N_3520,In_3037,In_253);
or U3521 (N_3521,In_2277,In_2245);
and U3522 (N_3522,In_3130,In_1872);
and U3523 (N_3523,In_3483,In_3148);
xor U3524 (N_3524,In_83,In_3975);
and U3525 (N_3525,In_3289,In_1034);
nand U3526 (N_3526,In_2519,In_3534);
nor U3527 (N_3527,In_4709,In_2046);
and U3528 (N_3528,In_3973,In_4953);
or U3529 (N_3529,In_847,In_4664);
and U3530 (N_3530,In_1338,In_2761);
and U3531 (N_3531,In_2495,In_1899);
xor U3532 (N_3532,In_4334,In_1175);
or U3533 (N_3533,In_247,In_1635);
nand U3534 (N_3534,In_1803,In_3168);
nand U3535 (N_3535,In_3334,In_275);
or U3536 (N_3536,In_1398,In_2524);
nor U3537 (N_3537,In_3091,In_4594);
xnor U3538 (N_3538,In_719,In_1025);
nor U3539 (N_3539,In_1032,In_230);
nor U3540 (N_3540,In_4780,In_3424);
or U3541 (N_3541,In_1535,In_29);
nor U3542 (N_3542,In_801,In_774);
or U3543 (N_3543,In_3599,In_704);
and U3544 (N_3544,In_143,In_2888);
xor U3545 (N_3545,In_4446,In_1412);
nand U3546 (N_3546,In_4092,In_3671);
or U3547 (N_3547,In_4428,In_1950);
xnor U3548 (N_3548,In_1557,In_3283);
and U3549 (N_3549,In_3890,In_2029);
nor U3550 (N_3550,In_2181,In_4958);
and U3551 (N_3551,In_149,In_1312);
and U3552 (N_3552,In_2123,In_4839);
nor U3553 (N_3553,In_299,In_1595);
nand U3554 (N_3554,In_1693,In_2768);
xnor U3555 (N_3555,In_768,In_3266);
nand U3556 (N_3556,In_3609,In_4357);
or U3557 (N_3557,In_1310,In_1593);
or U3558 (N_3558,In_93,In_1601);
or U3559 (N_3559,In_2741,In_4428);
nor U3560 (N_3560,In_4787,In_4630);
nand U3561 (N_3561,In_2214,In_738);
and U3562 (N_3562,In_3233,In_4769);
or U3563 (N_3563,In_379,In_871);
nand U3564 (N_3564,In_1997,In_2459);
or U3565 (N_3565,In_2268,In_3806);
or U3566 (N_3566,In_4052,In_1325);
and U3567 (N_3567,In_4517,In_1891);
nand U3568 (N_3568,In_2221,In_3864);
nand U3569 (N_3569,In_3877,In_2167);
xnor U3570 (N_3570,In_4364,In_4664);
nor U3571 (N_3571,In_1809,In_1850);
nand U3572 (N_3572,In_792,In_4471);
nor U3573 (N_3573,In_2536,In_4083);
and U3574 (N_3574,In_4577,In_2972);
and U3575 (N_3575,In_65,In_3070);
nand U3576 (N_3576,In_334,In_3566);
or U3577 (N_3577,In_483,In_319);
and U3578 (N_3578,In_4086,In_4403);
and U3579 (N_3579,In_1996,In_1333);
or U3580 (N_3580,In_4278,In_3864);
nand U3581 (N_3581,In_1724,In_2240);
and U3582 (N_3582,In_4357,In_343);
nand U3583 (N_3583,In_15,In_351);
or U3584 (N_3584,In_4310,In_2410);
nor U3585 (N_3585,In_772,In_2636);
and U3586 (N_3586,In_3922,In_156);
and U3587 (N_3587,In_3002,In_601);
nand U3588 (N_3588,In_1520,In_774);
and U3589 (N_3589,In_621,In_4915);
and U3590 (N_3590,In_3421,In_2386);
nor U3591 (N_3591,In_4747,In_1526);
nor U3592 (N_3592,In_4408,In_854);
and U3593 (N_3593,In_1582,In_1818);
nand U3594 (N_3594,In_2965,In_2480);
nor U3595 (N_3595,In_3525,In_2974);
nand U3596 (N_3596,In_4914,In_2305);
nor U3597 (N_3597,In_3187,In_2642);
or U3598 (N_3598,In_1766,In_2229);
nor U3599 (N_3599,In_4461,In_3117);
or U3600 (N_3600,In_4511,In_1360);
and U3601 (N_3601,In_1557,In_4757);
or U3602 (N_3602,In_3679,In_1830);
nand U3603 (N_3603,In_2343,In_3254);
or U3604 (N_3604,In_2321,In_2852);
or U3605 (N_3605,In_973,In_3748);
or U3606 (N_3606,In_288,In_1640);
nand U3607 (N_3607,In_3022,In_4654);
and U3608 (N_3608,In_1453,In_495);
and U3609 (N_3609,In_4864,In_1238);
or U3610 (N_3610,In_2789,In_670);
nand U3611 (N_3611,In_1129,In_3879);
or U3612 (N_3612,In_3023,In_4504);
nand U3613 (N_3613,In_3483,In_3485);
and U3614 (N_3614,In_1257,In_537);
nor U3615 (N_3615,In_4322,In_355);
nand U3616 (N_3616,In_974,In_167);
and U3617 (N_3617,In_3107,In_3147);
or U3618 (N_3618,In_4080,In_384);
nor U3619 (N_3619,In_4232,In_3502);
nand U3620 (N_3620,In_515,In_1175);
and U3621 (N_3621,In_3994,In_2615);
or U3622 (N_3622,In_4918,In_3773);
and U3623 (N_3623,In_3135,In_574);
or U3624 (N_3624,In_931,In_3388);
nand U3625 (N_3625,In_4280,In_2566);
or U3626 (N_3626,In_2420,In_686);
and U3627 (N_3627,In_742,In_4206);
nor U3628 (N_3628,In_4933,In_706);
or U3629 (N_3629,In_2570,In_3087);
nand U3630 (N_3630,In_3148,In_153);
xor U3631 (N_3631,In_3081,In_4471);
xnor U3632 (N_3632,In_2577,In_3898);
nand U3633 (N_3633,In_152,In_3539);
or U3634 (N_3634,In_1151,In_3158);
or U3635 (N_3635,In_1797,In_3404);
or U3636 (N_3636,In_3897,In_3031);
and U3637 (N_3637,In_2608,In_1440);
nand U3638 (N_3638,In_1455,In_3797);
nand U3639 (N_3639,In_286,In_644);
nor U3640 (N_3640,In_2078,In_1860);
or U3641 (N_3641,In_628,In_548);
or U3642 (N_3642,In_3551,In_3502);
nand U3643 (N_3643,In_2157,In_1459);
nor U3644 (N_3644,In_2461,In_919);
nand U3645 (N_3645,In_662,In_2374);
nor U3646 (N_3646,In_3586,In_1043);
or U3647 (N_3647,In_2410,In_4513);
nand U3648 (N_3648,In_3971,In_1989);
and U3649 (N_3649,In_1173,In_4371);
and U3650 (N_3650,In_2349,In_2290);
and U3651 (N_3651,In_3455,In_1630);
xnor U3652 (N_3652,In_4975,In_200);
xnor U3653 (N_3653,In_3261,In_645);
nand U3654 (N_3654,In_4514,In_4813);
nand U3655 (N_3655,In_1857,In_3637);
or U3656 (N_3656,In_51,In_4282);
nand U3657 (N_3657,In_4209,In_492);
nand U3658 (N_3658,In_4125,In_1906);
or U3659 (N_3659,In_3289,In_1231);
or U3660 (N_3660,In_1113,In_4703);
nor U3661 (N_3661,In_1770,In_2327);
and U3662 (N_3662,In_2462,In_3555);
and U3663 (N_3663,In_4209,In_2129);
or U3664 (N_3664,In_3676,In_3387);
or U3665 (N_3665,In_3867,In_1498);
nor U3666 (N_3666,In_2006,In_1442);
or U3667 (N_3667,In_4270,In_427);
or U3668 (N_3668,In_4774,In_33);
or U3669 (N_3669,In_1583,In_4326);
or U3670 (N_3670,In_2723,In_3936);
and U3671 (N_3671,In_3285,In_3112);
xnor U3672 (N_3672,In_2186,In_3580);
nand U3673 (N_3673,In_1736,In_2271);
nand U3674 (N_3674,In_3422,In_2761);
and U3675 (N_3675,In_1202,In_596);
or U3676 (N_3676,In_3814,In_2196);
xor U3677 (N_3677,In_3318,In_2934);
or U3678 (N_3678,In_1905,In_2999);
or U3679 (N_3679,In_3932,In_2092);
and U3680 (N_3680,In_4694,In_1787);
or U3681 (N_3681,In_935,In_2534);
nand U3682 (N_3682,In_327,In_4236);
nand U3683 (N_3683,In_1458,In_4611);
or U3684 (N_3684,In_2621,In_1721);
nand U3685 (N_3685,In_2944,In_4476);
and U3686 (N_3686,In_182,In_3467);
nand U3687 (N_3687,In_1227,In_3434);
xnor U3688 (N_3688,In_2324,In_1673);
or U3689 (N_3689,In_3832,In_339);
nor U3690 (N_3690,In_1396,In_2075);
and U3691 (N_3691,In_3228,In_4588);
and U3692 (N_3692,In_4564,In_349);
xor U3693 (N_3693,In_2478,In_3389);
nor U3694 (N_3694,In_3736,In_969);
and U3695 (N_3695,In_2730,In_4560);
nand U3696 (N_3696,In_3014,In_2892);
and U3697 (N_3697,In_4205,In_3142);
or U3698 (N_3698,In_4360,In_4613);
nand U3699 (N_3699,In_2625,In_2435);
nand U3700 (N_3700,In_3997,In_3710);
xnor U3701 (N_3701,In_2623,In_1026);
nand U3702 (N_3702,In_1196,In_730);
and U3703 (N_3703,In_3452,In_3755);
nand U3704 (N_3704,In_3601,In_1424);
and U3705 (N_3705,In_3477,In_1736);
nor U3706 (N_3706,In_3118,In_3065);
nand U3707 (N_3707,In_748,In_557);
or U3708 (N_3708,In_795,In_3769);
and U3709 (N_3709,In_593,In_2352);
or U3710 (N_3710,In_3572,In_2096);
nand U3711 (N_3711,In_800,In_364);
and U3712 (N_3712,In_1229,In_3401);
nor U3713 (N_3713,In_460,In_974);
or U3714 (N_3714,In_2637,In_3351);
nand U3715 (N_3715,In_3549,In_360);
or U3716 (N_3716,In_2618,In_2317);
and U3717 (N_3717,In_4990,In_2768);
nand U3718 (N_3718,In_36,In_4220);
nor U3719 (N_3719,In_136,In_4370);
nor U3720 (N_3720,In_2895,In_2235);
nor U3721 (N_3721,In_3043,In_4302);
nor U3722 (N_3722,In_1247,In_3485);
xnor U3723 (N_3723,In_2019,In_4840);
and U3724 (N_3724,In_3516,In_3847);
nor U3725 (N_3725,In_3392,In_3840);
and U3726 (N_3726,In_3502,In_1640);
or U3727 (N_3727,In_2537,In_2456);
nand U3728 (N_3728,In_2664,In_4867);
nor U3729 (N_3729,In_3794,In_1073);
xnor U3730 (N_3730,In_331,In_2158);
or U3731 (N_3731,In_2981,In_2755);
nand U3732 (N_3732,In_4151,In_548);
nand U3733 (N_3733,In_182,In_479);
or U3734 (N_3734,In_2220,In_2839);
and U3735 (N_3735,In_3752,In_1028);
nand U3736 (N_3736,In_258,In_3107);
nor U3737 (N_3737,In_1922,In_2090);
or U3738 (N_3738,In_1452,In_12);
and U3739 (N_3739,In_3321,In_4090);
nor U3740 (N_3740,In_1452,In_783);
nor U3741 (N_3741,In_3649,In_4687);
or U3742 (N_3742,In_2285,In_3688);
nand U3743 (N_3743,In_1699,In_387);
nand U3744 (N_3744,In_2990,In_89);
and U3745 (N_3745,In_2729,In_3080);
nor U3746 (N_3746,In_1537,In_4499);
nand U3747 (N_3747,In_1485,In_2237);
or U3748 (N_3748,In_4002,In_2877);
xor U3749 (N_3749,In_4434,In_1719);
nand U3750 (N_3750,In_1631,In_2985);
xor U3751 (N_3751,In_4355,In_1011);
xnor U3752 (N_3752,In_3915,In_4236);
or U3753 (N_3753,In_2341,In_4227);
nor U3754 (N_3754,In_2005,In_4981);
and U3755 (N_3755,In_3622,In_4390);
nor U3756 (N_3756,In_2689,In_2366);
xor U3757 (N_3757,In_3458,In_4329);
or U3758 (N_3758,In_1556,In_1778);
and U3759 (N_3759,In_826,In_637);
or U3760 (N_3760,In_1428,In_3043);
and U3761 (N_3761,In_4250,In_1525);
or U3762 (N_3762,In_233,In_3592);
and U3763 (N_3763,In_1683,In_3930);
and U3764 (N_3764,In_1855,In_1513);
nor U3765 (N_3765,In_163,In_4134);
nand U3766 (N_3766,In_1506,In_3967);
nand U3767 (N_3767,In_3656,In_1111);
and U3768 (N_3768,In_4878,In_2110);
nor U3769 (N_3769,In_4899,In_607);
nand U3770 (N_3770,In_2808,In_2300);
and U3771 (N_3771,In_138,In_2876);
or U3772 (N_3772,In_4515,In_2429);
nand U3773 (N_3773,In_1515,In_2367);
and U3774 (N_3774,In_4566,In_41);
or U3775 (N_3775,In_1706,In_4024);
or U3776 (N_3776,In_1346,In_4688);
nor U3777 (N_3777,In_831,In_1070);
xnor U3778 (N_3778,In_4740,In_3559);
or U3779 (N_3779,In_2258,In_4612);
nor U3780 (N_3780,In_3304,In_4625);
nor U3781 (N_3781,In_297,In_4517);
nor U3782 (N_3782,In_4617,In_3278);
nand U3783 (N_3783,In_1539,In_4086);
xor U3784 (N_3784,In_2064,In_971);
nor U3785 (N_3785,In_707,In_1550);
or U3786 (N_3786,In_492,In_2381);
and U3787 (N_3787,In_2586,In_2091);
nand U3788 (N_3788,In_2464,In_4792);
xor U3789 (N_3789,In_1744,In_3323);
or U3790 (N_3790,In_4471,In_3684);
and U3791 (N_3791,In_1741,In_4673);
xor U3792 (N_3792,In_1055,In_1520);
nand U3793 (N_3793,In_4886,In_1286);
xnor U3794 (N_3794,In_907,In_4450);
and U3795 (N_3795,In_3091,In_317);
and U3796 (N_3796,In_3491,In_1526);
nand U3797 (N_3797,In_3302,In_4263);
nor U3798 (N_3798,In_1321,In_3343);
xor U3799 (N_3799,In_4142,In_839);
or U3800 (N_3800,In_3646,In_961);
nor U3801 (N_3801,In_4498,In_4437);
xnor U3802 (N_3802,In_2047,In_3637);
nand U3803 (N_3803,In_130,In_2666);
or U3804 (N_3804,In_4815,In_264);
or U3805 (N_3805,In_1472,In_907);
nand U3806 (N_3806,In_4712,In_1472);
xor U3807 (N_3807,In_3784,In_2222);
nor U3808 (N_3808,In_2275,In_4783);
nand U3809 (N_3809,In_1530,In_207);
nand U3810 (N_3810,In_1133,In_1189);
and U3811 (N_3811,In_2329,In_4532);
and U3812 (N_3812,In_397,In_4685);
nand U3813 (N_3813,In_427,In_4632);
nand U3814 (N_3814,In_250,In_3945);
nand U3815 (N_3815,In_4342,In_3308);
nand U3816 (N_3816,In_3286,In_4714);
and U3817 (N_3817,In_3013,In_3999);
nand U3818 (N_3818,In_4403,In_2832);
or U3819 (N_3819,In_3220,In_2510);
nor U3820 (N_3820,In_922,In_4333);
nand U3821 (N_3821,In_2476,In_2399);
nor U3822 (N_3822,In_258,In_2097);
or U3823 (N_3823,In_3789,In_3036);
nand U3824 (N_3824,In_2121,In_4577);
and U3825 (N_3825,In_1274,In_1110);
and U3826 (N_3826,In_3529,In_70);
or U3827 (N_3827,In_4653,In_4389);
and U3828 (N_3828,In_3415,In_345);
and U3829 (N_3829,In_3679,In_149);
nor U3830 (N_3830,In_2241,In_2719);
xor U3831 (N_3831,In_3116,In_2168);
nand U3832 (N_3832,In_1747,In_2411);
or U3833 (N_3833,In_3730,In_1736);
and U3834 (N_3834,In_4793,In_1397);
nor U3835 (N_3835,In_232,In_221);
or U3836 (N_3836,In_3803,In_1886);
and U3837 (N_3837,In_3690,In_1104);
xor U3838 (N_3838,In_373,In_79);
or U3839 (N_3839,In_3204,In_2708);
nor U3840 (N_3840,In_4102,In_3534);
xnor U3841 (N_3841,In_2564,In_1000);
nand U3842 (N_3842,In_1267,In_1406);
or U3843 (N_3843,In_839,In_1623);
nand U3844 (N_3844,In_194,In_1601);
and U3845 (N_3845,In_929,In_4198);
or U3846 (N_3846,In_2013,In_736);
and U3847 (N_3847,In_1186,In_364);
and U3848 (N_3848,In_3818,In_3162);
nand U3849 (N_3849,In_1070,In_1855);
nand U3850 (N_3850,In_3376,In_2457);
or U3851 (N_3851,In_3335,In_3431);
and U3852 (N_3852,In_1218,In_4086);
xnor U3853 (N_3853,In_2671,In_3014);
nor U3854 (N_3854,In_520,In_1696);
or U3855 (N_3855,In_1090,In_2056);
and U3856 (N_3856,In_1508,In_1894);
or U3857 (N_3857,In_4949,In_3658);
or U3858 (N_3858,In_1345,In_2781);
or U3859 (N_3859,In_3158,In_1621);
nand U3860 (N_3860,In_1408,In_4072);
and U3861 (N_3861,In_1327,In_4377);
and U3862 (N_3862,In_1255,In_3661);
xor U3863 (N_3863,In_2763,In_2230);
nand U3864 (N_3864,In_3396,In_2738);
xnor U3865 (N_3865,In_1549,In_4970);
and U3866 (N_3866,In_4597,In_646);
nand U3867 (N_3867,In_439,In_240);
and U3868 (N_3868,In_2710,In_4669);
nor U3869 (N_3869,In_2348,In_2350);
xor U3870 (N_3870,In_1606,In_4150);
and U3871 (N_3871,In_4471,In_290);
nand U3872 (N_3872,In_1721,In_1325);
and U3873 (N_3873,In_257,In_325);
or U3874 (N_3874,In_3941,In_2510);
xnor U3875 (N_3875,In_2001,In_2248);
nor U3876 (N_3876,In_4283,In_870);
nand U3877 (N_3877,In_1316,In_4845);
nor U3878 (N_3878,In_738,In_4473);
nand U3879 (N_3879,In_2237,In_1912);
nand U3880 (N_3880,In_446,In_485);
xor U3881 (N_3881,In_3991,In_1319);
nand U3882 (N_3882,In_2033,In_4857);
nand U3883 (N_3883,In_4529,In_4024);
and U3884 (N_3884,In_4526,In_1713);
or U3885 (N_3885,In_2898,In_2995);
or U3886 (N_3886,In_2260,In_3678);
nand U3887 (N_3887,In_1606,In_3618);
nand U3888 (N_3888,In_779,In_3064);
nor U3889 (N_3889,In_4986,In_3708);
nand U3890 (N_3890,In_69,In_4215);
or U3891 (N_3891,In_4345,In_3866);
and U3892 (N_3892,In_3346,In_4768);
and U3893 (N_3893,In_2469,In_3548);
nor U3894 (N_3894,In_1097,In_883);
or U3895 (N_3895,In_1955,In_4265);
or U3896 (N_3896,In_1003,In_2857);
nor U3897 (N_3897,In_2483,In_204);
and U3898 (N_3898,In_3077,In_4901);
nor U3899 (N_3899,In_3003,In_4836);
xnor U3900 (N_3900,In_187,In_4918);
nor U3901 (N_3901,In_4526,In_2014);
nand U3902 (N_3902,In_537,In_2102);
and U3903 (N_3903,In_3704,In_1293);
nor U3904 (N_3904,In_3984,In_3851);
and U3905 (N_3905,In_1795,In_4594);
nand U3906 (N_3906,In_594,In_3548);
nor U3907 (N_3907,In_4469,In_3057);
or U3908 (N_3908,In_1529,In_4630);
xor U3909 (N_3909,In_1260,In_4506);
xnor U3910 (N_3910,In_3553,In_3628);
and U3911 (N_3911,In_4715,In_1239);
and U3912 (N_3912,In_1093,In_1393);
nor U3913 (N_3913,In_2626,In_2716);
and U3914 (N_3914,In_44,In_411);
and U3915 (N_3915,In_51,In_2663);
nor U3916 (N_3916,In_952,In_1548);
or U3917 (N_3917,In_2911,In_1724);
and U3918 (N_3918,In_2636,In_986);
or U3919 (N_3919,In_4771,In_3717);
and U3920 (N_3920,In_3552,In_191);
or U3921 (N_3921,In_3481,In_683);
nand U3922 (N_3922,In_321,In_896);
nor U3923 (N_3923,In_3020,In_874);
and U3924 (N_3924,In_4024,In_426);
and U3925 (N_3925,In_2066,In_495);
nand U3926 (N_3926,In_443,In_3690);
and U3927 (N_3927,In_2047,In_1246);
nor U3928 (N_3928,In_2706,In_1759);
or U3929 (N_3929,In_4152,In_1179);
nor U3930 (N_3930,In_2818,In_2961);
nand U3931 (N_3931,In_1325,In_395);
nor U3932 (N_3932,In_963,In_2668);
nand U3933 (N_3933,In_1827,In_1228);
nor U3934 (N_3934,In_4031,In_3178);
nor U3935 (N_3935,In_1890,In_448);
nand U3936 (N_3936,In_3980,In_2069);
nand U3937 (N_3937,In_2510,In_2297);
nor U3938 (N_3938,In_4357,In_1339);
or U3939 (N_3939,In_2106,In_2661);
or U3940 (N_3940,In_1651,In_3928);
nand U3941 (N_3941,In_2926,In_2664);
xnor U3942 (N_3942,In_4640,In_247);
or U3943 (N_3943,In_2580,In_2418);
and U3944 (N_3944,In_3629,In_1155);
nand U3945 (N_3945,In_1419,In_3497);
nor U3946 (N_3946,In_2335,In_4061);
nand U3947 (N_3947,In_4800,In_3546);
and U3948 (N_3948,In_3563,In_1521);
or U3949 (N_3949,In_4714,In_1848);
nor U3950 (N_3950,In_3423,In_3615);
or U3951 (N_3951,In_1196,In_3367);
and U3952 (N_3952,In_1445,In_405);
xor U3953 (N_3953,In_1931,In_721);
and U3954 (N_3954,In_4519,In_3258);
xor U3955 (N_3955,In_1911,In_3986);
xnor U3956 (N_3956,In_2237,In_2328);
or U3957 (N_3957,In_4751,In_3637);
nor U3958 (N_3958,In_2970,In_4837);
xnor U3959 (N_3959,In_1190,In_317);
nor U3960 (N_3960,In_779,In_1988);
or U3961 (N_3961,In_850,In_756);
nor U3962 (N_3962,In_2079,In_1755);
nand U3963 (N_3963,In_3879,In_2832);
nand U3964 (N_3964,In_3036,In_679);
or U3965 (N_3965,In_4317,In_4307);
or U3966 (N_3966,In_3516,In_2136);
xor U3967 (N_3967,In_469,In_4471);
and U3968 (N_3968,In_3615,In_2536);
or U3969 (N_3969,In_1167,In_2432);
nor U3970 (N_3970,In_175,In_280);
or U3971 (N_3971,In_3220,In_3599);
nor U3972 (N_3972,In_221,In_2358);
nor U3973 (N_3973,In_1683,In_4683);
xor U3974 (N_3974,In_4865,In_4882);
nor U3975 (N_3975,In_2620,In_3350);
and U3976 (N_3976,In_884,In_2420);
and U3977 (N_3977,In_2998,In_2930);
nor U3978 (N_3978,In_4739,In_2);
nor U3979 (N_3979,In_1141,In_4328);
nand U3980 (N_3980,In_3943,In_4525);
nor U3981 (N_3981,In_2783,In_2265);
nand U3982 (N_3982,In_528,In_3193);
and U3983 (N_3983,In_2355,In_3055);
nor U3984 (N_3984,In_819,In_2113);
and U3985 (N_3985,In_3739,In_4630);
nand U3986 (N_3986,In_4557,In_1080);
xor U3987 (N_3987,In_1242,In_145);
nor U3988 (N_3988,In_3571,In_4057);
nor U3989 (N_3989,In_828,In_2186);
nand U3990 (N_3990,In_2172,In_2747);
or U3991 (N_3991,In_1694,In_4794);
or U3992 (N_3992,In_3835,In_4147);
and U3993 (N_3993,In_3971,In_3594);
nor U3994 (N_3994,In_2278,In_2888);
and U3995 (N_3995,In_3867,In_947);
nand U3996 (N_3996,In_2347,In_4896);
xnor U3997 (N_3997,In_2528,In_264);
or U3998 (N_3998,In_2399,In_518);
or U3999 (N_3999,In_700,In_1667);
nor U4000 (N_4000,In_3675,In_1279);
and U4001 (N_4001,In_601,In_4611);
nor U4002 (N_4002,In_4422,In_4530);
and U4003 (N_4003,In_409,In_3695);
nor U4004 (N_4004,In_3820,In_31);
xor U4005 (N_4005,In_1970,In_4071);
nand U4006 (N_4006,In_2793,In_3869);
nor U4007 (N_4007,In_2270,In_1234);
nand U4008 (N_4008,In_39,In_4453);
xnor U4009 (N_4009,In_987,In_3018);
nor U4010 (N_4010,In_976,In_2127);
and U4011 (N_4011,In_4417,In_2755);
and U4012 (N_4012,In_1065,In_3448);
xnor U4013 (N_4013,In_4164,In_870);
nand U4014 (N_4014,In_1687,In_4474);
nor U4015 (N_4015,In_3927,In_3264);
nand U4016 (N_4016,In_4789,In_4042);
nor U4017 (N_4017,In_581,In_2365);
nand U4018 (N_4018,In_874,In_3140);
or U4019 (N_4019,In_2229,In_307);
nand U4020 (N_4020,In_3300,In_155);
or U4021 (N_4021,In_2367,In_2589);
or U4022 (N_4022,In_3783,In_106);
and U4023 (N_4023,In_296,In_1671);
xnor U4024 (N_4024,In_4974,In_4888);
or U4025 (N_4025,In_1738,In_581);
and U4026 (N_4026,In_2510,In_4702);
nand U4027 (N_4027,In_3848,In_2866);
xor U4028 (N_4028,In_4283,In_1557);
and U4029 (N_4029,In_161,In_2738);
nand U4030 (N_4030,In_1834,In_4404);
nor U4031 (N_4031,In_753,In_3304);
nor U4032 (N_4032,In_1100,In_529);
and U4033 (N_4033,In_4566,In_2500);
and U4034 (N_4034,In_607,In_4807);
nand U4035 (N_4035,In_1526,In_4104);
nand U4036 (N_4036,In_2548,In_4911);
or U4037 (N_4037,In_2810,In_2887);
nand U4038 (N_4038,In_333,In_3103);
or U4039 (N_4039,In_1082,In_2451);
or U4040 (N_4040,In_3571,In_1881);
or U4041 (N_4041,In_1721,In_2422);
and U4042 (N_4042,In_2347,In_1728);
and U4043 (N_4043,In_931,In_2333);
or U4044 (N_4044,In_2577,In_3713);
nor U4045 (N_4045,In_2525,In_4850);
or U4046 (N_4046,In_3068,In_981);
and U4047 (N_4047,In_2515,In_2982);
nor U4048 (N_4048,In_757,In_1196);
or U4049 (N_4049,In_4623,In_1787);
nor U4050 (N_4050,In_2026,In_4181);
and U4051 (N_4051,In_3164,In_125);
nand U4052 (N_4052,In_4735,In_370);
or U4053 (N_4053,In_2995,In_2831);
or U4054 (N_4054,In_2300,In_1305);
nor U4055 (N_4055,In_4237,In_115);
or U4056 (N_4056,In_4266,In_1204);
nor U4057 (N_4057,In_139,In_304);
nand U4058 (N_4058,In_3548,In_1279);
nand U4059 (N_4059,In_1105,In_4096);
nand U4060 (N_4060,In_1281,In_3190);
xnor U4061 (N_4061,In_1431,In_2245);
and U4062 (N_4062,In_576,In_848);
or U4063 (N_4063,In_2809,In_365);
nor U4064 (N_4064,In_1259,In_3789);
nor U4065 (N_4065,In_4803,In_250);
nor U4066 (N_4066,In_3986,In_3414);
nor U4067 (N_4067,In_1844,In_3312);
or U4068 (N_4068,In_2069,In_2625);
or U4069 (N_4069,In_928,In_2762);
nand U4070 (N_4070,In_288,In_3912);
nor U4071 (N_4071,In_4657,In_4274);
nand U4072 (N_4072,In_1406,In_3535);
nand U4073 (N_4073,In_176,In_4185);
xnor U4074 (N_4074,In_4627,In_3462);
and U4075 (N_4075,In_3793,In_2947);
nor U4076 (N_4076,In_4662,In_4149);
or U4077 (N_4077,In_1469,In_213);
nor U4078 (N_4078,In_2029,In_2275);
nand U4079 (N_4079,In_3858,In_1);
and U4080 (N_4080,In_4918,In_4429);
or U4081 (N_4081,In_3272,In_370);
nor U4082 (N_4082,In_1231,In_3086);
nor U4083 (N_4083,In_3366,In_4033);
or U4084 (N_4084,In_603,In_1447);
nor U4085 (N_4085,In_1059,In_4284);
and U4086 (N_4086,In_2248,In_3344);
nor U4087 (N_4087,In_3226,In_2429);
and U4088 (N_4088,In_2288,In_789);
nor U4089 (N_4089,In_2217,In_4478);
and U4090 (N_4090,In_4949,In_676);
and U4091 (N_4091,In_4132,In_1954);
and U4092 (N_4092,In_2139,In_3073);
and U4093 (N_4093,In_2798,In_4896);
nor U4094 (N_4094,In_3998,In_4117);
nor U4095 (N_4095,In_3217,In_2930);
nand U4096 (N_4096,In_743,In_3030);
xnor U4097 (N_4097,In_1018,In_255);
or U4098 (N_4098,In_3693,In_1611);
xor U4099 (N_4099,In_4250,In_2693);
or U4100 (N_4100,In_3677,In_1861);
nor U4101 (N_4101,In_4524,In_4848);
nor U4102 (N_4102,In_3675,In_3508);
nor U4103 (N_4103,In_1120,In_4583);
and U4104 (N_4104,In_4116,In_733);
nor U4105 (N_4105,In_2855,In_4356);
nand U4106 (N_4106,In_967,In_3678);
and U4107 (N_4107,In_2399,In_314);
nor U4108 (N_4108,In_4724,In_2080);
and U4109 (N_4109,In_1757,In_1804);
nor U4110 (N_4110,In_1246,In_4053);
or U4111 (N_4111,In_1445,In_133);
nor U4112 (N_4112,In_3826,In_1747);
or U4113 (N_4113,In_1096,In_4680);
nand U4114 (N_4114,In_2126,In_3551);
and U4115 (N_4115,In_4360,In_1219);
nor U4116 (N_4116,In_3178,In_2678);
or U4117 (N_4117,In_1383,In_2300);
nand U4118 (N_4118,In_3057,In_3448);
xor U4119 (N_4119,In_4832,In_2743);
and U4120 (N_4120,In_2628,In_384);
or U4121 (N_4121,In_3607,In_3318);
nand U4122 (N_4122,In_2020,In_3010);
and U4123 (N_4123,In_4746,In_910);
or U4124 (N_4124,In_2778,In_256);
or U4125 (N_4125,In_3275,In_4975);
and U4126 (N_4126,In_1408,In_322);
nand U4127 (N_4127,In_1639,In_1814);
and U4128 (N_4128,In_4168,In_3506);
and U4129 (N_4129,In_273,In_2052);
xor U4130 (N_4130,In_1934,In_3223);
nand U4131 (N_4131,In_3395,In_2753);
or U4132 (N_4132,In_694,In_3458);
nor U4133 (N_4133,In_1656,In_295);
or U4134 (N_4134,In_754,In_243);
or U4135 (N_4135,In_3089,In_2244);
nand U4136 (N_4136,In_3950,In_4324);
and U4137 (N_4137,In_1749,In_919);
xor U4138 (N_4138,In_45,In_2744);
xnor U4139 (N_4139,In_3157,In_2214);
or U4140 (N_4140,In_1154,In_2400);
and U4141 (N_4141,In_4416,In_4290);
nor U4142 (N_4142,In_4191,In_898);
and U4143 (N_4143,In_3684,In_1777);
nand U4144 (N_4144,In_896,In_2374);
and U4145 (N_4145,In_4875,In_2598);
nand U4146 (N_4146,In_1579,In_2829);
xor U4147 (N_4147,In_2460,In_1626);
nand U4148 (N_4148,In_3234,In_800);
xor U4149 (N_4149,In_1416,In_2137);
and U4150 (N_4150,In_4864,In_3629);
nor U4151 (N_4151,In_1529,In_2619);
and U4152 (N_4152,In_135,In_2037);
xnor U4153 (N_4153,In_2424,In_707);
nand U4154 (N_4154,In_4617,In_1568);
or U4155 (N_4155,In_247,In_2189);
nand U4156 (N_4156,In_2384,In_922);
xnor U4157 (N_4157,In_4353,In_4514);
or U4158 (N_4158,In_977,In_4366);
nor U4159 (N_4159,In_2602,In_538);
nor U4160 (N_4160,In_362,In_666);
and U4161 (N_4161,In_4149,In_2320);
nand U4162 (N_4162,In_4936,In_1531);
xnor U4163 (N_4163,In_253,In_1091);
nand U4164 (N_4164,In_3834,In_553);
xor U4165 (N_4165,In_1999,In_2373);
nand U4166 (N_4166,In_3338,In_4242);
and U4167 (N_4167,In_51,In_457);
and U4168 (N_4168,In_2227,In_4389);
nand U4169 (N_4169,In_1309,In_3797);
xnor U4170 (N_4170,In_3325,In_1116);
xnor U4171 (N_4171,In_1028,In_2825);
or U4172 (N_4172,In_2040,In_3708);
nand U4173 (N_4173,In_2317,In_3044);
nand U4174 (N_4174,In_3457,In_2948);
xnor U4175 (N_4175,In_88,In_252);
and U4176 (N_4176,In_234,In_2992);
nand U4177 (N_4177,In_1047,In_1298);
xnor U4178 (N_4178,In_134,In_1281);
or U4179 (N_4179,In_1045,In_2344);
and U4180 (N_4180,In_2277,In_2492);
nand U4181 (N_4181,In_778,In_2946);
or U4182 (N_4182,In_3387,In_1938);
nand U4183 (N_4183,In_1529,In_1111);
nor U4184 (N_4184,In_3578,In_585);
nand U4185 (N_4185,In_1086,In_503);
and U4186 (N_4186,In_888,In_3099);
nor U4187 (N_4187,In_908,In_4673);
and U4188 (N_4188,In_3839,In_2183);
or U4189 (N_4189,In_1189,In_4902);
nor U4190 (N_4190,In_1530,In_2754);
and U4191 (N_4191,In_2901,In_4207);
and U4192 (N_4192,In_2896,In_3449);
and U4193 (N_4193,In_4243,In_2310);
and U4194 (N_4194,In_4157,In_1469);
nand U4195 (N_4195,In_4147,In_854);
nand U4196 (N_4196,In_3425,In_3322);
and U4197 (N_4197,In_2218,In_3085);
and U4198 (N_4198,In_840,In_3603);
xor U4199 (N_4199,In_1672,In_4232);
nand U4200 (N_4200,In_2538,In_2423);
nand U4201 (N_4201,In_1782,In_386);
or U4202 (N_4202,In_3548,In_4722);
or U4203 (N_4203,In_3990,In_1608);
and U4204 (N_4204,In_4219,In_2682);
nand U4205 (N_4205,In_2913,In_3367);
or U4206 (N_4206,In_249,In_3380);
or U4207 (N_4207,In_3366,In_2102);
or U4208 (N_4208,In_31,In_3453);
nand U4209 (N_4209,In_3473,In_1243);
xor U4210 (N_4210,In_2617,In_1895);
nor U4211 (N_4211,In_3991,In_1620);
and U4212 (N_4212,In_600,In_1299);
nand U4213 (N_4213,In_722,In_910);
xor U4214 (N_4214,In_4084,In_2686);
or U4215 (N_4215,In_167,In_3883);
nor U4216 (N_4216,In_1792,In_1773);
and U4217 (N_4217,In_2588,In_3889);
xor U4218 (N_4218,In_3984,In_4881);
nand U4219 (N_4219,In_3446,In_2797);
or U4220 (N_4220,In_3271,In_2995);
xor U4221 (N_4221,In_1877,In_1996);
nand U4222 (N_4222,In_4707,In_4467);
xor U4223 (N_4223,In_4183,In_2825);
xor U4224 (N_4224,In_2917,In_3622);
nor U4225 (N_4225,In_1295,In_749);
or U4226 (N_4226,In_4045,In_319);
nand U4227 (N_4227,In_3438,In_1104);
and U4228 (N_4228,In_4493,In_4189);
and U4229 (N_4229,In_4181,In_3350);
or U4230 (N_4230,In_795,In_1790);
and U4231 (N_4231,In_3096,In_745);
nor U4232 (N_4232,In_3870,In_4365);
and U4233 (N_4233,In_136,In_848);
or U4234 (N_4234,In_898,In_430);
nor U4235 (N_4235,In_795,In_1794);
nor U4236 (N_4236,In_804,In_3478);
and U4237 (N_4237,In_3470,In_1484);
and U4238 (N_4238,In_2414,In_4478);
and U4239 (N_4239,In_1136,In_4861);
xnor U4240 (N_4240,In_3015,In_3627);
nand U4241 (N_4241,In_4375,In_851);
or U4242 (N_4242,In_2213,In_1633);
or U4243 (N_4243,In_4220,In_2250);
nor U4244 (N_4244,In_1678,In_757);
xor U4245 (N_4245,In_411,In_999);
nor U4246 (N_4246,In_3309,In_4365);
nand U4247 (N_4247,In_4672,In_1107);
nand U4248 (N_4248,In_3219,In_3566);
or U4249 (N_4249,In_224,In_4936);
or U4250 (N_4250,In_1020,In_2587);
or U4251 (N_4251,In_3677,In_431);
and U4252 (N_4252,In_2210,In_2268);
or U4253 (N_4253,In_4295,In_4708);
nor U4254 (N_4254,In_941,In_2825);
nand U4255 (N_4255,In_4346,In_3272);
or U4256 (N_4256,In_2324,In_3546);
nand U4257 (N_4257,In_1183,In_4347);
or U4258 (N_4258,In_2546,In_1744);
nor U4259 (N_4259,In_2302,In_3826);
nand U4260 (N_4260,In_2509,In_1853);
and U4261 (N_4261,In_4662,In_4932);
nand U4262 (N_4262,In_1509,In_1542);
xnor U4263 (N_4263,In_3247,In_4456);
xor U4264 (N_4264,In_4013,In_3138);
nor U4265 (N_4265,In_3232,In_1469);
nor U4266 (N_4266,In_4416,In_94);
nand U4267 (N_4267,In_3486,In_1847);
nor U4268 (N_4268,In_3480,In_3065);
or U4269 (N_4269,In_2060,In_302);
nand U4270 (N_4270,In_1732,In_1491);
or U4271 (N_4271,In_4994,In_4007);
and U4272 (N_4272,In_2181,In_2178);
nand U4273 (N_4273,In_4058,In_1434);
and U4274 (N_4274,In_1593,In_1901);
nor U4275 (N_4275,In_4730,In_2264);
nor U4276 (N_4276,In_4831,In_943);
nand U4277 (N_4277,In_2338,In_299);
nor U4278 (N_4278,In_3754,In_3414);
and U4279 (N_4279,In_903,In_2622);
and U4280 (N_4280,In_2802,In_3898);
nor U4281 (N_4281,In_2628,In_3801);
xnor U4282 (N_4282,In_4159,In_4874);
nand U4283 (N_4283,In_2320,In_4590);
or U4284 (N_4284,In_4367,In_2842);
xnor U4285 (N_4285,In_1337,In_4399);
nor U4286 (N_4286,In_2107,In_3345);
nor U4287 (N_4287,In_4980,In_4854);
or U4288 (N_4288,In_3135,In_2167);
nand U4289 (N_4289,In_3330,In_3222);
nor U4290 (N_4290,In_4039,In_3660);
nand U4291 (N_4291,In_749,In_1861);
or U4292 (N_4292,In_1656,In_2057);
nor U4293 (N_4293,In_3415,In_21);
and U4294 (N_4294,In_1503,In_1656);
or U4295 (N_4295,In_4598,In_3486);
nor U4296 (N_4296,In_2708,In_3780);
nor U4297 (N_4297,In_4092,In_1215);
or U4298 (N_4298,In_469,In_174);
or U4299 (N_4299,In_1785,In_1770);
xor U4300 (N_4300,In_580,In_905);
nand U4301 (N_4301,In_199,In_2110);
xnor U4302 (N_4302,In_2436,In_926);
or U4303 (N_4303,In_3516,In_3245);
nor U4304 (N_4304,In_1564,In_771);
nor U4305 (N_4305,In_1007,In_1663);
nand U4306 (N_4306,In_1533,In_3166);
or U4307 (N_4307,In_4313,In_1440);
and U4308 (N_4308,In_1659,In_405);
and U4309 (N_4309,In_3280,In_2573);
and U4310 (N_4310,In_3545,In_4945);
or U4311 (N_4311,In_4599,In_2190);
nor U4312 (N_4312,In_4419,In_3764);
and U4313 (N_4313,In_4851,In_4001);
or U4314 (N_4314,In_1216,In_4114);
or U4315 (N_4315,In_4935,In_2955);
and U4316 (N_4316,In_152,In_471);
and U4317 (N_4317,In_3096,In_4459);
nand U4318 (N_4318,In_109,In_4141);
nand U4319 (N_4319,In_3895,In_3116);
nand U4320 (N_4320,In_1829,In_278);
or U4321 (N_4321,In_1,In_1920);
and U4322 (N_4322,In_3859,In_4369);
nand U4323 (N_4323,In_207,In_896);
or U4324 (N_4324,In_601,In_1506);
nand U4325 (N_4325,In_4395,In_3922);
nand U4326 (N_4326,In_4646,In_2977);
nand U4327 (N_4327,In_1096,In_3813);
and U4328 (N_4328,In_4069,In_4665);
and U4329 (N_4329,In_4037,In_1892);
and U4330 (N_4330,In_1636,In_4428);
and U4331 (N_4331,In_2913,In_2071);
nand U4332 (N_4332,In_497,In_2515);
nor U4333 (N_4333,In_1355,In_615);
and U4334 (N_4334,In_2638,In_2159);
xor U4335 (N_4335,In_1121,In_2410);
xnor U4336 (N_4336,In_1559,In_1162);
or U4337 (N_4337,In_703,In_244);
or U4338 (N_4338,In_3608,In_3706);
nor U4339 (N_4339,In_4599,In_2772);
or U4340 (N_4340,In_4772,In_1273);
or U4341 (N_4341,In_4279,In_2868);
nor U4342 (N_4342,In_1728,In_2728);
and U4343 (N_4343,In_4455,In_1943);
nor U4344 (N_4344,In_3195,In_1730);
nand U4345 (N_4345,In_3110,In_3147);
or U4346 (N_4346,In_585,In_1015);
and U4347 (N_4347,In_429,In_460);
nand U4348 (N_4348,In_2461,In_2529);
or U4349 (N_4349,In_3453,In_1087);
and U4350 (N_4350,In_285,In_2571);
xnor U4351 (N_4351,In_219,In_4905);
nor U4352 (N_4352,In_473,In_3808);
or U4353 (N_4353,In_4669,In_3372);
and U4354 (N_4354,In_4293,In_4811);
or U4355 (N_4355,In_3662,In_3370);
xor U4356 (N_4356,In_2031,In_425);
nand U4357 (N_4357,In_3361,In_2673);
and U4358 (N_4358,In_99,In_4229);
or U4359 (N_4359,In_1183,In_4995);
or U4360 (N_4360,In_2150,In_4624);
nand U4361 (N_4361,In_54,In_3995);
nand U4362 (N_4362,In_2747,In_1517);
nand U4363 (N_4363,In_1099,In_2576);
and U4364 (N_4364,In_3432,In_672);
nor U4365 (N_4365,In_3260,In_2255);
and U4366 (N_4366,In_4798,In_4339);
or U4367 (N_4367,In_3581,In_3950);
and U4368 (N_4368,In_1371,In_842);
nand U4369 (N_4369,In_3193,In_3982);
xnor U4370 (N_4370,In_2981,In_2132);
nor U4371 (N_4371,In_4195,In_2004);
xor U4372 (N_4372,In_3699,In_4872);
or U4373 (N_4373,In_3943,In_4727);
nand U4374 (N_4374,In_3956,In_1925);
and U4375 (N_4375,In_376,In_3054);
xor U4376 (N_4376,In_3971,In_2543);
nand U4377 (N_4377,In_3177,In_2060);
nand U4378 (N_4378,In_4638,In_3137);
nand U4379 (N_4379,In_457,In_1587);
nand U4380 (N_4380,In_3150,In_1169);
nor U4381 (N_4381,In_3252,In_3711);
or U4382 (N_4382,In_366,In_3681);
or U4383 (N_4383,In_4246,In_2624);
nor U4384 (N_4384,In_3357,In_4886);
nand U4385 (N_4385,In_1136,In_4912);
nor U4386 (N_4386,In_3772,In_504);
or U4387 (N_4387,In_102,In_2900);
nor U4388 (N_4388,In_156,In_4486);
nand U4389 (N_4389,In_2786,In_4394);
or U4390 (N_4390,In_2597,In_2582);
nand U4391 (N_4391,In_1682,In_1838);
nor U4392 (N_4392,In_4521,In_1215);
nand U4393 (N_4393,In_4217,In_3074);
and U4394 (N_4394,In_2956,In_4295);
nor U4395 (N_4395,In_4610,In_436);
and U4396 (N_4396,In_1687,In_1002);
xor U4397 (N_4397,In_2846,In_3571);
nand U4398 (N_4398,In_1556,In_1734);
or U4399 (N_4399,In_3887,In_4783);
xor U4400 (N_4400,In_3144,In_3699);
nand U4401 (N_4401,In_2187,In_3919);
nor U4402 (N_4402,In_1383,In_2820);
and U4403 (N_4403,In_1391,In_3894);
nor U4404 (N_4404,In_3172,In_1351);
xnor U4405 (N_4405,In_597,In_1379);
or U4406 (N_4406,In_870,In_601);
xnor U4407 (N_4407,In_1405,In_2471);
and U4408 (N_4408,In_230,In_1076);
and U4409 (N_4409,In_742,In_2357);
nand U4410 (N_4410,In_2950,In_3264);
nand U4411 (N_4411,In_4719,In_307);
and U4412 (N_4412,In_2972,In_730);
and U4413 (N_4413,In_207,In_2776);
nand U4414 (N_4414,In_3721,In_4691);
and U4415 (N_4415,In_1651,In_3818);
xor U4416 (N_4416,In_1338,In_1517);
and U4417 (N_4417,In_3460,In_693);
nand U4418 (N_4418,In_120,In_820);
and U4419 (N_4419,In_3967,In_4942);
and U4420 (N_4420,In_490,In_1154);
xnor U4421 (N_4421,In_3787,In_4504);
nor U4422 (N_4422,In_2424,In_2436);
or U4423 (N_4423,In_1558,In_3424);
and U4424 (N_4424,In_2718,In_421);
nor U4425 (N_4425,In_1406,In_4324);
nor U4426 (N_4426,In_3488,In_4394);
xnor U4427 (N_4427,In_264,In_1276);
nand U4428 (N_4428,In_4123,In_372);
nor U4429 (N_4429,In_2193,In_1139);
and U4430 (N_4430,In_1419,In_3983);
xnor U4431 (N_4431,In_4776,In_996);
and U4432 (N_4432,In_2109,In_2402);
nor U4433 (N_4433,In_2728,In_1451);
and U4434 (N_4434,In_1846,In_1468);
or U4435 (N_4435,In_4019,In_660);
and U4436 (N_4436,In_4407,In_709);
or U4437 (N_4437,In_502,In_2302);
and U4438 (N_4438,In_1101,In_2002);
nand U4439 (N_4439,In_2343,In_3447);
nor U4440 (N_4440,In_1181,In_3135);
nor U4441 (N_4441,In_3371,In_4693);
nor U4442 (N_4442,In_2471,In_3692);
and U4443 (N_4443,In_2034,In_242);
or U4444 (N_4444,In_767,In_4151);
and U4445 (N_4445,In_4727,In_4334);
nand U4446 (N_4446,In_4001,In_4068);
or U4447 (N_4447,In_3361,In_1278);
nand U4448 (N_4448,In_2408,In_483);
and U4449 (N_4449,In_1594,In_624);
nor U4450 (N_4450,In_4467,In_1487);
or U4451 (N_4451,In_1058,In_4405);
nand U4452 (N_4452,In_480,In_786);
nand U4453 (N_4453,In_1738,In_4044);
and U4454 (N_4454,In_1466,In_3294);
nand U4455 (N_4455,In_1777,In_1139);
and U4456 (N_4456,In_2705,In_50);
nor U4457 (N_4457,In_726,In_3656);
nand U4458 (N_4458,In_3521,In_4656);
nor U4459 (N_4459,In_2026,In_471);
or U4460 (N_4460,In_1134,In_4442);
nor U4461 (N_4461,In_175,In_3407);
nand U4462 (N_4462,In_310,In_2965);
and U4463 (N_4463,In_32,In_2044);
or U4464 (N_4464,In_1987,In_1050);
nand U4465 (N_4465,In_2692,In_3727);
nor U4466 (N_4466,In_2523,In_4013);
xnor U4467 (N_4467,In_4363,In_178);
nor U4468 (N_4468,In_3877,In_2737);
xor U4469 (N_4469,In_1753,In_294);
or U4470 (N_4470,In_960,In_1139);
nor U4471 (N_4471,In_1360,In_169);
nand U4472 (N_4472,In_3881,In_665);
nor U4473 (N_4473,In_201,In_2303);
xnor U4474 (N_4474,In_2107,In_3398);
nand U4475 (N_4475,In_551,In_278);
or U4476 (N_4476,In_3574,In_2480);
xor U4477 (N_4477,In_872,In_3290);
or U4478 (N_4478,In_4196,In_1223);
nor U4479 (N_4479,In_3853,In_448);
and U4480 (N_4480,In_2886,In_4723);
xor U4481 (N_4481,In_3785,In_2098);
xor U4482 (N_4482,In_943,In_1797);
nor U4483 (N_4483,In_4685,In_2573);
xnor U4484 (N_4484,In_335,In_2371);
nor U4485 (N_4485,In_3269,In_475);
nand U4486 (N_4486,In_1173,In_2986);
nand U4487 (N_4487,In_3806,In_1316);
xnor U4488 (N_4488,In_2418,In_1492);
nand U4489 (N_4489,In_1138,In_594);
and U4490 (N_4490,In_1873,In_4566);
or U4491 (N_4491,In_1666,In_3354);
nor U4492 (N_4492,In_4554,In_4885);
or U4493 (N_4493,In_2375,In_4972);
and U4494 (N_4494,In_620,In_776);
xor U4495 (N_4495,In_4472,In_2153);
or U4496 (N_4496,In_4837,In_1039);
or U4497 (N_4497,In_2310,In_2125);
nor U4498 (N_4498,In_1074,In_2009);
nor U4499 (N_4499,In_4405,In_4671);
xor U4500 (N_4500,In_2155,In_1654);
nor U4501 (N_4501,In_2158,In_296);
and U4502 (N_4502,In_3982,In_3902);
nor U4503 (N_4503,In_4195,In_3624);
or U4504 (N_4504,In_955,In_1161);
nor U4505 (N_4505,In_3893,In_4944);
xnor U4506 (N_4506,In_530,In_2709);
nand U4507 (N_4507,In_4896,In_567);
nand U4508 (N_4508,In_3859,In_3485);
or U4509 (N_4509,In_1339,In_2861);
xor U4510 (N_4510,In_1193,In_1748);
and U4511 (N_4511,In_2055,In_1713);
xnor U4512 (N_4512,In_4656,In_848);
or U4513 (N_4513,In_975,In_3663);
nor U4514 (N_4514,In_633,In_1418);
or U4515 (N_4515,In_2481,In_3459);
and U4516 (N_4516,In_2310,In_4276);
nand U4517 (N_4517,In_2230,In_2775);
and U4518 (N_4518,In_3894,In_4575);
or U4519 (N_4519,In_1288,In_3550);
xnor U4520 (N_4520,In_3665,In_1437);
or U4521 (N_4521,In_3887,In_635);
and U4522 (N_4522,In_1171,In_622);
nor U4523 (N_4523,In_915,In_3478);
and U4524 (N_4524,In_2539,In_4076);
and U4525 (N_4525,In_2819,In_1633);
nand U4526 (N_4526,In_3930,In_898);
xor U4527 (N_4527,In_4430,In_4185);
or U4528 (N_4528,In_3660,In_4076);
and U4529 (N_4529,In_228,In_4354);
or U4530 (N_4530,In_4324,In_4838);
and U4531 (N_4531,In_1725,In_1275);
nand U4532 (N_4532,In_4082,In_3103);
nor U4533 (N_4533,In_1710,In_45);
xor U4534 (N_4534,In_2831,In_1314);
xor U4535 (N_4535,In_1818,In_2039);
or U4536 (N_4536,In_590,In_3407);
xor U4537 (N_4537,In_1986,In_2239);
or U4538 (N_4538,In_1627,In_1582);
nor U4539 (N_4539,In_2260,In_342);
nand U4540 (N_4540,In_4292,In_4528);
and U4541 (N_4541,In_4932,In_1989);
nor U4542 (N_4542,In_1155,In_4618);
and U4543 (N_4543,In_3733,In_1023);
xnor U4544 (N_4544,In_3767,In_3282);
nand U4545 (N_4545,In_1853,In_2770);
nand U4546 (N_4546,In_4349,In_3778);
nand U4547 (N_4547,In_1855,In_885);
and U4548 (N_4548,In_2049,In_2699);
nand U4549 (N_4549,In_2056,In_2519);
nand U4550 (N_4550,In_2004,In_1148);
nor U4551 (N_4551,In_2706,In_121);
xnor U4552 (N_4552,In_4425,In_2639);
or U4553 (N_4553,In_1745,In_2756);
and U4554 (N_4554,In_3920,In_4578);
and U4555 (N_4555,In_1054,In_4472);
and U4556 (N_4556,In_1716,In_4168);
nor U4557 (N_4557,In_1997,In_4338);
nor U4558 (N_4558,In_516,In_1860);
and U4559 (N_4559,In_3339,In_3906);
or U4560 (N_4560,In_2938,In_3225);
and U4561 (N_4561,In_842,In_3558);
or U4562 (N_4562,In_1613,In_4587);
nor U4563 (N_4563,In_4800,In_3309);
nand U4564 (N_4564,In_1832,In_359);
nor U4565 (N_4565,In_593,In_4530);
or U4566 (N_4566,In_2981,In_78);
or U4567 (N_4567,In_4223,In_850);
and U4568 (N_4568,In_4672,In_4023);
or U4569 (N_4569,In_4325,In_1949);
nand U4570 (N_4570,In_2316,In_3852);
and U4571 (N_4571,In_2204,In_1087);
nand U4572 (N_4572,In_3441,In_3687);
nand U4573 (N_4573,In_1380,In_4483);
nor U4574 (N_4574,In_3425,In_455);
and U4575 (N_4575,In_419,In_1428);
nor U4576 (N_4576,In_3637,In_2854);
nor U4577 (N_4577,In_3219,In_2408);
or U4578 (N_4578,In_4165,In_4363);
or U4579 (N_4579,In_3399,In_3896);
xor U4580 (N_4580,In_149,In_1334);
xnor U4581 (N_4581,In_1327,In_779);
nor U4582 (N_4582,In_2474,In_2741);
or U4583 (N_4583,In_652,In_3493);
xor U4584 (N_4584,In_2023,In_2110);
or U4585 (N_4585,In_4590,In_170);
nand U4586 (N_4586,In_644,In_212);
or U4587 (N_4587,In_52,In_2022);
xor U4588 (N_4588,In_780,In_2200);
xnor U4589 (N_4589,In_634,In_3804);
xnor U4590 (N_4590,In_617,In_4909);
or U4591 (N_4591,In_4782,In_2746);
xnor U4592 (N_4592,In_60,In_4967);
and U4593 (N_4593,In_2319,In_957);
or U4594 (N_4594,In_2586,In_1154);
or U4595 (N_4595,In_72,In_1747);
or U4596 (N_4596,In_2848,In_1770);
nand U4597 (N_4597,In_3282,In_4634);
xor U4598 (N_4598,In_3845,In_3276);
xor U4599 (N_4599,In_2470,In_1121);
and U4600 (N_4600,In_2933,In_2681);
nor U4601 (N_4601,In_2260,In_3750);
nand U4602 (N_4602,In_3553,In_4188);
nand U4603 (N_4603,In_153,In_250);
nor U4604 (N_4604,In_4593,In_1717);
and U4605 (N_4605,In_550,In_424);
and U4606 (N_4606,In_3647,In_2892);
nor U4607 (N_4607,In_4531,In_266);
and U4608 (N_4608,In_4865,In_1166);
nand U4609 (N_4609,In_4185,In_2814);
and U4610 (N_4610,In_1608,In_4805);
xnor U4611 (N_4611,In_4886,In_1325);
nor U4612 (N_4612,In_4315,In_1565);
and U4613 (N_4613,In_57,In_1477);
nor U4614 (N_4614,In_3206,In_3981);
nand U4615 (N_4615,In_3365,In_1373);
nor U4616 (N_4616,In_1027,In_2414);
nor U4617 (N_4617,In_2417,In_445);
xnor U4618 (N_4618,In_4747,In_562);
nand U4619 (N_4619,In_1976,In_158);
nor U4620 (N_4620,In_3409,In_4910);
nand U4621 (N_4621,In_4271,In_3750);
and U4622 (N_4622,In_1387,In_4274);
xnor U4623 (N_4623,In_3351,In_1918);
nand U4624 (N_4624,In_3505,In_4814);
nand U4625 (N_4625,In_1445,In_4654);
nor U4626 (N_4626,In_3636,In_4300);
and U4627 (N_4627,In_4664,In_4505);
nand U4628 (N_4628,In_410,In_1362);
xor U4629 (N_4629,In_1328,In_2500);
or U4630 (N_4630,In_134,In_217);
and U4631 (N_4631,In_4113,In_2411);
nor U4632 (N_4632,In_4319,In_3084);
nor U4633 (N_4633,In_162,In_2040);
nand U4634 (N_4634,In_4515,In_802);
or U4635 (N_4635,In_3845,In_1175);
and U4636 (N_4636,In_729,In_4501);
nor U4637 (N_4637,In_4807,In_4624);
and U4638 (N_4638,In_2410,In_1717);
nand U4639 (N_4639,In_4694,In_1565);
and U4640 (N_4640,In_3354,In_4510);
nor U4641 (N_4641,In_920,In_2351);
nor U4642 (N_4642,In_473,In_2829);
and U4643 (N_4643,In_4440,In_68);
nand U4644 (N_4644,In_3578,In_122);
nor U4645 (N_4645,In_3078,In_4344);
nand U4646 (N_4646,In_647,In_1761);
nor U4647 (N_4647,In_2667,In_1430);
nor U4648 (N_4648,In_590,In_4760);
or U4649 (N_4649,In_253,In_3638);
and U4650 (N_4650,In_3268,In_4382);
xnor U4651 (N_4651,In_4392,In_539);
and U4652 (N_4652,In_3935,In_1462);
xnor U4653 (N_4653,In_1052,In_106);
and U4654 (N_4654,In_2998,In_4768);
nor U4655 (N_4655,In_1282,In_3128);
or U4656 (N_4656,In_1375,In_2301);
nand U4657 (N_4657,In_1763,In_1178);
nor U4658 (N_4658,In_149,In_4494);
and U4659 (N_4659,In_4512,In_2555);
nor U4660 (N_4660,In_3544,In_939);
xor U4661 (N_4661,In_4410,In_1039);
and U4662 (N_4662,In_861,In_4898);
nor U4663 (N_4663,In_1592,In_3998);
and U4664 (N_4664,In_857,In_4317);
nand U4665 (N_4665,In_2607,In_4144);
nor U4666 (N_4666,In_1760,In_2899);
xnor U4667 (N_4667,In_4474,In_552);
xnor U4668 (N_4668,In_450,In_4892);
nor U4669 (N_4669,In_1856,In_2104);
nor U4670 (N_4670,In_4463,In_4034);
nor U4671 (N_4671,In_4795,In_1308);
and U4672 (N_4672,In_749,In_4853);
nor U4673 (N_4673,In_1913,In_4467);
and U4674 (N_4674,In_2957,In_1807);
and U4675 (N_4675,In_1081,In_2605);
xnor U4676 (N_4676,In_1616,In_1546);
xnor U4677 (N_4677,In_4735,In_2638);
and U4678 (N_4678,In_2140,In_3937);
and U4679 (N_4679,In_2858,In_4433);
and U4680 (N_4680,In_4951,In_59);
nand U4681 (N_4681,In_4064,In_2724);
nand U4682 (N_4682,In_4408,In_157);
or U4683 (N_4683,In_686,In_2096);
or U4684 (N_4684,In_3059,In_1476);
and U4685 (N_4685,In_1521,In_1925);
and U4686 (N_4686,In_1633,In_4859);
or U4687 (N_4687,In_2765,In_1816);
nand U4688 (N_4688,In_4058,In_4942);
nand U4689 (N_4689,In_2227,In_2272);
or U4690 (N_4690,In_250,In_1426);
xnor U4691 (N_4691,In_4959,In_1150);
nor U4692 (N_4692,In_2510,In_1948);
nand U4693 (N_4693,In_3748,In_1530);
or U4694 (N_4694,In_2953,In_1841);
and U4695 (N_4695,In_2852,In_764);
or U4696 (N_4696,In_1550,In_198);
or U4697 (N_4697,In_3644,In_1854);
and U4698 (N_4698,In_1040,In_2388);
nor U4699 (N_4699,In_1433,In_4254);
or U4700 (N_4700,In_4863,In_3333);
and U4701 (N_4701,In_257,In_3548);
and U4702 (N_4702,In_1777,In_4666);
or U4703 (N_4703,In_3454,In_3992);
nor U4704 (N_4704,In_1881,In_179);
and U4705 (N_4705,In_4392,In_852);
xor U4706 (N_4706,In_1687,In_3109);
nand U4707 (N_4707,In_1170,In_4866);
or U4708 (N_4708,In_4818,In_4888);
nor U4709 (N_4709,In_2786,In_4755);
and U4710 (N_4710,In_2077,In_4654);
or U4711 (N_4711,In_2341,In_4988);
or U4712 (N_4712,In_4340,In_4030);
nor U4713 (N_4713,In_1952,In_262);
nor U4714 (N_4714,In_3564,In_2710);
xor U4715 (N_4715,In_3068,In_1143);
or U4716 (N_4716,In_4293,In_4946);
nand U4717 (N_4717,In_2013,In_460);
or U4718 (N_4718,In_950,In_4025);
or U4719 (N_4719,In_4063,In_4568);
and U4720 (N_4720,In_2824,In_187);
and U4721 (N_4721,In_3954,In_3757);
or U4722 (N_4722,In_348,In_2401);
nor U4723 (N_4723,In_1954,In_1133);
nand U4724 (N_4724,In_4494,In_1682);
xor U4725 (N_4725,In_816,In_3776);
nand U4726 (N_4726,In_2279,In_2528);
or U4727 (N_4727,In_3603,In_4964);
xnor U4728 (N_4728,In_472,In_2248);
and U4729 (N_4729,In_585,In_1848);
or U4730 (N_4730,In_2621,In_3566);
and U4731 (N_4731,In_150,In_431);
nor U4732 (N_4732,In_4383,In_1347);
nand U4733 (N_4733,In_1950,In_705);
or U4734 (N_4734,In_924,In_4792);
nand U4735 (N_4735,In_4597,In_3394);
nor U4736 (N_4736,In_2052,In_435);
nand U4737 (N_4737,In_4689,In_398);
and U4738 (N_4738,In_3316,In_4266);
xor U4739 (N_4739,In_2176,In_1323);
or U4740 (N_4740,In_3052,In_2657);
or U4741 (N_4741,In_3786,In_164);
or U4742 (N_4742,In_1927,In_3023);
nor U4743 (N_4743,In_485,In_4985);
nand U4744 (N_4744,In_4125,In_4997);
and U4745 (N_4745,In_1835,In_1935);
and U4746 (N_4746,In_3197,In_1128);
nor U4747 (N_4747,In_2899,In_4895);
or U4748 (N_4748,In_2589,In_2931);
and U4749 (N_4749,In_3771,In_878);
nand U4750 (N_4750,In_3107,In_4399);
nand U4751 (N_4751,In_2989,In_759);
nor U4752 (N_4752,In_4523,In_4087);
and U4753 (N_4753,In_198,In_4831);
and U4754 (N_4754,In_4979,In_620);
or U4755 (N_4755,In_4011,In_4014);
or U4756 (N_4756,In_2083,In_3836);
nand U4757 (N_4757,In_3878,In_966);
and U4758 (N_4758,In_22,In_2286);
nor U4759 (N_4759,In_4334,In_1436);
and U4760 (N_4760,In_3295,In_1709);
and U4761 (N_4761,In_4064,In_3360);
nor U4762 (N_4762,In_468,In_2532);
nand U4763 (N_4763,In_1289,In_3379);
nand U4764 (N_4764,In_852,In_1628);
xor U4765 (N_4765,In_1311,In_1208);
nand U4766 (N_4766,In_938,In_543);
nor U4767 (N_4767,In_3986,In_3304);
xor U4768 (N_4768,In_167,In_3958);
nor U4769 (N_4769,In_2319,In_291);
and U4770 (N_4770,In_3412,In_4945);
nand U4771 (N_4771,In_1714,In_712);
xnor U4772 (N_4772,In_3986,In_4901);
nand U4773 (N_4773,In_3835,In_1066);
xor U4774 (N_4774,In_3888,In_4959);
nor U4775 (N_4775,In_760,In_3266);
or U4776 (N_4776,In_3870,In_42);
nand U4777 (N_4777,In_2242,In_2469);
nor U4778 (N_4778,In_1068,In_2042);
nand U4779 (N_4779,In_2833,In_1899);
or U4780 (N_4780,In_557,In_4530);
nand U4781 (N_4781,In_4971,In_2241);
nor U4782 (N_4782,In_3180,In_2604);
nand U4783 (N_4783,In_2706,In_1685);
and U4784 (N_4784,In_767,In_782);
nand U4785 (N_4785,In_4188,In_3753);
or U4786 (N_4786,In_2759,In_4536);
nand U4787 (N_4787,In_1778,In_2236);
nand U4788 (N_4788,In_3683,In_1333);
or U4789 (N_4789,In_2774,In_2706);
and U4790 (N_4790,In_1924,In_3521);
and U4791 (N_4791,In_4735,In_819);
or U4792 (N_4792,In_1073,In_636);
nor U4793 (N_4793,In_22,In_1316);
nand U4794 (N_4794,In_3236,In_819);
nor U4795 (N_4795,In_2950,In_3134);
xnor U4796 (N_4796,In_3003,In_3958);
and U4797 (N_4797,In_3457,In_3668);
or U4798 (N_4798,In_2585,In_2890);
xor U4799 (N_4799,In_2563,In_232);
nand U4800 (N_4800,In_2111,In_3935);
or U4801 (N_4801,In_2873,In_537);
or U4802 (N_4802,In_3465,In_4560);
nand U4803 (N_4803,In_1372,In_3659);
or U4804 (N_4804,In_3186,In_1261);
nor U4805 (N_4805,In_912,In_4327);
and U4806 (N_4806,In_4872,In_4392);
nor U4807 (N_4807,In_2020,In_4519);
nand U4808 (N_4808,In_2574,In_1194);
nor U4809 (N_4809,In_1854,In_3130);
and U4810 (N_4810,In_3377,In_4365);
and U4811 (N_4811,In_4710,In_412);
nor U4812 (N_4812,In_1362,In_4348);
or U4813 (N_4813,In_3965,In_1852);
or U4814 (N_4814,In_2363,In_3631);
or U4815 (N_4815,In_4070,In_1073);
or U4816 (N_4816,In_2349,In_984);
or U4817 (N_4817,In_4281,In_3871);
or U4818 (N_4818,In_4845,In_3392);
nand U4819 (N_4819,In_4666,In_4548);
or U4820 (N_4820,In_70,In_1992);
nor U4821 (N_4821,In_1023,In_1360);
or U4822 (N_4822,In_2192,In_953);
nand U4823 (N_4823,In_4673,In_3610);
or U4824 (N_4824,In_1011,In_3965);
and U4825 (N_4825,In_4514,In_4354);
and U4826 (N_4826,In_3565,In_1951);
or U4827 (N_4827,In_2020,In_1702);
nor U4828 (N_4828,In_2857,In_3277);
nand U4829 (N_4829,In_314,In_2839);
nor U4830 (N_4830,In_773,In_2196);
nand U4831 (N_4831,In_3969,In_717);
nor U4832 (N_4832,In_3939,In_3494);
and U4833 (N_4833,In_4182,In_1017);
xor U4834 (N_4834,In_371,In_3094);
nor U4835 (N_4835,In_2094,In_835);
xor U4836 (N_4836,In_4400,In_2668);
or U4837 (N_4837,In_463,In_1548);
nand U4838 (N_4838,In_1539,In_618);
and U4839 (N_4839,In_3796,In_1469);
nor U4840 (N_4840,In_486,In_4919);
nor U4841 (N_4841,In_1368,In_3729);
or U4842 (N_4842,In_1575,In_324);
nor U4843 (N_4843,In_4536,In_951);
and U4844 (N_4844,In_4331,In_4759);
nand U4845 (N_4845,In_1645,In_1709);
nand U4846 (N_4846,In_4969,In_12);
and U4847 (N_4847,In_3771,In_1296);
nor U4848 (N_4848,In_1603,In_4192);
nor U4849 (N_4849,In_4757,In_1665);
nor U4850 (N_4850,In_4328,In_3267);
or U4851 (N_4851,In_757,In_1465);
nand U4852 (N_4852,In_4179,In_4934);
and U4853 (N_4853,In_1524,In_3405);
and U4854 (N_4854,In_2987,In_772);
nor U4855 (N_4855,In_794,In_2471);
nor U4856 (N_4856,In_1270,In_2749);
nand U4857 (N_4857,In_3647,In_242);
nor U4858 (N_4858,In_1463,In_1665);
nor U4859 (N_4859,In_4124,In_3533);
or U4860 (N_4860,In_3906,In_1747);
nand U4861 (N_4861,In_2628,In_2558);
and U4862 (N_4862,In_4374,In_2688);
and U4863 (N_4863,In_1285,In_1068);
nor U4864 (N_4864,In_2568,In_3853);
nor U4865 (N_4865,In_1365,In_3469);
and U4866 (N_4866,In_3850,In_1549);
nor U4867 (N_4867,In_4205,In_3157);
or U4868 (N_4868,In_3459,In_2115);
and U4869 (N_4869,In_1059,In_4411);
or U4870 (N_4870,In_4214,In_1241);
or U4871 (N_4871,In_1243,In_2708);
nand U4872 (N_4872,In_4393,In_796);
and U4873 (N_4873,In_4635,In_2204);
or U4874 (N_4874,In_1898,In_750);
xnor U4875 (N_4875,In_448,In_3519);
nor U4876 (N_4876,In_580,In_1028);
and U4877 (N_4877,In_317,In_2358);
and U4878 (N_4878,In_4948,In_565);
nor U4879 (N_4879,In_3087,In_2365);
nor U4880 (N_4880,In_2799,In_1067);
and U4881 (N_4881,In_2052,In_533);
nand U4882 (N_4882,In_3756,In_3877);
nand U4883 (N_4883,In_1486,In_3167);
nor U4884 (N_4884,In_4307,In_1382);
or U4885 (N_4885,In_3947,In_3241);
or U4886 (N_4886,In_2182,In_3302);
nand U4887 (N_4887,In_128,In_160);
nand U4888 (N_4888,In_574,In_3756);
nand U4889 (N_4889,In_3964,In_4237);
and U4890 (N_4890,In_4857,In_2534);
nor U4891 (N_4891,In_1450,In_193);
xor U4892 (N_4892,In_4904,In_3505);
nand U4893 (N_4893,In_27,In_3732);
and U4894 (N_4894,In_872,In_1618);
nor U4895 (N_4895,In_4189,In_2535);
nand U4896 (N_4896,In_487,In_4769);
nor U4897 (N_4897,In_2200,In_2008);
or U4898 (N_4898,In_207,In_4790);
nand U4899 (N_4899,In_1289,In_2745);
nor U4900 (N_4900,In_2165,In_4620);
and U4901 (N_4901,In_4238,In_3937);
nand U4902 (N_4902,In_229,In_2261);
nor U4903 (N_4903,In_3279,In_954);
and U4904 (N_4904,In_3356,In_1605);
nand U4905 (N_4905,In_3376,In_554);
nand U4906 (N_4906,In_4848,In_517);
and U4907 (N_4907,In_4608,In_906);
xnor U4908 (N_4908,In_4023,In_3054);
nor U4909 (N_4909,In_4655,In_1745);
xnor U4910 (N_4910,In_415,In_2703);
xnor U4911 (N_4911,In_1418,In_1289);
or U4912 (N_4912,In_2424,In_4412);
or U4913 (N_4913,In_87,In_4118);
nor U4914 (N_4914,In_947,In_2560);
and U4915 (N_4915,In_2929,In_3195);
and U4916 (N_4916,In_3939,In_4221);
xnor U4917 (N_4917,In_1825,In_772);
nand U4918 (N_4918,In_2516,In_1431);
and U4919 (N_4919,In_2017,In_3047);
nand U4920 (N_4920,In_2661,In_2493);
or U4921 (N_4921,In_2065,In_2152);
nor U4922 (N_4922,In_2827,In_2806);
and U4923 (N_4923,In_4608,In_4243);
and U4924 (N_4924,In_1276,In_1239);
nor U4925 (N_4925,In_1243,In_1859);
nand U4926 (N_4926,In_2323,In_386);
nor U4927 (N_4927,In_3768,In_2775);
xnor U4928 (N_4928,In_2360,In_4825);
nand U4929 (N_4929,In_1206,In_4373);
and U4930 (N_4930,In_2377,In_1589);
and U4931 (N_4931,In_443,In_891);
and U4932 (N_4932,In_3645,In_169);
and U4933 (N_4933,In_1902,In_751);
xnor U4934 (N_4934,In_3819,In_225);
and U4935 (N_4935,In_3332,In_507);
nor U4936 (N_4936,In_4251,In_2366);
or U4937 (N_4937,In_4231,In_1522);
and U4938 (N_4938,In_2843,In_1836);
nand U4939 (N_4939,In_1142,In_125);
xnor U4940 (N_4940,In_4815,In_1834);
or U4941 (N_4941,In_4146,In_4504);
and U4942 (N_4942,In_133,In_1821);
xor U4943 (N_4943,In_1293,In_2619);
nor U4944 (N_4944,In_1724,In_4893);
and U4945 (N_4945,In_2847,In_3504);
or U4946 (N_4946,In_4954,In_2077);
and U4947 (N_4947,In_1338,In_4931);
or U4948 (N_4948,In_2736,In_2840);
or U4949 (N_4949,In_4490,In_4175);
nand U4950 (N_4950,In_2764,In_3359);
nand U4951 (N_4951,In_3747,In_3835);
and U4952 (N_4952,In_332,In_54);
xor U4953 (N_4953,In_4293,In_4457);
nor U4954 (N_4954,In_4979,In_3565);
nand U4955 (N_4955,In_42,In_4041);
or U4956 (N_4956,In_1943,In_4713);
nor U4957 (N_4957,In_2613,In_297);
or U4958 (N_4958,In_3770,In_960);
and U4959 (N_4959,In_243,In_3831);
or U4960 (N_4960,In_4706,In_4419);
or U4961 (N_4961,In_1463,In_1142);
nor U4962 (N_4962,In_1569,In_3270);
xnor U4963 (N_4963,In_335,In_1166);
xor U4964 (N_4964,In_1612,In_3069);
nand U4965 (N_4965,In_615,In_1225);
and U4966 (N_4966,In_91,In_3658);
or U4967 (N_4967,In_4120,In_961);
and U4968 (N_4968,In_1063,In_4550);
or U4969 (N_4969,In_304,In_1621);
nor U4970 (N_4970,In_1506,In_4037);
nand U4971 (N_4971,In_348,In_2721);
nand U4972 (N_4972,In_2594,In_4781);
or U4973 (N_4973,In_537,In_168);
nand U4974 (N_4974,In_3365,In_4523);
xnor U4975 (N_4975,In_3240,In_4151);
nand U4976 (N_4976,In_535,In_1345);
nor U4977 (N_4977,In_3251,In_2517);
nor U4978 (N_4978,In_4138,In_104);
nor U4979 (N_4979,In_690,In_1753);
or U4980 (N_4980,In_3495,In_2754);
nor U4981 (N_4981,In_1998,In_3182);
and U4982 (N_4982,In_3312,In_3116);
and U4983 (N_4983,In_3759,In_2509);
nor U4984 (N_4984,In_4946,In_1800);
xor U4985 (N_4985,In_493,In_3406);
nor U4986 (N_4986,In_2597,In_1593);
nand U4987 (N_4987,In_1025,In_3885);
and U4988 (N_4988,In_2099,In_243);
and U4989 (N_4989,In_574,In_28);
xnor U4990 (N_4990,In_783,In_580);
or U4991 (N_4991,In_3274,In_2344);
nand U4992 (N_4992,In_2260,In_3079);
or U4993 (N_4993,In_1234,In_4953);
nand U4994 (N_4994,In_2672,In_3288);
and U4995 (N_4995,In_4807,In_4477);
nor U4996 (N_4996,In_4112,In_332);
or U4997 (N_4997,In_1341,In_4556);
nor U4998 (N_4998,In_1373,In_3427);
xor U4999 (N_4999,In_845,In_2353);
nor U5000 (N_5000,N_3401,N_89);
nand U5001 (N_5001,N_4375,N_3920);
nor U5002 (N_5002,N_1397,N_4533);
and U5003 (N_5003,N_2733,N_2388);
nor U5004 (N_5004,N_2176,N_901);
nor U5005 (N_5005,N_2321,N_2629);
nand U5006 (N_5006,N_4300,N_3666);
nor U5007 (N_5007,N_3693,N_885);
nand U5008 (N_5008,N_2583,N_61);
or U5009 (N_5009,N_2868,N_1552);
and U5010 (N_5010,N_4723,N_393);
nor U5011 (N_5011,N_2762,N_3671);
or U5012 (N_5012,N_4,N_2823);
or U5013 (N_5013,N_806,N_2230);
and U5014 (N_5014,N_3446,N_3362);
and U5015 (N_5015,N_2455,N_4271);
and U5016 (N_5016,N_2094,N_1752);
nand U5017 (N_5017,N_4553,N_3252);
and U5018 (N_5018,N_4036,N_4909);
and U5019 (N_5019,N_1271,N_2200);
or U5020 (N_5020,N_2579,N_2298);
and U5021 (N_5021,N_4076,N_68);
and U5022 (N_5022,N_4401,N_4492);
nand U5023 (N_5023,N_1347,N_3155);
nand U5024 (N_5024,N_2711,N_3239);
xor U5025 (N_5025,N_2128,N_1656);
and U5026 (N_5026,N_3686,N_421);
and U5027 (N_5027,N_4333,N_1555);
nor U5028 (N_5028,N_4319,N_1612);
and U5029 (N_5029,N_2165,N_4833);
and U5030 (N_5030,N_2995,N_3115);
xor U5031 (N_5031,N_4911,N_1162);
nor U5032 (N_5032,N_3278,N_445);
nor U5033 (N_5033,N_2991,N_3489);
or U5034 (N_5034,N_942,N_657);
nor U5035 (N_5035,N_2704,N_4211);
or U5036 (N_5036,N_3809,N_1796);
nand U5037 (N_5037,N_4924,N_1222);
or U5038 (N_5038,N_4470,N_3325);
or U5039 (N_5039,N_3476,N_3586);
xnor U5040 (N_5040,N_589,N_1866);
or U5041 (N_5041,N_695,N_1813);
nor U5042 (N_5042,N_1539,N_4937);
and U5043 (N_5043,N_4193,N_4528);
nor U5044 (N_5044,N_4860,N_3684);
or U5045 (N_5045,N_2047,N_166);
or U5046 (N_5046,N_3991,N_1589);
nor U5047 (N_5047,N_4108,N_4182);
nor U5048 (N_5048,N_3166,N_411);
or U5049 (N_5049,N_4186,N_1158);
and U5050 (N_5050,N_4985,N_3378);
and U5051 (N_5051,N_746,N_4517);
and U5052 (N_5052,N_3199,N_2319);
nor U5053 (N_5053,N_3936,N_298);
nand U5054 (N_5054,N_532,N_1319);
and U5055 (N_5055,N_4745,N_1764);
xor U5056 (N_5056,N_4897,N_2138);
xnor U5057 (N_5057,N_3929,N_4145);
or U5058 (N_5058,N_4825,N_3122);
nor U5059 (N_5059,N_302,N_3086);
nand U5060 (N_5060,N_2233,N_440);
and U5061 (N_5061,N_3396,N_1938);
nand U5062 (N_5062,N_4586,N_3546);
and U5063 (N_5063,N_3738,N_2724);
nand U5064 (N_5064,N_4596,N_3363);
nand U5065 (N_5065,N_4709,N_1123);
and U5066 (N_5066,N_1226,N_878);
nor U5067 (N_5067,N_307,N_4231);
nand U5068 (N_5068,N_4432,N_3604);
nand U5069 (N_5069,N_4336,N_1543);
or U5070 (N_5070,N_1521,N_3903);
and U5071 (N_5071,N_356,N_3949);
or U5072 (N_5072,N_311,N_737);
nand U5073 (N_5073,N_4419,N_289);
nor U5074 (N_5074,N_4625,N_1779);
nand U5075 (N_5075,N_2734,N_3273);
or U5076 (N_5076,N_3358,N_3424);
xnor U5077 (N_5077,N_221,N_2433);
and U5078 (N_5078,N_716,N_937);
nand U5079 (N_5079,N_1522,N_3970);
or U5080 (N_5080,N_1704,N_799);
nand U5081 (N_5081,N_4240,N_2098);
and U5082 (N_5082,N_2637,N_596);
and U5083 (N_5083,N_15,N_818);
and U5084 (N_5084,N_4565,N_2745);
nor U5085 (N_5085,N_3963,N_519);
nor U5086 (N_5086,N_826,N_4755);
and U5087 (N_5087,N_830,N_1223);
nor U5088 (N_5088,N_3771,N_2067);
xnor U5089 (N_5089,N_2025,N_4244);
or U5090 (N_5090,N_814,N_2702);
nor U5091 (N_5091,N_1044,N_4578);
nand U5092 (N_5092,N_3876,N_1959);
xnor U5093 (N_5093,N_531,N_4526);
or U5094 (N_5094,N_3416,N_668);
nor U5095 (N_5095,N_4576,N_2761);
nand U5096 (N_5096,N_1056,N_3973);
or U5097 (N_5097,N_1942,N_4437);
nor U5098 (N_5098,N_4953,N_2006);
and U5099 (N_5099,N_1182,N_3573);
xor U5100 (N_5100,N_3966,N_908);
nand U5101 (N_5101,N_1117,N_190);
and U5102 (N_5102,N_3770,N_2195);
nor U5103 (N_5103,N_3701,N_4888);
and U5104 (N_5104,N_2982,N_754);
and U5105 (N_5105,N_861,N_2719);
nor U5106 (N_5106,N_4201,N_2521);
or U5107 (N_5107,N_4352,N_4091);
nand U5108 (N_5108,N_4129,N_3326);
and U5109 (N_5109,N_400,N_4136);
or U5110 (N_5110,N_4612,N_269);
or U5111 (N_5111,N_2698,N_280);
nand U5112 (N_5112,N_1885,N_4637);
and U5113 (N_5113,N_1253,N_4621);
xnor U5114 (N_5114,N_344,N_1105);
nand U5115 (N_5115,N_2616,N_1677);
or U5116 (N_5116,N_40,N_859);
or U5117 (N_5117,N_1301,N_562);
or U5118 (N_5118,N_2595,N_4908);
and U5119 (N_5119,N_643,N_499);
or U5120 (N_5120,N_1024,N_3948);
and U5121 (N_5121,N_392,N_4701);
or U5122 (N_5122,N_3387,N_1623);
nand U5123 (N_5123,N_4534,N_1619);
or U5124 (N_5124,N_3612,N_148);
nor U5125 (N_5125,N_4183,N_996);
nor U5126 (N_5126,N_4384,N_4007);
or U5127 (N_5127,N_1459,N_1815);
nor U5128 (N_5128,N_3514,N_225);
or U5129 (N_5129,N_4281,N_1549);
and U5130 (N_5130,N_28,N_2207);
nand U5131 (N_5131,N_3825,N_3411);
nand U5132 (N_5132,N_187,N_3370);
or U5133 (N_5133,N_4964,N_1432);
xor U5134 (N_5134,N_4799,N_181);
or U5135 (N_5135,N_3008,N_2366);
and U5136 (N_5136,N_2679,N_13);
and U5137 (N_5137,N_3529,N_2948);
xnor U5138 (N_5138,N_70,N_4498);
nand U5139 (N_5139,N_1978,N_1348);
nand U5140 (N_5140,N_4077,N_1682);
or U5141 (N_5141,N_2665,N_4486);
or U5142 (N_5142,N_3403,N_3822);
and U5143 (N_5143,N_481,N_4125);
nand U5144 (N_5144,N_1931,N_2785);
nand U5145 (N_5145,N_4503,N_2820);
nor U5146 (N_5146,N_3608,N_2383);
nor U5147 (N_5147,N_4259,N_2531);
and U5148 (N_5148,N_4017,N_2456);
nand U5149 (N_5149,N_1402,N_3862);
or U5150 (N_5150,N_4624,N_2282);
nor U5151 (N_5151,N_970,N_2143);
and U5152 (N_5152,N_1523,N_1136);
nand U5153 (N_5153,N_2895,N_525);
nand U5154 (N_5154,N_154,N_2569);
or U5155 (N_5155,N_3906,N_4782);
nor U5156 (N_5156,N_1040,N_2580);
xor U5157 (N_5157,N_3860,N_47);
nor U5158 (N_5158,N_3961,N_1016);
and U5159 (N_5159,N_4542,N_3430);
or U5160 (N_5160,N_4960,N_1644);
nand U5161 (N_5161,N_4121,N_3742);
nand U5162 (N_5162,N_2986,N_1374);
nor U5163 (N_5163,N_3481,N_1037);
nor U5164 (N_5164,N_3164,N_4758);
or U5165 (N_5165,N_4887,N_3210);
and U5166 (N_5166,N_1786,N_4010);
or U5167 (N_5167,N_808,N_3734);
and U5168 (N_5168,N_2317,N_1287);
nand U5169 (N_5169,N_4824,N_2381);
and U5170 (N_5170,N_3540,N_950);
or U5171 (N_5171,N_2299,N_1944);
nor U5172 (N_5172,N_599,N_3275);
xnor U5173 (N_5173,N_3957,N_3756);
and U5174 (N_5174,N_123,N_1715);
nand U5175 (N_5175,N_4390,N_2337);
nand U5176 (N_5176,N_748,N_636);
and U5177 (N_5177,N_1110,N_3972);
or U5178 (N_5178,N_3369,N_881);
and U5179 (N_5179,N_1538,N_4223);
nor U5180 (N_5180,N_4163,N_4307);
and U5181 (N_5181,N_4254,N_536);
and U5182 (N_5182,N_2744,N_981);
nor U5183 (N_5183,N_353,N_2707);
nand U5184 (N_5184,N_2286,N_1964);
nor U5185 (N_5185,N_2812,N_4350);
nand U5186 (N_5186,N_483,N_3640);
nor U5187 (N_5187,N_2426,N_1603);
nand U5188 (N_5188,N_555,N_734);
and U5189 (N_5189,N_3627,N_1751);
nor U5190 (N_5190,N_2396,N_1932);
xnor U5191 (N_5191,N_4731,N_2210);
nand U5192 (N_5192,N_3533,N_1683);
nand U5193 (N_5193,N_4872,N_4198);
nand U5194 (N_5194,N_87,N_468);
nand U5195 (N_5195,N_3786,N_823);
and U5196 (N_5196,N_4722,N_3209);
or U5197 (N_5197,N_2803,N_3266);
nor U5198 (N_5198,N_4312,N_1621);
nor U5199 (N_5199,N_4740,N_2221);
or U5200 (N_5200,N_731,N_1205);
nor U5201 (N_5201,N_2493,N_658);
nand U5202 (N_5202,N_4316,N_407);
or U5203 (N_5203,N_3421,N_3993);
xor U5204 (N_5204,N_2652,N_3260);
nor U5205 (N_5205,N_309,N_3);
nor U5206 (N_5206,N_3933,N_1022);
or U5207 (N_5207,N_3519,N_4795);
nand U5208 (N_5208,N_3685,N_1741);
or U5209 (N_5209,N_3212,N_3160);
and U5210 (N_5210,N_1719,N_3934);
nor U5211 (N_5211,N_3784,N_3832);
and U5212 (N_5212,N_3617,N_378);
nor U5213 (N_5213,N_3391,N_4761);
or U5214 (N_5214,N_3538,N_2093);
and U5215 (N_5215,N_240,N_4836);
nand U5216 (N_5216,N_3690,N_3333);
nor U5217 (N_5217,N_3074,N_3301);
nor U5218 (N_5218,N_4792,N_2326);
or U5219 (N_5219,N_4355,N_3642);
nor U5220 (N_5220,N_2065,N_2754);
nand U5221 (N_5221,N_4631,N_4410);
nor U5222 (N_5222,N_2671,N_1785);
or U5223 (N_5223,N_1470,N_3023);
and U5224 (N_5224,N_1924,N_4233);
or U5225 (N_5225,N_503,N_2100);
nor U5226 (N_5226,N_2348,N_2229);
xnor U5227 (N_5227,N_215,N_2749);
and U5228 (N_5228,N_3073,N_2979);
and U5229 (N_5229,N_2750,N_2550);
and U5230 (N_5230,N_4383,N_3549);
nor U5231 (N_5231,N_432,N_433);
and U5232 (N_5232,N_1987,N_3726);
nor U5233 (N_5233,N_1661,N_3480);
nor U5234 (N_5234,N_2778,N_4510);
nor U5235 (N_5235,N_3217,N_3835);
or U5236 (N_5236,N_3276,N_2071);
xnor U5237 (N_5237,N_1339,N_4008);
xor U5238 (N_5238,N_165,N_3950);
nor U5239 (N_5239,N_4747,N_2187);
nor U5240 (N_5240,N_2101,N_745);
nand U5241 (N_5241,N_4327,N_2809);
nor U5242 (N_5242,N_2320,N_4192);
and U5243 (N_5243,N_1586,N_771);
or U5244 (N_5244,N_963,N_4828);
and U5245 (N_5245,N_4177,N_592);
nor U5246 (N_5246,N_2048,N_2873);
nand U5247 (N_5247,N_3114,N_1191);
nor U5248 (N_5248,N_4770,N_4680);
and U5249 (N_5249,N_2329,N_3758);
and U5250 (N_5250,N_1714,N_2136);
nor U5251 (N_5251,N_3094,N_2377);
and U5252 (N_5252,N_3465,N_4870);
nand U5253 (N_5253,N_1579,N_2607);
nor U5254 (N_5254,N_2180,N_2590);
and U5255 (N_5255,N_1650,N_2014);
nand U5256 (N_5256,N_1377,N_2919);
nor U5257 (N_5257,N_418,N_2597);
and U5258 (N_5258,N_313,N_3989);
nor U5259 (N_5259,N_4942,N_4907);
nor U5260 (N_5260,N_4839,N_1150);
nand U5261 (N_5261,N_1312,N_565);
or U5262 (N_5262,N_1230,N_3352);
nor U5263 (N_5263,N_1986,N_4055);
or U5264 (N_5264,N_4948,N_394);
and U5265 (N_5265,N_17,N_2027);
xor U5266 (N_5266,N_3940,N_2837);
and U5267 (N_5267,N_266,N_3850);
or U5268 (N_5268,N_1132,N_417);
and U5269 (N_5269,N_516,N_4049);
or U5270 (N_5270,N_1531,N_2677);
nand U5271 (N_5271,N_728,N_4242);
nand U5272 (N_5272,N_497,N_2821);
nor U5273 (N_5273,N_522,N_2256);
nor U5274 (N_5274,N_3737,N_195);
nor U5275 (N_5275,N_778,N_3222);
or U5276 (N_5276,N_1357,N_4850);
nor U5277 (N_5277,N_4629,N_1121);
and U5278 (N_5278,N_2680,N_4998);
nor U5279 (N_5279,N_3389,N_4377);
xnor U5280 (N_5280,N_1581,N_2389);
and U5281 (N_5281,N_3556,N_1439);
nand U5282 (N_5282,N_4563,N_1845);
nor U5283 (N_5283,N_366,N_3852);
or U5284 (N_5284,N_1266,N_1088);
and U5285 (N_5285,N_4321,N_3995);
and U5286 (N_5286,N_1332,N_2227);
xnor U5287 (N_5287,N_4015,N_176);
nor U5288 (N_5288,N_1179,N_988);
nand U5289 (N_5289,N_4651,N_2118);
and U5290 (N_5290,N_3081,N_3682);
nor U5291 (N_5291,N_705,N_3547);
and U5292 (N_5292,N_3909,N_4944);
nor U5293 (N_5293,N_1052,N_4171);
or U5294 (N_5294,N_4222,N_3557);
xor U5295 (N_5295,N_3808,N_1091);
and U5296 (N_5296,N_1697,N_3512);
nor U5297 (N_5297,N_2892,N_2205);
nor U5298 (N_5298,N_2738,N_4243);
nand U5299 (N_5299,N_3169,N_1535);
nand U5300 (N_5300,N_3196,N_4704);
nor U5301 (N_5301,N_858,N_446);
nor U5302 (N_5302,N_974,N_4575);
nor U5303 (N_5303,N_2281,N_4979);
nand U5304 (N_5304,N_2474,N_2368);
nor U5305 (N_5305,N_794,N_569);
and U5306 (N_5306,N_3354,N_3555);
nor U5307 (N_5307,N_4078,N_3576);
xor U5308 (N_5308,N_2942,N_3853);
xnor U5309 (N_5309,N_3486,N_4769);
nor U5310 (N_5310,N_1240,N_1074);
or U5311 (N_5311,N_2601,N_3721);
or U5312 (N_5312,N_655,N_2782);
and U5313 (N_5313,N_1283,N_1277);
or U5314 (N_5314,N_3807,N_2984);
and U5315 (N_5315,N_4956,N_4464);
nor U5316 (N_5316,N_2507,N_1901);
or U5317 (N_5317,N_1429,N_3603);
xnor U5318 (N_5318,N_682,N_4019);
and U5319 (N_5319,N_4739,N_3998);
and U5320 (N_5320,N_1562,N_2797);
or U5321 (N_5321,N_1310,N_4277);
xnor U5322 (N_5322,N_188,N_2675);
nand U5323 (N_5323,N_2324,N_4139);
nand U5324 (N_5324,N_4212,N_3788);
and U5325 (N_5325,N_837,N_4245);
nand U5326 (N_5326,N_1126,N_472);
xnor U5327 (N_5327,N_4516,N_4142);
or U5328 (N_5328,N_4028,N_1524);
nor U5329 (N_5329,N_1078,N_2503);
or U5330 (N_5330,N_4706,N_3648);
or U5331 (N_5331,N_800,N_1920);
and U5332 (N_5332,N_1810,N_4905);
or U5333 (N_5333,N_926,N_2560);
nand U5334 (N_5334,N_485,N_2032);
and U5335 (N_5335,N_4204,N_3413);
or U5336 (N_5336,N_2311,N_1560);
nor U5337 (N_5337,N_4362,N_4591);
and U5338 (N_5338,N_372,N_3031);
nand U5339 (N_5339,N_4021,N_3660);
nand U5340 (N_5340,N_2844,N_2107);
xor U5341 (N_5341,N_4144,N_3955);
nand U5342 (N_5342,N_3543,N_1527);
and U5343 (N_5343,N_2046,N_1009);
nor U5344 (N_5344,N_2646,N_3818);
and U5345 (N_5345,N_2384,N_4646);
or U5346 (N_5346,N_141,N_3708);
nor U5347 (N_5347,N_2917,N_2472);
and U5348 (N_5348,N_4230,N_2886);
or U5349 (N_5349,N_3040,N_345);
nor U5350 (N_5350,N_4499,N_3602);
and U5351 (N_5351,N_4034,N_1163);
nand U5352 (N_5352,N_3028,N_2385);
and U5353 (N_5353,N_412,N_2218);
and U5354 (N_5354,N_4974,N_2272);
or U5355 (N_5355,N_1992,N_3651);
nand U5356 (N_5356,N_1567,N_4086);
xor U5357 (N_5357,N_2747,N_554);
and U5358 (N_5358,N_96,N_4149);
nor U5359 (N_5359,N_649,N_1280);
or U5360 (N_5360,N_545,N_3058);
and U5361 (N_5361,N_3975,N_706);
and U5362 (N_5362,N_3505,N_1834);
nand U5363 (N_5363,N_320,N_2113);
and U5364 (N_5364,N_3134,N_887);
xor U5365 (N_5365,N_3639,N_1977);
nor U5366 (N_5366,N_2374,N_1138);
nor U5367 (N_5367,N_3675,N_350);
or U5368 (N_5368,N_291,N_3819);
nor U5369 (N_5369,N_1300,N_3441);
xor U5370 (N_5370,N_1371,N_3865);
or U5371 (N_5371,N_2131,N_92);
nand U5372 (N_5372,N_130,N_1392);
nand U5373 (N_5373,N_151,N_1058);
and U5374 (N_5374,N_2692,N_2386);
or U5375 (N_5375,N_3945,N_3451);
nand U5376 (N_5376,N_4675,N_2875);
and U5377 (N_5377,N_4527,N_3235);
and U5378 (N_5378,N_1500,N_2732);
nor U5379 (N_5379,N_1968,N_4800);
or U5380 (N_5380,N_84,N_2087);
nor U5381 (N_5381,N_4508,N_3131);
nand U5382 (N_5382,N_2520,N_3118);
nor U5383 (N_5383,N_2859,N_1829);
or U5384 (N_5384,N_3716,N_495);
nor U5385 (N_5385,N_4750,N_4634);
nor U5386 (N_5386,N_4536,N_1703);
nor U5387 (N_5387,N_2572,N_664);
or U5388 (N_5388,N_4644,N_1791);
nand U5389 (N_5389,N_3712,N_4376);
nor U5390 (N_5390,N_4718,N_1745);
nand U5391 (N_5391,N_3921,N_1216);
or U5392 (N_5392,N_1828,N_4609);
and U5393 (N_5393,N_4100,N_3080);
xnor U5394 (N_5394,N_3152,N_2408);
nand U5395 (N_5395,N_3834,N_3774);
nand U5396 (N_5396,N_162,N_4524);
or U5397 (N_5397,N_3587,N_1613);
nand U5398 (N_5398,N_890,N_3676);
nand U5399 (N_5399,N_822,N_1943);
nand U5400 (N_5400,N_325,N_3200);
nor U5401 (N_5401,N_52,N_1636);
nor U5402 (N_5402,N_2526,N_767);
nand U5403 (N_5403,N_23,N_352);
nor U5404 (N_5404,N_2043,N_899);
xor U5405 (N_5405,N_2565,N_3915);
or U5406 (N_5406,N_488,N_798);
nand U5407 (N_5407,N_817,N_4000);
or U5408 (N_5408,N_1072,N_924);
and U5409 (N_5409,N_1444,N_2713);
xnor U5410 (N_5410,N_4673,N_3601);
nor U5411 (N_5411,N_2751,N_2602);
nand U5412 (N_5412,N_4848,N_2954);
and U5413 (N_5413,N_3637,N_218);
and U5414 (N_5414,N_1647,N_3475);
nor U5415 (N_5415,N_4730,N_4988);
nand U5416 (N_5416,N_4054,N_3702);
nor U5417 (N_5417,N_1750,N_500);
nand U5418 (N_5418,N_146,N_4950);
nand U5419 (N_5419,N_399,N_2716);
and U5420 (N_5420,N_4681,N_1219);
nand U5421 (N_5421,N_2097,N_4270);
or U5422 (N_5422,N_4959,N_3075);
nand U5423 (N_5423,N_3051,N_178);
and U5424 (N_5424,N_2694,N_3733);
nor U5425 (N_5425,N_4405,N_3242);
xnor U5426 (N_5426,N_2807,N_3705);
nor U5427 (N_5427,N_2814,N_4299);
nand U5428 (N_5428,N_634,N_4594);
and U5429 (N_5429,N_2613,N_3683);
nor U5430 (N_5430,N_4398,N_2708);
nor U5431 (N_5431,N_2029,N_3673);
or U5432 (N_5432,N_223,N_4153);
and U5433 (N_5433,N_879,N_4184);
and U5434 (N_5434,N_290,N_4386);
nand U5435 (N_5435,N_4518,N_3012);
nor U5436 (N_5436,N_3553,N_1012);
and U5437 (N_5437,N_1166,N_2040);
xor U5438 (N_5438,N_907,N_4018);
and U5439 (N_5439,N_1454,N_2805);
xnor U5440 (N_5440,N_4643,N_920);
nand U5441 (N_5441,N_2042,N_4278);
or U5442 (N_5442,N_951,N_3959);
nor U5443 (N_5443,N_1995,N_4031);
nand U5444 (N_5444,N_3965,N_2335);
nand U5445 (N_5445,N_4345,N_2973);
or U5446 (N_5446,N_3307,N_949);
or U5447 (N_5447,N_2276,N_1611);
or U5448 (N_5448,N_1506,N_3285);
nor U5449 (N_5449,N_3232,N_1934);
nor U5450 (N_5450,N_1398,N_4232);
nor U5451 (N_5451,N_2208,N_676);
nor U5452 (N_5452,N_4991,N_2501);
nor U5453 (N_5453,N_2467,N_2354);
nand U5454 (N_5454,N_2416,N_1876);
nand U5455 (N_5455,N_1853,N_83);
or U5456 (N_5456,N_1125,N_3219);
or U5457 (N_5457,N_1869,N_4048);
or U5458 (N_5458,N_3054,N_4147);
and U5459 (N_5459,N_3518,N_2648);
nor U5460 (N_5460,N_465,N_4691);
and U5461 (N_5461,N_275,N_560);
or U5462 (N_5462,N_54,N_2031);
or U5463 (N_5463,N_250,N_4784);
nand U5464 (N_5464,N_892,N_4306);
nand U5465 (N_5465,N_2285,N_1727);
and U5466 (N_5466,N_3725,N_2792);
nand U5467 (N_5467,N_1178,N_2075);
nor U5468 (N_5468,N_3142,N_2663);
or U5469 (N_5469,N_3605,N_316);
nand U5470 (N_5470,N_1858,N_1237);
nand U5471 (N_5471,N_470,N_1143);
and U5472 (N_5472,N_4209,N_2905);
or U5473 (N_5473,N_2280,N_2454);
or U5474 (N_5474,N_1900,N_4678);
nand U5475 (N_5475,N_638,N_1015);
and U5476 (N_5476,N_2573,N_1627);
or U5477 (N_5477,N_747,N_2400);
xor U5478 (N_5478,N_2666,N_4549);
or U5479 (N_5479,N_3703,N_1090);
and U5480 (N_5480,N_3607,N_6);
or U5481 (N_5481,N_2273,N_3806);
nand U5482 (N_5482,N_1462,N_2793);
nand U5483 (N_5483,N_2668,N_2604);
and U5484 (N_5484,N_2452,N_2206);
nor U5485 (N_5485,N_3718,N_1605);
or U5486 (N_5486,N_3952,N_4666);
and U5487 (N_5487,N_810,N_2307);
nand U5488 (N_5488,N_4554,N_2336);
and U5489 (N_5489,N_1440,N_4463);
nand U5490 (N_5490,N_1193,N_850);
nor U5491 (N_5491,N_170,N_4496);
or U5492 (N_5492,N_3125,N_3063);
nor U5493 (N_5493,N_4173,N_2955);
and U5494 (N_5494,N_3049,N_2904);
and U5495 (N_5495,N_3029,N_4005);
or U5496 (N_5496,N_478,N_39);
nand U5497 (N_5497,N_733,N_925);
nor U5498 (N_5498,N_2164,N_3107);
and U5499 (N_5499,N_2081,N_4568);
nor U5500 (N_5500,N_4200,N_915);
and U5501 (N_5501,N_4558,N_1945);
or U5502 (N_5502,N_4235,N_2391);
or U5503 (N_5503,N_2158,N_3007);
or U5504 (N_5504,N_1311,N_3971);
nand U5505 (N_5505,N_1267,N_3014);
nand U5506 (N_5506,N_1218,N_2978);
nor U5507 (N_5507,N_2735,N_670);
xnor U5508 (N_5508,N_2784,N_4817);
nand U5509 (N_5509,N_3292,N_3377);
nand U5510 (N_5510,N_4272,N_3414);
nand U5511 (N_5511,N_3748,N_4325);
or U5512 (N_5512,N_783,N_524);
and U5513 (N_5513,N_1115,N_1485);
nor U5514 (N_5514,N_2558,N_3159);
nand U5515 (N_5515,N_4255,N_1114);
nor U5516 (N_5516,N_2152,N_3531);
nand U5517 (N_5517,N_4214,N_1585);
or U5518 (N_5518,N_3388,N_410);
and U5519 (N_5519,N_4241,N_567);
or U5520 (N_5520,N_1382,N_4379);
and U5521 (N_5521,N_62,N_1973);
xor U5522 (N_5522,N_3709,N_1278);
nor U5523 (N_5523,N_2951,N_2527);
and U5524 (N_5524,N_4435,N_34);
nor U5525 (N_5525,N_238,N_1477);
nor U5526 (N_5526,N_2302,N_911);
and U5527 (N_5527,N_2072,N_3195);
or U5528 (N_5528,N_1344,N_3093);
or U5529 (N_5529,N_4290,N_1767);
and U5530 (N_5530,N_1825,N_438);
and U5531 (N_5531,N_3224,N_2549);
and U5532 (N_5532,N_444,N_2634);
xnor U5533 (N_5533,N_3994,N_1846);
or U5534 (N_5534,N_3535,N_4038);
xor U5535 (N_5535,N_3308,N_2849);
nand U5536 (N_5536,N_1046,N_1602);
and U5537 (N_5537,N_3847,N_1783);
nor U5538 (N_5538,N_1087,N_1122);
or U5539 (N_5539,N_511,N_1529);
or U5540 (N_5540,N_3590,N_340);
and U5541 (N_5541,N_928,N_2191);
nand U5542 (N_5542,N_3385,N_3532);
and U5543 (N_5543,N_1687,N_3887);
nand U5544 (N_5544,N_261,N_3977);
nand U5545 (N_5545,N_3306,N_155);
or U5546 (N_5546,N_3470,N_624);
nor U5547 (N_5547,N_2684,N_4685);
and U5548 (N_5548,N_2949,N_1980);
and U5549 (N_5549,N_4148,N_4943);
and U5550 (N_5550,N_3667,N_2994);
and U5551 (N_5551,N_2980,N_9);
nand U5552 (N_5552,N_1584,N_3947);
nand U5553 (N_5553,N_587,N_1060);
nor U5554 (N_5554,N_1568,N_3541);
or U5555 (N_5555,N_3041,N_1547);
xnor U5556 (N_5556,N_339,N_4892);
and U5557 (N_5557,N_3816,N_1097);
nand U5558 (N_5558,N_2127,N_867);
or U5559 (N_5559,N_1517,N_546);
or U5560 (N_5560,N_4116,N_902);
or U5561 (N_5561,N_3513,N_1606);
or U5562 (N_5562,N_4289,N_998);
nand U5563 (N_5563,N_1084,N_4543);
xnor U5564 (N_5564,N_1383,N_3630);
nand U5565 (N_5565,N_1553,N_105);
nand U5566 (N_5566,N_1597,N_3905);
nand U5567 (N_5567,N_693,N_4427);
and U5568 (N_5568,N_4202,N_4921);
nand U5569 (N_5569,N_2404,N_66);
nand U5570 (N_5570,N_4227,N_3119);
or U5571 (N_5571,N_2288,N_543);
xnor U5572 (N_5572,N_4579,N_3309);
nor U5573 (N_5573,N_4583,N_422);
nor U5574 (N_5574,N_2655,N_1307);
nand U5575 (N_5575,N_725,N_2612);
xnor U5576 (N_5576,N_326,N_3508);
or U5577 (N_5577,N_2674,N_4459);
or U5578 (N_5578,N_588,N_4716);
or U5579 (N_5579,N_3104,N_943);
nor U5580 (N_5580,N_121,N_164);
nand U5581 (N_5581,N_999,N_994);
nand U5582 (N_5582,N_1499,N_1755);
nand U5583 (N_5583,N_4642,N_742);
and U5584 (N_5584,N_622,N_4861);
nand U5585 (N_5585,N_3582,N_3374);
nor U5586 (N_5586,N_3942,N_2274);
and U5587 (N_5587,N_1991,N_227);
nand U5588 (N_5588,N_2283,N_1837);
and U5589 (N_5589,N_611,N_124);
nor U5590 (N_5590,N_116,N_3001);
or U5591 (N_5591,N_2940,N_1967);
nor U5592 (N_5592,N_4927,N_1578);
nor U5593 (N_5593,N_4249,N_2216);
nor U5594 (N_5594,N_4343,N_3048);
and U5595 (N_5595,N_1415,N_2470);
and U5596 (N_5596,N_508,N_4687);
nor U5597 (N_5597,N_1190,N_35);
or U5598 (N_5598,N_2293,N_41);
xor U5599 (N_5599,N_3875,N_3606);
nor U5600 (N_5600,N_4951,N_3393);
nor U5601 (N_5601,N_4097,N_2035);
nor U5602 (N_5602,N_4157,N_3979);
or U5603 (N_5603,N_1161,N_2913);
nor U5604 (N_5604,N_3581,N_2936);
and U5605 (N_5605,N_3394,N_4689);
nand U5606 (N_5606,N_1358,N_2727);
nor U5607 (N_5607,N_1147,N_1430);
xor U5608 (N_5608,N_464,N_2442);
nand U5609 (N_5609,N_3801,N_4067);
and U5610 (N_5610,N_912,N_3892);
nand U5611 (N_5611,N_138,N_3641);
and U5612 (N_5612,N_4205,N_4751);
nor U5613 (N_5613,N_3528,N_4367);
or U5614 (N_5614,N_2292,N_3752);
nor U5615 (N_5615,N_1782,N_2045);
nor U5616 (N_5616,N_4357,N_2162);
and U5617 (N_5617,N_4416,N_3849);
nor U5618 (N_5618,N_801,N_909);
and U5619 (N_5619,N_172,N_505);
or U5620 (N_5620,N_3677,N_4721);
or U5621 (N_5621,N_4228,N_1194);
and U5622 (N_5622,N_933,N_3539);
or U5623 (N_5623,N_3208,N_1575);
and U5624 (N_5624,N_2016,N_3365);
nor U5625 (N_5625,N_3953,N_3302);
or U5626 (N_5626,N_2907,N_2439);
xnor U5627 (N_5627,N_4368,N_1684);
nor U5628 (N_5628,N_234,N_1906);
and U5629 (N_5629,N_4009,N_2395);
xnor U5630 (N_5630,N_2870,N_3980);
and U5631 (N_5631,N_2869,N_4555);
nor U5632 (N_5632,N_1706,N_2630);
or U5633 (N_5633,N_4471,N_3679);
nor U5634 (N_5634,N_108,N_1718);
and U5635 (N_5635,N_182,N_4922);
nand U5636 (N_5636,N_3678,N_3968);
or U5637 (N_5637,N_4364,N_3739);
and U5638 (N_5638,N_2872,N_2952);
nand U5639 (N_5639,N_797,N_600);
and U5640 (N_5640,N_2878,N_3511);
and U5641 (N_5641,N_4674,N_1789);
and U5642 (N_5642,N_4226,N_1850);
nor U5643 (N_5643,N_11,N_979);
xnor U5644 (N_5644,N_4589,N_3317);
and U5645 (N_5645,N_2105,N_48);
nand U5646 (N_5646,N_945,N_3415);
nand U5647 (N_5647,N_2748,N_1426);
or U5648 (N_5648,N_3085,N_2073);
nand U5649 (N_5649,N_373,N_4652);
nand U5650 (N_5650,N_3255,N_370);
xnor U5651 (N_5651,N_1183,N_2861);
or U5652 (N_5652,N_496,N_276);
and U5653 (N_5653,N_2810,N_4841);
nor U5654 (N_5654,N_60,N_3941);
or U5655 (N_5655,N_95,N_1614);
or U5656 (N_5656,N_3813,N_4074);
and U5657 (N_5657,N_700,N_4303);
nand U5658 (N_5658,N_2997,N_2881);
nand U5659 (N_5659,N_3880,N_1378);
nand U5660 (N_5660,N_4360,N_3579);
and U5661 (N_5661,N_729,N_1364);
nor U5662 (N_5662,N_3468,N_917);
and U5663 (N_5663,N_601,N_3450);
nand U5664 (N_5664,N_2356,N_2971);
or U5665 (N_5665,N_1151,N_3907);
and U5666 (N_5666,N_3567,N_3088);
nor U5667 (N_5667,N_206,N_4777);
nand U5668 (N_5668,N_4089,N_1221);
nand U5669 (N_5669,N_2996,N_1849);
nand U5670 (N_5670,N_4620,N_4441);
and U5671 (N_5671,N_2141,N_2357);
or U5672 (N_5672,N_2833,N_1327);
nand U5673 (N_5673,N_1561,N_3916);
nor U5674 (N_5674,N_1804,N_3379);
xnor U5675 (N_5675,N_374,N_3698);
nor U5676 (N_5676,N_1497,N_3904);
nand U5677 (N_5677,N_4632,N_3599);
nor U5678 (N_5678,N_1413,N_1495);
xnor U5679 (N_5679,N_173,N_4668);
nor U5680 (N_5680,N_1481,N_3167);
and U5681 (N_5681,N_619,N_4900);
or U5682 (N_5682,N_2561,N_3409);
and U5683 (N_5683,N_4152,N_1963);
or U5684 (N_5684,N_1411,N_2974);
nor U5685 (N_5685,N_1545,N_574);
nor U5686 (N_5686,N_1051,N_512);
nor U5687 (N_5687,N_1646,N_1152);
nand U5688 (N_5688,N_2514,N_3759);
and U5689 (N_5689,N_840,N_4679);
and U5690 (N_5690,N_94,N_2963);
nand U5691 (N_5691,N_4865,N_2968);
nand U5692 (N_5692,N_4256,N_713);
nor U5693 (N_5693,N_694,N_4891);
or U5694 (N_5694,N_1565,N_3149);
nand U5695 (N_5695,N_255,N_4775);
nand U5696 (N_5696,N_3802,N_4340);
nor U5697 (N_5697,N_4311,N_4531);
and U5698 (N_5698,N_1588,N_97);
or U5699 (N_5699,N_4901,N_3672);
and U5700 (N_5700,N_2414,N_591);
or U5701 (N_5701,N_3580,N_4285);
or U5702 (N_5702,N_4995,N_1102);
and U5703 (N_5703,N_1532,N_262);
and U5704 (N_5704,N_993,N_2226);
nor U5705 (N_5705,N_2421,N_3783);
and U5706 (N_5706,N_502,N_1353);
and U5707 (N_5707,N_3699,N_4274);
or U5708 (N_5708,N_3342,N_1442);
nand U5709 (N_5709,N_1038,N_2847);
and U5710 (N_5710,N_3132,N_1270);
or U5711 (N_5711,N_4693,N_1880);
or U5712 (N_5712,N_80,N_2961);
xnor U5713 (N_5713,N_1419,N_3037);
or U5714 (N_5714,N_2928,N_4912);
and U5715 (N_5715,N_1314,N_4837);
nand U5716 (N_5716,N_2908,N_1493);
nor U5717 (N_5717,N_86,N_2108);
or U5718 (N_5718,N_2806,N_4765);
nand U5719 (N_5719,N_4296,N_2920);
nand U5720 (N_5720,N_2323,N_3175);
or U5721 (N_5721,N_277,N_4396);
xor U5722 (N_5722,N_3349,N_1546);
xor U5723 (N_5723,N_2415,N_2159);
nand U5724 (N_5724,N_4046,N_2538);
nor U5725 (N_5725,N_3402,N_12);
or U5726 (N_5726,N_1922,N_1975);
or U5727 (N_5727,N_3141,N_1424);
or U5728 (N_5728,N_1171,N_3331);
nand U5729 (N_5729,N_3127,N_1423);
and U5730 (N_5730,N_4073,N_328);
nor U5731 (N_5731,N_3992,N_4502);
nor U5732 (N_5732,N_1663,N_3644);
and U5733 (N_5733,N_4059,N_1870);
or U5734 (N_5734,N_2678,N_2092);
nand U5735 (N_5735,N_3656,N_4037);
nor U5736 (N_5736,N_1212,N_1590);
or U5737 (N_5737,N_4874,N_4699);
and U5738 (N_5738,N_2379,N_3883);
xnor U5739 (N_5739,N_2842,N_2372);
nand U5740 (N_5740,N_2509,N_4354);
nand U5741 (N_5741,N_3572,N_1690);
and U5742 (N_5742,N_2193,N_1410);
or U5743 (N_5743,N_3958,N_336);
or U5744 (N_5744,N_4972,N_785);
nor U5745 (N_5745,N_2053,N_3749);
nor U5746 (N_5746,N_1817,N_1707);
xor U5747 (N_5747,N_3778,N_1536);
or U5748 (N_5748,N_660,N_2360);
or U5749 (N_5749,N_3408,N_1185);
and U5750 (N_5750,N_3002,N_4932);
nand U5751 (N_5751,N_2964,N_448);
or U5752 (N_5752,N_4422,N_2213);
nor U5753 (N_5753,N_873,N_3527);
nor U5754 (N_5754,N_3382,N_535);
nand U5755 (N_5755,N_2468,N_1366);
nor U5756 (N_5756,N_1335,N_4969);
nand U5757 (N_5757,N_646,N_1775);
nor U5758 (N_5758,N_3493,N_1197);
nor U5759 (N_5759,N_3803,N_2768);
or U5760 (N_5760,N_3240,N_1983);
nor U5761 (N_5761,N_3741,N_527);
or U5762 (N_5762,N_4489,N_4447);
xor U5763 (N_5763,N_3615,N_168);
nand U5764 (N_5764,N_884,N_2672);
xnor U5765 (N_5765,N_1473,N_1023);
and U5766 (N_5766,N_1998,N_405);
xor U5767 (N_5767,N_207,N_228);
xnor U5768 (N_5768,N_1338,N_3189);
or U5769 (N_5769,N_3982,N_4635);
nand U5770 (N_5770,N_2464,N_1050);
xor U5771 (N_5771,N_1847,N_1351);
xnor U5772 (N_5772,N_3130,N_2611);
or U5773 (N_5773,N_4433,N_836);
nor U5774 (N_5774,N_1550,N_1490);
and U5775 (N_5775,N_3985,N_1106);
nand U5776 (N_5776,N_1908,N_2038);
or U5777 (N_5777,N_2709,N_3375);
xnor U5778 (N_5778,N_4638,N_3584);
and U5779 (N_5779,N_3569,N_3171);
nor U5780 (N_5780,N_1372,N_833);
or U5781 (N_5781,N_4628,N_3121);
and U5782 (N_5782,N_3700,N_1359);
or U5783 (N_5783,N_3272,N_2287);
nand U5784 (N_5784,N_2945,N_1824);
or U5785 (N_5785,N_1450,N_1373);
nand U5786 (N_5786,N_4356,N_1245);
nand U5787 (N_5787,N_424,N_605);
and U5788 (N_5788,N_819,N_117);
or U5789 (N_5789,N_3223,N_3600);
or U5790 (N_5790,N_4657,N_4529);
and U5791 (N_5791,N_921,N_4759);
and U5792 (N_5792,N_3123,N_3767);
and U5793 (N_5793,N_1744,N_613);
or U5794 (N_5794,N_3890,N_4439);
nor U5795 (N_5795,N_3449,N_4547);
nor U5796 (N_5796,N_4963,N_4925);
nor U5797 (N_5797,N_2911,N_2901);
nor U5798 (N_5798,N_2412,N_1881);
and U5799 (N_5799,N_1049,N_375);
nor U5800 (N_5800,N_2953,N_2893);
nor U5801 (N_5801,N_1976,N_4882);
nor U5802 (N_5802,N_1962,N_93);
and U5803 (N_5803,N_3564,N_3264);
or U5804 (N_5804,N_4649,N_1073);
nand U5805 (N_5805,N_3148,N_4790);
and U5806 (N_5806,N_904,N_2828);
or U5807 (N_5807,N_2532,N_4744);
or U5808 (N_5808,N_651,N_1557);
or U5809 (N_5809,N_3868,N_688);
nor U5810 (N_5810,N_2078,N_4484);
nor U5811 (N_5811,N_578,N_2011);
nand U5812 (N_5812,N_1019,N_453);
or U5813 (N_5813,N_4916,N_371);
nor U5814 (N_5814,N_2826,N_1302);
nor U5815 (N_5815,N_4849,N_1840);
xnor U5816 (N_5816,N_409,N_2451);
nand U5817 (N_5817,N_2300,N_3932);
and U5818 (N_5818,N_1294,N_1214);
nand U5819 (N_5819,N_3633,N_2882);
xnor U5820 (N_5820,N_1693,N_938);
and U5821 (N_5821,N_3146,N_4856);
and U5822 (N_5822,N_91,N_4160);
and U5823 (N_5823,N_2899,N_4798);
nand U5824 (N_5824,N_2638,N_4483);
nor U5825 (N_5825,N_4934,N_376);
and U5826 (N_5826,N_3597,N_3856);
or U5827 (N_5827,N_3763,N_299);
and U5828 (N_5828,N_2462,N_2361);
or U5829 (N_5829,N_3895,N_3491);
or U5830 (N_5830,N_1298,N_2628);
or U5831 (N_5831,N_4816,N_385);
xnor U5832 (N_5832,N_1844,N_160);
nand U5833 (N_5833,N_2513,N_4613);
and U5834 (N_5834,N_1008,N_1966);
or U5835 (N_5835,N_3318,N_4151);
nor U5836 (N_5836,N_3324,N_1814);
nor U5837 (N_5837,N_948,N_3078);
or U5838 (N_5838,N_4472,N_1672);
xor U5839 (N_5839,N_2717,N_4904);
xnor U5840 (N_5840,N_2765,N_630);
or U5841 (N_5841,N_1762,N_1518);
xnor U5842 (N_5842,N_3020,N_869);
or U5843 (N_5843,N_3482,N_4295);
nor U5844 (N_5844,N_4611,N_813);
nor U5845 (N_5845,N_1747,N_2714);
xor U5846 (N_5846,N_4002,N_2938);
nor U5847 (N_5847,N_1431,N_666);
xnor U5848 (N_5848,N_4164,N_1735);
nand U5849 (N_5849,N_1912,N_2236);
nor U5850 (N_5850,N_718,N_2327);
xnor U5851 (N_5851,N_1509,N_1658);
or U5852 (N_5852,N_351,N_4676);
nor U5853 (N_5853,N_3151,N_358);
nand U5854 (N_5854,N_1000,N_3635);
or U5855 (N_5855,N_3188,N_1256);
or U5856 (N_5856,N_2498,N_4365);
xor U5857 (N_5857,N_3594,N_4101);
nor U5858 (N_5858,N_3471,N_3286);
nor U5859 (N_5859,N_197,N_644);
and U5860 (N_5860,N_2375,N_1808);
xnor U5861 (N_5861,N_3003,N_2988);
nand U5862 (N_5862,N_1362,N_2260);
or U5863 (N_5863,N_3202,N_53);
nor U5864 (N_5864,N_4707,N_402);
nand U5865 (N_5865,N_3311,N_758);
nor U5866 (N_5866,N_4975,N_415);
nand U5867 (N_5867,N_3254,N_2528);
and U5868 (N_5868,N_685,N_341);
nand U5869 (N_5869,N_1769,N_2480);
or U5870 (N_5870,N_242,N_4879);
nand U5871 (N_5871,N_98,N_1759);
and U5872 (N_5872,N_3831,N_1345);
or U5873 (N_5873,N_1877,N_3912);
nor U5874 (N_5874,N_2458,N_633);
nand U5875 (N_5875,N_2083,N_2898);
xor U5876 (N_5876,N_2983,N_3727);
nand U5877 (N_5877,N_3751,N_2008);
or U5878 (N_5878,N_2202,N_4626);
nor U5879 (N_5879,N_2786,N_1195);
or U5880 (N_5880,N_4339,N_3762);
and U5881 (N_5881,N_380,N_2787);
nor U5882 (N_5882,N_1801,N_4541);
or U5883 (N_5883,N_1576,N_936);
nand U5884 (N_5884,N_4767,N_1577);
or U5885 (N_5885,N_4029,N_3872);
or U5886 (N_5886,N_1921,N_3779);
or U5887 (N_5887,N_473,N_4273);
nand U5888 (N_5888,N_3598,N_990);
and U5889 (N_5889,N_3997,N_4062);
and U5890 (N_5890,N_724,N_2650);
and U5891 (N_5891,N_2056,N_910);
nor U5892 (N_5892,N_3053,N_2203);
or U5893 (N_5893,N_662,N_1464);
and U5894 (N_5894,N_3420,N_4293);
or U5895 (N_5895,N_4167,N_3542);
or U5896 (N_5896,N_2696,N_515);
and U5897 (N_5897,N_2824,N_2535);
xnor U5898 (N_5898,N_4570,N_4334);
and U5899 (N_5899,N_528,N_1520);
or U5900 (N_5900,N_1069,N_547);
and U5901 (N_5901,N_874,N_4338);
or U5902 (N_5902,N_805,N_2592);
nand U5903 (N_5903,N_4443,N_1935);
or U5904 (N_5904,N_122,N_2972);
nand U5905 (N_5905,N_968,N_1239);
nand U5906 (N_5906,N_391,N_2811);
nor U5907 (N_5907,N_3072,N_3346);
and U5908 (N_5908,N_2618,N_3344);
nand U5909 (N_5909,N_2960,N_1026);
and U5910 (N_5910,N_2536,N_4406);
and U5911 (N_5911,N_3503,N_1795);
and U5912 (N_5912,N_3263,N_3177);
or U5913 (N_5913,N_1063,N_553);
nor U5914 (N_5914,N_930,N_1181);
nand U5915 (N_5915,N_2021,N_3844);
or U5916 (N_5916,N_452,N_201);
nor U5917 (N_5917,N_1939,N_1438);
xnor U5918 (N_5918,N_1955,N_3099);
nor U5919 (N_5919,N_4698,N_628);
nand U5920 (N_5920,N_3462,N_3395);
nor U5921 (N_5921,N_3536,N_3026);
or U5922 (N_5922,N_3366,N_2957);
nand U5923 (N_5923,N_1139,N_2587);
nand U5924 (N_5924,N_2333,N_1622);
and U5925 (N_5925,N_4917,N_1264);
nor U5926 (N_5926,N_3207,N_3372);
nand U5927 (N_5927,N_4627,N_2114);
nand U5928 (N_5928,N_484,N_2147);
or U5929 (N_5929,N_471,N_1699);
or U5930 (N_5930,N_4618,N_965);
nor U5931 (N_5931,N_2012,N_1036);
nand U5932 (N_5932,N_586,N_1133);
nand U5933 (N_5933,N_1208,N_4003);
or U5934 (N_5934,N_824,N_7);
or U5935 (N_5935,N_4252,N_1196);
nand U5936 (N_5936,N_3206,N_4663);
nand U5937 (N_5937,N_2962,N_2063);
or U5938 (N_5938,N_3330,N_1308);
nor U5939 (N_5939,N_3855,N_4738);
nand U5940 (N_5940,N_3231,N_4491);
and U5941 (N_5941,N_3214,N_147);
nand U5942 (N_5942,N_2295,N_3496);
or U5943 (N_5943,N_969,N_2268);
or U5944 (N_5944,N_3400,N_625);
or U5945 (N_5945,N_3610,N_4719);
nor U5946 (N_5946,N_2422,N_248);
and U5947 (N_5947,N_1910,N_1766);
and U5948 (N_5948,N_2989,N_2044);
and U5949 (N_5949,N_1128,N_3417);
nand U5950 (N_5950,N_2515,N_3488);
nor U5951 (N_5951,N_4525,N_306);
and U5952 (N_5952,N_2902,N_1476);
xor U5953 (N_5953,N_4349,N_4781);
nand U5954 (N_5954,N_918,N_3249);
nor U5955 (N_5955,N_1748,N_4363);
nand U5956 (N_5956,N_3688,N_631);
nor U5957 (N_5957,N_2689,N_1691);
xnor U5958 (N_5958,N_2516,N_4462);
and U5959 (N_5959,N_726,N_1254);
xor U5960 (N_5960,N_3247,N_2392);
nand U5961 (N_5961,N_4999,N_1443);
or U5962 (N_5962,N_4684,N_893);
or U5963 (N_5963,N_1790,N_4424);
or U5964 (N_5964,N_847,N_2039);
nand U5965 (N_5965,N_3357,N_2540);
nand U5966 (N_5966,N_841,N_1809);
or U5967 (N_5967,N_4400,N_4538);
nor U5968 (N_5968,N_4686,N_210);
or U5969 (N_5969,N_3859,N_580);
nand U5970 (N_5970,N_684,N_3900);
and U5971 (N_5971,N_3410,N_4923);
nor U5972 (N_5972,N_796,N_1805);
and U5973 (N_5973,N_2344,N_1842);
or U5974 (N_5974,N_1957,N_4871);
nor U5975 (N_5975,N_3034,N_3713);
or U5976 (N_5976,N_359,N_3918);
or U5977 (N_5977,N_2249,N_701);
nor U5978 (N_5978,N_829,N_2903);
or U5979 (N_5979,N_4898,N_2855);
and U5980 (N_5980,N_3433,N_4712);
nand U5981 (N_5981,N_4515,N_870);
and U5982 (N_5982,N_2351,N_2475);
nand U5983 (N_5983,N_296,N_315);
nor U5984 (N_5984,N_2013,N_1563);
or U5985 (N_5985,N_537,N_1120);
nand U5986 (N_5986,N_1712,N_282);
nor U5987 (N_5987,N_809,N_2606);
and U5988 (N_5988,N_2393,N_2756);
or U5989 (N_5989,N_1863,N_4965);
and U5990 (N_5990,N_3244,N_179);
and U5991 (N_5991,N_3024,N_426);
xor U5992 (N_5992,N_2002,N_3291);
nor U5993 (N_5993,N_1841,N_552);
or U5994 (N_5994,N_1108,N_1685);
or U5995 (N_5995,N_191,N_3879);
and U5996 (N_5996,N_4936,N_3238);
nor U5997 (N_5997,N_2495,N_2330);
and U5998 (N_5998,N_3760,N_287);
nand U5999 (N_5999,N_4702,N_4158);
and U6000 (N_6000,N_4504,N_1600);
nor U6001 (N_6001,N_3516,N_2346);
and U6002 (N_6002,N_3864,N_3661);
nor U6003 (N_6003,N_2918,N_459);
or U6004 (N_6004,N_2322,N_1331);
nand U6005 (N_6005,N_1210,N_4446);
nor U6006 (N_6006,N_679,N_2499);
nand U6007 (N_6007,N_501,N_3797);
xnor U6008 (N_6008,N_1763,N_506);
or U6009 (N_6009,N_167,N_2649);
nor U6010 (N_6010,N_4710,N_1594);
nand U6011 (N_6011,N_2220,N_2500);
or U6012 (N_6012,N_2577,N_2715);
nor U6013 (N_6013,N_461,N_434);
and U6014 (N_6014,N_2066,N_781);
and U6015 (N_6015,N_2240,N_1919);
nand U6016 (N_6016,N_3670,N_1376);
xnor U6017 (N_6017,N_3506,N_2453);
and U6018 (N_6018,N_3562,N_844);
nand U6019 (N_6019,N_4480,N_2817);
or U6020 (N_6020,N_1215,N_51);
and U6021 (N_6021,N_1421,N_510);
and U6022 (N_6022,N_1228,N_145);
nand U6023 (N_6023,N_442,N_260);
nor U6024 (N_6024,N_2741,N_3938);
or U6025 (N_6025,N_3201,N_4434);
nand U6026 (N_6026,N_3150,N_4473);
or U6027 (N_6027,N_2586,N_59);
nand U6028 (N_6028,N_4081,N_2977);
and U6029 (N_6029,N_2835,N_4485);
or U6030 (N_6030,N_3293,N_3636);
or U6031 (N_6031,N_983,N_3566);
nand U6032 (N_6032,N_2460,N_1742);
or U6033 (N_6033,N_623,N_8);
nor U6034 (N_6034,N_2659,N_4347);
and U6035 (N_6035,N_3005,N_3351);
nor U6036 (N_6036,N_3198,N_1489);
or U6037 (N_6037,N_2508,N_2764);
xnor U6038 (N_6038,N_3559,N_1889);
nand U6039 (N_6039,N_991,N_2897);
nand U6040 (N_6040,N_539,N_419);
nor U6041 (N_6041,N_786,N_4743);
nand U6042 (N_6042,N_4537,N_1933);
nand U6043 (N_6043,N_2089,N_386);
xnor U6044 (N_6044,N_3545,N_4027);
xor U6045 (N_6045,N_27,N_1717);
xor U6046 (N_6046,N_161,N_1394);
and U6047 (N_6047,N_2865,N_1232);
nand U6048 (N_6048,N_4601,N_1369);
and U6049 (N_6049,N_347,N_3447);
and U6050 (N_6050,N_4827,N_4793);
or U6051 (N_6051,N_1710,N_3893);
nor U6052 (N_6052,N_2058,N_2593);
or U6053 (N_6053,N_3857,N_2776);
xnor U6054 (N_6054,N_3561,N_330);
nand U6055 (N_6055,N_2290,N_1914);
and U6056 (N_6056,N_1064,N_4218);
or U6057 (N_6057,N_530,N_3147);
nor U6058 (N_6058,N_463,N_4835);
and U6059 (N_6059,N_1765,N_4683);
nor U6060 (N_6060,N_4134,N_3548);
or U6061 (N_6061,N_2449,N_2699);
nor U6062 (N_6062,N_4513,N_2596);
nor U6063 (N_6063,N_4682,N_3866);
or U6064 (N_6064,N_677,N_4788);
nand U6065 (N_6065,N_523,N_3459);
or U6066 (N_6066,N_2250,N_2900);
xnor U6067 (N_6067,N_37,N_3719);
and U6068 (N_6068,N_2054,N_2255);
nor U6069 (N_6069,N_1420,N_4174);
nand U6070 (N_6070,N_115,N_2076);
or U6071 (N_6071,N_3460,N_4786);
and U6072 (N_6072,N_1149,N_1632);
or U6073 (N_6073,N_3228,N_2605);
nor U6074 (N_6074,N_1007,N_952);
nand U6075 (N_6075,N_3091,N_401);
nand U6076 (N_6076,N_4190,N_2910);
nor U6077 (N_6077,N_4708,N_3521);
nand U6078 (N_6078,N_736,N_3258);
nand U6079 (N_6079,N_521,N_3371);
nor U6080 (N_6080,N_2022,N_4215);
nor U6081 (N_6081,N_2091,N_4179);
or U6082 (N_6082,N_3795,N_2617);
nor U6083 (N_6083,N_984,N_4677);
and U6084 (N_6084,N_1928,N_4811);
or U6085 (N_6085,N_3274,N_1832);
nand U6086 (N_6086,N_3793,N_3425);
or U6087 (N_6087,N_3740,N_2115);
nand U6088 (N_6088,N_757,N_1268);
or U6089 (N_6089,N_38,N_3343);
nor U6090 (N_6090,N_2033,N_1501);
and U6091 (N_6091,N_67,N_1686);
and U6092 (N_6092,N_4746,N_1836);
and U6093 (N_6093,N_1507,N_3837);
xnor U6094 (N_6094,N_2387,N_3336);
and U6095 (N_6095,N_3109,N_106);
and U6096 (N_6096,N_308,N_1740);
nand U6097 (N_6097,N_4728,N_288);
xor U6098 (N_6098,N_2278,N_3426);
and U6099 (N_6099,N_2843,N_1167);
nor U6100 (N_6100,N_3455,N_1954);
nand U6101 (N_6101,N_3964,N_2214);
nand U6102 (N_6102,N_2993,N_1062);
nand U6103 (N_6103,N_213,N_125);
xnor U6104 (N_6104,N_1574,N_43);
nor U6105 (N_6105,N_2247,N_2340);
nor U6106 (N_6106,N_4581,N_4185);
or U6107 (N_6107,N_3565,N_1515);
and U6108 (N_6108,N_4854,N_4863);
nand U6109 (N_6109,N_1466,N_3924);
and U6110 (N_6110,N_2641,N_1890);
xor U6111 (N_6111,N_2581,N_4335);
xor U6112 (N_6112,N_3650,N_4458);
nand U6113 (N_6113,N_1315,N_4426);
xnor U6114 (N_6114,N_3083,N_1488);
or U6115 (N_6115,N_2269,N_3213);
nand U6116 (N_6116,N_2270,N_1720);
nand U6117 (N_6117,N_1678,N_3084);
xor U6118 (N_6118,N_1048,N_3172);
or U6119 (N_6119,N_868,N_4615);
nand U6120 (N_6120,N_2457,N_4315);
and U6121 (N_6121,N_2156,N_1159);
nand U6122 (N_6122,N_3775,N_4475);
nor U6123 (N_6123,N_3498,N_2888);
and U6124 (N_6124,N_3218,N_2469);
xnor U6125 (N_6125,N_4606,N_4451);
nor U6126 (N_6126,N_711,N_3181);
and U6127 (N_6127,N_2308,N_618);
and U6128 (N_6128,N_2234,N_1961);
and U6129 (N_6129,N_1989,N_1071);
xor U6130 (N_6130,N_1184,N_953);
and U6131 (N_6131,N_1839,N_1170);
or U6132 (N_6132,N_2157,N_4246);
and U6133 (N_6133,N_4732,N_2755);
xnor U6134 (N_6134,N_3746,N_65);
and U6135 (N_6135,N_513,N_2095);
nor U6136 (N_6136,N_4978,N_2624);
nor U6137 (N_6137,N_1852,N_2796);
nand U6138 (N_6138,N_1981,N_803);
and U6139 (N_6139,N_1281,N_2096);
or U6140 (N_6140,N_1494,N_1318);
or U6141 (N_6141,N_576,N_4656);
or U6142 (N_6142,N_4264,N_2621);
xor U6143 (N_6143,N_355,N_4203);
nor U6144 (N_6144,N_571,N_2705);
xnor U6145 (N_6145,N_126,N_958);
or U6146 (N_6146,N_1172,N_4342);
nor U6147 (N_6147,N_3036,N_2552);
and U6148 (N_6148,N_4947,N_4207);
xor U6149 (N_6149,N_2813,N_2987);
and U6150 (N_6150,N_1918,N_2160);
nand U6151 (N_6151,N_1911,N_1272);
nor U6152 (N_6152,N_4088,N_3225);
or U6153 (N_6153,N_1260,N_2769);
and U6154 (N_6154,N_4079,N_2730);
or U6155 (N_6155,N_3723,N_4658);
or U6156 (N_6156,N_1618,N_3241);
nand U6157 (N_6157,N_653,N_667);
nor U6158 (N_6158,N_72,N_3474);
or U6159 (N_6159,N_2237,N_3359);
nand U6160 (N_6160,N_2005,N_462);
nand U6161 (N_6161,N_3339,N_3744);
and U6162 (N_6162,N_467,N_2841);
nand U6163 (N_6163,N_1304,N_254);
nand U6164 (N_6164,N_2530,N_626);
nand U6165 (N_6165,N_927,N_4952);
and U6166 (N_6166,N_3485,N_2519);
nand U6167 (N_6167,N_4220,N_157);
or U6168 (N_6168,N_1994,N_1367);
nor U6169 (N_6169,N_4990,N_727);
xor U6170 (N_6170,N_3479,N_1213);
nand U6171 (N_6171,N_3946,N_3140);
or U6172 (N_6172,N_245,N_4022);
nand U6173 (N_6173,N_2019,N_4457);
xnor U6174 (N_6174,N_665,N_77);
or U6175 (N_6175,N_883,N_3515);
and U6176 (N_6176,N_1604,N_3360);
and U6177 (N_6177,N_1483,N_955);
nand U6178 (N_6178,N_529,N_1259);
nand U6179 (N_6179,N_750,N_2876);
and U6180 (N_6180,N_2950,N_1021);
xnor U6181 (N_6181,N_2069,N_1969);
nand U6182 (N_6182,N_4809,N_629);
nand U6183 (N_6183,N_3101,N_4989);
nor U6184 (N_6184,N_3454,N_1381);
and U6185 (N_6185,N_278,N_1781);
nand U6186 (N_6186,N_1251,N_3059);
and U6187 (N_6187,N_2192,N_2830);
nor U6188 (N_6188,N_815,N_3338);
and U6189 (N_6189,N_1556,N_4420);
nand U6190 (N_6190,N_1333,N_1337);
and U6191 (N_6191,N_2334,N_4280);
xnor U6192 (N_6192,N_2542,N_1503);
and U6193 (N_6193,N_4785,N_959);
nand U6194 (N_6194,N_1666,N_4361);
nand U6195 (N_6195,N_1140,N_3170);
nand U6196 (N_6196,N_1878,N_4326);
and U6197 (N_6197,N_1638,N_2197);
nand U6198 (N_6198,N_294,N_4772);
nor U6199 (N_6199,N_3833,N_1958);
nor U6200 (N_6200,N_2874,N_163);
nor U6201 (N_6201,N_3609,N_200);
or U6202 (N_6202,N_4283,N_1275);
and U6203 (N_6203,N_1802,N_838);
nor U6204 (N_6204,N_4763,N_2068);
nand U6205 (N_6205,N_2614,N_3799);
and U6206 (N_6206,N_321,N_1077);
and U6207 (N_6207,N_3111,N_2304);
nand U6208 (N_6208,N_4001,N_2305);
and U6209 (N_6209,N_2264,N_1516);
nor U6210 (N_6210,N_4519,N_1391);
nand U6211 (N_6211,N_4111,N_1843);
nand U6212 (N_6212,N_621,N_1329);
and U6213 (N_6213,N_3500,N_789);
nand U6214 (N_6214,N_3279,N_3032);
or U6215 (N_6215,N_1433,N_2504);
nand U6216 (N_6216,N_2564,N_1458);
and U6217 (N_6217,N_674,N_4135);
nand U6218 (N_6218,N_2822,N_4840);
nor U6219 (N_6219,N_2438,N_3898);
and U6220 (N_6220,N_450,N_3435);
nor U6221 (N_6221,N_2529,N_361);
and U6222 (N_6222,N_4700,N_189);
nand U6223 (N_6223,N_2496,N_2966);
and U6224 (N_6224,N_1269,N_4843);
nor U6225 (N_6225,N_4216,N_2051);
nor U6226 (N_6226,N_4713,N_312);
nor U6227 (N_6227,N_455,N_56);
and U6228 (N_6228,N_323,N_3692);
or U6229 (N_6229,N_961,N_3097);
or U6230 (N_6230,N_4973,N_4671);
or U6231 (N_6231,N_2518,N_4468);
and U6232 (N_6232,N_715,N_2825);
nor U6233 (N_6233,N_862,N_540);
nand U6234 (N_6234,N_2199,N_3015);
nand U6235 (N_6235,N_2566,N_1164);
and U6236 (N_6236,N_149,N_3593);
nand U6237 (N_6237,N_3913,N_2838);
and U6238 (N_6238,N_1160,N_4894);
nor U6239 (N_6239,N_2819,N_305);
or U6240 (N_6240,N_1418,N_159);
or U6241 (N_6241,N_1778,N_4168);
or U6242 (N_6242,N_4430,N_1384);
nand U6243 (N_6243,N_639,N_2946);
or U6244 (N_6244,N_3261,N_2642);
nand U6245 (N_6245,N_2263,N_4093);
or U6246 (N_6246,N_784,N_1774);
nand U6247 (N_6247,N_1370,N_111);
and U6248 (N_6248,N_2916,N_4970);
nand U6249 (N_6249,N_14,N_1985);
nor U6250 (N_6250,N_4291,N_4083);
nand U6251 (N_6251,N_1733,N_835);
nor U6252 (N_6252,N_3785,N_3495);
or U6253 (N_6253,N_1587,N_3773);
nor U6254 (N_6254,N_2690,N_3444);
nor U6255 (N_6255,N_196,N_1947);
nand U6256 (N_6256,N_2090,N_3355);
or U6257 (N_6257,N_1279,N_2992);
nor U6258 (N_6258,N_2551,N_1);
nand U6259 (N_6259,N_2783,N_2840);
nand U6260 (N_6260,N_582,N_2103);
or U6261 (N_6261,N_2975,N_1180);
xnor U6262 (N_6262,N_4314,N_4366);
nand U6263 (N_6263,N_494,N_454);
nor U6264 (N_6264,N_741,N_3453);
nor U6265 (N_6265,N_4331,N_1711);
nand U6266 (N_6266,N_4789,N_1096);
and U6267 (N_6267,N_3314,N_1784);
nor U6268 (N_6268,N_2478,N_3284);
nand U6269 (N_6269,N_3017,N_4132);
or U6270 (N_6270,N_285,N_603);
and U6271 (N_6271,N_4199,N_4572);
and U6272 (N_6272,N_2126,N_4453);
or U6273 (N_6273,N_3571,N_4225);
nor U6274 (N_6274,N_1303,N_2635);
xnor U6275 (N_6275,N_384,N_1234);
nand U6276 (N_6276,N_617,N_2753);
nor U6277 (N_6277,N_4913,N_2070);
or U6278 (N_6278,N_3380,N_895);
nand U6279 (N_6279,N_3299,N_2600);
and U6280 (N_6280,N_4976,N_3390);
or U6281 (N_6281,N_4734,N_3988);
nor U6282 (N_6282,N_1083,N_1580);
or U6283 (N_6283,N_3658,N_3510);
nand U6284 (N_6284,N_3484,N_204);
xnor U6285 (N_6285,N_1388,N_2758);
or U6286 (N_6286,N_4095,N_740);
and U6287 (N_6287,N_474,N_4717);
nor U6288 (N_6288,N_2145,N_184);
or U6289 (N_6289,N_4431,N_1262);
nor U6290 (N_6290,N_348,N_2687);
xor U6291 (N_6291,N_3070,N_2623);
xor U6292 (N_6292,N_387,N_42);
nor U6293 (N_6293,N_230,N_1695);
and U6294 (N_6294,N_4403,N_4412);
xnor U6295 (N_6295,N_3502,N_404);
nand U6296 (N_6296,N_1768,N_558);
nor U6297 (N_6297,N_648,N_1812);
or U6298 (N_6298,N_4720,N_3657);
xnor U6299 (N_6299,N_3009,N_4346);
or U6300 (N_6300,N_1250,N_257);
and U6301 (N_6301,N_437,N_1098);
nor U6302 (N_6302,N_2224,N_751);
xor U6303 (N_6303,N_1101,N_956);
nand U6304 (N_6304,N_3618,N_3996);
and U6305 (N_6305,N_3854,N_1540);
nor U6306 (N_6306,N_2481,N_79);
nand U6307 (N_6307,N_3884,N_3158);
nand U6308 (N_6308,N_2277,N_4593);
nor U6309 (N_6309,N_1709,N_3729);
nor U6310 (N_6310,N_1800,N_4004);
nand U6311 (N_6311,N_4239,N_4040);
nor U6312 (N_6312,N_1484,N_2555);
nand U6313 (N_6313,N_112,N_3765);
or U6314 (N_6314,N_4667,N_131);
and U6315 (N_6315,N_3364,N_4859);
nand U6316 (N_6316,N_3437,N_3524);
and U6317 (N_6317,N_3838,N_3467);
nand U6318 (N_6318,N_2483,N_3653);
nor U6319 (N_6319,N_2436,N_2119);
xor U6320 (N_6320,N_2183,N_310);
nand U6321 (N_6321,N_898,N_3944);
nand U6322 (N_6322,N_3303,N_1773);
nor U6323 (N_6323,N_1806,N_4844);
nand U6324 (N_6324,N_3668,N_3332);
and U6325 (N_6325,N_2173,N_4928);
nand U6326 (N_6326,N_4106,N_4322);
or U6327 (N_6327,N_2658,N_1907);
or U6328 (N_6328,N_4899,N_3429);
nor U6329 (N_6329,N_2001,N_2289);
nand U6330 (N_6330,N_2151,N_2673);
nand U6331 (N_6331,N_3035,N_4221);
nor U6332 (N_6332,N_2017,N_88);
and U6333 (N_6333,N_3823,N_1244);
nor U6334 (N_6334,N_3983,N_1425);
nand U6335 (N_6335,N_4213,N_3270);
nand U6336 (N_6336,N_431,N_1320);
nand U6337 (N_6337,N_1153,N_2559);
and U6338 (N_6338,N_1820,N_2409);
nand U6339 (N_6339,N_3969,N_851);
nand U6340 (N_6340,N_1289,N_4766);
nand U6341 (N_6341,N_2267,N_3499);
nand U6342 (N_6342,N_1660,N_2941);
or U6343 (N_6343,N_4633,N_3724);
nand U6344 (N_6344,N_4655,N_4103);
nor U6345 (N_6345,N_698,N_216);
and U6346 (N_6346,N_3757,N_3870);
xnor U6347 (N_6347,N_4358,N_397);
or U6348 (N_6348,N_2656,N_4323);
and U6349 (N_6349,N_2238,N_1209);
nand U6350 (N_6350,N_4562,N_1882);
nand U6351 (N_6351,N_2568,N_211);
nand U6352 (N_6352,N_2934,N_1902);
xor U6353 (N_6353,N_957,N_4208);
nand U6354 (N_6354,N_3731,N_1352);
nand U6355 (N_6355,N_3962,N_3623);
nor U6356 (N_6356,N_303,N_3570);
and U6357 (N_6357,N_3190,N_3923);
nand U6358 (N_6358,N_1798,N_2461);
nand U6359 (N_6359,N_2037,N_1203);
xnor U6360 (N_6360,N_2482,N_498);
xor U6361 (N_6361,N_2251,N_2390);
xor U6362 (N_6362,N_964,N_4085);
or U6363 (N_6363,N_2365,N_3552);
nand U6364 (N_6364,N_50,N_1776);
xnor U6365 (N_6365,N_4818,N_654);
or U6366 (N_6366,N_1794,N_1202);
and U6367 (N_6367,N_3245,N_2688);
nand U6368 (N_6368,N_4715,N_1615);
nand U6369 (N_6369,N_2306,N_4234);
and U6370 (N_6370,N_4938,N_3162);
nand U6371 (N_6371,N_335,N_723);
nor U6372 (N_6372,N_3861,N_4736);
nor U6373 (N_6373,N_2010,N_3157);
or U6374 (N_6374,N_4919,N_2358);
or U6375 (N_6375,N_854,N_1113);
nor U6376 (N_6376,N_1220,N_4248);
xnor U6377 (N_6377,N_4159,N_4261);
xnor U6378 (N_6378,N_1502,N_2248);
or U6379 (N_6379,N_533,N_1633);
nor U6380 (N_6380,N_4460,N_1971);
nor U6381 (N_6381,N_2567,N_3466);
and U6382 (N_6382,N_4949,N_2169);
and U6383 (N_6383,N_4752,N_1990);
nand U6384 (N_6384,N_2405,N_1177);
nor U6385 (N_6385,N_4986,N_3211);
nor U6386 (N_6386,N_4348,N_913);
nor U6387 (N_6387,N_2430,N_3796);
xor U6388 (N_6388,N_2219,N_2347);
or U6389 (N_6389,N_1452,N_4063);
or U6390 (N_6390,N_3522,N_4868);
nand U6391 (N_6391,N_1157,N_4016);
or U6392 (N_6392,N_2297,N_2773);
and U6393 (N_6393,N_144,N_2378);
nor U6394 (N_6394,N_4600,N_2086);
nand U6395 (N_6395,N_4328,N_256);
and U6396 (N_6396,N_1999,N_3422);
or U6397 (N_6397,N_2654,N_989);
or U6398 (N_6398,N_1135,N_2829);
nand U6399 (N_6399,N_4414,N_1317);
or U6400 (N_6400,N_538,N_416);
or U6401 (N_6401,N_1566,N_4599);
nor U6402 (N_6402,N_4584,N_1896);
and U6403 (N_6403,N_3877,N_3841);
nor U6404 (N_6404,N_2459,N_4665);
or U6405 (N_6405,N_3137,N_1792);
nand U6406 (N_6406,N_2171,N_4382);
nor U6407 (N_6407,N_1554,N_2752);
nor U6408 (N_6408,N_1681,N_3501);
and U6409 (N_6409,N_2887,N_2450);
or U6410 (N_6410,N_1460,N_443);
and U6411 (N_6411,N_4268,N_4166);
nor U6412 (N_6412,N_4450,N_4830);
and U6413 (N_6413,N_3858,N_4694);
or U6414 (N_6414,N_4104,N_2944);
or U6415 (N_6415,N_4110,N_2168);
nor U6416 (N_6416,N_929,N_1827);
and U6417 (N_6417,N_2757,N_1937);
nor U6418 (N_6418,N_369,N_1094);
and U6419 (N_6419,N_103,N_4476);
nand U6420 (N_6420,N_4224,N_680);
nand U6421 (N_6421,N_710,N_3691);
nand U6422 (N_6422,N_2110,N_1570);
or U6423 (N_6423,N_1799,N_4695);
and U6424 (N_6424,N_1243,N_2492);
or U6425 (N_6425,N_768,N_3755);
or U6426 (N_6426,N_171,N_4714);
nand U6427 (N_6427,N_2889,N_3310);
nor U6428 (N_6428,N_1713,N_1227);
nand U6429 (N_6429,N_109,N_22);
nor U6430 (N_6430,N_2254,N_3812);
nand U6431 (N_6431,N_4045,N_1142);
or U6432 (N_6432,N_1206,N_3914);
xnor U6433 (N_6433,N_1498,N_2487);
nor U6434 (N_6434,N_2194,N_4359);
nor U6435 (N_6435,N_2133,N_2185);
nor U6436 (N_6436,N_1696,N_2479);
or U6437 (N_6437,N_2161,N_104);
nand U6438 (N_6438,N_1200,N_490);
and U6439 (N_6439,N_2632,N_4013);
nand U6440 (N_6440,N_57,N_4968);
or U6441 (N_6441,N_3504,N_3473);
and U6442 (N_6442,N_3016,N_2777);
nor U6443 (N_6443,N_1003,N_4154);
and U6444 (N_6444,N_4025,N_4057);
xor U6445 (N_6445,N_2712,N_4391);
nor U6446 (N_6446,N_3102,N_1297);
and U6447 (N_6447,N_905,N_4690);
and U6448 (N_6448,N_1826,N_1465);
or U6449 (N_6449,N_3830,N_2781);
nor U6450 (N_6450,N_4821,N_820);
nand U6451 (N_6451,N_3136,N_3384);
nor U6452 (N_6452,N_722,N_107);
and U6453 (N_6453,N_3193,N_3820);
nand U6454 (N_6454,N_2155,N_3381);
and U6455 (N_6455,N_2261,N_3006);
or U6456 (N_6456,N_2790,N_2144);
nand U6457 (N_6457,N_4308,N_2537);
nand U6458 (N_6458,N_99,N_3622);
and U6459 (N_6459,N_916,N_2275);
and U6460 (N_6460,N_4197,N_3554);
nand U6461 (N_6461,N_3824,N_3781);
or U6462 (N_6462,N_102,N_1952);
or U6463 (N_6463,N_2312,N_2325);
xor U6464 (N_6464,N_337,N_2373);
and U6465 (N_6465,N_4757,N_349);
or U6466 (N_6466,N_114,N_4556);
nand U6467 (N_6467,N_2284,N_1070);
nand U6468 (N_6468,N_763,N_4645);
and U6469 (N_6469,N_3227,N_134);
nand U6470 (N_6470,N_441,N_2681);
nor U6471 (N_6471,N_1086,N_2510);
or U6472 (N_6472,N_4195,N_595);
nand U6473 (N_6473,N_1640,N_101);
nand U6474 (N_6474,N_3987,N_4815);
or U6475 (N_6475,N_4229,N_4161);
and U6476 (N_6476,N_3178,N_1436);
nand U6477 (N_6477,N_1861,N_3321);
nor U6478 (N_6478,N_4880,N_4026);
or U6479 (N_6479,N_2609,N_4436);
xor U6480 (N_6480,N_1897,N_1385);
and U6481 (N_6481,N_4838,N_1165);
nand U6482 (N_6482,N_1970,N_4418);
or U6483 (N_6483,N_3065,N_33);
nor U6484 (N_6484,N_1903,N_3442);
or U6485 (N_6485,N_1608,N_3507);
nand U6486 (N_6486,N_1899,N_3071);
or U6487 (N_6487,N_4939,N_4068);
nand U6488 (N_6488,N_258,N_1916);
nor U6489 (N_6489,N_3076,N_4466);
xor U6490 (N_6490,N_44,N_3457);
xnor U6491 (N_6491,N_2722,N_504);
nand U6492 (N_6492,N_4669,N_2884);
or U6493 (N_6493,N_3896,N_842);
nor U6494 (N_6494,N_379,N_1404);
and U6495 (N_6495,N_3312,N_1035);
nand U6496 (N_6496,N_1787,N_3288);
nand U6497 (N_6497,N_2407,N_2985);
nor U6498 (N_6498,N_3000,N_2502);
or U6499 (N_6499,N_2402,N_3316);
nand U6500 (N_6500,N_2170,N_1573);
or U6501 (N_6501,N_3687,N_663);
nor U6502 (N_6502,N_3204,N_1505);
nor U6503 (N_6503,N_2780,N_113);
nor U6504 (N_6504,N_3092,N_1637);
nand U6505 (N_6505,N_3619,N_886);
xor U6506 (N_6506,N_3694,N_1700);
nor U6507 (N_6507,N_2380,N_1449);
nand U6508 (N_6508,N_4421,N_2178);
nor U6509 (N_6509,N_4653,N_365);
or U6510 (N_6510,N_1360,N_4566);
or U6511 (N_6511,N_3925,N_1093);
and U6512 (N_6512,N_4257,N_1386);
nor U6513 (N_6513,N_3899,N_863);
and U6514 (N_6514,N_4117,N_4194);
and U6515 (N_6515,N_3464,N_575);
nand U6516 (N_6516,N_4639,N_408);
nand U6517 (N_6517,N_1504,N_4392);
or U6518 (N_6518,N_2506,N_3348);
nand U6519 (N_6519,N_2890,N_4647);
or U6520 (N_6520,N_4903,N_4065);
or U6521 (N_6521,N_4791,N_3294);
nor U6522 (N_6522,N_1887,N_2697);
and U6523 (N_6523,N_2556,N_139);
and U6524 (N_6524,N_396,N_449);
and U6525 (N_6525,N_2534,N_1130);
nor U6526 (N_6526,N_509,N_4501);
and U6527 (N_6527,N_1628,N_1662);
nand U6528 (N_6528,N_413,N_3625);
and U6529 (N_6529,N_1447,N_3334);
nand U6530 (N_6530,N_4906,N_2789);
and U6531 (N_6531,N_3163,N_251);
and U6532 (N_6532,N_4660,N_2217);
or U6533 (N_6533,N_697,N_1821);
or U6534 (N_6534,N_2059,N_1823);
or U6535 (N_6535,N_3439,N_3935);
xnor U6536 (N_6536,N_2728,N_24);
nor U6537 (N_6537,N_292,N_2932);
xnor U6538 (N_6538,N_1708,N_1265);
and U6539 (N_6539,N_1334,N_1407);
nand U6540 (N_6540,N_1513,N_3087);
and U6541 (N_6541,N_3064,N_1322);
nand U6542 (N_6542,N_4370,N_49);
nand U6543 (N_6543,N_2352,N_2622);
nand U6544 (N_6544,N_4196,N_2124);
or U6545 (N_6545,N_2184,N_3722);
and U6546 (N_6546,N_4175,N_2691);
and U6547 (N_6547,N_20,N_1112);
xnor U6548 (N_6548,N_4852,N_1734);
and U6549 (N_6549,N_4902,N_4552);
nor U6550 (N_6550,N_2061,N_4044);
nand U6551 (N_6551,N_1610,N_4276);
nand U6552 (N_6552,N_1754,N_1956);
or U6553 (N_6553,N_4138,N_1972);
and U6554 (N_6554,N_1731,N_594);
and U6555 (N_6555,N_2175,N_3419);
xor U6556 (N_6556,N_46,N_1446);
and U6557 (N_6557,N_3497,N_1241);
nor U6558 (N_6558,N_4877,N_1030);
nand U6559 (N_6559,N_2879,N_793);
nand U6560 (N_6560,N_563,N_194);
or U6561 (N_6561,N_2643,N_2891);
nor U6562 (N_6562,N_4050,N_3611);
nand U6563 (N_6563,N_3728,N_2080);
or U6564 (N_6564,N_1997,N_2432);
nor U6565 (N_6565,N_1032,N_3361);
nand U6566 (N_6566,N_4893,N_1187);
nand U6567 (N_6567,N_3215,N_4914);
or U6568 (N_6568,N_720,N_2591);
xor U6569 (N_6569,N_3277,N_1045);
and U6570 (N_6570,N_2570,N_1186);
and U6571 (N_6571,N_300,N_1328);
or U6572 (N_6572,N_3943,N_2924);
xor U6573 (N_6573,N_906,N_1085);
and U6574 (N_6574,N_4505,N_721);
nand U6575 (N_6575,N_2644,N_3179);
and U6576 (N_6576,N_3418,N_1399);
nand U6577 (N_6577,N_2661,N_3984);
nor U6578 (N_6578,N_3010,N_4330);
and U6579 (N_6579,N_237,N_1305);
nor U6580 (N_6580,N_4210,N_175);
and U6581 (N_6581,N_1010,N_1380);
xor U6582 (N_6582,N_3745,N_3295);
and U6583 (N_6583,N_3423,N_3674);
or U6584 (N_6584,N_4511,N_3589);
and U6585 (N_6585,N_4607,N_2018);
nand U6586 (N_6586,N_3289,N_3736);
nor U6587 (N_6587,N_4094,N_1025);
nand U6588 (N_6588,N_4585,N_1757);
and U6589 (N_6589,N_1224,N_2533);
or U6590 (N_6590,N_1467,N_2883);
and U6591 (N_6591,N_3230,N_2000);
or U6592 (N_6592,N_360,N_2245);
nand U6593 (N_6593,N_877,N_3523);
nand U6594 (N_6594,N_4429,N_1292);
or U6595 (N_6595,N_4140,N_4217);
nand U6596 (N_6596,N_4602,N_941);
xor U6597 (N_6597,N_1865,N_1204);
xnor U6598 (N_6598,N_985,N_1406);
nand U6599 (N_6599,N_3999,N_2939);
nand U6600 (N_6600,N_743,N_4754);
or U6601 (N_6601,N_3710,N_3383);
nand U6602 (N_6602,N_3297,N_3030);
nand U6603 (N_6603,N_2315,N_3680);
nand U6604 (N_6604,N_3404,N_342);
nand U6605 (N_6605,N_2137,N_2242);
nor U6606 (N_6606,N_606,N_1316);
nor U6607 (N_6607,N_739,N_3664);
nor U6608 (N_6608,N_3477,N_2418);
nor U6609 (N_6609,N_2544,N_367);
nor U6610 (N_6610,N_4082,N_3353);
nand U6611 (N_6611,N_2223,N_1629);
or U6612 (N_6612,N_1356,N_177);
or U6613 (N_6613,N_3836,N_1617);
or U6614 (N_6614,N_4380,N_2791);
or U6615 (N_6615,N_2225,N_4981);
or U6616 (N_6616,N_3440,N_1926);
and U6617 (N_6617,N_4753,N_2598);
and U6618 (N_6618,N_3937,N_1340);
xnor U6619 (N_6619,N_3792,N_2222);
nand U6620 (N_6620,N_1851,N_4456);
or U6621 (N_6621,N_2332,N_3082);
nor U6622 (N_6622,N_2857,N_4573);
and U6623 (N_6623,N_127,N_1625);
nor U6624 (N_6624,N_3747,N_2802);
and U6625 (N_6625,N_4479,N_4561);
or U6626 (N_6626,N_4648,N_2403);
nand U6627 (N_6627,N_4402,N_2111);
nand U6628 (N_6628,N_673,N_678);
nand U6629 (N_6629,N_2239,N_686);
xnor U6630 (N_6630,N_1080,N_607);
and U6631 (N_6631,N_3090,N_222);
nor U6632 (N_6632,N_4084,N_3320);
nor U6633 (N_6633,N_327,N_333);
nor U6634 (N_6634,N_3250,N_857);
and U6635 (N_6635,N_1898,N_74);
nand U6636 (N_6636,N_2052,N_3780);
nor U6637 (N_6637,N_2922,N_2774);
and U6638 (N_6638,N_272,N_1657);
nand U6639 (N_6639,N_982,N_4532);
and U6640 (N_6640,N_4012,N_1109);
or U6641 (N_6641,N_4408,N_2153);
xor U6642 (N_6642,N_482,N_1726);
and U6643 (N_6643,N_1676,N_4385);
nor U6644 (N_6644,N_1830,N_1043);
nand U6645 (N_6645,N_1118,N_507);
nand U6646 (N_6646,N_2419,N_4035);
nand U6647 (N_6647,N_2434,N_1743);
nor U6648 (N_6648,N_978,N_2394);
nor U6649 (N_6649,N_2444,N_919);
or U6650 (N_6650,N_1412,N_314);
nand U6651 (N_6651,N_1569,N_2880);
and U6652 (N_6652,N_26,N_4819);
nand U6653 (N_6653,N_120,N_110);
xnor U6654 (N_6654,N_4381,N_4292);
xnor U6655 (N_6655,N_980,N_3117);
nand U6656 (N_6656,N_2179,N_4332);
nor U6657 (N_6657,N_1679,N_16);
and U6658 (N_6658,N_559,N_232);
or U6659 (N_6659,N_564,N_4550);
xor U6660 (N_6660,N_2525,N_752);
or U6661 (N_6661,N_3926,N_4014);
or U6662 (N_6662,N_4051,N_2742);
and U6663 (N_6663,N_2314,N_4047);
and U6664 (N_6664,N_198,N_3062);
nor U6665 (N_6665,N_3828,N_3156);
or U6666 (N_6666,N_2959,N_4162);
nand U6667 (N_6667,N_2406,N_2779);
nor U6668 (N_6668,N_615,N_133);
nand U6669 (N_6669,N_4250,N_3243);
nor U6670 (N_6670,N_3350,N_3154);
nor U6671 (N_6671,N_1144,N_4069);
nand U6672 (N_6672,N_3039,N_1107);
xor U6673 (N_6673,N_2074,N_428);
and U6674 (N_6674,N_790,N_4748);
or U6675 (N_6675,N_2990,N_2425);
or U6676 (N_6676,N_3790,N_301);
and U6677 (N_6677,N_4107,N_4282);
and U6678 (N_6678,N_1276,N_811);
nor U6679 (N_6679,N_3897,N_458);
xnor U6680 (N_6680,N_3047,N_3990);
nand U6681 (N_6681,N_3183,N_4187);
or U6682 (N_6682,N_1005,N_1496);
xnor U6683 (N_6683,N_4237,N_1486);
and U6684 (N_6684,N_3287,N_236);
nor U6685 (N_6685,N_971,N_1868);
nand U6686 (N_6686,N_1753,N_2585);
and U6687 (N_6687,N_973,N_150);
nand U6688 (N_6688,N_4590,N_2041);
xnor U6689 (N_6689,N_4075,N_3695);
nor U6690 (N_6690,N_2921,N_2446);
xnor U6691 (N_6691,N_4474,N_2106);
nor U6692 (N_6692,N_2512,N_583);
xor U6693 (N_6693,N_4661,N_3621);
nor U6694 (N_6694,N_4387,N_1951);
nor U6695 (N_6695,N_2186,N_2125);
nand U6696 (N_6696,N_284,N_4329);
nand U6697 (N_6697,N_383,N_4984);
or U6698 (N_6698,N_1027,N_669);
nor U6699 (N_6699,N_152,N_4188);
or U6700 (N_6700,N_2121,N_4109);
and U6701 (N_6701,N_3626,N_3829);
nor U6702 (N_6702,N_2198,N_4545);
and U6703 (N_6703,N_2703,N_541);
nor U6704 (N_6704,N_1771,N_1417);
xnor U6705 (N_6705,N_3267,N_3096);
or U6706 (N_6706,N_2201,N_2296);
nand U6707 (N_6707,N_3798,N_2915);
nor U6708 (N_6708,N_3056,N_3133);
xnor U6709 (N_6709,N_1930,N_2411);
or U6710 (N_6710,N_3910,N_252);
nand U6711 (N_6711,N_3487,N_1780);
nor U6712 (N_6712,N_1480,N_4574);
and U6713 (N_6713,N_4423,N_1041);
xor U6714 (N_6714,N_2582,N_2831);
nand U6715 (N_6715,N_3233,N_2856);
nor U6716 (N_6716,N_3591,N_4056);
and U6717 (N_6717,N_1673,N_3445);
or U6718 (N_6718,N_75,N_4449);
xor U6719 (N_6719,N_1649,N_707);
nor U6720 (N_6720,N_3800,N_3550);
nand U6721 (N_6721,N_3124,N_4454);
or U6722 (N_6722,N_2371,N_3089);
xor U6723 (N_6723,N_202,N_2667);
or U6724 (N_6724,N_3537,N_2523);
or U6725 (N_6725,N_1455,N_872);
and U6726 (N_6726,N_2030,N_3399);
or U6727 (N_6727,N_2477,N_4597);
and U6728 (N_6728,N_2123,N_2428);
nor U6729 (N_6729,N_3077,N_3456);
and U6730 (N_6730,N_3438,N_3614);
nor U6731 (N_6731,N_286,N_4801);
and U6732 (N_6732,N_2930,N_1838);
xor U6733 (N_6733,N_2763,N_3103);
or U6734 (N_6734,N_2116,N_2057);
and U6735 (N_6735,N_2228,N_1886);
and U6736 (N_6736,N_3095,N_4756);
nor U6737 (N_6737,N_4992,N_58);
and U6738 (N_6738,N_4371,N_3192);
or U6739 (N_6739,N_4389,N_1803);
nand U6740 (N_6740,N_2188,N_3696);
xor U6741 (N_6741,N_2023,N_3878);
and U6742 (N_6742,N_598,N_3791);
and U6743 (N_6743,N_787,N_2359);
nand U6744 (N_6744,N_4805,N_825);
nor U6745 (N_6745,N_2189,N_2547);
or U6746 (N_6746,N_3560,N_2369);
nand U6747 (N_6747,N_477,N_2816);
nor U6748 (N_6748,N_2466,N_975);
or U6749 (N_6749,N_3432,N_3405);
nand U6750 (N_6750,N_3954,N_3113);
nand U6751 (N_6751,N_2246,N_1641);
or U6752 (N_6752,N_2036,N_1033);
nor U6753 (N_6753,N_4741,N_1929);
nand U6754 (N_6754,N_4155,N_1014);
nand U6755 (N_6755,N_1379,N_259);
nor U6756 (N_6756,N_4726,N_73);
nor U6757 (N_6757,N_2345,N_3817);
and U6758 (N_6758,N_2647,N_3110);
or U6759 (N_6759,N_1039,N_947);
or U6760 (N_6760,N_549,N_3492);
or U6761 (N_6761,N_4878,N_4455);
or U6762 (N_6762,N_1675,N_1879);
or U6763 (N_6763,N_4983,N_1749);
nor U6764 (N_6764,N_4269,N_4853);
or U6765 (N_6765,N_3269,N_2553);
xor U6766 (N_6766,N_1692,N_2545);
and U6767 (N_6767,N_2662,N_866);
xnor U6768 (N_6768,N_1670,N_4445);
or U6769 (N_6769,N_556,N_2441);
nor U6770 (N_6770,N_4918,N_1722);
xor U6771 (N_6771,N_620,N_1601);
nor U6772 (N_6772,N_2166,N_1057);
nor U6773 (N_6773,N_1475,N_1909);
or U6774 (N_6774,N_4654,N_3874);
nand U6775 (N_6775,N_1816,N_4595);
or U6776 (N_6776,N_3730,N_1422);
and U6777 (N_6777,N_4945,N_447);
and U6778 (N_6778,N_1525,N_1534);
or U6779 (N_6779,N_2241,N_3628);
nor U6780 (N_6780,N_90,N_1211);
or U6781 (N_6781,N_140,N_4711);
nor U6782 (N_6782,N_4559,N_2129);
and U6783 (N_6783,N_4206,N_997);
nand U6784 (N_6784,N_1341,N_3290);
xnor U6785 (N_6785,N_2102,N_557);
or U6786 (N_6786,N_1729,N_3271);
nand U6787 (N_6787,N_1343,N_338);
nor U6788 (N_6788,N_1680,N_709);
nor U6789 (N_6789,N_4039,N_3577);
nand U6790 (N_6790,N_4664,N_1533);
nand U6791 (N_6791,N_3659,N_3431);
nor U6792 (N_6792,N_1453,N_3814);
nor U6793 (N_6793,N_3315,N_3777);
and U6794 (N_6794,N_923,N_590);
nand U6795 (N_6795,N_764,N_4309);
xnor U6796 (N_6796,N_2894,N_4369);
nand U6797 (N_6797,N_1408,N_1544);
nand U6798 (N_6798,N_4191,N_4301);
nand U6799 (N_6799,N_548,N_4287);
nand U6800 (N_6800,N_2148,N_2906);
nand U6801 (N_6801,N_4881,N_2163);
or U6802 (N_6802,N_129,N_3902);
nand U6803 (N_6803,N_64,N_891);
and U6804 (N_6804,N_1336,N_1746);
nand U6805 (N_6805,N_1701,N_4958);
nor U6806 (N_6806,N_4165,N_831);
or U6807 (N_6807,N_4407,N_1065);
or U6808 (N_6808,N_1061,N_967);
or U6809 (N_6809,N_4260,N_2085);
or U6810 (N_6810,N_4438,N_3840);
and U6811 (N_6811,N_2877,N_4540);
nor U6812 (N_6812,N_1129,N_3143);
nand U6813 (N_6813,N_2766,N_761);
and U6814 (N_6814,N_4617,N_4033);
nand U6815 (N_6815,N_570,N_788);
or U6816 (N_6816,N_4662,N_2437);
nor U6817 (N_6817,N_2117,N_3236);
and U6818 (N_6818,N_3768,N_4884);
nand U6819 (N_6819,N_4053,N_779);
or U6820 (N_6820,N_436,N_4064);
or U6821 (N_6821,N_922,N_2122);
and U6822 (N_6822,N_1996,N_1572);
or U6823 (N_6823,N_935,N_4832);
nor U6824 (N_6824,N_2235,N_2933);
nand U6825 (N_6825,N_4577,N_1273);
nand U6826 (N_6826,N_3753,N_3769);
and U6827 (N_6827,N_2146,N_71);
nand U6828 (N_6828,N_4966,N_1634);
and U6829 (N_6829,N_3347,N_845);
nor U6830 (N_6830,N_3406,N_2718);
and U6831 (N_6831,N_3112,N_1389);
or U6832 (N_6832,N_2653,N_864);
nor U6833 (N_6833,N_3313,N_4831);
and U6834 (N_6834,N_2135,N_293);
nand U6835 (N_6835,N_4247,N_1478);
xor U6836 (N_6836,N_4967,N_4826);
and U6837 (N_6837,N_192,N_1199);
and U6838 (N_6838,N_4178,N_2370);
nor U6839 (N_6839,N_1469,N_2851);
xnor U6840 (N_6840,N_749,N_585);
and U6841 (N_6841,N_1403,N_1246);
nor U6842 (N_6842,N_2546,N_1659);
or U6843 (N_6843,N_1857,N_4845);
and U6844 (N_6844,N_2120,N_4941);
xnor U6845 (N_6845,N_4098,N_1511);
nor U6846 (N_6846,N_2182,N_4886);
nor U6847 (N_6847,N_3069,N_4764);
and U6848 (N_6848,N_3259,N_4760);
nor U6849 (N_6849,N_865,N_4417);
nand U6850 (N_6850,N_1435,N_3981);
or U6851 (N_6851,N_3262,N_986);
and U6852 (N_6852,N_4940,N_4614);
and U6853 (N_6853,N_4866,N_744);
or U6854 (N_6854,N_708,N_381);
nor U6855 (N_6855,N_3100,N_76);
nand U6856 (N_6856,N_3689,N_3873);
and U6857 (N_6857,N_2294,N_4619);
and U6858 (N_6858,N_4512,N_63);
nand U6859 (N_6859,N_1321,N_2291);
nor U6860 (N_6860,N_4351,N_2349);
and U6861 (N_6861,N_19,N_3574);
nor U6862 (N_6862,N_212,N_2524);
nor U6863 (N_6863,N_1639,N_3226);
and U6864 (N_6864,N_3956,N_2313);
or U6865 (N_6865,N_791,N_2420);
nand U6866 (N_6866,N_2885,N_3304);
xnor U6867 (N_6867,N_1689,N_2215);
and U6868 (N_6868,N_493,N_304);
nor U6869 (N_6869,N_4933,N_2931);
nand U6870 (N_6870,N_1811,N_2575);
nor U6871 (N_6871,N_4258,N_224);
nand U6872 (N_6872,N_2836,N_2112);
xnor U6873 (N_6873,N_3472,N_616);
and U6874 (N_6874,N_4783,N_3043);
nor U6875 (N_6875,N_1645,N_4994);
or U6876 (N_6876,N_3229,N_4172);
nor U6877 (N_6877,N_609,N_1651);
nor U6878 (N_6878,N_3407,N_4284);
nand U6879 (N_6879,N_4588,N_3463);
xnor U6880 (N_6880,N_566,N_1368);
nor U6881 (N_6881,N_2134,N_1913);
and U6882 (N_6882,N_4344,N_268);
nor U6883 (N_6883,N_466,N_2801);
or U6884 (N_6884,N_1441,N_476);
nor U6885 (N_6885,N_2760,N_1648);
and U6886 (N_6886,N_2376,N_4006);
and U6887 (N_6887,N_219,N_2266);
nor U6888 (N_6888,N_719,N_4127);
or U6889 (N_6889,N_1819,N_2929);
xnor U6890 (N_6890,N_3894,N_153);
xor U6891 (N_6891,N_2710,N_4768);
and U6892 (N_6892,N_3715,N_2795);
or U6893 (N_6893,N_940,N_4946);
and U6894 (N_6894,N_762,N_3067);
and U6895 (N_6895,N_2003,N_4428);
xor U6896 (N_6896,N_766,N_4133);
and U6897 (N_6897,N_246,N_1888);
and U6898 (N_6898,N_3368,N_1871);
nor U6899 (N_6899,N_4522,N_4096);
xor U6900 (N_6900,N_3645,N_3754);
and U6901 (N_6901,N_2845,N_2858);
and U6902 (N_6902,N_3298,N_18);
and U6903 (N_6903,N_2860,N_2548);
nor U6904 (N_6904,N_4803,N_2050);
nor U6905 (N_6905,N_1066,N_1542);
or U6906 (N_6906,N_2484,N_377);
nor U6907 (N_6907,N_183,N_2541);
or U6908 (N_6908,N_3534,N_2443);
nor U6909 (N_6909,N_640,N_1818);
nand U6910 (N_6910,N_1355,N_4869);
and U6911 (N_6911,N_3248,N_4310);
xor U6912 (N_6912,N_2554,N_1173);
nand U6913 (N_6913,N_4842,N_3662);
and U6914 (N_6914,N_2788,N_2435);
or U6915 (N_6915,N_2651,N_972);
and U6916 (N_6916,N_4982,N_1474);
nand U6917 (N_6917,N_3917,N_1510);
and U6918 (N_6918,N_2154,N_1387);
or U6919 (N_6919,N_852,N_457);
xnor U6920 (N_6920,N_4935,N_2486);
nand U6921 (N_6921,N_1326,N_1883);
nor U6922 (N_6922,N_4802,N_3021);
and U6923 (N_6923,N_1448,N_4807);
and U6924 (N_6924,N_3794,N_1950);
nor U6925 (N_6925,N_2620,N_4776);
or U6926 (N_6926,N_427,N_3305);
and U6927 (N_6927,N_3221,N_2476);
nand U6928 (N_6928,N_4955,N_977);
nand U6929 (N_6929,N_3776,N_894);
xor U6930 (N_6930,N_2815,N_3138);
and U6931 (N_6931,N_3810,N_3649);
nor U6932 (N_6932,N_3782,N_2309);
or U6933 (N_6933,N_802,N_3256);
or U6934 (N_6934,N_203,N_2862);
nand U6935 (N_6935,N_1875,N_2132);
nor U6936 (N_6936,N_581,N_3356);
nor U6937 (N_6937,N_4181,N_1894);
and U6938 (N_6938,N_656,N_1396);
nor U6939 (N_6939,N_3011,N_1346);
xor U6940 (N_6940,N_1409,N_2139);
or U6941 (N_6941,N_1309,N_702);
nor U6942 (N_6942,N_843,N_1293);
nand U6943 (N_6943,N_3165,N_1089);
xnor U6944 (N_6944,N_1508,N_270);
nor U6945 (N_6945,N_3126,N_1285);
or U6946 (N_6946,N_4452,N_1519);
xor U6947 (N_6947,N_398,N_2576);
xnor U6948 (N_6948,N_3469,N_3282);
xor U6949 (N_6949,N_3205,N_1067);
nand U6950 (N_6950,N_2631,N_1238);
or U6951 (N_6951,N_2259,N_451);
nand U6952 (N_6952,N_4253,N_2700);
xnor U6953 (N_6953,N_2077,N_3842);
nor U6954 (N_6954,N_4487,N_550);
nor U6955 (N_6955,N_1146,N_514);
nor U6956 (N_6956,N_4813,N_2401);
or U6957 (N_6957,N_931,N_672);
and U6958 (N_6958,N_3525,N_1609);
or U6959 (N_6959,N_4477,N_3145);
or U6960 (N_6960,N_3116,N_772);
xnor U6961 (N_6961,N_4931,N_4176);
nor U6962 (N_6962,N_3281,N_717);
or U6963 (N_6963,N_3986,N_4448);
xor U6964 (N_6964,N_2771,N_4725);
nor U6965 (N_6965,N_4696,N_1217);
nor U6966 (N_6966,N_4411,N_2445);
and U6967 (N_6967,N_1993,N_1174);
and U6968 (N_6968,N_4796,N_1248);
xor U6969 (N_6969,N_1893,N_2232);
or U6970 (N_6970,N_3182,N_3881);
nand U6971 (N_6971,N_2448,N_730);
xor U6972 (N_6972,N_526,N_4304);
or U6973 (N_6973,N_81,N_821);
nand U6974 (N_6974,N_1468,N_1076);
nand U6975 (N_6975,N_792,N_1528);
nand U6976 (N_6976,N_1029,N_1760);
nor U6977 (N_6977,N_880,N_2909);
and U6978 (N_6978,N_2998,N_4011);
xor U6979 (N_6979,N_3328,N_1512);
xnor U6980 (N_6980,N_3928,N_2706);
nand U6981 (N_6981,N_1822,N_3575);
or U6982 (N_6982,N_2004,N_1940);
nor U6983 (N_6983,N_3743,N_579);
and U6984 (N_6984,N_1068,N_2867);
nand U6985 (N_6985,N_4847,N_3592);
and U6986 (N_6986,N_2463,N_4042);
nand U6987 (N_6987,N_4742,N_1004);
nand U6988 (N_6988,N_4774,N_1313);
nor U6989 (N_6989,N_2935,N_4481);
xor U6990 (N_6990,N_1702,N_932);
xor U6991 (N_6991,N_4640,N_4514);
and U6992 (N_6992,N_3717,N_759);
nor U6993 (N_6993,N_2489,N_395);
or U6994 (N_6994,N_1176,N_2852);
xor U6995 (N_6995,N_4313,N_1738);
and U6996 (N_6996,N_2608,N_4551);
xnor U6997 (N_6997,N_3246,N_1859);
and U6998 (N_6998,N_2660,N_1665);
nor U6999 (N_6999,N_363,N_2543);
or U7000 (N_7000,N_1047,N_1848);
and U7001 (N_7001,N_2937,N_934);
nand U7002 (N_7002,N_4762,N_2399);
nor U7003 (N_7003,N_4650,N_1723);
nand U7004 (N_7004,N_1075,N_1905);
nand U7005 (N_7005,N_1698,N_2342);
and U7006 (N_7006,N_4507,N_960);
and U7007 (N_7007,N_3922,N_1482);
nand U7008 (N_7008,N_243,N_1941);
nand U7009 (N_7009,N_2999,N_683);
or U7010 (N_7010,N_2610,N_2669);
xor U7011 (N_7011,N_2912,N_2172);
nand U7012 (N_7012,N_4130,N_3613);
nand U7013 (N_7013,N_4399,N_3888);
or U7014 (N_7014,N_2410,N_4890);
xor U7015 (N_7015,N_4862,N_2832);
and U7016 (N_7016,N_3624,N_3098);
or U7017 (N_7017,N_1405,N_4324);
nand U7018 (N_7018,N_4598,N_4052);
xnor U7019 (N_7019,N_1593,N_690);
and U7020 (N_7020,N_3978,N_3340);
nand U7021 (N_7021,N_4864,N_180);
nand U7022 (N_7022,N_3544,N_69);
nor U7023 (N_7023,N_4670,N_4023);
nand U7024 (N_7024,N_2947,N_4113);
and U7025 (N_7025,N_1104,N_329);
or U7026 (N_7026,N_1296,N_3106);
and U7027 (N_7027,N_2686,N_1154);
nand U7028 (N_7028,N_776,N_3843);
and U7029 (N_7029,N_3646,N_4126);
nand U7030 (N_7030,N_889,N_2413);
nor U7031 (N_7031,N_1233,N_1249);
and U7032 (N_7032,N_795,N_816);
xor U7033 (N_7033,N_4263,N_2009);
or U7034 (N_7034,N_3578,N_4697);
nor U7035 (N_7035,N_3173,N_3013);
and U7036 (N_7036,N_3187,N_1793);
and U7037 (N_7037,N_3478,N_3811);
and U7038 (N_7038,N_1872,N_3960);
nor U7039 (N_7039,N_2701,N_3706);
nand U7040 (N_7040,N_414,N_4705);
and U7041 (N_7041,N_4493,N_3526);
nor U7042 (N_7042,N_3558,N_1395);
and U7043 (N_7043,N_4442,N_1988);
nor U7044 (N_7044,N_849,N_602);
or U7045 (N_7045,N_4883,N_1188);
nand U7046 (N_7046,N_4808,N_4564);
nand U7047 (N_7047,N_1095,N_1664);
nor U7048 (N_7048,N_3629,N_2079);
nand U7049 (N_7049,N_2683,N_281);
and U7050 (N_7050,N_82,N_4189);
xor U7051 (N_7051,N_1626,N_3750);
or U7052 (N_7052,N_4971,N_610);
xor U7053 (N_7053,N_1652,N_2150);
nand U7054 (N_7054,N_1001,N_2431);
xor U7055 (N_7055,N_4672,N_518);
nor U7056 (N_7056,N_4288,N_4544);
or U7057 (N_7057,N_2563,N_946);
or U7058 (N_7058,N_2034,N_4378);
nand U7059 (N_7059,N_3882,N_1984);
and U7060 (N_7060,N_3634,N_1917);
or U7061 (N_7061,N_765,N_322);
or U7062 (N_7062,N_4659,N_3397);
nor U7063 (N_7063,N_4569,N_2574);
nand U7064 (N_7064,N_2853,N_4467);
nand U7065 (N_7065,N_1668,N_209);
nor U7066 (N_7066,N_241,N_2084);
or U7067 (N_7067,N_1054,N_4279);
and U7068 (N_7068,N_1974,N_3885);
or U7069 (N_7069,N_319,N_1042);
nand U7070 (N_7070,N_2244,N_1855);
nor U7071 (N_7071,N_1948,N_1583);
and U7072 (N_7072,N_604,N_1598);
and U7073 (N_7073,N_2088,N_3185);
nand U7074 (N_7074,N_283,N_572);
nand U7075 (N_7075,N_4341,N_3616);
nor U7076 (N_7076,N_1013,N_3563);
or U7077 (N_7077,N_273,N_100);
nand U7078 (N_7078,N_45,N_4582);
nand U7079 (N_7079,N_712,N_3867);
and U7080 (N_7080,N_3976,N_4961);
and U7081 (N_7081,N_1643,N_362);
nand U7082 (N_7082,N_4238,N_4823);
and U7083 (N_7083,N_2424,N_4610);
nor U7084 (N_7084,N_1119,N_1936);
or U7085 (N_7085,N_388,N_3186);
or U7086 (N_7086,N_249,N_2721);
or U7087 (N_7087,N_855,N_4810);
nor U7088 (N_7088,N_2318,N_853);
nor U7089 (N_7089,N_3050,N_645);
nand U7090 (N_7090,N_2204,N_3234);
or U7091 (N_7091,N_1492,N_4889);
nor U7092 (N_7092,N_593,N_1653);
xnor U7093 (N_7093,N_3027,N_3665);
or U7094 (N_7094,N_2362,N_1414);
nor U7095 (N_7095,N_4873,N_3042);
xnor U7096 (N_7096,N_3025,N_324);
nand U7097 (N_7097,N_2099,N_687);
nor U7098 (N_7098,N_882,N_4478);
and U7099 (N_7099,N_2695,N_118);
or U7100 (N_7100,N_1982,N_4557);
nor U7101 (N_7101,N_1116,N_1011);
nor U7102 (N_7102,N_4374,N_573);
and U7103 (N_7103,N_517,N_1915);
nor U7104 (N_7104,N_4469,N_875);
nor U7105 (N_7105,N_4993,N_2682);
nand U7106 (N_7106,N_3663,N_1235);
nand U7107 (N_7107,N_3764,N_2664);
nand U7108 (N_7108,N_456,N_1111);
nor U7109 (N_7109,N_3804,N_659);
nand U7110 (N_7110,N_1596,N_425);
and U7111 (N_7111,N_475,N_4060);
or U7112 (N_7112,N_205,N_962);
and U7113 (N_7113,N_4286,N_995);
and U7114 (N_7114,N_2028,N_681);
or U7115 (N_7115,N_2627,N_3720);
or U7116 (N_7116,N_780,N_1053);
and U7117 (N_7117,N_3341,N_769);
and U7118 (N_7118,N_492,N_839);
nor U7119 (N_7119,N_1169,N_4521);
nor U7120 (N_7120,N_3863,N_420);
and U7121 (N_7121,N_3367,N_3596);
nand U7122 (N_7122,N_390,N_2740);
or U7123 (N_7123,N_2670,N_1736);
nor U7124 (N_7124,N_1342,N_2571);
nand U7125 (N_7125,N_4814,N_3889);
nor U7126 (N_7126,N_1263,N_3319);
nor U7127 (N_7127,N_3153,N_3018);
and U7128 (N_7128,N_4251,N_4915);
or U7129 (N_7129,N_382,N_2926);
xor U7130 (N_7130,N_4373,N_1564);
nor U7131 (N_7131,N_770,N_2243);
or U7132 (N_7132,N_3588,N_3520);
and U7133 (N_7133,N_2491,N_3869);
nor U7134 (N_7134,N_3412,N_1375);
and U7135 (N_7135,N_2896,N_4929);
nand U7136 (N_7136,N_2440,N_1299);
and U7137 (N_7137,N_136,N_2104);
and U7138 (N_7138,N_2015,N_1737);
nand U7139 (N_7139,N_486,N_1124);
and U7140 (N_7140,N_1630,N_4560);
nor U7141 (N_7141,N_279,N_3066);
and U7142 (N_7142,N_856,N_1028);
nor U7143 (N_7143,N_346,N_4834);
nand U7144 (N_7144,N_4114,N_3300);
xor U7145 (N_7145,N_3632,N_4024);
nor U7146 (N_7146,N_3191,N_2211);
nor U7147 (N_7147,N_4020,N_3494);
xor U7148 (N_7148,N_1349,N_4954);
or U7149 (N_7149,N_2382,N_732);
nor U7150 (N_7150,N_534,N_4636);
and U7151 (N_7151,N_185,N_233);
nor U7152 (N_7152,N_3919,N_1229);
and U7153 (N_7153,N_1558,N_1127);
nand U7154 (N_7154,N_1002,N_900);
and U7155 (N_7155,N_1716,N_1134);
xor U7156 (N_7156,N_1103,N_364);
and U7157 (N_7157,N_2338,N_3927);
nand U7158 (N_7158,N_4820,N_429);
nand U7159 (N_7159,N_3652,N_480);
and U7160 (N_7160,N_1457,N_1261);
or U7161 (N_7161,N_3443,N_4535);
xnor U7162 (N_7162,N_650,N_1018);
nor U7163 (N_7163,N_208,N_3376);
nand U7164 (N_7164,N_4987,N_317);
and U7165 (N_7165,N_2594,N_3583);
nor U7166 (N_7166,N_4506,N_760);
nor U7167 (N_7167,N_4267,N_4829);
and U7168 (N_7168,N_641,N_3461);
nand U7169 (N_7169,N_689,N_1156);
nor U7170 (N_7170,N_439,N_2854);
nor U7171 (N_7171,N_4058,N_2);
nor U7172 (N_7172,N_4804,N_1671);
and U7173 (N_7173,N_297,N_10);
or U7174 (N_7174,N_3323,N_4858);
and U7175 (N_7175,N_3638,N_1079);
and U7176 (N_7176,N_2064,N_244);
nor U7177 (N_7177,N_1537,N_1616);
nand U7178 (N_7178,N_3373,N_4262);
or U7179 (N_7179,N_703,N_1867);
and U7180 (N_7180,N_4616,N_2633);
nand U7181 (N_7181,N_3620,N_156);
nand U7182 (N_7182,N_1862,N_1231);
nand U7183 (N_7183,N_2142,N_976);
or U7184 (N_7184,N_2231,N_4851);
and U7185 (N_7185,N_1225,N_318);
nor U7186 (N_7186,N_3669,N_2743);
nor U7187 (N_7187,N_1020,N_1728);
or U7188 (N_7188,N_1100,N_782);
nor U7189 (N_7189,N_1284,N_1595);
and U7190 (N_7190,N_357,N_1247);
nand U7191 (N_7191,N_1654,N_1437);
nand U7192 (N_7192,N_4092,N_1168);
and U7193 (N_7193,N_2331,N_263);
nand U7194 (N_7194,N_2804,N_3045);
nor U7195 (N_7195,N_143,N_1400);
and U7196 (N_7196,N_2328,N_1155);
nor U7197 (N_7197,N_3851,N_4317);
and U7198 (N_7198,N_4605,N_1059);
xnor U7199 (N_7199,N_2367,N_4302);
nor U7200 (N_7200,N_1669,N_3398);
nand U7201 (N_7201,N_4393,N_2020);
nand U7202 (N_7202,N_295,N_3908);
nand U7203 (N_7203,N_4957,N_4122);
nor U7204 (N_7204,N_756,N_4488);
nor U7205 (N_7205,N_4580,N_520);
nor U7206 (N_7206,N_403,N_4265);
or U7207 (N_7207,N_3038,N_4461);
nand U7208 (N_7208,N_4735,N_1777);
or U7209 (N_7209,N_334,N_3732);
nand U7210 (N_7210,N_4592,N_3436);
and U7211 (N_7211,N_3144,N_2871);
nor U7212 (N_7212,N_4118,N_1895);
nor U7213 (N_7213,N_1624,N_2427);
and U7214 (N_7214,N_2578,N_2488);
nand U7215 (N_7215,N_4490,N_1831);
and U7216 (N_7216,N_3392,N_3257);
nand U7217 (N_7217,N_2645,N_1949);
nor U7218 (N_7218,N_1092,N_568);
nor U7219 (N_7219,N_4780,N_487);
nand U7220 (N_7220,N_4733,N_4571);
or U7221 (N_7221,N_2864,N_2759);
xnor U7222 (N_7222,N_1642,N_4072);
xor U7223 (N_7223,N_1607,N_4112);
and U7224 (N_7224,N_3735,N_4622);
nand U7225 (N_7225,N_1252,N_4425);
and U7226 (N_7226,N_229,N_3704);
or U7227 (N_7227,N_1674,N_4297);
and U7228 (N_7228,N_4787,N_3327);
or U7229 (N_7229,N_3194,N_1137);
and U7230 (N_7230,N_3220,N_4090);
and U7231 (N_7231,N_4895,N_3283);
or U7232 (N_7232,N_4131,N_2965);
nor U7233 (N_7233,N_4170,N_3180);
and U7234 (N_7234,N_4141,N_903);
and U7235 (N_7235,N_4603,N_137);
and U7236 (N_7236,N_4298,N_939);
and U7237 (N_7237,N_0,N_3458);
nor U7238 (N_7238,N_4372,N_4099);
nor U7239 (N_7239,N_435,N_132);
or U7240 (N_7240,N_4520,N_544);
nor U7241 (N_7241,N_584,N_661);
and U7242 (N_7242,N_3845,N_30);
nor U7243 (N_7243,N_3044,N_1694);
and U7244 (N_7244,N_3595,N_1965);
and U7245 (N_7245,N_2341,N_3647);
nor U7246 (N_7246,N_804,N_2174);
or U7247 (N_7247,N_4749,N_4102);
or U7248 (N_7248,N_2739,N_1807);
nand U7249 (N_7249,N_2808,N_966);
nor U7250 (N_7250,N_239,N_2417);
or U7251 (N_7251,N_226,N_4066);
nor U7252 (N_7252,N_1286,N_2746);
nand U7253 (N_7253,N_4724,N_3821);
and U7254 (N_7254,N_2866,N_551);
nor U7255 (N_7255,N_4703,N_4394);
xnor U7256 (N_7256,N_3930,N_954);
or U7257 (N_7257,N_235,N_3848);
nor U7258 (N_7258,N_2190,N_1393);
and U7259 (N_7259,N_265,N_3337);
nand U7260 (N_7260,N_3772,N_4885);
and U7261 (N_7261,N_2640,N_4143);
nor U7262 (N_7262,N_4641,N_1772);
nand U7263 (N_7263,N_4773,N_777);
nand U7264 (N_7264,N_4119,N_4771);
and U7265 (N_7265,N_2794,N_4509);
and U7266 (N_7266,N_4337,N_4497);
and U7267 (N_7267,N_469,N_4855);
xnor U7268 (N_7268,N_888,N_1559);
or U7269 (N_7269,N_3901,N_3129);
nor U7270 (N_7270,N_1833,N_1291);
nor U7271 (N_7271,N_2800,N_4876);
xnor U7272 (N_7272,N_247,N_4729);
nand U7273 (N_7273,N_4105,N_3951);
nor U7274 (N_7274,N_1891,N_627);
nand U7275 (N_7275,N_774,N_479);
or U7276 (N_7276,N_2958,N_4727);
and U7277 (N_7277,N_2343,N_2657);
or U7278 (N_7278,N_3631,N_735);
and U7279 (N_7279,N_3886,N_992);
nand U7280 (N_7280,N_1099,N_614);
xnor U7281 (N_7281,N_406,N_1461);
nor U7282 (N_7282,N_1434,N_2271);
or U7283 (N_7283,N_3707,N_612);
and U7284 (N_7284,N_1631,N_2636);
and U7285 (N_7285,N_1034,N_1148);
and U7286 (N_7286,N_1591,N_4608);
nor U7287 (N_7287,N_2562,N_1548);
nor U7288 (N_7288,N_3681,N_3197);
nand U7289 (N_7289,N_460,N_2693);
and U7290 (N_7290,N_1892,N_1330);
or U7291 (N_7291,N_2511,N_561);
and U7292 (N_7292,N_332,N_3176);
nand U7293 (N_7293,N_632,N_3004);
or U7294 (N_7294,N_1324,N_1946);
or U7295 (N_7295,N_3128,N_2818);
or U7296 (N_7296,N_389,N_2923);
or U7297 (N_7297,N_2720,N_1739);
nor U7298 (N_7298,N_2967,N_4080);
nor U7299 (N_7299,N_1445,N_1472);
nor U7300 (N_7300,N_1514,N_343);
nor U7301 (N_7301,N_3296,N_186);
and U7302 (N_7302,N_1479,N_3805);
and U7303 (N_7303,N_4482,N_1874);
nor U7304 (N_7304,N_1599,N_812);
or U7305 (N_7305,N_1207,N_1923);
and U7306 (N_7306,N_846,N_78);
nand U7307 (N_7307,N_2265,N_4318);
nor U7308 (N_7308,N_1463,N_1323);
and U7309 (N_7309,N_4587,N_3766);
and U7310 (N_7310,N_2398,N_4494);
or U7311 (N_7311,N_331,N_3448);
nand U7312 (N_7312,N_2262,N_3061);
and U7313 (N_7313,N_135,N_642);
or U7314 (N_7314,N_4806,N_2925);
nor U7315 (N_7315,N_1451,N_3789);
and U7316 (N_7316,N_4070,N_1189);
nor U7317 (N_7317,N_4910,N_1732);
nor U7318 (N_7318,N_1756,N_1761);
and U7319 (N_7319,N_4061,N_1175);
or U7320 (N_7320,N_542,N_704);
and U7321 (N_7321,N_1960,N_1325);
or U7322 (N_7322,N_3655,N_4219);
and U7323 (N_7323,N_2505,N_3509);
or U7324 (N_7324,N_1582,N_1864);
nand U7325 (N_7325,N_4977,N_2557);
xnor U7326 (N_7326,N_4087,N_3280);
or U7327 (N_7327,N_423,N_1770);
nand U7328 (N_7328,N_4822,N_4440);
nand U7329 (N_7329,N_85,N_3022);
or U7330 (N_7330,N_3055,N_3161);
and U7331 (N_7331,N_3046,N_2839);
and U7332 (N_7332,N_220,N_2196);
nand U7333 (N_7333,N_2914,N_4567);
or U7334 (N_7334,N_3839,N_4546);
or U7335 (N_7335,N_3714,N_3551);
and U7336 (N_7336,N_1541,N_3974);
nand U7337 (N_7337,N_3216,N_4530);
nor U7338 (N_7338,N_2258,N_4409);
nor U7339 (N_7339,N_3967,N_3057);
or U7340 (N_7340,N_2209,N_1979);
xnor U7341 (N_7341,N_4778,N_635);
nand U7342 (N_7342,N_3871,N_264);
and U7343 (N_7343,N_3654,N_3060);
nor U7344 (N_7344,N_5,N_2303);
and U7345 (N_7345,N_4623,N_775);
or U7346 (N_7346,N_2599,N_3483);
or U7347 (N_7347,N_1236,N_4523);
nor U7348 (N_7348,N_2177,N_354);
or U7349 (N_7349,N_4857,N_274);
nand U7350 (N_7350,N_2834,N_4030);
nor U7351 (N_7351,N_1361,N_1471);
and U7352 (N_7352,N_4353,N_2799);
nor U7353 (N_7353,N_692,N_4930);
nor U7354 (N_7354,N_2485,N_4875);
nand U7355 (N_7355,N_1288,N_1487);
nand U7356 (N_7356,N_2615,N_1427);
nor U7357 (N_7357,N_1904,N_1927);
nand U7358 (N_7358,N_1953,N_1198);
and U7359 (N_7359,N_4926,N_1456);
nand U7360 (N_7360,N_4797,N_4156);
xor U7361 (N_7361,N_3711,N_4962);
and U7362 (N_7362,N_1255,N_1141);
and U7363 (N_7363,N_2253,N_3135);
nor U7364 (N_7364,N_4137,N_871);
and U7365 (N_7365,N_3891,N_4920);
nand U7366 (N_7366,N_3568,N_169);
or U7367 (N_7367,N_828,N_3033);
or U7368 (N_7368,N_36,N_699);
nor U7369 (N_7369,N_2731,N_2465);
xor U7370 (N_7370,N_3939,N_691);
xnor U7371 (N_7371,N_2943,N_2140);
nand U7372 (N_7372,N_944,N_1201);
nor U7373 (N_7373,N_31,N_4500);
nand U7374 (N_7374,N_2109,N_2490);
nand U7375 (N_7375,N_3105,N_897);
or U7376 (N_7376,N_2736,N_3911);
nor U7377 (N_7377,N_4980,N_3237);
or U7378 (N_7378,N_1721,N_4495);
and U7379 (N_7379,N_4404,N_4320);
nor U7380 (N_7380,N_652,N_4465);
nand U7381 (N_7381,N_876,N_1081);
or U7382 (N_7382,N_671,N_4896);
or U7383 (N_7383,N_834,N_1365);
nor U7384 (N_7384,N_2167,N_2725);
and U7385 (N_7385,N_2976,N_738);
or U7386 (N_7386,N_1145,N_2363);
and U7387 (N_7387,N_1797,N_4123);
or U7388 (N_7388,N_4630,N_914);
or U7389 (N_7389,N_2729,N_3697);
or U7390 (N_7390,N_832,N_1416);
nand U7391 (N_7391,N_827,N_2339);
or U7392 (N_7392,N_193,N_2863);
and U7393 (N_7393,N_4388,N_3203);
xor U7394 (N_7394,N_1282,N_3139);
xor U7395 (N_7395,N_1006,N_1290);
or U7396 (N_7396,N_4120,N_577);
or U7397 (N_7397,N_2026,N_1655);
xor U7398 (N_7398,N_2350,N_753);
nand U7399 (N_7399,N_4539,N_1873);
or U7400 (N_7400,N_2619,N_3585);
nand U7401 (N_7401,N_2584,N_1835);
xnor U7402 (N_7402,N_4997,N_1526);
or U7403 (N_7403,N_2737,N_2497);
and U7404 (N_7404,N_1031,N_2473);
nor U7405 (N_7405,N_3386,N_896);
nand U7406 (N_7406,N_1925,N_4169);
nand U7407 (N_7407,N_2252,N_4071);
nor U7408 (N_7408,N_489,N_3787);
xor U7409 (N_7409,N_4604,N_1017);
and U7410 (N_7410,N_1688,N_2130);
or U7411 (N_7411,N_2494,N_1788);
nand U7412 (N_7412,N_3265,N_3322);
and U7413 (N_7413,N_2429,N_637);
nor U7414 (N_7414,N_1082,N_3826);
and U7415 (N_7415,N_2676,N_2310);
nor U7416 (N_7416,N_1192,N_3052);
and U7417 (N_7417,N_2770,N_2517);
and U7418 (N_7418,N_2969,N_3434);
nor U7419 (N_7419,N_1242,N_696);
nor U7420 (N_7420,N_1667,N_2423);
xnor U7421 (N_7421,N_55,N_2397);
nand U7422 (N_7422,N_1530,N_3068);
and U7423 (N_7423,N_3452,N_158);
and U7424 (N_7424,N_4688,N_2846);
or U7425 (N_7425,N_2970,N_3079);
or U7426 (N_7426,N_2848,N_3517);
nand U7427 (N_7427,N_2279,N_4128);
or U7428 (N_7428,N_29,N_2726);
nand U7429 (N_7429,N_2447,N_4779);
or U7430 (N_7430,N_1884,N_4115);
nand U7431 (N_7431,N_3530,N_2850);
nand U7432 (N_7432,N_4150,N_25);
or U7433 (N_7433,N_675,N_3827);
nand U7434 (N_7434,N_1620,N_2626);
and U7435 (N_7435,N_4236,N_1592);
nand U7436 (N_7436,N_1354,N_773);
xnor U7437 (N_7437,N_2723,N_271);
or U7438 (N_7438,N_3761,N_3253);
and U7439 (N_7439,N_597,N_1491);
nor U7440 (N_7440,N_1295,N_4794);
or U7441 (N_7441,N_2956,N_199);
nand U7442 (N_7442,N_491,N_1724);
nor U7443 (N_7443,N_1131,N_174);
or U7444 (N_7444,N_4548,N_32);
or U7445 (N_7445,N_3428,N_807);
and U7446 (N_7446,N_21,N_3168);
and U7447 (N_7447,N_1725,N_4180);
nand U7448 (N_7448,N_2212,N_4146);
or U7449 (N_7449,N_3643,N_3345);
nor U7450 (N_7450,N_3019,N_3120);
and U7451 (N_7451,N_4395,N_2471);
nor U7452 (N_7452,N_1635,N_3931);
nor U7453 (N_7453,N_2316,N_1363);
and U7454 (N_7454,N_714,N_142);
nand U7455 (N_7455,N_4737,N_2603);
xor U7456 (N_7456,N_2588,N_4032);
xor U7457 (N_7457,N_2981,N_2639);
nor U7458 (N_7458,N_4413,N_2625);
or U7459 (N_7459,N_4266,N_2353);
nor U7460 (N_7460,N_430,N_1428);
or U7461 (N_7461,N_217,N_1758);
xor U7462 (N_7462,N_4812,N_4124);
nand U7463 (N_7463,N_2522,N_2060);
nor U7464 (N_7464,N_755,N_128);
or U7465 (N_7465,N_2775,N_2007);
and U7466 (N_7466,N_2927,N_1705);
nand U7467 (N_7467,N_4305,N_1551);
nand U7468 (N_7468,N_2767,N_860);
or U7469 (N_7469,N_214,N_4275);
nand U7470 (N_7470,N_2772,N_4415);
and U7471 (N_7471,N_4996,N_4867);
and U7472 (N_7472,N_1055,N_1860);
nor U7473 (N_7473,N_987,N_267);
nand U7474 (N_7474,N_4041,N_3490);
xnor U7475 (N_7475,N_2355,N_2049);
xor U7476 (N_7476,N_1390,N_608);
or U7477 (N_7477,N_2827,N_2364);
nand U7478 (N_7478,N_848,N_253);
or U7479 (N_7479,N_1258,N_3427);
nor U7480 (N_7480,N_4692,N_1257);
nor U7481 (N_7481,N_2539,N_3846);
nor U7482 (N_7482,N_2082,N_1274);
nand U7483 (N_7483,N_647,N_2024);
nand U7484 (N_7484,N_4444,N_1401);
or U7485 (N_7485,N_2181,N_2055);
or U7486 (N_7486,N_4043,N_1854);
nand U7487 (N_7487,N_3174,N_4397);
xnor U7488 (N_7488,N_3184,N_1730);
nor U7489 (N_7489,N_2301,N_2062);
nand U7490 (N_7490,N_231,N_4846);
nor U7491 (N_7491,N_1350,N_3251);
xor U7492 (N_7492,N_3329,N_1571);
nand U7493 (N_7493,N_2589,N_2798);
nand U7494 (N_7494,N_4294,N_2149);
or U7495 (N_7495,N_1306,N_119);
or U7496 (N_7496,N_3815,N_3335);
or U7497 (N_7497,N_3108,N_3268);
and U7498 (N_7498,N_368,N_1856);
nor U7499 (N_7499,N_2257,N_2685);
or U7500 (N_7500,N_1474,N_1246);
nand U7501 (N_7501,N_4070,N_162);
and U7502 (N_7502,N_992,N_2899);
xnor U7503 (N_7503,N_3429,N_4859);
and U7504 (N_7504,N_4711,N_477);
or U7505 (N_7505,N_404,N_2621);
and U7506 (N_7506,N_3569,N_575);
nor U7507 (N_7507,N_167,N_1146);
and U7508 (N_7508,N_801,N_2098);
xnor U7509 (N_7509,N_3384,N_1829);
or U7510 (N_7510,N_4895,N_3731);
or U7511 (N_7511,N_508,N_2997);
and U7512 (N_7512,N_1608,N_2572);
and U7513 (N_7513,N_2744,N_1569);
nand U7514 (N_7514,N_2660,N_940);
nand U7515 (N_7515,N_301,N_4234);
nand U7516 (N_7516,N_891,N_4493);
and U7517 (N_7517,N_4315,N_3948);
and U7518 (N_7518,N_1309,N_3578);
and U7519 (N_7519,N_2854,N_2166);
or U7520 (N_7520,N_4633,N_2682);
nor U7521 (N_7521,N_925,N_4968);
and U7522 (N_7522,N_1904,N_3568);
nand U7523 (N_7523,N_2809,N_1510);
or U7524 (N_7524,N_4418,N_3166);
nor U7525 (N_7525,N_1086,N_2162);
nand U7526 (N_7526,N_1332,N_2657);
or U7527 (N_7527,N_3732,N_192);
nand U7528 (N_7528,N_500,N_926);
nor U7529 (N_7529,N_2652,N_3250);
nor U7530 (N_7530,N_3648,N_978);
nor U7531 (N_7531,N_3080,N_606);
or U7532 (N_7532,N_1419,N_544);
and U7533 (N_7533,N_1262,N_857);
nand U7534 (N_7534,N_4227,N_698);
or U7535 (N_7535,N_3311,N_3260);
and U7536 (N_7536,N_3111,N_720);
and U7537 (N_7537,N_3756,N_2085);
nor U7538 (N_7538,N_3227,N_32);
nor U7539 (N_7539,N_2682,N_2801);
and U7540 (N_7540,N_408,N_1481);
nand U7541 (N_7541,N_4230,N_2430);
nand U7542 (N_7542,N_2795,N_3140);
or U7543 (N_7543,N_2870,N_243);
nand U7544 (N_7544,N_52,N_683);
or U7545 (N_7545,N_1684,N_1013);
or U7546 (N_7546,N_2735,N_600);
or U7547 (N_7547,N_3101,N_929);
nand U7548 (N_7548,N_1351,N_3149);
nand U7549 (N_7549,N_664,N_1111);
nor U7550 (N_7550,N_4837,N_1702);
and U7551 (N_7551,N_577,N_1719);
nand U7552 (N_7552,N_3131,N_2100);
nor U7553 (N_7553,N_1691,N_4867);
nand U7554 (N_7554,N_699,N_3443);
and U7555 (N_7555,N_3431,N_725);
and U7556 (N_7556,N_141,N_490);
and U7557 (N_7557,N_745,N_4639);
and U7558 (N_7558,N_1577,N_367);
or U7559 (N_7559,N_2223,N_1706);
nor U7560 (N_7560,N_2782,N_2713);
and U7561 (N_7561,N_358,N_2240);
xnor U7562 (N_7562,N_1225,N_3890);
nor U7563 (N_7563,N_2590,N_1040);
nand U7564 (N_7564,N_3382,N_1993);
nor U7565 (N_7565,N_1622,N_4715);
or U7566 (N_7566,N_849,N_478);
nand U7567 (N_7567,N_3400,N_4994);
nor U7568 (N_7568,N_4345,N_3938);
nor U7569 (N_7569,N_1836,N_4516);
nand U7570 (N_7570,N_1509,N_474);
xor U7571 (N_7571,N_3069,N_1805);
and U7572 (N_7572,N_632,N_4384);
and U7573 (N_7573,N_851,N_2527);
and U7574 (N_7574,N_4442,N_979);
nor U7575 (N_7575,N_678,N_39);
nor U7576 (N_7576,N_2566,N_520);
nor U7577 (N_7577,N_3217,N_4450);
or U7578 (N_7578,N_3968,N_4245);
and U7579 (N_7579,N_4834,N_4348);
xor U7580 (N_7580,N_1489,N_434);
or U7581 (N_7581,N_4849,N_90);
xnor U7582 (N_7582,N_2021,N_1372);
or U7583 (N_7583,N_3770,N_4937);
and U7584 (N_7584,N_2778,N_1233);
or U7585 (N_7585,N_2578,N_1048);
nand U7586 (N_7586,N_1086,N_803);
nor U7587 (N_7587,N_1439,N_4652);
and U7588 (N_7588,N_1243,N_2629);
nor U7589 (N_7589,N_338,N_316);
nand U7590 (N_7590,N_1526,N_2674);
nor U7591 (N_7591,N_1032,N_3278);
nand U7592 (N_7592,N_489,N_1013);
or U7593 (N_7593,N_1502,N_4525);
nand U7594 (N_7594,N_4771,N_418);
nand U7595 (N_7595,N_1493,N_1476);
and U7596 (N_7596,N_2181,N_292);
and U7597 (N_7597,N_4437,N_4543);
xnor U7598 (N_7598,N_427,N_2684);
xnor U7599 (N_7599,N_1710,N_2048);
xor U7600 (N_7600,N_4247,N_344);
and U7601 (N_7601,N_1441,N_2871);
nand U7602 (N_7602,N_3717,N_2239);
nor U7603 (N_7603,N_3369,N_3293);
nor U7604 (N_7604,N_1346,N_4083);
or U7605 (N_7605,N_1848,N_526);
or U7606 (N_7606,N_2608,N_4912);
nor U7607 (N_7607,N_2406,N_3267);
nand U7608 (N_7608,N_1846,N_3360);
or U7609 (N_7609,N_3789,N_625);
and U7610 (N_7610,N_2271,N_2460);
or U7611 (N_7611,N_1229,N_1010);
nor U7612 (N_7612,N_3147,N_2647);
and U7613 (N_7613,N_3199,N_4413);
nor U7614 (N_7614,N_4024,N_1509);
nand U7615 (N_7615,N_4016,N_3150);
or U7616 (N_7616,N_2507,N_1685);
or U7617 (N_7617,N_4533,N_3124);
xor U7618 (N_7618,N_4811,N_4376);
or U7619 (N_7619,N_2447,N_170);
or U7620 (N_7620,N_1893,N_3468);
nor U7621 (N_7621,N_1753,N_2424);
nor U7622 (N_7622,N_829,N_1289);
nor U7623 (N_7623,N_30,N_2801);
nor U7624 (N_7624,N_1586,N_4751);
nor U7625 (N_7625,N_922,N_4857);
and U7626 (N_7626,N_3691,N_1010);
and U7627 (N_7627,N_1914,N_3041);
nand U7628 (N_7628,N_2809,N_4053);
and U7629 (N_7629,N_2534,N_2754);
and U7630 (N_7630,N_3929,N_4984);
nand U7631 (N_7631,N_448,N_1927);
and U7632 (N_7632,N_741,N_2467);
or U7633 (N_7633,N_4862,N_3826);
and U7634 (N_7634,N_3289,N_4824);
nor U7635 (N_7635,N_4547,N_4966);
nor U7636 (N_7636,N_2361,N_4522);
and U7637 (N_7637,N_3526,N_3383);
and U7638 (N_7638,N_362,N_2415);
or U7639 (N_7639,N_4566,N_1393);
nor U7640 (N_7640,N_2045,N_4976);
nand U7641 (N_7641,N_2338,N_3988);
nor U7642 (N_7642,N_4788,N_3895);
nand U7643 (N_7643,N_2471,N_867);
nor U7644 (N_7644,N_1421,N_2376);
nand U7645 (N_7645,N_819,N_3929);
or U7646 (N_7646,N_3974,N_4913);
nand U7647 (N_7647,N_2709,N_2645);
or U7648 (N_7648,N_1804,N_2655);
nor U7649 (N_7649,N_4590,N_3416);
nand U7650 (N_7650,N_4262,N_3520);
or U7651 (N_7651,N_3753,N_3999);
nor U7652 (N_7652,N_733,N_2768);
and U7653 (N_7653,N_1184,N_317);
and U7654 (N_7654,N_3835,N_223);
nor U7655 (N_7655,N_1579,N_3435);
xnor U7656 (N_7656,N_4562,N_82);
nand U7657 (N_7657,N_4477,N_852);
nand U7658 (N_7658,N_608,N_602);
nand U7659 (N_7659,N_1146,N_299);
nand U7660 (N_7660,N_1039,N_1252);
xor U7661 (N_7661,N_256,N_3905);
nand U7662 (N_7662,N_991,N_2716);
xor U7663 (N_7663,N_1266,N_297);
nor U7664 (N_7664,N_4764,N_832);
nand U7665 (N_7665,N_983,N_4128);
nand U7666 (N_7666,N_122,N_541);
and U7667 (N_7667,N_626,N_1179);
xnor U7668 (N_7668,N_1806,N_2675);
nand U7669 (N_7669,N_1470,N_928);
or U7670 (N_7670,N_3368,N_4264);
nand U7671 (N_7671,N_71,N_3452);
and U7672 (N_7672,N_2998,N_2070);
nor U7673 (N_7673,N_3331,N_876);
or U7674 (N_7674,N_1661,N_2861);
nor U7675 (N_7675,N_1567,N_124);
nor U7676 (N_7676,N_2483,N_3574);
or U7677 (N_7677,N_3859,N_336);
and U7678 (N_7678,N_1017,N_1067);
or U7679 (N_7679,N_2108,N_3661);
and U7680 (N_7680,N_4058,N_2893);
and U7681 (N_7681,N_3720,N_4961);
and U7682 (N_7682,N_4460,N_1817);
or U7683 (N_7683,N_1461,N_4063);
and U7684 (N_7684,N_4155,N_4078);
nor U7685 (N_7685,N_3996,N_949);
nand U7686 (N_7686,N_2026,N_3432);
and U7687 (N_7687,N_1142,N_3346);
and U7688 (N_7688,N_2116,N_4748);
nand U7689 (N_7689,N_1433,N_844);
nand U7690 (N_7690,N_4622,N_3883);
nand U7691 (N_7691,N_3647,N_2915);
nand U7692 (N_7692,N_904,N_781);
nand U7693 (N_7693,N_4194,N_522);
nor U7694 (N_7694,N_1830,N_4961);
nand U7695 (N_7695,N_2551,N_2832);
or U7696 (N_7696,N_4792,N_3157);
nor U7697 (N_7697,N_3032,N_3557);
nor U7698 (N_7698,N_1364,N_4397);
xor U7699 (N_7699,N_4297,N_1591);
and U7700 (N_7700,N_684,N_3163);
nand U7701 (N_7701,N_767,N_1982);
nor U7702 (N_7702,N_1958,N_4441);
and U7703 (N_7703,N_4442,N_4230);
xor U7704 (N_7704,N_551,N_3431);
nand U7705 (N_7705,N_1498,N_721);
or U7706 (N_7706,N_4957,N_3908);
nand U7707 (N_7707,N_352,N_4406);
xor U7708 (N_7708,N_1793,N_2860);
and U7709 (N_7709,N_90,N_1334);
nand U7710 (N_7710,N_3991,N_2298);
xnor U7711 (N_7711,N_2478,N_4447);
nor U7712 (N_7712,N_3733,N_1033);
and U7713 (N_7713,N_2926,N_628);
and U7714 (N_7714,N_740,N_3154);
or U7715 (N_7715,N_741,N_2789);
or U7716 (N_7716,N_1219,N_1882);
nand U7717 (N_7717,N_800,N_2488);
nor U7718 (N_7718,N_3709,N_2538);
nand U7719 (N_7719,N_2681,N_12);
nand U7720 (N_7720,N_4896,N_4549);
or U7721 (N_7721,N_3117,N_3131);
and U7722 (N_7722,N_4221,N_754);
and U7723 (N_7723,N_3668,N_1544);
nand U7724 (N_7724,N_1998,N_2623);
and U7725 (N_7725,N_3339,N_3939);
xnor U7726 (N_7726,N_4502,N_402);
and U7727 (N_7727,N_2410,N_4530);
and U7728 (N_7728,N_3611,N_815);
nor U7729 (N_7729,N_237,N_3475);
and U7730 (N_7730,N_3265,N_3409);
or U7731 (N_7731,N_1384,N_4946);
and U7732 (N_7732,N_3552,N_1051);
or U7733 (N_7733,N_658,N_2177);
or U7734 (N_7734,N_2123,N_4381);
nor U7735 (N_7735,N_1245,N_1125);
and U7736 (N_7736,N_3513,N_1058);
nand U7737 (N_7737,N_3236,N_4830);
xnor U7738 (N_7738,N_1244,N_461);
nor U7739 (N_7739,N_1242,N_3308);
nor U7740 (N_7740,N_571,N_3457);
and U7741 (N_7741,N_4029,N_3206);
or U7742 (N_7742,N_4510,N_3430);
or U7743 (N_7743,N_1822,N_1034);
and U7744 (N_7744,N_369,N_2871);
xnor U7745 (N_7745,N_3893,N_2943);
or U7746 (N_7746,N_4947,N_2380);
or U7747 (N_7747,N_883,N_4849);
or U7748 (N_7748,N_120,N_3704);
nor U7749 (N_7749,N_139,N_2348);
and U7750 (N_7750,N_4321,N_1393);
xor U7751 (N_7751,N_1897,N_3703);
and U7752 (N_7752,N_4345,N_4157);
nand U7753 (N_7753,N_646,N_4295);
nand U7754 (N_7754,N_3958,N_1822);
or U7755 (N_7755,N_1843,N_2576);
xnor U7756 (N_7756,N_4763,N_884);
xor U7757 (N_7757,N_4565,N_3625);
nor U7758 (N_7758,N_2131,N_3067);
or U7759 (N_7759,N_1043,N_3103);
nand U7760 (N_7760,N_4075,N_3718);
nand U7761 (N_7761,N_1555,N_2507);
or U7762 (N_7762,N_2695,N_4777);
nor U7763 (N_7763,N_38,N_2920);
nand U7764 (N_7764,N_4360,N_1892);
xnor U7765 (N_7765,N_1149,N_4123);
xnor U7766 (N_7766,N_734,N_1521);
or U7767 (N_7767,N_4736,N_1575);
and U7768 (N_7768,N_3831,N_219);
xor U7769 (N_7769,N_1290,N_1265);
and U7770 (N_7770,N_4214,N_4795);
or U7771 (N_7771,N_3318,N_3339);
and U7772 (N_7772,N_2908,N_4957);
nor U7773 (N_7773,N_2601,N_2106);
or U7774 (N_7774,N_4865,N_2440);
nor U7775 (N_7775,N_4415,N_2648);
xor U7776 (N_7776,N_115,N_3811);
nand U7777 (N_7777,N_4017,N_2661);
xnor U7778 (N_7778,N_3563,N_353);
nand U7779 (N_7779,N_4633,N_823);
or U7780 (N_7780,N_1152,N_4231);
nor U7781 (N_7781,N_387,N_3065);
or U7782 (N_7782,N_1355,N_645);
xor U7783 (N_7783,N_1931,N_1797);
and U7784 (N_7784,N_2412,N_3677);
nor U7785 (N_7785,N_4116,N_1762);
or U7786 (N_7786,N_3426,N_1642);
nand U7787 (N_7787,N_2285,N_1761);
nand U7788 (N_7788,N_1460,N_4120);
xnor U7789 (N_7789,N_739,N_3454);
nand U7790 (N_7790,N_4703,N_860);
and U7791 (N_7791,N_1370,N_892);
nand U7792 (N_7792,N_3031,N_1414);
or U7793 (N_7793,N_672,N_3311);
nand U7794 (N_7794,N_4041,N_1457);
nand U7795 (N_7795,N_328,N_1877);
xor U7796 (N_7796,N_1012,N_4601);
or U7797 (N_7797,N_1007,N_406);
and U7798 (N_7798,N_4013,N_503);
nand U7799 (N_7799,N_3640,N_4324);
xor U7800 (N_7800,N_3515,N_3709);
nor U7801 (N_7801,N_2817,N_1268);
or U7802 (N_7802,N_3191,N_3479);
nand U7803 (N_7803,N_1361,N_701);
or U7804 (N_7804,N_4319,N_4555);
nor U7805 (N_7805,N_3884,N_2445);
nor U7806 (N_7806,N_3228,N_4807);
nand U7807 (N_7807,N_531,N_964);
nor U7808 (N_7808,N_3250,N_2015);
xnor U7809 (N_7809,N_355,N_3096);
or U7810 (N_7810,N_4353,N_3000);
nor U7811 (N_7811,N_4110,N_2493);
and U7812 (N_7812,N_1197,N_479);
xor U7813 (N_7813,N_4469,N_2001);
or U7814 (N_7814,N_4338,N_488);
or U7815 (N_7815,N_983,N_2538);
xor U7816 (N_7816,N_85,N_2978);
or U7817 (N_7817,N_2159,N_439);
nor U7818 (N_7818,N_2431,N_3520);
nor U7819 (N_7819,N_192,N_2739);
or U7820 (N_7820,N_4974,N_843);
xor U7821 (N_7821,N_1738,N_368);
xor U7822 (N_7822,N_852,N_1877);
or U7823 (N_7823,N_4090,N_3442);
and U7824 (N_7824,N_1000,N_1916);
and U7825 (N_7825,N_169,N_753);
and U7826 (N_7826,N_1954,N_2454);
nand U7827 (N_7827,N_2885,N_948);
or U7828 (N_7828,N_4053,N_3219);
and U7829 (N_7829,N_1735,N_419);
nor U7830 (N_7830,N_140,N_1241);
or U7831 (N_7831,N_2925,N_2857);
or U7832 (N_7832,N_711,N_958);
nor U7833 (N_7833,N_286,N_369);
and U7834 (N_7834,N_2558,N_2857);
nand U7835 (N_7835,N_4261,N_3262);
nor U7836 (N_7836,N_55,N_2882);
nor U7837 (N_7837,N_3512,N_3106);
or U7838 (N_7838,N_328,N_3849);
nand U7839 (N_7839,N_2845,N_3295);
xor U7840 (N_7840,N_4948,N_2662);
or U7841 (N_7841,N_233,N_4755);
nor U7842 (N_7842,N_1455,N_2514);
nand U7843 (N_7843,N_290,N_1129);
and U7844 (N_7844,N_818,N_1842);
or U7845 (N_7845,N_2223,N_4582);
nor U7846 (N_7846,N_3678,N_399);
nor U7847 (N_7847,N_4917,N_2847);
nor U7848 (N_7848,N_2494,N_2865);
nor U7849 (N_7849,N_1991,N_2801);
nor U7850 (N_7850,N_84,N_4603);
nor U7851 (N_7851,N_2728,N_3690);
or U7852 (N_7852,N_344,N_4931);
xnor U7853 (N_7853,N_1966,N_1504);
or U7854 (N_7854,N_2998,N_2812);
nor U7855 (N_7855,N_3196,N_3572);
nor U7856 (N_7856,N_1817,N_1911);
nor U7857 (N_7857,N_2569,N_577);
or U7858 (N_7858,N_120,N_2873);
or U7859 (N_7859,N_86,N_4197);
xnor U7860 (N_7860,N_3657,N_761);
and U7861 (N_7861,N_4284,N_533);
nor U7862 (N_7862,N_3080,N_851);
or U7863 (N_7863,N_1476,N_4790);
and U7864 (N_7864,N_2471,N_3498);
and U7865 (N_7865,N_424,N_2475);
nor U7866 (N_7866,N_1852,N_964);
and U7867 (N_7867,N_4940,N_4386);
nand U7868 (N_7868,N_164,N_1185);
and U7869 (N_7869,N_1015,N_834);
and U7870 (N_7870,N_2693,N_4997);
or U7871 (N_7871,N_11,N_4068);
nand U7872 (N_7872,N_870,N_2829);
nor U7873 (N_7873,N_1722,N_3375);
or U7874 (N_7874,N_2021,N_659);
and U7875 (N_7875,N_2496,N_947);
nand U7876 (N_7876,N_151,N_508);
nor U7877 (N_7877,N_663,N_4405);
and U7878 (N_7878,N_3415,N_1589);
and U7879 (N_7879,N_883,N_3100);
nor U7880 (N_7880,N_2502,N_2284);
nand U7881 (N_7881,N_2638,N_185);
nor U7882 (N_7882,N_1900,N_4798);
nand U7883 (N_7883,N_3412,N_4365);
nand U7884 (N_7884,N_1991,N_3547);
and U7885 (N_7885,N_4296,N_1314);
nor U7886 (N_7886,N_463,N_978);
and U7887 (N_7887,N_2743,N_582);
nand U7888 (N_7888,N_1567,N_238);
nand U7889 (N_7889,N_4052,N_4040);
nand U7890 (N_7890,N_2472,N_3515);
and U7891 (N_7891,N_416,N_679);
or U7892 (N_7892,N_4705,N_3306);
xnor U7893 (N_7893,N_4801,N_4470);
nor U7894 (N_7894,N_1051,N_4691);
or U7895 (N_7895,N_26,N_180);
nand U7896 (N_7896,N_500,N_4901);
or U7897 (N_7897,N_1308,N_2392);
and U7898 (N_7898,N_4896,N_4834);
and U7899 (N_7899,N_3396,N_1421);
nor U7900 (N_7900,N_3335,N_1100);
and U7901 (N_7901,N_1643,N_1835);
and U7902 (N_7902,N_2294,N_3041);
or U7903 (N_7903,N_3533,N_1076);
nand U7904 (N_7904,N_1059,N_2709);
and U7905 (N_7905,N_4234,N_318);
xnor U7906 (N_7906,N_4818,N_182);
nor U7907 (N_7907,N_2678,N_2908);
nor U7908 (N_7908,N_414,N_56);
nor U7909 (N_7909,N_2670,N_2397);
nor U7910 (N_7910,N_2174,N_2477);
nor U7911 (N_7911,N_3623,N_3936);
nand U7912 (N_7912,N_1527,N_721);
and U7913 (N_7913,N_2570,N_2054);
xor U7914 (N_7914,N_2053,N_3529);
and U7915 (N_7915,N_1960,N_4399);
and U7916 (N_7916,N_322,N_840);
nand U7917 (N_7917,N_722,N_1780);
xor U7918 (N_7918,N_2792,N_2267);
and U7919 (N_7919,N_3923,N_1597);
or U7920 (N_7920,N_928,N_2287);
nand U7921 (N_7921,N_3547,N_1015);
or U7922 (N_7922,N_3430,N_1272);
nor U7923 (N_7923,N_4363,N_282);
or U7924 (N_7924,N_3835,N_13);
nor U7925 (N_7925,N_4460,N_482);
and U7926 (N_7926,N_1872,N_4166);
nor U7927 (N_7927,N_4079,N_4593);
nand U7928 (N_7928,N_2981,N_2590);
or U7929 (N_7929,N_4056,N_4080);
or U7930 (N_7930,N_690,N_3762);
nand U7931 (N_7931,N_4285,N_1608);
nand U7932 (N_7932,N_2041,N_2393);
nor U7933 (N_7933,N_4825,N_2392);
or U7934 (N_7934,N_3448,N_4973);
and U7935 (N_7935,N_3726,N_2455);
or U7936 (N_7936,N_1536,N_1440);
or U7937 (N_7937,N_3281,N_3309);
nor U7938 (N_7938,N_1188,N_1245);
or U7939 (N_7939,N_4945,N_4253);
and U7940 (N_7940,N_4641,N_1017);
and U7941 (N_7941,N_3890,N_4346);
nand U7942 (N_7942,N_2811,N_1);
xnor U7943 (N_7943,N_3971,N_3273);
nor U7944 (N_7944,N_4368,N_2965);
or U7945 (N_7945,N_142,N_3843);
nand U7946 (N_7946,N_1480,N_970);
nand U7947 (N_7947,N_796,N_3623);
nor U7948 (N_7948,N_1976,N_2832);
xnor U7949 (N_7949,N_2909,N_2417);
nor U7950 (N_7950,N_1425,N_575);
and U7951 (N_7951,N_4934,N_445);
xor U7952 (N_7952,N_1136,N_2656);
or U7953 (N_7953,N_4984,N_953);
and U7954 (N_7954,N_2902,N_1831);
nor U7955 (N_7955,N_2796,N_2020);
and U7956 (N_7956,N_2440,N_2487);
nand U7957 (N_7957,N_2648,N_87);
nor U7958 (N_7958,N_1831,N_3432);
nor U7959 (N_7959,N_885,N_142);
or U7960 (N_7960,N_4210,N_3647);
nor U7961 (N_7961,N_1007,N_821);
nor U7962 (N_7962,N_3809,N_3308);
nor U7963 (N_7963,N_3844,N_1830);
or U7964 (N_7964,N_1524,N_2965);
nor U7965 (N_7965,N_4153,N_3339);
and U7966 (N_7966,N_2601,N_3062);
and U7967 (N_7967,N_3169,N_3150);
xnor U7968 (N_7968,N_386,N_2786);
and U7969 (N_7969,N_3016,N_565);
nand U7970 (N_7970,N_1653,N_1502);
nor U7971 (N_7971,N_2904,N_3404);
and U7972 (N_7972,N_324,N_1449);
and U7973 (N_7973,N_3419,N_4993);
nor U7974 (N_7974,N_240,N_1769);
and U7975 (N_7975,N_4436,N_530);
and U7976 (N_7976,N_347,N_2388);
xor U7977 (N_7977,N_730,N_2709);
or U7978 (N_7978,N_829,N_415);
and U7979 (N_7979,N_4076,N_3755);
and U7980 (N_7980,N_484,N_4603);
nor U7981 (N_7981,N_2443,N_2454);
xor U7982 (N_7982,N_1415,N_4973);
xor U7983 (N_7983,N_2757,N_4224);
nor U7984 (N_7984,N_4312,N_3373);
nor U7985 (N_7985,N_1886,N_1055);
and U7986 (N_7986,N_3172,N_1397);
or U7987 (N_7987,N_2584,N_2060);
nand U7988 (N_7988,N_946,N_3774);
or U7989 (N_7989,N_4104,N_4899);
nand U7990 (N_7990,N_611,N_3826);
or U7991 (N_7991,N_4961,N_4380);
or U7992 (N_7992,N_2009,N_2392);
nand U7993 (N_7993,N_1532,N_1685);
or U7994 (N_7994,N_4663,N_4725);
nand U7995 (N_7995,N_1484,N_1195);
nand U7996 (N_7996,N_583,N_2014);
and U7997 (N_7997,N_3814,N_1152);
nand U7998 (N_7998,N_4218,N_1718);
nand U7999 (N_7999,N_349,N_4855);
nor U8000 (N_8000,N_2947,N_398);
or U8001 (N_8001,N_2734,N_3603);
xnor U8002 (N_8002,N_4047,N_3965);
xnor U8003 (N_8003,N_1060,N_92);
and U8004 (N_8004,N_4195,N_1389);
nand U8005 (N_8005,N_1092,N_1621);
nand U8006 (N_8006,N_4173,N_331);
or U8007 (N_8007,N_1759,N_2889);
or U8008 (N_8008,N_1249,N_4774);
nand U8009 (N_8009,N_4196,N_4298);
nand U8010 (N_8010,N_3979,N_4650);
nand U8011 (N_8011,N_1517,N_2822);
or U8012 (N_8012,N_886,N_3506);
or U8013 (N_8013,N_2716,N_3763);
nor U8014 (N_8014,N_1132,N_493);
nor U8015 (N_8015,N_1884,N_886);
nand U8016 (N_8016,N_2528,N_323);
and U8017 (N_8017,N_1527,N_3474);
or U8018 (N_8018,N_2162,N_4696);
nand U8019 (N_8019,N_4684,N_75);
or U8020 (N_8020,N_1147,N_1538);
nor U8021 (N_8021,N_282,N_4873);
nand U8022 (N_8022,N_1670,N_2019);
and U8023 (N_8023,N_2957,N_2257);
or U8024 (N_8024,N_235,N_3468);
nor U8025 (N_8025,N_162,N_1663);
and U8026 (N_8026,N_2820,N_22);
nand U8027 (N_8027,N_2882,N_388);
xnor U8028 (N_8028,N_3690,N_3943);
or U8029 (N_8029,N_3751,N_3171);
nand U8030 (N_8030,N_2831,N_4083);
and U8031 (N_8031,N_2218,N_92);
nand U8032 (N_8032,N_4082,N_2491);
nor U8033 (N_8033,N_4781,N_1373);
nand U8034 (N_8034,N_791,N_2403);
nor U8035 (N_8035,N_1618,N_4970);
nand U8036 (N_8036,N_4034,N_3632);
and U8037 (N_8037,N_2295,N_2533);
nand U8038 (N_8038,N_3959,N_1047);
and U8039 (N_8039,N_1585,N_3913);
nor U8040 (N_8040,N_332,N_3993);
and U8041 (N_8041,N_3996,N_3825);
nor U8042 (N_8042,N_3360,N_2446);
nand U8043 (N_8043,N_2487,N_3494);
nor U8044 (N_8044,N_4964,N_4010);
nand U8045 (N_8045,N_664,N_688);
and U8046 (N_8046,N_4230,N_4600);
or U8047 (N_8047,N_1908,N_3661);
or U8048 (N_8048,N_323,N_2573);
nor U8049 (N_8049,N_2102,N_2086);
and U8050 (N_8050,N_3937,N_4194);
or U8051 (N_8051,N_1288,N_4997);
xnor U8052 (N_8052,N_3157,N_4900);
or U8053 (N_8053,N_4387,N_1544);
or U8054 (N_8054,N_3,N_156);
nand U8055 (N_8055,N_1869,N_2156);
and U8056 (N_8056,N_1089,N_292);
nor U8057 (N_8057,N_4312,N_3569);
nor U8058 (N_8058,N_2009,N_3194);
nand U8059 (N_8059,N_4641,N_1416);
or U8060 (N_8060,N_550,N_2963);
nor U8061 (N_8061,N_4702,N_592);
and U8062 (N_8062,N_2411,N_3429);
nand U8063 (N_8063,N_1197,N_3188);
or U8064 (N_8064,N_4677,N_2839);
and U8065 (N_8065,N_1607,N_1981);
and U8066 (N_8066,N_722,N_3591);
nor U8067 (N_8067,N_1405,N_2505);
and U8068 (N_8068,N_4333,N_3587);
nor U8069 (N_8069,N_3004,N_491);
nand U8070 (N_8070,N_1739,N_3811);
nor U8071 (N_8071,N_1942,N_3847);
nor U8072 (N_8072,N_3395,N_4385);
and U8073 (N_8073,N_3966,N_1298);
nor U8074 (N_8074,N_4757,N_125);
nand U8075 (N_8075,N_1418,N_4291);
nor U8076 (N_8076,N_4113,N_4157);
and U8077 (N_8077,N_2295,N_4749);
or U8078 (N_8078,N_3985,N_4091);
nand U8079 (N_8079,N_674,N_2958);
nand U8080 (N_8080,N_4381,N_3440);
and U8081 (N_8081,N_1444,N_3304);
or U8082 (N_8082,N_3422,N_991);
nand U8083 (N_8083,N_2386,N_3484);
or U8084 (N_8084,N_3946,N_270);
nor U8085 (N_8085,N_9,N_4133);
nand U8086 (N_8086,N_1221,N_1900);
nor U8087 (N_8087,N_3435,N_348);
nand U8088 (N_8088,N_3582,N_3497);
nand U8089 (N_8089,N_3495,N_614);
nand U8090 (N_8090,N_4720,N_2378);
nand U8091 (N_8091,N_2633,N_453);
or U8092 (N_8092,N_735,N_1421);
nor U8093 (N_8093,N_4211,N_754);
nand U8094 (N_8094,N_935,N_1192);
nor U8095 (N_8095,N_2840,N_1567);
and U8096 (N_8096,N_3722,N_1219);
nand U8097 (N_8097,N_916,N_3848);
xnor U8098 (N_8098,N_1135,N_1897);
and U8099 (N_8099,N_2174,N_4596);
nor U8100 (N_8100,N_676,N_605);
and U8101 (N_8101,N_562,N_866);
nor U8102 (N_8102,N_2389,N_972);
nand U8103 (N_8103,N_584,N_851);
nand U8104 (N_8104,N_1892,N_1818);
nand U8105 (N_8105,N_150,N_2597);
nor U8106 (N_8106,N_1319,N_836);
or U8107 (N_8107,N_3246,N_13);
and U8108 (N_8108,N_1894,N_3748);
or U8109 (N_8109,N_595,N_721);
nor U8110 (N_8110,N_1864,N_169);
and U8111 (N_8111,N_2856,N_1839);
xor U8112 (N_8112,N_693,N_3838);
or U8113 (N_8113,N_4754,N_1911);
nor U8114 (N_8114,N_4612,N_631);
and U8115 (N_8115,N_4567,N_3656);
or U8116 (N_8116,N_403,N_1091);
nor U8117 (N_8117,N_142,N_3037);
nor U8118 (N_8118,N_1161,N_1303);
nand U8119 (N_8119,N_4492,N_333);
and U8120 (N_8120,N_386,N_4505);
and U8121 (N_8121,N_4906,N_388);
nand U8122 (N_8122,N_4228,N_503);
nand U8123 (N_8123,N_271,N_1990);
and U8124 (N_8124,N_3974,N_2719);
and U8125 (N_8125,N_2647,N_3831);
or U8126 (N_8126,N_1212,N_4386);
nor U8127 (N_8127,N_1277,N_1971);
xor U8128 (N_8128,N_4798,N_4234);
and U8129 (N_8129,N_2585,N_825);
xnor U8130 (N_8130,N_4792,N_2539);
and U8131 (N_8131,N_1512,N_4386);
nor U8132 (N_8132,N_2554,N_3865);
nand U8133 (N_8133,N_2398,N_2638);
xor U8134 (N_8134,N_1402,N_624);
and U8135 (N_8135,N_1299,N_3253);
or U8136 (N_8136,N_3975,N_3595);
nand U8137 (N_8137,N_3172,N_4529);
nand U8138 (N_8138,N_4404,N_1483);
nand U8139 (N_8139,N_3764,N_577);
and U8140 (N_8140,N_1971,N_2688);
or U8141 (N_8141,N_4207,N_480);
xor U8142 (N_8142,N_1897,N_2635);
or U8143 (N_8143,N_1664,N_3228);
nor U8144 (N_8144,N_2320,N_4204);
nor U8145 (N_8145,N_3898,N_352);
nor U8146 (N_8146,N_2466,N_383);
nand U8147 (N_8147,N_4342,N_4205);
or U8148 (N_8148,N_3261,N_1385);
and U8149 (N_8149,N_1929,N_4635);
or U8150 (N_8150,N_2581,N_4908);
and U8151 (N_8151,N_2237,N_4802);
nor U8152 (N_8152,N_3724,N_1788);
nor U8153 (N_8153,N_1671,N_349);
or U8154 (N_8154,N_1250,N_3125);
or U8155 (N_8155,N_743,N_3885);
and U8156 (N_8156,N_1666,N_2201);
nand U8157 (N_8157,N_1573,N_4223);
or U8158 (N_8158,N_4850,N_1944);
or U8159 (N_8159,N_1237,N_901);
and U8160 (N_8160,N_3211,N_3304);
xnor U8161 (N_8161,N_4552,N_2273);
and U8162 (N_8162,N_1409,N_4848);
nand U8163 (N_8163,N_2013,N_3257);
or U8164 (N_8164,N_1807,N_313);
or U8165 (N_8165,N_2922,N_2549);
and U8166 (N_8166,N_2284,N_4248);
or U8167 (N_8167,N_935,N_2285);
or U8168 (N_8168,N_2391,N_1643);
xnor U8169 (N_8169,N_2384,N_1830);
nor U8170 (N_8170,N_2755,N_1618);
and U8171 (N_8171,N_37,N_1627);
and U8172 (N_8172,N_221,N_3422);
nand U8173 (N_8173,N_1460,N_3601);
nor U8174 (N_8174,N_4401,N_666);
and U8175 (N_8175,N_2294,N_2488);
xor U8176 (N_8176,N_4302,N_2807);
or U8177 (N_8177,N_583,N_3889);
or U8178 (N_8178,N_4263,N_3537);
and U8179 (N_8179,N_1044,N_2357);
nor U8180 (N_8180,N_4631,N_3883);
xor U8181 (N_8181,N_2866,N_144);
or U8182 (N_8182,N_2238,N_3580);
or U8183 (N_8183,N_104,N_4912);
nor U8184 (N_8184,N_2297,N_2513);
or U8185 (N_8185,N_4195,N_1339);
and U8186 (N_8186,N_1501,N_680);
nor U8187 (N_8187,N_3192,N_4386);
nand U8188 (N_8188,N_213,N_2094);
nand U8189 (N_8189,N_1826,N_901);
xor U8190 (N_8190,N_657,N_908);
or U8191 (N_8191,N_3334,N_4922);
and U8192 (N_8192,N_1294,N_3693);
nor U8193 (N_8193,N_571,N_1112);
nor U8194 (N_8194,N_495,N_2087);
nand U8195 (N_8195,N_299,N_3876);
nand U8196 (N_8196,N_4007,N_4846);
nor U8197 (N_8197,N_3450,N_3867);
or U8198 (N_8198,N_306,N_3331);
or U8199 (N_8199,N_1587,N_1885);
and U8200 (N_8200,N_4093,N_2996);
or U8201 (N_8201,N_114,N_3730);
or U8202 (N_8202,N_999,N_36);
nor U8203 (N_8203,N_3951,N_1902);
or U8204 (N_8204,N_1575,N_4264);
xor U8205 (N_8205,N_4547,N_3785);
or U8206 (N_8206,N_4863,N_802);
xnor U8207 (N_8207,N_2431,N_4997);
or U8208 (N_8208,N_4284,N_4596);
nand U8209 (N_8209,N_4497,N_1138);
or U8210 (N_8210,N_4726,N_1549);
and U8211 (N_8211,N_1803,N_446);
and U8212 (N_8212,N_4317,N_4601);
nor U8213 (N_8213,N_4049,N_1817);
nand U8214 (N_8214,N_1210,N_3916);
and U8215 (N_8215,N_1319,N_166);
nand U8216 (N_8216,N_1594,N_4732);
or U8217 (N_8217,N_1725,N_1625);
or U8218 (N_8218,N_4871,N_237);
xnor U8219 (N_8219,N_3781,N_1829);
xnor U8220 (N_8220,N_3789,N_1773);
nor U8221 (N_8221,N_3428,N_1044);
nand U8222 (N_8222,N_909,N_1863);
nand U8223 (N_8223,N_3571,N_42);
or U8224 (N_8224,N_1348,N_3818);
or U8225 (N_8225,N_223,N_729);
and U8226 (N_8226,N_1571,N_24);
and U8227 (N_8227,N_107,N_168);
xnor U8228 (N_8228,N_2028,N_2385);
nand U8229 (N_8229,N_1557,N_1931);
and U8230 (N_8230,N_2053,N_3448);
and U8231 (N_8231,N_776,N_1529);
or U8232 (N_8232,N_1482,N_4023);
nor U8233 (N_8233,N_2515,N_2623);
nand U8234 (N_8234,N_580,N_466);
and U8235 (N_8235,N_2581,N_1906);
or U8236 (N_8236,N_2289,N_206);
or U8237 (N_8237,N_3445,N_332);
and U8238 (N_8238,N_4420,N_1675);
and U8239 (N_8239,N_2682,N_2685);
nand U8240 (N_8240,N_3878,N_3770);
or U8241 (N_8241,N_656,N_2287);
xnor U8242 (N_8242,N_4084,N_1870);
and U8243 (N_8243,N_4114,N_378);
xor U8244 (N_8244,N_4655,N_1528);
xnor U8245 (N_8245,N_4003,N_2976);
and U8246 (N_8246,N_2943,N_4620);
nand U8247 (N_8247,N_2209,N_698);
xor U8248 (N_8248,N_4173,N_2987);
xor U8249 (N_8249,N_2883,N_275);
nand U8250 (N_8250,N_1245,N_4673);
nor U8251 (N_8251,N_3782,N_1256);
nor U8252 (N_8252,N_3906,N_1339);
or U8253 (N_8253,N_760,N_1027);
nand U8254 (N_8254,N_1632,N_945);
nor U8255 (N_8255,N_576,N_4844);
and U8256 (N_8256,N_4692,N_2240);
and U8257 (N_8257,N_1895,N_4749);
nor U8258 (N_8258,N_3169,N_4742);
nand U8259 (N_8259,N_3866,N_4052);
and U8260 (N_8260,N_4181,N_2500);
or U8261 (N_8261,N_4996,N_867);
nand U8262 (N_8262,N_3119,N_1541);
or U8263 (N_8263,N_336,N_3942);
and U8264 (N_8264,N_4923,N_3795);
nand U8265 (N_8265,N_3851,N_1120);
nor U8266 (N_8266,N_1440,N_3916);
xnor U8267 (N_8267,N_264,N_1564);
or U8268 (N_8268,N_3251,N_3655);
nand U8269 (N_8269,N_3334,N_4503);
nand U8270 (N_8270,N_4378,N_2207);
or U8271 (N_8271,N_3126,N_3570);
nand U8272 (N_8272,N_3796,N_4265);
and U8273 (N_8273,N_2374,N_28);
xor U8274 (N_8274,N_3268,N_3302);
or U8275 (N_8275,N_3932,N_1999);
nand U8276 (N_8276,N_3403,N_3197);
or U8277 (N_8277,N_4428,N_3941);
or U8278 (N_8278,N_625,N_264);
or U8279 (N_8279,N_156,N_3706);
nor U8280 (N_8280,N_2033,N_642);
or U8281 (N_8281,N_3723,N_4881);
nand U8282 (N_8282,N_3955,N_1187);
xnor U8283 (N_8283,N_699,N_479);
and U8284 (N_8284,N_3588,N_991);
or U8285 (N_8285,N_3098,N_2658);
or U8286 (N_8286,N_308,N_3429);
or U8287 (N_8287,N_4283,N_4492);
or U8288 (N_8288,N_775,N_2492);
nand U8289 (N_8289,N_4184,N_1498);
nor U8290 (N_8290,N_1252,N_798);
nor U8291 (N_8291,N_4906,N_1751);
nand U8292 (N_8292,N_394,N_3674);
and U8293 (N_8293,N_1595,N_133);
nand U8294 (N_8294,N_2523,N_3875);
or U8295 (N_8295,N_4453,N_1076);
and U8296 (N_8296,N_244,N_3243);
nor U8297 (N_8297,N_2691,N_1923);
and U8298 (N_8298,N_3786,N_2726);
or U8299 (N_8299,N_391,N_1232);
nor U8300 (N_8300,N_4673,N_687);
nor U8301 (N_8301,N_1427,N_4444);
nor U8302 (N_8302,N_3200,N_44);
and U8303 (N_8303,N_3867,N_3827);
or U8304 (N_8304,N_1837,N_1247);
nand U8305 (N_8305,N_3719,N_4437);
or U8306 (N_8306,N_2296,N_668);
and U8307 (N_8307,N_2834,N_606);
or U8308 (N_8308,N_3331,N_1050);
and U8309 (N_8309,N_1062,N_1021);
nor U8310 (N_8310,N_3504,N_154);
or U8311 (N_8311,N_4629,N_3509);
nor U8312 (N_8312,N_4121,N_1394);
nor U8313 (N_8313,N_3295,N_753);
or U8314 (N_8314,N_3204,N_2273);
or U8315 (N_8315,N_1392,N_615);
nand U8316 (N_8316,N_4202,N_4201);
and U8317 (N_8317,N_3300,N_4760);
or U8318 (N_8318,N_1430,N_1876);
or U8319 (N_8319,N_4525,N_1376);
nand U8320 (N_8320,N_4725,N_4439);
nor U8321 (N_8321,N_3105,N_1657);
nor U8322 (N_8322,N_4185,N_3);
and U8323 (N_8323,N_2904,N_3088);
or U8324 (N_8324,N_724,N_556);
or U8325 (N_8325,N_3781,N_58);
nor U8326 (N_8326,N_1839,N_118);
and U8327 (N_8327,N_4864,N_3109);
nand U8328 (N_8328,N_3523,N_2056);
nor U8329 (N_8329,N_2777,N_2872);
nand U8330 (N_8330,N_3989,N_3418);
nor U8331 (N_8331,N_2718,N_4587);
nor U8332 (N_8332,N_4491,N_286);
xnor U8333 (N_8333,N_2852,N_4660);
or U8334 (N_8334,N_1721,N_520);
nand U8335 (N_8335,N_4687,N_3729);
and U8336 (N_8336,N_3065,N_1208);
and U8337 (N_8337,N_2528,N_2362);
or U8338 (N_8338,N_118,N_2459);
and U8339 (N_8339,N_2764,N_1062);
and U8340 (N_8340,N_1123,N_2835);
nand U8341 (N_8341,N_686,N_3927);
nor U8342 (N_8342,N_3537,N_34);
and U8343 (N_8343,N_2273,N_1703);
or U8344 (N_8344,N_4418,N_1539);
nor U8345 (N_8345,N_554,N_408);
or U8346 (N_8346,N_3767,N_833);
nor U8347 (N_8347,N_1769,N_843);
nand U8348 (N_8348,N_2426,N_1654);
and U8349 (N_8349,N_2235,N_306);
and U8350 (N_8350,N_3741,N_4039);
nand U8351 (N_8351,N_4862,N_4637);
and U8352 (N_8352,N_2719,N_2125);
xor U8353 (N_8353,N_1562,N_433);
nand U8354 (N_8354,N_2763,N_4560);
and U8355 (N_8355,N_3207,N_4844);
or U8356 (N_8356,N_928,N_3933);
nor U8357 (N_8357,N_3160,N_1206);
and U8358 (N_8358,N_1720,N_4421);
xnor U8359 (N_8359,N_3271,N_1337);
nor U8360 (N_8360,N_2532,N_2271);
and U8361 (N_8361,N_2061,N_2716);
nand U8362 (N_8362,N_1731,N_4982);
nand U8363 (N_8363,N_317,N_3056);
nand U8364 (N_8364,N_4537,N_2606);
nand U8365 (N_8365,N_94,N_4998);
xor U8366 (N_8366,N_4431,N_500);
and U8367 (N_8367,N_475,N_165);
and U8368 (N_8368,N_2760,N_2607);
and U8369 (N_8369,N_1450,N_2275);
nand U8370 (N_8370,N_2440,N_3294);
nor U8371 (N_8371,N_3024,N_2860);
or U8372 (N_8372,N_4451,N_2709);
or U8373 (N_8373,N_63,N_2345);
nand U8374 (N_8374,N_3386,N_1921);
xor U8375 (N_8375,N_2339,N_1913);
and U8376 (N_8376,N_4723,N_4951);
nand U8377 (N_8377,N_1006,N_1477);
nand U8378 (N_8378,N_2994,N_1313);
nand U8379 (N_8379,N_604,N_144);
or U8380 (N_8380,N_4235,N_2639);
xor U8381 (N_8381,N_4023,N_3570);
or U8382 (N_8382,N_1547,N_1351);
nand U8383 (N_8383,N_168,N_4905);
and U8384 (N_8384,N_3684,N_1555);
nand U8385 (N_8385,N_2721,N_1526);
nand U8386 (N_8386,N_4110,N_3288);
nor U8387 (N_8387,N_1915,N_4166);
nor U8388 (N_8388,N_1955,N_1538);
or U8389 (N_8389,N_1837,N_3280);
and U8390 (N_8390,N_471,N_4436);
nand U8391 (N_8391,N_2579,N_946);
nand U8392 (N_8392,N_1656,N_1278);
or U8393 (N_8393,N_2164,N_2658);
nand U8394 (N_8394,N_4581,N_176);
or U8395 (N_8395,N_1610,N_1314);
or U8396 (N_8396,N_2487,N_2769);
nand U8397 (N_8397,N_4824,N_464);
and U8398 (N_8398,N_4129,N_3925);
nor U8399 (N_8399,N_1992,N_1166);
xor U8400 (N_8400,N_1461,N_359);
nor U8401 (N_8401,N_4012,N_2811);
and U8402 (N_8402,N_4804,N_3023);
xor U8403 (N_8403,N_1089,N_1162);
or U8404 (N_8404,N_2866,N_2685);
nand U8405 (N_8405,N_1190,N_326);
and U8406 (N_8406,N_939,N_2106);
xor U8407 (N_8407,N_4818,N_1462);
nor U8408 (N_8408,N_2278,N_3404);
nor U8409 (N_8409,N_4489,N_2000);
or U8410 (N_8410,N_4361,N_922);
xor U8411 (N_8411,N_2469,N_3518);
or U8412 (N_8412,N_1939,N_2529);
nand U8413 (N_8413,N_1855,N_152);
and U8414 (N_8414,N_539,N_1552);
or U8415 (N_8415,N_3596,N_1530);
nor U8416 (N_8416,N_3363,N_335);
nand U8417 (N_8417,N_1761,N_3710);
and U8418 (N_8418,N_1888,N_549);
nand U8419 (N_8419,N_2919,N_462);
nand U8420 (N_8420,N_372,N_2151);
and U8421 (N_8421,N_4600,N_1309);
xnor U8422 (N_8422,N_2994,N_1675);
xnor U8423 (N_8423,N_2623,N_2819);
xnor U8424 (N_8424,N_4080,N_1614);
or U8425 (N_8425,N_1008,N_3583);
xor U8426 (N_8426,N_1326,N_3234);
nor U8427 (N_8427,N_2932,N_2275);
and U8428 (N_8428,N_3042,N_2816);
nand U8429 (N_8429,N_2018,N_1282);
and U8430 (N_8430,N_398,N_2874);
nor U8431 (N_8431,N_2952,N_4778);
and U8432 (N_8432,N_1746,N_2470);
or U8433 (N_8433,N_3918,N_3133);
nor U8434 (N_8434,N_4504,N_4532);
nand U8435 (N_8435,N_3018,N_268);
and U8436 (N_8436,N_2505,N_833);
and U8437 (N_8437,N_4840,N_942);
and U8438 (N_8438,N_1671,N_2708);
nand U8439 (N_8439,N_390,N_2848);
or U8440 (N_8440,N_4641,N_3429);
or U8441 (N_8441,N_4878,N_2023);
nand U8442 (N_8442,N_670,N_1559);
nor U8443 (N_8443,N_544,N_4142);
nand U8444 (N_8444,N_4966,N_2645);
xor U8445 (N_8445,N_641,N_3655);
nand U8446 (N_8446,N_3413,N_4785);
and U8447 (N_8447,N_1560,N_2975);
or U8448 (N_8448,N_4790,N_3410);
or U8449 (N_8449,N_658,N_1224);
nor U8450 (N_8450,N_2330,N_3024);
or U8451 (N_8451,N_3009,N_4484);
nand U8452 (N_8452,N_3248,N_4648);
and U8453 (N_8453,N_739,N_4645);
xor U8454 (N_8454,N_14,N_3518);
nor U8455 (N_8455,N_4024,N_4310);
nand U8456 (N_8456,N_448,N_534);
or U8457 (N_8457,N_887,N_2050);
xnor U8458 (N_8458,N_799,N_2424);
nor U8459 (N_8459,N_4746,N_4988);
nand U8460 (N_8460,N_1651,N_1240);
or U8461 (N_8461,N_2337,N_1130);
or U8462 (N_8462,N_3349,N_3140);
or U8463 (N_8463,N_4165,N_3703);
nor U8464 (N_8464,N_2234,N_2537);
nand U8465 (N_8465,N_2006,N_1589);
xnor U8466 (N_8466,N_4478,N_4974);
and U8467 (N_8467,N_494,N_3965);
nand U8468 (N_8468,N_4171,N_3096);
xor U8469 (N_8469,N_4442,N_4768);
and U8470 (N_8470,N_2253,N_4962);
nor U8471 (N_8471,N_4606,N_4915);
and U8472 (N_8472,N_3157,N_203);
and U8473 (N_8473,N_2660,N_4820);
or U8474 (N_8474,N_2796,N_2379);
nand U8475 (N_8475,N_3205,N_35);
and U8476 (N_8476,N_1857,N_852);
nor U8477 (N_8477,N_4933,N_2425);
nand U8478 (N_8478,N_1778,N_1734);
nand U8479 (N_8479,N_1491,N_2598);
or U8480 (N_8480,N_3450,N_2514);
nand U8481 (N_8481,N_4640,N_1506);
or U8482 (N_8482,N_4420,N_4133);
or U8483 (N_8483,N_4857,N_2295);
and U8484 (N_8484,N_4923,N_2375);
and U8485 (N_8485,N_852,N_2739);
and U8486 (N_8486,N_4602,N_3549);
nor U8487 (N_8487,N_1153,N_2611);
nand U8488 (N_8488,N_4327,N_2021);
xor U8489 (N_8489,N_2965,N_4769);
nor U8490 (N_8490,N_1423,N_3512);
nand U8491 (N_8491,N_3587,N_1844);
nor U8492 (N_8492,N_748,N_1468);
nor U8493 (N_8493,N_3677,N_3950);
nor U8494 (N_8494,N_2317,N_4371);
nor U8495 (N_8495,N_3978,N_2967);
or U8496 (N_8496,N_3249,N_2853);
nand U8497 (N_8497,N_569,N_2080);
nand U8498 (N_8498,N_3703,N_2092);
nand U8499 (N_8499,N_2094,N_281);
and U8500 (N_8500,N_4990,N_3874);
xnor U8501 (N_8501,N_3497,N_1649);
nor U8502 (N_8502,N_3369,N_1711);
and U8503 (N_8503,N_103,N_2468);
and U8504 (N_8504,N_3913,N_4531);
nand U8505 (N_8505,N_4412,N_2069);
nand U8506 (N_8506,N_1631,N_4916);
and U8507 (N_8507,N_3986,N_4547);
nor U8508 (N_8508,N_1663,N_772);
nand U8509 (N_8509,N_4190,N_4482);
xnor U8510 (N_8510,N_4599,N_4642);
and U8511 (N_8511,N_2550,N_3986);
or U8512 (N_8512,N_891,N_2123);
nand U8513 (N_8513,N_1125,N_1572);
nand U8514 (N_8514,N_1442,N_3186);
or U8515 (N_8515,N_3042,N_1638);
or U8516 (N_8516,N_4799,N_1298);
nand U8517 (N_8517,N_62,N_3287);
or U8518 (N_8518,N_2710,N_1514);
nand U8519 (N_8519,N_2867,N_1550);
nand U8520 (N_8520,N_4912,N_124);
or U8521 (N_8521,N_4973,N_848);
and U8522 (N_8522,N_92,N_4322);
and U8523 (N_8523,N_3722,N_1501);
and U8524 (N_8524,N_4994,N_2131);
nand U8525 (N_8525,N_4852,N_1258);
and U8526 (N_8526,N_2120,N_4381);
and U8527 (N_8527,N_4614,N_4269);
nor U8528 (N_8528,N_3136,N_1842);
and U8529 (N_8529,N_1045,N_530);
and U8530 (N_8530,N_10,N_1135);
and U8531 (N_8531,N_1057,N_751);
or U8532 (N_8532,N_2988,N_3080);
and U8533 (N_8533,N_2109,N_2068);
xor U8534 (N_8534,N_997,N_3793);
or U8535 (N_8535,N_1933,N_2653);
nor U8536 (N_8536,N_2281,N_2323);
and U8537 (N_8537,N_3960,N_3361);
or U8538 (N_8538,N_1055,N_3288);
and U8539 (N_8539,N_4007,N_3927);
nor U8540 (N_8540,N_423,N_2917);
xor U8541 (N_8541,N_3956,N_3750);
and U8542 (N_8542,N_1418,N_4104);
and U8543 (N_8543,N_3636,N_2770);
nor U8544 (N_8544,N_642,N_655);
or U8545 (N_8545,N_2227,N_719);
nor U8546 (N_8546,N_4456,N_2354);
or U8547 (N_8547,N_861,N_2659);
nor U8548 (N_8548,N_1672,N_1668);
and U8549 (N_8549,N_3254,N_1150);
nor U8550 (N_8550,N_613,N_644);
nor U8551 (N_8551,N_4538,N_1996);
nor U8552 (N_8552,N_3493,N_3983);
nand U8553 (N_8553,N_4392,N_2375);
or U8554 (N_8554,N_873,N_2769);
nand U8555 (N_8555,N_4609,N_1471);
and U8556 (N_8556,N_4529,N_2959);
and U8557 (N_8557,N_2676,N_4721);
and U8558 (N_8558,N_1615,N_548);
and U8559 (N_8559,N_4950,N_1531);
xor U8560 (N_8560,N_853,N_629);
and U8561 (N_8561,N_2430,N_3219);
or U8562 (N_8562,N_4362,N_4484);
and U8563 (N_8563,N_2336,N_142);
and U8564 (N_8564,N_3957,N_2739);
nand U8565 (N_8565,N_3973,N_2401);
nor U8566 (N_8566,N_3770,N_394);
or U8567 (N_8567,N_1719,N_3291);
nand U8568 (N_8568,N_4115,N_3147);
nor U8569 (N_8569,N_3389,N_87);
nor U8570 (N_8570,N_4388,N_1911);
or U8571 (N_8571,N_229,N_3481);
and U8572 (N_8572,N_1269,N_3026);
and U8573 (N_8573,N_1563,N_526);
and U8574 (N_8574,N_712,N_2801);
and U8575 (N_8575,N_3974,N_2818);
and U8576 (N_8576,N_1059,N_3637);
nand U8577 (N_8577,N_1221,N_2053);
nor U8578 (N_8578,N_4179,N_2982);
or U8579 (N_8579,N_2197,N_1596);
and U8580 (N_8580,N_4357,N_3672);
nand U8581 (N_8581,N_3124,N_2856);
and U8582 (N_8582,N_185,N_3750);
and U8583 (N_8583,N_4053,N_3450);
xor U8584 (N_8584,N_2100,N_4035);
xor U8585 (N_8585,N_4421,N_4219);
or U8586 (N_8586,N_2947,N_2460);
or U8587 (N_8587,N_4953,N_4555);
xnor U8588 (N_8588,N_3566,N_534);
and U8589 (N_8589,N_4386,N_3273);
and U8590 (N_8590,N_3837,N_357);
and U8591 (N_8591,N_433,N_2108);
nor U8592 (N_8592,N_303,N_1972);
or U8593 (N_8593,N_3357,N_3806);
xnor U8594 (N_8594,N_4296,N_4203);
nand U8595 (N_8595,N_3262,N_4814);
nand U8596 (N_8596,N_4013,N_3608);
nand U8597 (N_8597,N_2479,N_1687);
and U8598 (N_8598,N_2669,N_1794);
and U8599 (N_8599,N_2721,N_3041);
nor U8600 (N_8600,N_2606,N_4145);
and U8601 (N_8601,N_3604,N_789);
and U8602 (N_8602,N_2233,N_2755);
xor U8603 (N_8603,N_2786,N_1763);
nor U8604 (N_8604,N_1961,N_4865);
and U8605 (N_8605,N_295,N_1932);
xnor U8606 (N_8606,N_4904,N_4760);
nand U8607 (N_8607,N_1103,N_1562);
nand U8608 (N_8608,N_4521,N_3216);
and U8609 (N_8609,N_2010,N_3057);
or U8610 (N_8610,N_4569,N_426);
nand U8611 (N_8611,N_3617,N_368);
nand U8612 (N_8612,N_4380,N_558);
xor U8613 (N_8613,N_626,N_4751);
or U8614 (N_8614,N_4462,N_2580);
and U8615 (N_8615,N_2907,N_3882);
nand U8616 (N_8616,N_456,N_4828);
or U8617 (N_8617,N_2406,N_2980);
nand U8618 (N_8618,N_1852,N_1255);
and U8619 (N_8619,N_1208,N_2148);
or U8620 (N_8620,N_4253,N_3659);
nor U8621 (N_8621,N_3825,N_1385);
nand U8622 (N_8622,N_139,N_4880);
nor U8623 (N_8623,N_4995,N_4354);
and U8624 (N_8624,N_2164,N_1236);
or U8625 (N_8625,N_3043,N_1995);
nand U8626 (N_8626,N_2824,N_3636);
nand U8627 (N_8627,N_2450,N_142);
nand U8628 (N_8628,N_2241,N_1587);
nor U8629 (N_8629,N_2341,N_4908);
xor U8630 (N_8630,N_2673,N_635);
nor U8631 (N_8631,N_4532,N_487);
or U8632 (N_8632,N_1390,N_4357);
or U8633 (N_8633,N_3652,N_3195);
or U8634 (N_8634,N_4291,N_2575);
or U8635 (N_8635,N_407,N_175);
or U8636 (N_8636,N_1955,N_551);
nand U8637 (N_8637,N_2502,N_3835);
or U8638 (N_8638,N_4943,N_1850);
nor U8639 (N_8639,N_135,N_1061);
and U8640 (N_8640,N_519,N_4497);
and U8641 (N_8641,N_3683,N_3304);
and U8642 (N_8642,N_3660,N_2445);
nand U8643 (N_8643,N_2733,N_3030);
nand U8644 (N_8644,N_3143,N_4352);
or U8645 (N_8645,N_4042,N_3584);
or U8646 (N_8646,N_4340,N_3196);
nand U8647 (N_8647,N_4064,N_383);
xor U8648 (N_8648,N_3453,N_3518);
nand U8649 (N_8649,N_2754,N_4180);
nor U8650 (N_8650,N_2045,N_3357);
xor U8651 (N_8651,N_1400,N_4990);
nor U8652 (N_8652,N_2118,N_2244);
nor U8653 (N_8653,N_4756,N_1579);
and U8654 (N_8654,N_113,N_2279);
and U8655 (N_8655,N_3039,N_690);
nor U8656 (N_8656,N_4649,N_4567);
or U8657 (N_8657,N_1449,N_2196);
or U8658 (N_8658,N_2170,N_2339);
and U8659 (N_8659,N_812,N_1280);
or U8660 (N_8660,N_3141,N_2200);
xnor U8661 (N_8661,N_2589,N_2812);
and U8662 (N_8662,N_4013,N_3176);
or U8663 (N_8663,N_3028,N_4403);
and U8664 (N_8664,N_592,N_4797);
and U8665 (N_8665,N_1400,N_3594);
xor U8666 (N_8666,N_3231,N_1218);
nand U8667 (N_8667,N_1960,N_3529);
nor U8668 (N_8668,N_2037,N_4719);
nor U8669 (N_8669,N_3978,N_2207);
nor U8670 (N_8670,N_835,N_1131);
and U8671 (N_8671,N_780,N_4386);
and U8672 (N_8672,N_4806,N_2616);
nor U8673 (N_8673,N_23,N_1222);
or U8674 (N_8674,N_767,N_2350);
or U8675 (N_8675,N_436,N_1078);
nor U8676 (N_8676,N_1530,N_3399);
nand U8677 (N_8677,N_2472,N_3099);
or U8678 (N_8678,N_4022,N_1660);
and U8679 (N_8679,N_3237,N_1270);
or U8680 (N_8680,N_3019,N_1945);
nand U8681 (N_8681,N_4035,N_1491);
or U8682 (N_8682,N_3396,N_4123);
and U8683 (N_8683,N_2525,N_628);
and U8684 (N_8684,N_407,N_3132);
and U8685 (N_8685,N_3037,N_1897);
nand U8686 (N_8686,N_2080,N_741);
and U8687 (N_8687,N_1329,N_3574);
nor U8688 (N_8688,N_4812,N_3315);
nor U8689 (N_8689,N_4297,N_4712);
nor U8690 (N_8690,N_1214,N_4314);
and U8691 (N_8691,N_1476,N_2392);
and U8692 (N_8692,N_1075,N_962);
nor U8693 (N_8693,N_3607,N_4094);
and U8694 (N_8694,N_2204,N_3434);
and U8695 (N_8695,N_3827,N_2931);
xor U8696 (N_8696,N_1407,N_3987);
nand U8697 (N_8697,N_1481,N_2057);
xnor U8698 (N_8698,N_1776,N_3122);
and U8699 (N_8699,N_2493,N_3359);
and U8700 (N_8700,N_1677,N_1654);
nand U8701 (N_8701,N_438,N_346);
and U8702 (N_8702,N_1903,N_3633);
or U8703 (N_8703,N_3932,N_2208);
nand U8704 (N_8704,N_3597,N_4122);
and U8705 (N_8705,N_4136,N_2110);
or U8706 (N_8706,N_3869,N_2338);
nor U8707 (N_8707,N_715,N_4505);
nand U8708 (N_8708,N_2983,N_3729);
nor U8709 (N_8709,N_2576,N_1650);
and U8710 (N_8710,N_329,N_3941);
or U8711 (N_8711,N_4597,N_3006);
and U8712 (N_8712,N_2720,N_750);
and U8713 (N_8713,N_4195,N_1840);
or U8714 (N_8714,N_3738,N_3392);
or U8715 (N_8715,N_3857,N_423);
or U8716 (N_8716,N_4104,N_4807);
and U8717 (N_8717,N_3170,N_4580);
and U8718 (N_8718,N_1150,N_1929);
nor U8719 (N_8719,N_4223,N_3869);
or U8720 (N_8720,N_3348,N_67);
xnor U8721 (N_8721,N_143,N_1120);
nor U8722 (N_8722,N_2068,N_3353);
and U8723 (N_8723,N_2820,N_1825);
or U8724 (N_8724,N_1775,N_1064);
nand U8725 (N_8725,N_1438,N_1923);
or U8726 (N_8726,N_4697,N_2063);
nand U8727 (N_8727,N_1454,N_2947);
nand U8728 (N_8728,N_2822,N_2536);
xnor U8729 (N_8729,N_754,N_1180);
nand U8730 (N_8730,N_1407,N_1985);
nand U8731 (N_8731,N_54,N_51);
and U8732 (N_8732,N_1206,N_3729);
or U8733 (N_8733,N_3621,N_1388);
nor U8734 (N_8734,N_4290,N_1790);
or U8735 (N_8735,N_532,N_4916);
or U8736 (N_8736,N_249,N_4749);
xor U8737 (N_8737,N_3343,N_2733);
and U8738 (N_8738,N_2740,N_4453);
nand U8739 (N_8739,N_508,N_3162);
nor U8740 (N_8740,N_2955,N_503);
and U8741 (N_8741,N_2835,N_3232);
nand U8742 (N_8742,N_1289,N_3790);
xor U8743 (N_8743,N_4719,N_553);
or U8744 (N_8744,N_358,N_1820);
and U8745 (N_8745,N_2444,N_3619);
xnor U8746 (N_8746,N_3586,N_1137);
or U8747 (N_8747,N_3214,N_112);
or U8748 (N_8748,N_4699,N_3053);
nor U8749 (N_8749,N_1630,N_1632);
or U8750 (N_8750,N_632,N_564);
and U8751 (N_8751,N_297,N_4196);
nor U8752 (N_8752,N_4704,N_2966);
and U8753 (N_8753,N_2446,N_2950);
and U8754 (N_8754,N_3872,N_1963);
and U8755 (N_8755,N_2023,N_4700);
nor U8756 (N_8756,N_4744,N_4360);
or U8757 (N_8757,N_3476,N_378);
nand U8758 (N_8758,N_3306,N_4476);
nor U8759 (N_8759,N_2101,N_314);
nand U8760 (N_8760,N_2795,N_3989);
nand U8761 (N_8761,N_4133,N_2257);
and U8762 (N_8762,N_860,N_2914);
nor U8763 (N_8763,N_1116,N_581);
or U8764 (N_8764,N_2019,N_698);
xor U8765 (N_8765,N_757,N_177);
nand U8766 (N_8766,N_2163,N_3434);
nand U8767 (N_8767,N_1596,N_390);
nor U8768 (N_8768,N_3955,N_4671);
and U8769 (N_8769,N_2721,N_951);
or U8770 (N_8770,N_3345,N_1270);
or U8771 (N_8771,N_289,N_3795);
nand U8772 (N_8772,N_1123,N_3733);
or U8773 (N_8773,N_590,N_4904);
nand U8774 (N_8774,N_3034,N_1152);
nand U8775 (N_8775,N_2485,N_1921);
nand U8776 (N_8776,N_3095,N_1868);
xnor U8777 (N_8777,N_4661,N_3356);
or U8778 (N_8778,N_2077,N_250);
nand U8779 (N_8779,N_1157,N_1024);
or U8780 (N_8780,N_3128,N_361);
or U8781 (N_8781,N_2380,N_2911);
and U8782 (N_8782,N_2567,N_1519);
nor U8783 (N_8783,N_1378,N_2907);
and U8784 (N_8784,N_3053,N_1087);
xnor U8785 (N_8785,N_1407,N_2325);
or U8786 (N_8786,N_2840,N_914);
nor U8787 (N_8787,N_2040,N_3685);
and U8788 (N_8788,N_963,N_3750);
and U8789 (N_8789,N_942,N_3077);
nor U8790 (N_8790,N_2297,N_4116);
and U8791 (N_8791,N_516,N_4732);
nand U8792 (N_8792,N_239,N_4129);
nand U8793 (N_8793,N_2898,N_665);
or U8794 (N_8794,N_3990,N_511);
nand U8795 (N_8795,N_3825,N_1222);
and U8796 (N_8796,N_1888,N_494);
nor U8797 (N_8797,N_1338,N_2617);
nor U8798 (N_8798,N_4993,N_4664);
xor U8799 (N_8799,N_799,N_93);
xor U8800 (N_8800,N_1009,N_1339);
nand U8801 (N_8801,N_2272,N_597);
and U8802 (N_8802,N_1081,N_3242);
xnor U8803 (N_8803,N_624,N_2976);
nand U8804 (N_8804,N_116,N_2439);
xnor U8805 (N_8805,N_493,N_2618);
nand U8806 (N_8806,N_4107,N_4801);
nand U8807 (N_8807,N_1619,N_4712);
nor U8808 (N_8808,N_1188,N_1987);
nor U8809 (N_8809,N_2496,N_4260);
and U8810 (N_8810,N_1646,N_1396);
nand U8811 (N_8811,N_3946,N_688);
nor U8812 (N_8812,N_4382,N_2750);
or U8813 (N_8813,N_2230,N_3672);
nor U8814 (N_8814,N_3294,N_1500);
nand U8815 (N_8815,N_4969,N_1787);
nand U8816 (N_8816,N_313,N_4774);
or U8817 (N_8817,N_4306,N_626);
and U8818 (N_8818,N_3897,N_841);
xnor U8819 (N_8819,N_2168,N_560);
or U8820 (N_8820,N_1824,N_2171);
and U8821 (N_8821,N_24,N_1931);
or U8822 (N_8822,N_4274,N_3124);
nand U8823 (N_8823,N_1690,N_356);
or U8824 (N_8824,N_1645,N_3928);
nor U8825 (N_8825,N_768,N_860);
nand U8826 (N_8826,N_2279,N_452);
or U8827 (N_8827,N_3803,N_66);
and U8828 (N_8828,N_583,N_2187);
or U8829 (N_8829,N_1348,N_2384);
or U8830 (N_8830,N_2987,N_1743);
nor U8831 (N_8831,N_4370,N_921);
and U8832 (N_8832,N_4964,N_2088);
and U8833 (N_8833,N_1291,N_3167);
and U8834 (N_8834,N_1672,N_1975);
or U8835 (N_8835,N_4569,N_1108);
and U8836 (N_8836,N_2230,N_3495);
nor U8837 (N_8837,N_4974,N_3331);
or U8838 (N_8838,N_3653,N_1732);
nand U8839 (N_8839,N_3966,N_3626);
and U8840 (N_8840,N_3471,N_1133);
nand U8841 (N_8841,N_3499,N_1351);
nor U8842 (N_8842,N_828,N_4269);
nor U8843 (N_8843,N_3717,N_2034);
nor U8844 (N_8844,N_4020,N_2218);
nor U8845 (N_8845,N_4651,N_4850);
nand U8846 (N_8846,N_4884,N_4303);
nor U8847 (N_8847,N_2953,N_1161);
nand U8848 (N_8848,N_1545,N_3831);
xor U8849 (N_8849,N_721,N_720);
nand U8850 (N_8850,N_2845,N_2874);
nor U8851 (N_8851,N_4375,N_1908);
nor U8852 (N_8852,N_2458,N_2638);
and U8853 (N_8853,N_4386,N_2843);
nand U8854 (N_8854,N_4699,N_733);
nand U8855 (N_8855,N_3712,N_4370);
or U8856 (N_8856,N_4144,N_3200);
or U8857 (N_8857,N_3945,N_385);
and U8858 (N_8858,N_2221,N_4337);
nand U8859 (N_8859,N_2488,N_3731);
nor U8860 (N_8860,N_126,N_146);
nand U8861 (N_8861,N_778,N_2190);
nor U8862 (N_8862,N_4903,N_1508);
nor U8863 (N_8863,N_4909,N_4212);
and U8864 (N_8864,N_976,N_2008);
and U8865 (N_8865,N_4687,N_159);
or U8866 (N_8866,N_3385,N_130);
or U8867 (N_8867,N_1833,N_1254);
nor U8868 (N_8868,N_2386,N_1586);
or U8869 (N_8869,N_1385,N_2314);
and U8870 (N_8870,N_4341,N_2087);
nor U8871 (N_8871,N_2052,N_2494);
nor U8872 (N_8872,N_4035,N_1788);
nor U8873 (N_8873,N_4837,N_3330);
nand U8874 (N_8874,N_2697,N_2744);
nor U8875 (N_8875,N_4617,N_4047);
and U8876 (N_8876,N_457,N_2884);
xor U8877 (N_8877,N_1517,N_3877);
and U8878 (N_8878,N_3277,N_3595);
and U8879 (N_8879,N_1920,N_650);
nor U8880 (N_8880,N_4167,N_3886);
nand U8881 (N_8881,N_4359,N_3855);
and U8882 (N_8882,N_2012,N_2329);
or U8883 (N_8883,N_703,N_4437);
nor U8884 (N_8884,N_4764,N_4947);
nor U8885 (N_8885,N_4169,N_332);
nand U8886 (N_8886,N_3317,N_3574);
and U8887 (N_8887,N_2568,N_6);
nand U8888 (N_8888,N_1714,N_297);
or U8889 (N_8889,N_2770,N_4887);
or U8890 (N_8890,N_2531,N_1316);
xor U8891 (N_8891,N_1926,N_1356);
nand U8892 (N_8892,N_3552,N_4083);
and U8893 (N_8893,N_3413,N_1226);
nor U8894 (N_8894,N_2717,N_23);
or U8895 (N_8895,N_239,N_4054);
xnor U8896 (N_8896,N_4755,N_3998);
or U8897 (N_8897,N_4543,N_22);
nor U8898 (N_8898,N_1035,N_460);
nand U8899 (N_8899,N_3657,N_1324);
and U8900 (N_8900,N_4604,N_306);
nor U8901 (N_8901,N_787,N_4270);
nor U8902 (N_8902,N_34,N_2157);
and U8903 (N_8903,N_4574,N_2696);
nor U8904 (N_8904,N_183,N_3016);
xnor U8905 (N_8905,N_3228,N_2668);
nor U8906 (N_8906,N_3615,N_1211);
nand U8907 (N_8907,N_502,N_1418);
or U8908 (N_8908,N_91,N_14);
or U8909 (N_8909,N_3154,N_3848);
nand U8910 (N_8910,N_1928,N_2620);
nand U8911 (N_8911,N_4025,N_1497);
or U8912 (N_8912,N_4145,N_3035);
xor U8913 (N_8913,N_1586,N_4957);
and U8914 (N_8914,N_2803,N_52);
nand U8915 (N_8915,N_541,N_2818);
nand U8916 (N_8916,N_3281,N_4113);
xnor U8917 (N_8917,N_844,N_217);
nand U8918 (N_8918,N_337,N_4093);
nand U8919 (N_8919,N_2773,N_4917);
or U8920 (N_8920,N_3617,N_2122);
nor U8921 (N_8921,N_1372,N_45);
and U8922 (N_8922,N_1155,N_756);
and U8923 (N_8923,N_213,N_1647);
and U8924 (N_8924,N_2488,N_2414);
nand U8925 (N_8925,N_4220,N_1594);
or U8926 (N_8926,N_1318,N_3524);
nor U8927 (N_8927,N_4897,N_2434);
xnor U8928 (N_8928,N_3616,N_2905);
and U8929 (N_8929,N_4786,N_3538);
nor U8930 (N_8930,N_1448,N_4815);
or U8931 (N_8931,N_3313,N_3469);
nand U8932 (N_8932,N_998,N_3730);
or U8933 (N_8933,N_2596,N_2322);
or U8934 (N_8934,N_4627,N_900);
nor U8935 (N_8935,N_3100,N_683);
nand U8936 (N_8936,N_3960,N_4104);
or U8937 (N_8937,N_1149,N_79);
or U8938 (N_8938,N_4198,N_4593);
nand U8939 (N_8939,N_2225,N_2738);
nand U8940 (N_8940,N_868,N_98);
or U8941 (N_8941,N_3022,N_3944);
nor U8942 (N_8942,N_77,N_1318);
nor U8943 (N_8943,N_2940,N_4724);
nor U8944 (N_8944,N_1254,N_2610);
or U8945 (N_8945,N_3657,N_2188);
or U8946 (N_8946,N_2921,N_831);
nor U8947 (N_8947,N_484,N_779);
or U8948 (N_8948,N_2531,N_1077);
and U8949 (N_8949,N_2928,N_459);
and U8950 (N_8950,N_3629,N_3634);
nor U8951 (N_8951,N_2643,N_4383);
and U8952 (N_8952,N_2916,N_3470);
nor U8953 (N_8953,N_2980,N_533);
nor U8954 (N_8954,N_1507,N_1362);
nand U8955 (N_8955,N_4281,N_1497);
and U8956 (N_8956,N_4488,N_379);
nand U8957 (N_8957,N_93,N_4463);
and U8958 (N_8958,N_1005,N_3805);
xnor U8959 (N_8959,N_858,N_3440);
or U8960 (N_8960,N_717,N_3903);
or U8961 (N_8961,N_619,N_333);
nor U8962 (N_8962,N_1644,N_2134);
or U8963 (N_8963,N_3035,N_3671);
nand U8964 (N_8964,N_2559,N_2392);
xnor U8965 (N_8965,N_823,N_3975);
or U8966 (N_8966,N_2164,N_4174);
nand U8967 (N_8967,N_4436,N_2770);
nor U8968 (N_8968,N_1149,N_1373);
or U8969 (N_8969,N_1308,N_2350);
xnor U8970 (N_8970,N_3249,N_125);
nand U8971 (N_8971,N_3998,N_1447);
nor U8972 (N_8972,N_3554,N_683);
nor U8973 (N_8973,N_3542,N_837);
or U8974 (N_8974,N_1568,N_3505);
xor U8975 (N_8975,N_842,N_3320);
or U8976 (N_8976,N_114,N_2920);
nor U8977 (N_8977,N_699,N_4652);
nand U8978 (N_8978,N_3963,N_4976);
and U8979 (N_8979,N_974,N_2);
nand U8980 (N_8980,N_3,N_2171);
or U8981 (N_8981,N_1105,N_99);
nor U8982 (N_8982,N_4928,N_4458);
nand U8983 (N_8983,N_2245,N_2805);
nand U8984 (N_8984,N_4156,N_3737);
or U8985 (N_8985,N_1442,N_1592);
nor U8986 (N_8986,N_2467,N_735);
and U8987 (N_8987,N_1129,N_4919);
or U8988 (N_8988,N_4044,N_2651);
xnor U8989 (N_8989,N_4926,N_1128);
nor U8990 (N_8990,N_2688,N_2402);
and U8991 (N_8991,N_890,N_4242);
nor U8992 (N_8992,N_1083,N_3079);
nand U8993 (N_8993,N_4590,N_4625);
xnor U8994 (N_8994,N_434,N_4744);
nand U8995 (N_8995,N_3195,N_2657);
or U8996 (N_8996,N_3035,N_1656);
nor U8997 (N_8997,N_3440,N_3363);
and U8998 (N_8998,N_4282,N_2199);
nand U8999 (N_8999,N_1573,N_505);
nor U9000 (N_9000,N_2662,N_2434);
or U9001 (N_9001,N_2525,N_1108);
nor U9002 (N_9002,N_2634,N_354);
or U9003 (N_9003,N_4570,N_2423);
or U9004 (N_9004,N_4094,N_2598);
nor U9005 (N_9005,N_2990,N_417);
or U9006 (N_9006,N_3294,N_4122);
and U9007 (N_9007,N_4526,N_2041);
or U9008 (N_9008,N_2770,N_966);
and U9009 (N_9009,N_796,N_1285);
xor U9010 (N_9010,N_2484,N_3083);
or U9011 (N_9011,N_872,N_3550);
nand U9012 (N_9012,N_463,N_231);
nor U9013 (N_9013,N_2678,N_3861);
and U9014 (N_9014,N_4001,N_3181);
or U9015 (N_9015,N_1413,N_1552);
xnor U9016 (N_9016,N_2763,N_1304);
nor U9017 (N_9017,N_216,N_2412);
nor U9018 (N_9018,N_4435,N_2398);
or U9019 (N_9019,N_1015,N_3627);
or U9020 (N_9020,N_1472,N_129);
or U9021 (N_9021,N_4113,N_2421);
or U9022 (N_9022,N_2089,N_3035);
or U9023 (N_9023,N_4463,N_830);
nor U9024 (N_9024,N_2418,N_1134);
or U9025 (N_9025,N_3522,N_4243);
and U9026 (N_9026,N_3968,N_4566);
or U9027 (N_9027,N_2089,N_2386);
nand U9028 (N_9028,N_1897,N_2814);
xor U9029 (N_9029,N_3079,N_487);
nor U9030 (N_9030,N_4014,N_2505);
nor U9031 (N_9031,N_1833,N_4006);
nor U9032 (N_9032,N_2783,N_1210);
nand U9033 (N_9033,N_3326,N_4573);
xnor U9034 (N_9034,N_15,N_4022);
nand U9035 (N_9035,N_46,N_2422);
or U9036 (N_9036,N_3813,N_3603);
or U9037 (N_9037,N_664,N_2499);
nand U9038 (N_9038,N_1648,N_349);
xor U9039 (N_9039,N_901,N_1018);
or U9040 (N_9040,N_1661,N_1181);
nand U9041 (N_9041,N_4458,N_766);
nor U9042 (N_9042,N_4087,N_1521);
or U9043 (N_9043,N_59,N_1856);
or U9044 (N_9044,N_3432,N_4931);
nand U9045 (N_9045,N_4667,N_2902);
and U9046 (N_9046,N_658,N_4929);
nor U9047 (N_9047,N_988,N_4501);
nor U9048 (N_9048,N_7,N_4285);
or U9049 (N_9049,N_2112,N_3849);
xor U9050 (N_9050,N_1019,N_3641);
xnor U9051 (N_9051,N_1243,N_4553);
or U9052 (N_9052,N_1117,N_899);
and U9053 (N_9053,N_1426,N_2152);
nor U9054 (N_9054,N_3385,N_4543);
nor U9055 (N_9055,N_3968,N_4483);
nor U9056 (N_9056,N_429,N_4256);
and U9057 (N_9057,N_4363,N_803);
and U9058 (N_9058,N_1977,N_2736);
xor U9059 (N_9059,N_3004,N_843);
nand U9060 (N_9060,N_551,N_1335);
and U9061 (N_9061,N_1129,N_1240);
or U9062 (N_9062,N_4542,N_2147);
and U9063 (N_9063,N_3781,N_3939);
nor U9064 (N_9064,N_4810,N_2372);
or U9065 (N_9065,N_722,N_3313);
nor U9066 (N_9066,N_3668,N_4997);
or U9067 (N_9067,N_1865,N_3411);
nand U9068 (N_9068,N_263,N_743);
or U9069 (N_9069,N_487,N_3719);
nand U9070 (N_9070,N_2037,N_1313);
nor U9071 (N_9071,N_3847,N_4412);
or U9072 (N_9072,N_4980,N_4984);
nor U9073 (N_9073,N_395,N_4630);
and U9074 (N_9074,N_2919,N_3616);
or U9075 (N_9075,N_1029,N_2685);
xnor U9076 (N_9076,N_2844,N_4741);
and U9077 (N_9077,N_3162,N_1724);
or U9078 (N_9078,N_902,N_736);
nor U9079 (N_9079,N_3948,N_4508);
nand U9080 (N_9080,N_2610,N_4683);
or U9081 (N_9081,N_1718,N_641);
nor U9082 (N_9082,N_4928,N_4865);
nand U9083 (N_9083,N_1769,N_4803);
and U9084 (N_9084,N_4753,N_2674);
or U9085 (N_9085,N_4421,N_796);
nand U9086 (N_9086,N_549,N_932);
nor U9087 (N_9087,N_2116,N_2943);
and U9088 (N_9088,N_476,N_2503);
or U9089 (N_9089,N_4502,N_1399);
nand U9090 (N_9090,N_3259,N_1371);
nand U9091 (N_9091,N_161,N_4974);
or U9092 (N_9092,N_844,N_1340);
nor U9093 (N_9093,N_958,N_1723);
and U9094 (N_9094,N_2348,N_2386);
nand U9095 (N_9095,N_4558,N_1188);
or U9096 (N_9096,N_3943,N_2242);
and U9097 (N_9097,N_77,N_4961);
or U9098 (N_9098,N_128,N_425);
nand U9099 (N_9099,N_3377,N_3490);
nand U9100 (N_9100,N_4539,N_4784);
and U9101 (N_9101,N_4732,N_3689);
nand U9102 (N_9102,N_1515,N_1207);
or U9103 (N_9103,N_1161,N_2874);
nor U9104 (N_9104,N_1526,N_3437);
or U9105 (N_9105,N_45,N_2848);
nor U9106 (N_9106,N_4694,N_293);
nand U9107 (N_9107,N_269,N_3493);
and U9108 (N_9108,N_149,N_416);
nor U9109 (N_9109,N_3107,N_1143);
xnor U9110 (N_9110,N_4539,N_1207);
or U9111 (N_9111,N_10,N_1592);
or U9112 (N_9112,N_1280,N_1757);
nor U9113 (N_9113,N_2868,N_715);
nand U9114 (N_9114,N_3619,N_3290);
nor U9115 (N_9115,N_2338,N_2957);
or U9116 (N_9116,N_4848,N_4939);
nand U9117 (N_9117,N_4805,N_3852);
xnor U9118 (N_9118,N_623,N_2793);
nand U9119 (N_9119,N_1709,N_1893);
nand U9120 (N_9120,N_2302,N_507);
or U9121 (N_9121,N_889,N_558);
or U9122 (N_9122,N_2313,N_3126);
nand U9123 (N_9123,N_1049,N_753);
and U9124 (N_9124,N_1455,N_893);
nor U9125 (N_9125,N_4542,N_1552);
and U9126 (N_9126,N_4300,N_1885);
xnor U9127 (N_9127,N_2022,N_3109);
nand U9128 (N_9128,N_837,N_4148);
or U9129 (N_9129,N_2423,N_1995);
nor U9130 (N_9130,N_2558,N_2270);
nor U9131 (N_9131,N_4273,N_1416);
xnor U9132 (N_9132,N_4918,N_2496);
nor U9133 (N_9133,N_3990,N_235);
nand U9134 (N_9134,N_2716,N_4820);
or U9135 (N_9135,N_46,N_1473);
xnor U9136 (N_9136,N_2664,N_4706);
and U9137 (N_9137,N_78,N_2069);
nand U9138 (N_9138,N_1619,N_951);
or U9139 (N_9139,N_849,N_4662);
nor U9140 (N_9140,N_2835,N_2698);
nor U9141 (N_9141,N_4400,N_4212);
and U9142 (N_9142,N_3726,N_4903);
nor U9143 (N_9143,N_746,N_2076);
and U9144 (N_9144,N_1196,N_140);
and U9145 (N_9145,N_4480,N_806);
xnor U9146 (N_9146,N_3929,N_1588);
or U9147 (N_9147,N_4867,N_4531);
or U9148 (N_9148,N_2601,N_1009);
nand U9149 (N_9149,N_1389,N_1443);
nand U9150 (N_9150,N_2783,N_3582);
nor U9151 (N_9151,N_4506,N_4361);
nand U9152 (N_9152,N_4738,N_2153);
nand U9153 (N_9153,N_4454,N_4695);
and U9154 (N_9154,N_1774,N_695);
nor U9155 (N_9155,N_1050,N_1329);
or U9156 (N_9156,N_1180,N_1209);
nand U9157 (N_9157,N_3347,N_2397);
and U9158 (N_9158,N_2957,N_2016);
or U9159 (N_9159,N_595,N_3389);
xnor U9160 (N_9160,N_1814,N_2525);
nand U9161 (N_9161,N_473,N_3508);
xor U9162 (N_9162,N_1998,N_1188);
and U9163 (N_9163,N_4360,N_246);
and U9164 (N_9164,N_4867,N_4891);
and U9165 (N_9165,N_4055,N_4758);
and U9166 (N_9166,N_4596,N_0);
and U9167 (N_9167,N_3954,N_2790);
nand U9168 (N_9168,N_4818,N_4400);
nor U9169 (N_9169,N_775,N_2399);
or U9170 (N_9170,N_422,N_4453);
nor U9171 (N_9171,N_4531,N_1258);
nor U9172 (N_9172,N_3709,N_1111);
xnor U9173 (N_9173,N_3256,N_3793);
nor U9174 (N_9174,N_4504,N_1841);
nand U9175 (N_9175,N_1368,N_537);
and U9176 (N_9176,N_4154,N_2346);
or U9177 (N_9177,N_4049,N_1671);
or U9178 (N_9178,N_37,N_3645);
xnor U9179 (N_9179,N_2112,N_1717);
or U9180 (N_9180,N_4009,N_3094);
or U9181 (N_9181,N_1478,N_2869);
and U9182 (N_9182,N_3514,N_3973);
nand U9183 (N_9183,N_339,N_4297);
xnor U9184 (N_9184,N_62,N_4668);
or U9185 (N_9185,N_395,N_262);
or U9186 (N_9186,N_4649,N_511);
nor U9187 (N_9187,N_71,N_394);
or U9188 (N_9188,N_3435,N_1848);
nand U9189 (N_9189,N_2520,N_4538);
nand U9190 (N_9190,N_2340,N_4516);
or U9191 (N_9191,N_1124,N_974);
nor U9192 (N_9192,N_3338,N_4539);
nor U9193 (N_9193,N_3872,N_4948);
nor U9194 (N_9194,N_455,N_4579);
nand U9195 (N_9195,N_1239,N_2302);
nand U9196 (N_9196,N_296,N_429);
nand U9197 (N_9197,N_390,N_1014);
nand U9198 (N_9198,N_1877,N_874);
nor U9199 (N_9199,N_1177,N_1287);
nor U9200 (N_9200,N_1828,N_257);
nand U9201 (N_9201,N_3342,N_1974);
or U9202 (N_9202,N_1353,N_1468);
nor U9203 (N_9203,N_1002,N_3536);
nor U9204 (N_9204,N_1598,N_1611);
and U9205 (N_9205,N_4681,N_3694);
nor U9206 (N_9206,N_4255,N_2552);
or U9207 (N_9207,N_3095,N_3230);
or U9208 (N_9208,N_4931,N_3867);
nor U9209 (N_9209,N_1505,N_1565);
xor U9210 (N_9210,N_1108,N_1215);
nor U9211 (N_9211,N_2080,N_3514);
or U9212 (N_9212,N_1500,N_4402);
nor U9213 (N_9213,N_2338,N_4472);
nand U9214 (N_9214,N_922,N_2613);
nor U9215 (N_9215,N_1450,N_3159);
nand U9216 (N_9216,N_1309,N_326);
xnor U9217 (N_9217,N_591,N_3548);
nor U9218 (N_9218,N_2843,N_4423);
and U9219 (N_9219,N_2393,N_4481);
or U9220 (N_9220,N_586,N_218);
nor U9221 (N_9221,N_64,N_387);
nand U9222 (N_9222,N_894,N_4473);
or U9223 (N_9223,N_2970,N_1895);
and U9224 (N_9224,N_4578,N_4357);
and U9225 (N_9225,N_3379,N_4188);
and U9226 (N_9226,N_4107,N_1704);
or U9227 (N_9227,N_2113,N_1372);
xor U9228 (N_9228,N_2398,N_4298);
nor U9229 (N_9229,N_2106,N_586);
or U9230 (N_9230,N_4427,N_754);
nor U9231 (N_9231,N_1024,N_17);
xnor U9232 (N_9232,N_3651,N_3836);
and U9233 (N_9233,N_4447,N_1514);
nand U9234 (N_9234,N_1368,N_801);
or U9235 (N_9235,N_216,N_4831);
or U9236 (N_9236,N_969,N_3773);
or U9237 (N_9237,N_4776,N_2655);
or U9238 (N_9238,N_3628,N_4308);
or U9239 (N_9239,N_4008,N_1961);
nand U9240 (N_9240,N_4831,N_2468);
nor U9241 (N_9241,N_2073,N_3625);
nor U9242 (N_9242,N_2538,N_3721);
and U9243 (N_9243,N_1553,N_1953);
nand U9244 (N_9244,N_4170,N_739);
nand U9245 (N_9245,N_173,N_4963);
nand U9246 (N_9246,N_4826,N_4295);
or U9247 (N_9247,N_666,N_4240);
nand U9248 (N_9248,N_1032,N_4164);
xor U9249 (N_9249,N_4731,N_608);
nand U9250 (N_9250,N_1662,N_3441);
nand U9251 (N_9251,N_420,N_2531);
nand U9252 (N_9252,N_2529,N_1436);
or U9253 (N_9253,N_1013,N_4946);
nand U9254 (N_9254,N_4674,N_1436);
or U9255 (N_9255,N_2768,N_4205);
nor U9256 (N_9256,N_1240,N_1848);
nand U9257 (N_9257,N_3236,N_1229);
xnor U9258 (N_9258,N_2398,N_1263);
and U9259 (N_9259,N_1399,N_741);
nor U9260 (N_9260,N_3780,N_570);
nor U9261 (N_9261,N_4210,N_1217);
nand U9262 (N_9262,N_377,N_2502);
and U9263 (N_9263,N_1098,N_2282);
and U9264 (N_9264,N_1421,N_4533);
or U9265 (N_9265,N_791,N_1703);
xor U9266 (N_9266,N_3312,N_4153);
and U9267 (N_9267,N_482,N_4752);
and U9268 (N_9268,N_1952,N_6);
nor U9269 (N_9269,N_3367,N_4519);
and U9270 (N_9270,N_4887,N_4564);
nand U9271 (N_9271,N_1904,N_1586);
nor U9272 (N_9272,N_4327,N_4554);
and U9273 (N_9273,N_281,N_736);
nor U9274 (N_9274,N_2299,N_4331);
nand U9275 (N_9275,N_4949,N_378);
or U9276 (N_9276,N_1615,N_1335);
nand U9277 (N_9277,N_2145,N_3180);
nand U9278 (N_9278,N_4642,N_782);
or U9279 (N_9279,N_4646,N_3328);
nor U9280 (N_9280,N_1714,N_2598);
and U9281 (N_9281,N_1970,N_485);
and U9282 (N_9282,N_2569,N_719);
nand U9283 (N_9283,N_4080,N_2795);
xor U9284 (N_9284,N_4314,N_2353);
and U9285 (N_9285,N_12,N_1552);
and U9286 (N_9286,N_4388,N_3437);
and U9287 (N_9287,N_4244,N_3087);
nor U9288 (N_9288,N_3291,N_793);
or U9289 (N_9289,N_27,N_1247);
and U9290 (N_9290,N_660,N_3635);
nand U9291 (N_9291,N_1508,N_578);
nor U9292 (N_9292,N_2782,N_1605);
xor U9293 (N_9293,N_1945,N_3145);
and U9294 (N_9294,N_2045,N_4870);
nand U9295 (N_9295,N_3130,N_4957);
and U9296 (N_9296,N_1266,N_247);
nor U9297 (N_9297,N_89,N_710);
or U9298 (N_9298,N_2006,N_1575);
and U9299 (N_9299,N_3729,N_1944);
or U9300 (N_9300,N_2850,N_3802);
nand U9301 (N_9301,N_3799,N_2759);
nand U9302 (N_9302,N_3862,N_4377);
nand U9303 (N_9303,N_1099,N_926);
or U9304 (N_9304,N_4455,N_2828);
nand U9305 (N_9305,N_3757,N_941);
xnor U9306 (N_9306,N_1585,N_3296);
nand U9307 (N_9307,N_4009,N_3624);
nor U9308 (N_9308,N_1901,N_2182);
nand U9309 (N_9309,N_3966,N_3854);
and U9310 (N_9310,N_2732,N_3207);
xor U9311 (N_9311,N_4380,N_1230);
nor U9312 (N_9312,N_3639,N_481);
nor U9313 (N_9313,N_31,N_3442);
or U9314 (N_9314,N_531,N_1213);
xnor U9315 (N_9315,N_1883,N_3676);
or U9316 (N_9316,N_1531,N_3767);
nand U9317 (N_9317,N_4093,N_144);
nor U9318 (N_9318,N_2525,N_2388);
or U9319 (N_9319,N_1286,N_926);
nor U9320 (N_9320,N_1478,N_2201);
and U9321 (N_9321,N_863,N_1049);
xnor U9322 (N_9322,N_787,N_3815);
nor U9323 (N_9323,N_2137,N_3044);
nand U9324 (N_9324,N_3191,N_3958);
nor U9325 (N_9325,N_4259,N_2876);
or U9326 (N_9326,N_4551,N_4871);
nand U9327 (N_9327,N_717,N_1943);
nand U9328 (N_9328,N_583,N_761);
xnor U9329 (N_9329,N_169,N_4363);
and U9330 (N_9330,N_1781,N_1920);
nand U9331 (N_9331,N_594,N_588);
nand U9332 (N_9332,N_581,N_1676);
nor U9333 (N_9333,N_1107,N_943);
or U9334 (N_9334,N_1395,N_1727);
or U9335 (N_9335,N_4390,N_3928);
and U9336 (N_9336,N_3987,N_4685);
nand U9337 (N_9337,N_2582,N_636);
nor U9338 (N_9338,N_1037,N_3953);
nor U9339 (N_9339,N_1507,N_1780);
and U9340 (N_9340,N_312,N_3254);
and U9341 (N_9341,N_4926,N_2116);
nor U9342 (N_9342,N_2917,N_3609);
nand U9343 (N_9343,N_2034,N_3120);
and U9344 (N_9344,N_1029,N_552);
nand U9345 (N_9345,N_1160,N_2780);
nor U9346 (N_9346,N_3811,N_2219);
and U9347 (N_9347,N_1635,N_1540);
and U9348 (N_9348,N_819,N_4840);
and U9349 (N_9349,N_1962,N_3135);
nand U9350 (N_9350,N_869,N_3155);
nand U9351 (N_9351,N_284,N_2723);
nor U9352 (N_9352,N_1656,N_819);
xnor U9353 (N_9353,N_1451,N_49);
nand U9354 (N_9354,N_4906,N_717);
and U9355 (N_9355,N_1452,N_2811);
and U9356 (N_9356,N_100,N_2411);
and U9357 (N_9357,N_1645,N_4464);
nor U9358 (N_9358,N_504,N_2596);
or U9359 (N_9359,N_2239,N_3629);
nor U9360 (N_9360,N_352,N_2670);
xor U9361 (N_9361,N_2605,N_2956);
nor U9362 (N_9362,N_3257,N_4190);
nand U9363 (N_9363,N_1429,N_2342);
xor U9364 (N_9364,N_3208,N_1038);
or U9365 (N_9365,N_144,N_1287);
and U9366 (N_9366,N_2379,N_1272);
and U9367 (N_9367,N_2543,N_3580);
nor U9368 (N_9368,N_2273,N_645);
and U9369 (N_9369,N_2949,N_2726);
nor U9370 (N_9370,N_3656,N_958);
or U9371 (N_9371,N_2451,N_4820);
xnor U9372 (N_9372,N_2827,N_4747);
and U9373 (N_9373,N_4191,N_4503);
and U9374 (N_9374,N_4541,N_1041);
nor U9375 (N_9375,N_1210,N_4807);
and U9376 (N_9376,N_1,N_1040);
or U9377 (N_9377,N_2074,N_3897);
nor U9378 (N_9378,N_4911,N_3684);
nor U9379 (N_9379,N_325,N_3481);
nor U9380 (N_9380,N_1238,N_1253);
and U9381 (N_9381,N_2835,N_3807);
or U9382 (N_9382,N_4333,N_4420);
xnor U9383 (N_9383,N_926,N_1927);
nor U9384 (N_9384,N_196,N_3698);
nor U9385 (N_9385,N_3378,N_106);
and U9386 (N_9386,N_4418,N_3264);
and U9387 (N_9387,N_338,N_3132);
xor U9388 (N_9388,N_3367,N_977);
nor U9389 (N_9389,N_4791,N_1730);
or U9390 (N_9390,N_3041,N_3937);
nand U9391 (N_9391,N_2824,N_3559);
or U9392 (N_9392,N_2749,N_1443);
nand U9393 (N_9393,N_1614,N_3374);
and U9394 (N_9394,N_3943,N_1734);
nand U9395 (N_9395,N_644,N_2971);
nand U9396 (N_9396,N_1113,N_3621);
or U9397 (N_9397,N_2546,N_4686);
nand U9398 (N_9398,N_773,N_3822);
or U9399 (N_9399,N_686,N_1966);
or U9400 (N_9400,N_2348,N_4868);
nand U9401 (N_9401,N_3882,N_3317);
nor U9402 (N_9402,N_3080,N_93);
nand U9403 (N_9403,N_3107,N_3222);
nor U9404 (N_9404,N_2011,N_3483);
and U9405 (N_9405,N_2515,N_2216);
nor U9406 (N_9406,N_234,N_204);
nor U9407 (N_9407,N_948,N_2313);
or U9408 (N_9408,N_3407,N_34);
nor U9409 (N_9409,N_4905,N_1872);
and U9410 (N_9410,N_957,N_4237);
nor U9411 (N_9411,N_4089,N_29);
xnor U9412 (N_9412,N_1640,N_1085);
nor U9413 (N_9413,N_2880,N_1306);
or U9414 (N_9414,N_3592,N_164);
xor U9415 (N_9415,N_1947,N_1217);
nand U9416 (N_9416,N_1533,N_4728);
nand U9417 (N_9417,N_2251,N_3434);
nand U9418 (N_9418,N_3473,N_1595);
and U9419 (N_9419,N_3543,N_3612);
nand U9420 (N_9420,N_1111,N_1083);
nor U9421 (N_9421,N_4138,N_521);
nand U9422 (N_9422,N_4456,N_2462);
or U9423 (N_9423,N_978,N_2141);
nor U9424 (N_9424,N_3310,N_4996);
nand U9425 (N_9425,N_4332,N_1932);
nor U9426 (N_9426,N_678,N_2869);
or U9427 (N_9427,N_1127,N_922);
or U9428 (N_9428,N_4029,N_2010);
and U9429 (N_9429,N_1027,N_1607);
nand U9430 (N_9430,N_2317,N_4469);
or U9431 (N_9431,N_1630,N_816);
and U9432 (N_9432,N_4590,N_1298);
xnor U9433 (N_9433,N_3296,N_837);
nand U9434 (N_9434,N_648,N_4694);
nor U9435 (N_9435,N_4133,N_4170);
nor U9436 (N_9436,N_3635,N_2236);
nand U9437 (N_9437,N_2028,N_4669);
and U9438 (N_9438,N_2012,N_252);
or U9439 (N_9439,N_3376,N_315);
nor U9440 (N_9440,N_3653,N_3512);
xnor U9441 (N_9441,N_3814,N_1458);
and U9442 (N_9442,N_2231,N_1722);
xor U9443 (N_9443,N_2401,N_894);
and U9444 (N_9444,N_2031,N_3466);
or U9445 (N_9445,N_3096,N_331);
nor U9446 (N_9446,N_616,N_3264);
nor U9447 (N_9447,N_1660,N_3617);
xnor U9448 (N_9448,N_1539,N_3057);
xor U9449 (N_9449,N_1261,N_4241);
nor U9450 (N_9450,N_2035,N_4106);
nand U9451 (N_9451,N_785,N_3338);
and U9452 (N_9452,N_2782,N_3421);
or U9453 (N_9453,N_4841,N_4660);
nor U9454 (N_9454,N_4413,N_4951);
nor U9455 (N_9455,N_2550,N_4069);
nand U9456 (N_9456,N_3769,N_4601);
or U9457 (N_9457,N_3199,N_3000);
xor U9458 (N_9458,N_2858,N_4235);
or U9459 (N_9459,N_1574,N_3634);
nand U9460 (N_9460,N_2330,N_1927);
and U9461 (N_9461,N_3425,N_2012);
or U9462 (N_9462,N_4686,N_199);
nand U9463 (N_9463,N_122,N_2517);
or U9464 (N_9464,N_2521,N_4995);
or U9465 (N_9465,N_2200,N_1807);
nand U9466 (N_9466,N_704,N_3602);
or U9467 (N_9467,N_910,N_3413);
or U9468 (N_9468,N_296,N_1691);
nand U9469 (N_9469,N_4453,N_2743);
nor U9470 (N_9470,N_2309,N_1239);
nand U9471 (N_9471,N_4751,N_2256);
or U9472 (N_9472,N_4452,N_4143);
and U9473 (N_9473,N_2304,N_2024);
and U9474 (N_9474,N_992,N_945);
nand U9475 (N_9475,N_2140,N_116);
or U9476 (N_9476,N_2494,N_535);
xor U9477 (N_9477,N_4562,N_3291);
and U9478 (N_9478,N_1869,N_3541);
nand U9479 (N_9479,N_3934,N_193);
xnor U9480 (N_9480,N_3381,N_1735);
and U9481 (N_9481,N_2494,N_4087);
and U9482 (N_9482,N_2571,N_157);
nand U9483 (N_9483,N_4608,N_1768);
xnor U9484 (N_9484,N_4250,N_3207);
or U9485 (N_9485,N_266,N_4410);
or U9486 (N_9486,N_791,N_4134);
or U9487 (N_9487,N_1681,N_4386);
nor U9488 (N_9488,N_1537,N_1572);
and U9489 (N_9489,N_4042,N_1042);
xnor U9490 (N_9490,N_2913,N_72);
xnor U9491 (N_9491,N_2972,N_4025);
nand U9492 (N_9492,N_1066,N_2290);
nor U9493 (N_9493,N_762,N_635);
and U9494 (N_9494,N_2553,N_2285);
nor U9495 (N_9495,N_744,N_4075);
and U9496 (N_9496,N_1419,N_3715);
nor U9497 (N_9497,N_4798,N_2462);
xor U9498 (N_9498,N_2857,N_2322);
and U9499 (N_9499,N_31,N_2394);
nor U9500 (N_9500,N_306,N_2136);
nor U9501 (N_9501,N_1103,N_4374);
and U9502 (N_9502,N_328,N_2964);
nor U9503 (N_9503,N_1088,N_831);
nand U9504 (N_9504,N_4228,N_807);
nand U9505 (N_9505,N_830,N_3941);
nand U9506 (N_9506,N_798,N_4198);
and U9507 (N_9507,N_2825,N_1923);
or U9508 (N_9508,N_4714,N_1863);
or U9509 (N_9509,N_1287,N_2626);
xnor U9510 (N_9510,N_3552,N_4165);
or U9511 (N_9511,N_3878,N_4546);
or U9512 (N_9512,N_1473,N_1414);
nand U9513 (N_9513,N_2146,N_3233);
and U9514 (N_9514,N_3367,N_3160);
xnor U9515 (N_9515,N_3495,N_1004);
nand U9516 (N_9516,N_772,N_348);
or U9517 (N_9517,N_938,N_4103);
nand U9518 (N_9518,N_2177,N_3720);
and U9519 (N_9519,N_4262,N_917);
xnor U9520 (N_9520,N_3029,N_3987);
nor U9521 (N_9521,N_2145,N_1923);
nand U9522 (N_9522,N_1851,N_1050);
nor U9523 (N_9523,N_670,N_4138);
and U9524 (N_9524,N_67,N_3541);
nand U9525 (N_9525,N_3201,N_3879);
or U9526 (N_9526,N_4236,N_1093);
xor U9527 (N_9527,N_2201,N_1183);
or U9528 (N_9528,N_4501,N_2530);
xnor U9529 (N_9529,N_2555,N_4195);
xor U9530 (N_9530,N_2157,N_4234);
nor U9531 (N_9531,N_1987,N_2070);
nand U9532 (N_9532,N_3934,N_4173);
xor U9533 (N_9533,N_73,N_4214);
nand U9534 (N_9534,N_2906,N_1971);
nor U9535 (N_9535,N_1643,N_3962);
nand U9536 (N_9536,N_158,N_3572);
nand U9537 (N_9537,N_1495,N_390);
and U9538 (N_9538,N_2610,N_949);
or U9539 (N_9539,N_3979,N_1723);
nand U9540 (N_9540,N_2273,N_3256);
or U9541 (N_9541,N_579,N_3728);
or U9542 (N_9542,N_305,N_2701);
or U9543 (N_9543,N_3510,N_910);
nor U9544 (N_9544,N_2664,N_2815);
nor U9545 (N_9545,N_2547,N_3175);
nor U9546 (N_9546,N_2298,N_1334);
nor U9547 (N_9547,N_324,N_3140);
xnor U9548 (N_9548,N_4479,N_849);
nor U9549 (N_9549,N_4228,N_995);
and U9550 (N_9550,N_2194,N_3790);
and U9551 (N_9551,N_1993,N_4651);
or U9552 (N_9552,N_993,N_3441);
nor U9553 (N_9553,N_6,N_4193);
xor U9554 (N_9554,N_2934,N_662);
and U9555 (N_9555,N_4146,N_4030);
nand U9556 (N_9556,N_4645,N_2754);
and U9557 (N_9557,N_678,N_327);
nor U9558 (N_9558,N_3236,N_619);
or U9559 (N_9559,N_166,N_3216);
and U9560 (N_9560,N_3782,N_1716);
or U9561 (N_9561,N_4340,N_3350);
or U9562 (N_9562,N_3409,N_2972);
and U9563 (N_9563,N_3686,N_1218);
and U9564 (N_9564,N_1336,N_263);
nor U9565 (N_9565,N_268,N_3611);
nand U9566 (N_9566,N_1063,N_4041);
or U9567 (N_9567,N_1352,N_4488);
xor U9568 (N_9568,N_3980,N_1215);
nand U9569 (N_9569,N_1980,N_3313);
nand U9570 (N_9570,N_4109,N_655);
nand U9571 (N_9571,N_849,N_2412);
or U9572 (N_9572,N_659,N_556);
and U9573 (N_9573,N_4368,N_2773);
or U9574 (N_9574,N_3388,N_1716);
nor U9575 (N_9575,N_831,N_1262);
and U9576 (N_9576,N_261,N_2848);
or U9577 (N_9577,N_2893,N_1515);
nand U9578 (N_9578,N_4634,N_2639);
nor U9579 (N_9579,N_3073,N_51);
xnor U9580 (N_9580,N_4534,N_4873);
xnor U9581 (N_9581,N_1544,N_3839);
or U9582 (N_9582,N_1568,N_2561);
and U9583 (N_9583,N_4329,N_2271);
or U9584 (N_9584,N_728,N_1618);
nand U9585 (N_9585,N_2049,N_315);
nand U9586 (N_9586,N_374,N_3764);
nor U9587 (N_9587,N_2263,N_4465);
and U9588 (N_9588,N_2321,N_2545);
xnor U9589 (N_9589,N_4075,N_2817);
and U9590 (N_9590,N_3672,N_3913);
nand U9591 (N_9591,N_534,N_585);
and U9592 (N_9592,N_2496,N_3059);
and U9593 (N_9593,N_20,N_2092);
or U9594 (N_9594,N_2693,N_2336);
or U9595 (N_9595,N_447,N_2947);
nand U9596 (N_9596,N_1297,N_2837);
and U9597 (N_9597,N_4755,N_4113);
or U9598 (N_9598,N_1561,N_4580);
and U9599 (N_9599,N_2227,N_4802);
nor U9600 (N_9600,N_503,N_712);
nand U9601 (N_9601,N_3619,N_1552);
nor U9602 (N_9602,N_2117,N_362);
nor U9603 (N_9603,N_2351,N_502);
nand U9604 (N_9604,N_1403,N_3752);
xnor U9605 (N_9605,N_2759,N_3565);
nand U9606 (N_9606,N_4958,N_4268);
nor U9607 (N_9607,N_3492,N_1109);
or U9608 (N_9608,N_1195,N_4242);
nand U9609 (N_9609,N_724,N_145);
and U9610 (N_9610,N_815,N_2688);
nand U9611 (N_9611,N_3271,N_3000);
or U9612 (N_9612,N_4221,N_297);
and U9613 (N_9613,N_4257,N_1437);
or U9614 (N_9614,N_2057,N_605);
nand U9615 (N_9615,N_4270,N_1778);
and U9616 (N_9616,N_3009,N_2034);
or U9617 (N_9617,N_344,N_671);
nand U9618 (N_9618,N_3561,N_1506);
nand U9619 (N_9619,N_3526,N_1807);
nor U9620 (N_9620,N_135,N_3947);
or U9621 (N_9621,N_796,N_1688);
nor U9622 (N_9622,N_4982,N_1891);
nand U9623 (N_9623,N_646,N_830);
nor U9624 (N_9624,N_3991,N_3599);
or U9625 (N_9625,N_2282,N_610);
and U9626 (N_9626,N_3671,N_3917);
or U9627 (N_9627,N_3441,N_2504);
and U9628 (N_9628,N_4888,N_744);
xor U9629 (N_9629,N_2740,N_3269);
and U9630 (N_9630,N_529,N_2193);
and U9631 (N_9631,N_4059,N_2959);
and U9632 (N_9632,N_2030,N_3310);
nand U9633 (N_9633,N_99,N_3103);
xnor U9634 (N_9634,N_4663,N_661);
and U9635 (N_9635,N_2688,N_1432);
nor U9636 (N_9636,N_3622,N_693);
nor U9637 (N_9637,N_694,N_2554);
or U9638 (N_9638,N_4647,N_4038);
or U9639 (N_9639,N_4236,N_156);
nor U9640 (N_9640,N_3107,N_1092);
nand U9641 (N_9641,N_3152,N_2315);
or U9642 (N_9642,N_144,N_4745);
or U9643 (N_9643,N_1327,N_2517);
nand U9644 (N_9644,N_161,N_4560);
nand U9645 (N_9645,N_3954,N_2191);
nand U9646 (N_9646,N_228,N_4493);
or U9647 (N_9647,N_3309,N_587);
nand U9648 (N_9648,N_1363,N_4141);
or U9649 (N_9649,N_3382,N_3791);
and U9650 (N_9650,N_349,N_3287);
or U9651 (N_9651,N_3150,N_1432);
nand U9652 (N_9652,N_2841,N_39);
nand U9653 (N_9653,N_1306,N_4237);
nand U9654 (N_9654,N_1956,N_1209);
nand U9655 (N_9655,N_2255,N_1440);
nand U9656 (N_9656,N_2810,N_4540);
or U9657 (N_9657,N_2899,N_3217);
or U9658 (N_9658,N_3475,N_1613);
and U9659 (N_9659,N_1266,N_4457);
nand U9660 (N_9660,N_4167,N_4324);
or U9661 (N_9661,N_1643,N_1353);
nor U9662 (N_9662,N_1580,N_2883);
nand U9663 (N_9663,N_1891,N_3297);
or U9664 (N_9664,N_2167,N_2422);
nor U9665 (N_9665,N_986,N_2965);
nand U9666 (N_9666,N_1670,N_1949);
or U9667 (N_9667,N_4012,N_362);
nor U9668 (N_9668,N_1313,N_3850);
nand U9669 (N_9669,N_2612,N_2796);
or U9670 (N_9670,N_1371,N_1283);
nor U9671 (N_9671,N_3205,N_3020);
nor U9672 (N_9672,N_13,N_3008);
and U9673 (N_9673,N_4471,N_3519);
nor U9674 (N_9674,N_579,N_2234);
nor U9675 (N_9675,N_4397,N_1067);
nand U9676 (N_9676,N_3828,N_717);
nand U9677 (N_9677,N_3732,N_407);
nor U9678 (N_9678,N_2046,N_2268);
nand U9679 (N_9679,N_1159,N_4352);
or U9680 (N_9680,N_3430,N_2031);
and U9681 (N_9681,N_4882,N_3763);
nor U9682 (N_9682,N_760,N_811);
and U9683 (N_9683,N_4709,N_1207);
nor U9684 (N_9684,N_3692,N_4424);
and U9685 (N_9685,N_728,N_3529);
and U9686 (N_9686,N_1610,N_1279);
nor U9687 (N_9687,N_2578,N_1453);
nand U9688 (N_9688,N_380,N_4257);
nand U9689 (N_9689,N_677,N_4480);
and U9690 (N_9690,N_1845,N_3580);
or U9691 (N_9691,N_4157,N_4072);
or U9692 (N_9692,N_3996,N_1045);
or U9693 (N_9693,N_1077,N_422);
nand U9694 (N_9694,N_1140,N_3099);
and U9695 (N_9695,N_1931,N_391);
or U9696 (N_9696,N_138,N_2402);
and U9697 (N_9697,N_1453,N_4977);
nand U9698 (N_9698,N_1504,N_1388);
and U9699 (N_9699,N_2867,N_1269);
or U9700 (N_9700,N_2841,N_1935);
or U9701 (N_9701,N_1867,N_2639);
and U9702 (N_9702,N_4694,N_4987);
xor U9703 (N_9703,N_1652,N_958);
or U9704 (N_9704,N_1679,N_3899);
and U9705 (N_9705,N_2759,N_2147);
or U9706 (N_9706,N_1158,N_1573);
and U9707 (N_9707,N_4416,N_4960);
or U9708 (N_9708,N_4978,N_1079);
nor U9709 (N_9709,N_4718,N_1674);
nand U9710 (N_9710,N_3595,N_3563);
xnor U9711 (N_9711,N_2143,N_2533);
nand U9712 (N_9712,N_432,N_283);
or U9713 (N_9713,N_3151,N_237);
xnor U9714 (N_9714,N_4673,N_2586);
xnor U9715 (N_9715,N_4466,N_1269);
nand U9716 (N_9716,N_746,N_617);
nand U9717 (N_9717,N_2397,N_2318);
and U9718 (N_9718,N_4922,N_3637);
or U9719 (N_9719,N_3975,N_3409);
nor U9720 (N_9720,N_2696,N_4099);
nand U9721 (N_9721,N_2913,N_965);
or U9722 (N_9722,N_4387,N_4022);
nor U9723 (N_9723,N_748,N_1956);
nor U9724 (N_9724,N_3618,N_698);
nor U9725 (N_9725,N_1902,N_1409);
nor U9726 (N_9726,N_3445,N_2877);
nor U9727 (N_9727,N_1755,N_2188);
and U9728 (N_9728,N_1408,N_1921);
nand U9729 (N_9729,N_4607,N_1686);
nand U9730 (N_9730,N_838,N_675);
or U9731 (N_9731,N_755,N_2203);
xnor U9732 (N_9732,N_1987,N_4734);
nor U9733 (N_9733,N_3943,N_4481);
or U9734 (N_9734,N_4006,N_2108);
and U9735 (N_9735,N_1670,N_1335);
or U9736 (N_9736,N_2406,N_4825);
nand U9737 (N_9737,N_3720,N_3519);
nand U9738 (N_9738,N_1273,N_4735);
and U9739 (N_9739,N_124,N_2939);
nand U9740 (N_9740,N_520,N_3506);
nor U9741 (N_9741,N_1397,N_3508);
or U9742 (N_9742,N_2520,N_543);
or U9743 (N_9743,N_4125,N_4050);
and U9744 (N_9744,N_4364,N_1753);
or U9745 (N_9745,N_3439,N_2817);
nand U9746 (N_9746,N_3331,N_1049);
nor U9747 (N_9747,N_567,N_1471);
nor U9748 (N_9748,N_2711,N_4495);
or U9749 (N_9749,N_3165,N_4009);
nand U9750 (N_9750,N_3204,N_3707);
xnor U9751 (N_9751,N_497,N_1760);
xnor U9752 (N_9752,N_1252,N_2673);
nand U9753 (N_9753,N_4602,N_4951);
nand U9754 (N_9754,N_4774,N_1901);
and U9755 (N_9755,N_640,N_2509);
or U9756 (N_9756,N_1092,N_3594);
nand U9757 (N_9757,N_2903,N_4854);
nand U9758 (N_9758,N_930,N_2138);
and U9759 (N_9759,N_3429,N_2097);
nor U9760 (N_9760,N_3344,N_4788);
xor U9761 (N_9761,N_907,N_2692);
or U9762 (N_9762,N_4510,N_1922);
nor U9763 (N_9763,N_902,N_4278);
nand U9764 (N_9764,N_4544,N_1217);
nor U9765 (N_9765,N_2853,N_4150);
nand U9766 (N_9766,N_441,N_4027);
nand U9767 (N_9767,N_3206,N_136);
and U9768 (N_9768,N_3776,N_529);
and U9769 (N_9769,N_1782,N_2918);
nor U9770 (N_9770,N_1507,N_954);
nor U9771 (N_9771,N_4537,N_1790);
or U9772 (N_9772,N_4810,N_3865);
or U9773 (N_9773,N_3782,N_2218);
xor U9774 (N_9774,N_109,N_2520);
nand U9775 (N_9775,N_4099,N_3579);
or U9776 (N_9776,N_667,N_1791);
xor U9777 (N_9777,N_3648,N_1329);
nor U9778 (N_9778,N_4734,N_1864);
nand U9779 (N_9779,N_2622,N_2214);
and U9780 (N_9780,N_1558,N_4187);
and U9781 (N_9781,N_713,N_3723);
and U9782 (N_9782,N_4854,N_4385);
or U9783 (N_9783,N_1409,N_2619);
nor U9784 (N_9784,N_2444,N_955);
nand U9785 (N_9785,N_715,N_314);
and U9786 (N_9786,N_1130,N_3383);
or U9787 (N_9787,N_3367,N_4023);
nor U9788 (N_9788,N_2448,N_3657);
nor U9789 (N_9789,N_257,N_2869);
and U9790 (N_9790,N_1922,N_3476);
nor U9791 (N_9791,N_374,N_4562);
xor U9792 (N_9792,N_1968,N_3185);
nor U9793 (N_9793,N_380,N_788);
and U9794 (N_9794,N_3539,N_2676);
xor U9795 (N_9795,N_2166,N_4071);
and U9796 (N_9796,N_4495,N_577);
and U9797 (N_9797,N_4561,N_1675);
nor U9798 (N_9798,N_3670,N_955);
or U9799 (N_9799,N_58,N_1820);
nand U9800 (N_9800,N_3838,N_3684);
and U9801 (N_9801,N_4661,N_3527);
or U9802 (N_9802,N_548,N_1861);
xor U9803 (N_9803,N_4017,N_192);
nand U9804 (N_9804,N_2511,N_4545);
or U9805 (N_9805,N_4452,N_2787);
nor U9806 (N_9806,N_3902,N_3032);
nor U9807 (N_9807,N_2492,N_1832);
and U9808 (N_9808,N_4829,N_4835);
or U9809 (N_9809,N_4503,N_644);
or U9810 (N_9810,N_2565,N_1633);
and U9811 (N_9811,N_3939,N_934);
nand U9812 (N_9812,N_2336,N_1051);
and U9813 (N_9813,N_1051,N_4995);
and U9814 (N_9814,N_4935,N_1637);
nand U9815 (N_9815,N_4849,N_494);
nand U9816 (N_9816,N_1269,N_2407);
nand U9817 (N_9817,N_1825,N_3691);
xor U9818 (N_9818,N_351,N_1690);
or U9819 (N_9819,N_4444,N_1886);
nand U9820 (N_9820,N_2171,N_1616);
and U9821 (N_9821,N_2908,N_4568);
nand U9822 (N_9822,N_2339,N_684);
and U9823 (N_9823,N_948,N_933);
or U9824 (N_9824,N_1570,N_2196);
nor U9825 (N_9825,N_536,N_381);
nor U9826 (N_9826,N_4446,N_2353);
nor U9827 (N_9827,N_4684,N_803);
and U9828 (N_9828,N_3565,N_783);
nand U9829 (N_9829,N_4281,N_2218);
or U9830 (N_9830,N_1255,N_2454);
nand U9831 (N_9831,N_660,N_4077);
or U9832 (N_9832,N_2039,N_4290);
nand U9833 (N_9833,N_1214,N_3044);
nor U9834 (N_9834,N_1031,N_4758);
or U9835 (N_9835,N_4234,N_4569);
and U9836 (N_9836,N_2670,N_2684);
nand U9837 (N_9837,N_4352,N_2405);
or U9838 (N_9838,N_621,N_3955);
nor U9839 (N_9839,N_2886,N_3770);
nor U9840 (N_9840,N_2917,N_1576);
xor U9841 (N_9841,N_1490,N_1478);
and U9842 (N_9842,N_1606,N_4844);
and U9843 (N_9843,N_2401,N_2295);
nand U9844 (N_9844,N_4717,N_2551);
nor U9845 (N_9845,N_1171,N_1324);
or U9846 (N_9846,N_2420,N_2803);
and U9847 (N_9847,N_2591,N_3240);
nand U9848 (N_9848,N_4619,N_4397);
nand U9849 (N_9849,N_2180,N_4697);
or U9850 (N_9850,N_3383,N_1324);
xor U9851 (N_9851,N_422,N_4316);
and U9852 (N_9852,N_4422,N_1630);
or U9853 (N_9853,N_4987,N_2570);
nand U9854 (N_9854,N_4238,N_1982);
xnor U9855 (N_9855,N_202,N_2594);
nor U9856 (N_9856,N_4296,N_4873);
and U9857 (N_9857,N_1129,N_2121);
xor U9858 (N_9858,N_756,N_4494);
nor U9859 (N_9859,N_2089,N_3709);
nand U9860 (N_9860,N_1879,N_3914);
and U9861 (N_9861,N_853,N_4030);
or U9862 (N_9862,N_2103,N_4863);
nand U9863 (N_9863,N_4027,N_2368);
or U9864 (N_9864,N_4300,N_3557);
nor U9865 (N_9865,N_3056,N_1523);
and U9866 (N_9866,N_274,N_4967);
nor U9867 (N_9867,N_1817,N_1133);
or U9868 (N_9868,N_336,N_3011);
nand U9869 (N_9869,N_468,N_2497);
and U9870 (N_9870,N_2847,N_2228);
or U9871 (N_9871,N_1697,N_872);
nor U9872 (N_9872,N_178,N_395);
xnor U9873 (N_9873,N_3525,N_2560);
nor U9874 (N_9874,N_4106,N_2636);
and U9875 (N_9875,N_2844,N_3514);
and U9876 (N_9876,N_613,N_1263);
nor U9877 (N_9877,N_2167,N_2918);
or U9878 (N_9878,N_80,N_1877);
nor U9879 (N_9879,N_4168,N_4129);
and U9880 (N_9880,N_2710,N_2031);
nand U9881 (N_9881,N_3261,N_4001);
or U9882 (N_9882,N_1030,N_2067);
and U9883 (N_9883,N_4073,N_4552);
nand U9884 (N_9884,N_3588,N_2934);
nand U9885 (N_9885,N_236,N_4745);
and U9886 (N_9886,N_2604,N_2750);
nor U9887 (N_9887,N_511,N_345);
and U9888 (N_9888,N_4136,N_4172);
nand U9889 (N_9889,N_1964,N_4933);
or U9890 (N_9890,N_4811,N_1545);
nor U9891 (N_9891,N_4772,N_1954);
nor U9892 (N_9892,N_1200,N_2813);
or U9893 (N_9893,N_647,N_504);
nor U9894 (N_9894,N_516,N_4677);
nand U9895 (N_9895,N_666,N_1798);
or U9896 (N_9896,N_396,N_1770);
xnor U9897 (N_9897,N_2314,N_4556);
xor U9898 (N_9898,N_2241,N_298);
xnor U9899 (N_9899,N_4328,N_2923);
and U9900 (N_9900,N_2746,N_4396);
nand U9901 (N_9901,N_4811,N_2681);
nand U9902 (N_9902,N_1551,N_223);
nand U9903 (N_9903,N_32,N_822);
or U9904 (N_9904,N_307,N_2207);
and U9905 (N_9905,N_3759,N_2409);
or U9906 (N_9906,N_2355,N_1065);
or U9907 (N_9907,N_4924,N_3563);
or U9908 (N_9908,N_2703,N_787);
and U9909 (N_9909,N_906,N_477);
xor U9910 (N_9910,N_547,N_3304);
nor U9911 (N_9911,N_3987,N_1943);
nor U9912 (N_9912,N_2927,N_3964);
xor U9913 (N_9913,N_530,N_3560);
nand U9914 (N_9914,N_97,N_1035);
or U9915 (N_9915,N_4225,N_3179);
nor U9916 (N_9916,N_799,N_2879);
nand U9917 (N_9917,N_3385,N_432);
xnor U9918 (N_9918,N_3006,N_3947);
nand U9919 (N_9919,N_1613,N_221);
nor U9920 (N_9920,N_2964,N_1660);
or U9921 (N_9921,N_2247,N_790);
and U9922 (N_9922,N_1120,N_4761);
and U9923 (N_9923,N_4168,N_1075);
nor U9924 (N_9924,N_2519,N_6);
or U9925 (N_9925,N_3560,N_3948);
nand U9926 (N_9926,N_4373,N_4593);
nand U9927 (N_9927,N_4157,N_2752);
and U9928 (N_9928,N_2128,N_3731);
or U9929 (N_9929,N_2092,N_1134);
or U9930 (N_9930,N_4030,N_4131);
or U9931 (N_9931,N_1718,N_3589);
nor U9932 (N_9932,N_2706,N_672);
and U9933 (N_9933,N_898,N_2209);
nor U9934 (N_9934,N_471,N_1107);
and U9935 (N_9935,N_3676,N_1453);
nor U9936 (N_9936,N_304,N_3271);
or U9937 (N_9937,N_4724,N_3922);
nor U9938 (N_9938,N_1785,N_2478);
nor U9939 (N_9939,N_4959,N_4605);
nand U9940 (N_9940,N_4088,N_2847);
or U9941 (N_9941,N_4545,N_750);
or U9942 (N_9942,N_1882,N_1727);
or U9943 (N_9943,N_4577,N_4360);
nor U9944 (N_9944,N_3052,N_3628);
and U9945 (N_9945,N_3961,N_4484);
nand U9946 (N_9946,N_3375,N_4621);
nor U9947 (N_9947,N_3004,N_299);
and U9948 (N_9948,N_3440,N_2342);
nand U9949 (N_9949,N_482,N_1330);
nor U9950 (N_9950,N_3243,N_3861);
or U9951 (N_9951,N_1380,N_2626);
or U9952 (N_9952,N_4350,N_1368);
or U9953 (N_9953,N_3511,N_1754);
xnor U9954 (N_9954,N_4542,N_919);
nand U9955 (N_9955,N_4336,N_4033);
xnor U9956 (N_9956,N_2797,N_11);
nor U9957 (N_9957,N_862,N_3603);
and U9958 (N_9958,N_3787,N_87);
nand U9959 (N_9959,N_1904,N_3639);
nand U9960 (N_9960,N_4292,N_1906);
xor U9961 (N_9961,N_956,N_4121);
or U9962 (N_9962,N_3404,N_3481);
or U9963 (N_9963,N_1646,N_4373);
or U9964 (N_9964,N_4507,N_2194);
xnor U9965 (N_9965,N_4893,N_3954);
xnor U9966 (N_9966,N_4071,N_2601);
nand U9967 (N_9967,N_2648,N_1959);
or U9968 (N_9968,N_346,N_581);
nor U9969 (N_9969,N_2445,N_1325);
and U9970 (N_9970,N_1800,N_2051);
and U9971 (N_9971,N_1447,N_535);
xnor U9972 (N_9972,N_4425,N_68);
and U9973 (N_9973,N_114,N_1498);
nor U9974 (N_9974,N_1070,N_2165);
nor U9975 (N_9975,N_2244,N_755);
or U9976 (N_9976,N_3086,N_3135);
xor U9977 (N_9977,N_1516,N_507);
and U9978 (N_9978,N_265,N_2983);
and U9979 (N_9979,N_1755,N_2998);
or U9980 (N_9980,N_2354,N_2902);
and U9981 (N_9981,N_3184,N_305);
nor U9982 (N_9982,N_1400,N_1465);
nor U9983 (N_9983,N_2815,N_4086);
nor U9984 (N_9984,N_3570,N_2952);
nor U9985 (N_9985,N_1040,N_4559);
xor U9986 (N_9986,N_4084,N_2719);
nand U9987 (N_9987,N_558,N_1154);
nor U9988 (N_9988,N_2888,N_3398);
nor U9989 (N_9989,N_2053,N_2549);
nor U9990 (N_9990,N_2299,N_958);
nor U9991 (N_9991,N_3311,N_3087);
or U9992 (N_9992,N_3259,N_3145);
and U9993 (N_9993,N_912,N_1394);
nand U9994 (N_9994,N_4535,N_1422);
and U9995 (N_9995,N_2027,N_4260);
nand U9996 (N_9996,N_3036,N_2664);
nand U9997 (N_9997,N_2813,N_4293);
or U9998 (N_9998,N_3111,N_1104);
nand U9999 (N_9999,N_712,N_2436);
nor U10000 (N_10000,N_5023,N_8284);
nor U10001 (N_10001,N_7874,N_5203);
and U10002 (N_10002,N_7959,N_5071);
or U10003 (N_10003,N_7102,N_8530);
or U10004 (N_10004,N_8133,N_9475);
and U10005 (N_10005,N_8107,N_6566);
nor U10006 (N_10006,N_5384,N_9008);
nor U10007 (N_10007,N_8891,N_8110);
or U10008 (N_10008,N_5753,N_8356);
nor U10009 (N_10009,N_7767,N_6807);
nand U10010 (N_10010,N_7296,N_8608);
nand U10011 (N_10011,N_6918,N_7036);
or U10012 (N_10012,N_6890,N_7809);
or U10013 (N_10013,N_9749,N_7508);
and U10014 (N_10014,N_9313,N_6838);
nor U10015 (N_10015,N_6555,N_8219);
and U10016 (N_10016,N_5837,N_9478);
and U10017 (N_10017,N_8248,N_7673);
and U10018 (N_10018,N_8402,N_9707);
nor U10019 (N_10019,N_5183,N_5665);
xnor U10020 (N_10020,N_7483,N_9738);
nor U10021 (N_10021,N_5504,N_9615);
nor U10022 (N_10022,N_9299,N_5977);
nand U10023 (N_10023,N_7780,N_9546);
and U10024 (N_10024,N_5114,N_6317);
nor U10025 (N_10025,N_7756,N_9332);
nand U10026 (N_10026,N_6028,N_6655);
xnor U10027 (N_10027,N_5637,N_6251);
and U10028 (N_10028,N_7880,N_5774);
and U10029 (N_10029,N_9335,N_7933);
nand U10030 (N_10030,N_7843,N_7311);
nor U10031 (N_10031,N_7157,N_7962);
xnor U10032 (N_10032,N_5802,N_7750);
nand U10033 (N_10033,N_5043,N_8411);
nand U10034 (N_10034,N_7680,N_7233);
and U10035 (N_10035,N_7377,N_9592);
or U10036 (N_10036,N_5271,N_5532);
and U10037 (N_10037,N_6642,N_8688);
or U10038 (N_10038,N_9722,N_9384);
nand U10039 (N_10039,N_7331,N_7453);
or U10040 (N_10040,N_6470,N_5938);
nor U10041 (N_10041,N_6177,N_5263);
nor U10042 (N_10042,N_8959,N_7869);
or U10043 (N_10043,N_6290,N_9044);
xnor U10044 (N_10044,N_6909,N_5266);
nand U10045 (N_10045,N_8626,N_8625);
and U10046 (N_10046,N_8311,N_5234);
and U10047 (N_10047,N_8423,N_9990);
nand U10048 (N_10048,N_7010,N_9046);
and U10049 (N_10049,N_8047,N_6079);
xnor U10050 (N_10050,N_8708,N_6204);
or U10051 (N_10051,N_7170,N_7626);
nand U10052 (N_10052,N_6243,N_5167);
and U10053 (N_10053,N_8194,N_7766);
nor U10054 (N_10054,N_9892,N_8798);
and U10055 (N_10055,N_7129,N_9355);
and U10056 (N_10056,N_9394,N_8200);
nand U10057 (N_10057,N_5590,N_7186);
xnor U10058 (N_10058,N_5654,N_6946);
nand U10059 (N_10059,N_8760,N_6007);
or U10060 (N_10060,N_8148,N_7642);
or U10061 (N_10061,N_7066,N_7524);
and U10062 (N_10062,N_8205,N_6161);
nand U10063 (N_10063,N_7449,N_6236);
nor U10064 (N_10064,N_8967,N_8266);
nand U10065 (N_10065,N_7250,N_7439);
nand U10066 (N_10066,N_6574,N_8880);
or U10067 (N_10067,N_5869,N_5566);
nand U10068 (N_10068,N_7747,N_9261);
or U10069 (N_10069,N_5691,N_9294);
nor U10070 (N_10070,N_6665,N_8113);
and U10071 (N_10071,N_7405,N_7204);
nor U10072 (N_10072,N_8671,N_6561);
and U10073 (N_10073,N_7293,N_5954);
nand U10074 (N_10074,N_6368,N_9543);
xor U10075 (N_10075,N_8337,N_8914);
nand U10076 (N_10076,N_6127,N_5685);
nor U10077 (N_10077,N_8464,N_7338);
xnor U10078 (N_10078,N_7344,N_5297);
and U10079 (N_10079,N_8268,N_5926);
and U10080 (N_10080,N_6657,N_9515);
and U10081 (N_10081,N_7165,N_5427);
xnor U10082 (N_10082,N_6463,N_5000);
xnor U10083 (N_10083,N_9727,N_7290);
and U10084 (N_10084,N_9582,N_5729);
xor U10085 (N_10085,N_8040,N_7238);
and U10086 (N_10086,N_9014,N_8218);
nor U10087 (N_10087,N_7523,N_6289);
nand U10088 (N_10088,N_8534,N_5188);
nand U10089 (N_10089,N_5990,N_5440);
xnor U10090 (N_10090,N_9288,N_6381);
or U10091 (N_10091,N_6851,N_8136);
and U10092 (N_10092,N_8640,N_5292);
nor U10093 (N_10093,N_9954,N_9520);
nand U10094 (N_10094,N_8463,N_8126);
nand U10095 (N_10095,N_9743,N_8397);
and U10096 (N_10096,N_8335,N_7949);
nor U10097 (N_10097,N_7878,N_6427);
and U10098 (N_10098,N_9759,N_5885);
nand U10099 (N_10099,N_6779,N_5048);
or U10100 (N_10100,N_6626,N_7635);
nor U10101 (N_10101,N_7676,N_8217);
nand U10102 (N_10102,N_9206,N_5128);
nor U10103 (N_10103,N_9870,N_9523);
or U10104 (N_10104,N_8233,N_8225);
or U10105 (N_10105,N_8135,N_5275);
or U10106 (N_10106,N_8869,N_5010);
nor U10107 (N_10107,N_7342,N_8257);
nand U10108 (N_10108,N_6213,N_7215);
nand U10109 (N_10109,N_5482,N_5195);
nand U10110 (N_10110,N_7340,N_7212);
nand U10111 (N_10111,N_9226,N_6706);
nor U10112 (N_10112,N_7113,N_5414);
xnor U10113 (N_10113,N_5904,N_6766);
nand U10114 (N_10114,N_7720,N_7663);
nand U10115 (N_10115,N_7814,N_8923);
nand U10116 (N_10116,N_9694,N_5830);
nor U10117 (N_10117,N_6420,N_5241);
xnor U10118 (N_10118,N_8836,N_9188);
nor U10119 (N_10119,N_7681,N_7650);
nand U10120 (N_10120,N_9279,N_7370);
or U10121 (N_10121,N_9302,N_5295);
xor U10122 (N_10122,N_9411,N_8554);
nand U10123 (N_10123,N_7435,N_5116);
xor U10124 (N_10124,N_8761,N_6187);
or U10125 (N_10125,N_6003,N_6349);
xor U10126 (N_10126,N_6682,N_9851);
or U10127 (N_10127,N_9361,N_5648);
nor U10128 (N_10128,N_8964,N_8473);
nor U10129 (N_10129,N_6728,N_8504);
or U10130 (N_10130,N_9522,N_7565);
or U10131 (N_10131,N_7777,N_9449);
or U10132 (N_10132,N_8030,N_5792);
or U10133 (N_10133,N_6501,N_5040);
nor U10134 (N_10134,N_7566,N_8446);
or U10135 (N_10135,N_6314,N_9060);
and U10136 (N_10136,N_9664,N_6060);
or U10137 (N_10137,N_7368,N_7132);
or U10138 (N_10138,N_8174,N_5528);
nor U10139 (N_10139,N_9252,N_5917);
and U10140 (N_10140,N_5335,N_6955);
nand U10141 (N_10141,N_7348,N_7306);
or U10142 (N_10142,N_9076,N_7028);
nor U10143 (N_10143,N_7828,N_9260);
or U10144 (N_10144,N_9048,N_8331);
or U10145 (N_10145,N_6016,N_9780);
nand U10146 (N_10146,N_5849,N_6661);
nor U10147 (N_10147,N_7572,N_8762);
and U10148 (N_10148,N_7854,N_8156);
or U10149 (N_10149,N_6577,N_7938);
nor U10150 (N_10150,N_8898,N_7522);
or U10151 (N_10151,N_8876,N_9812);
and U10152 (N_10152,N_5300,N_6302);
nand U10153 (N_10153,N_8661,N_5541);
nor U10154 (N_10154,N_5153,N_9640);
nor U10155 (N_10155,N_9340,N_6696);
nand U10156 (N_10156,N_8975,N_8306);
nand U10157 (N_10157,N_8336,N_7582);
xnor U10158 (N_10158,N_6552,N_7585);
and U10159 (N_10159,N_5896,N_6421);
nand U10160 (N_10160,N_9827,N_5616);
and U10161 (N_10161,N_5171,N_7805);
xor U10162 (N_10162,N_6892,N_6419);
and U10163 (N_10163,N_8817,N_5077);
or U10164 (N_10164,N_6369,N_5211);
nor U10165 (N_10165,N_8167,N_7425);
and U10166 (N_10166,N_8521,N_7622);
and U10167 (N_10167,N_5454,N_7471);
and U10168 (N_10168,N_5015,N_8084);
and U10169 (N_10169,N_7423,N_6708);
xor U10170 (N_10170,N_9562,N_9968);
and U10171 (N_10171,N_5923,N_6153);
and U10172 (N_10172,N_6698,N_6397);
and U10173 (N_10173,N_9276,N_5140);
nand U10174 (N_10174,N_7283,N_8339);
nand U10175 (N_10175,N_8827,N_7133);
or U10176 (N_10176,N_9835,N_8789);
nand U10177 (N_10177,N_7643,N_5582);
nand U10178 (N_10178,N_8855,N_9203);
xor U10179 (N_10179,N_8607,N_8104);
nand U10180 (N_10180,N_7893,N_7271);
nor U10181 (N_10181,N_6166,N_7817);
or U10182 (N_10182,N_5578,N_8856);
nor U10183 (N_10183,N_8777,N_6798);
or U10184 (N_10184,N_7083,N_6371);
and U10185 (N_10185,N_6796,N_5014);
or U10186 (N_10186,N_5137,N_8750);
xnor U10187 (N_10187,N_9671,N_7683);
nand U10188 (N_10188,N_7867,N_8875);
and U10189 (N_10189,N_9233,N_8332);
nor U10190 (N_10190,N_7070,N_8681);
and U10191 (N_10191,N_6754,N_7637);
xnor U10192 (N_10192,N_8187,N_7702);
nand U10193 (N_10193,N_8468,N_8531);
or U10194 (N_10194,N_7084,N_8064);
or U10195 (N_10195,N_9551,N_9825);
nand U10196 (N_10196,N_8757,N_8820);
nor U10197 (N_10197,N_8286,N_9366);
and U10198 (N_10198,N_9508,N_6171);
xor U10199 (N_10199,N_5945,N_5217);
nand U10200 (N_10200,N_9028,N_6925);
or U10201 (N_10201,N_7496,N_7154);
nand U10202 (N_10202,N_6418,N_7167);
and U10203 (N_10203,N_8570,N_6628);
nand U10204 (N_10204,N_8767,N_6509);
nor U10205 (N_10205,N_7755,N_5809);
nor U10206 (N_10206,N_7615,N_7833);
nand U10207 (N_10207,N_8497,N_6765);
and U10208 (N_10208,N_8229,N_7699);
or U10209 (N_10209,N_6639,N_9909);
xor U10210 (N_10210,N_8952,N_5035);
or U10211 (N_10211,N_5261,N_5121);
or U10212 (N_10212,N_9310,N_6582);
nand U10213 (N_10213,N_6319,N_5796);
nor U10214 (N_10214,N_6379,N_8621);
or U10215 (N_10215,N_8732,N_7601);
and U10216 (N_10216,N_7035,N_8153);
or U10217 (N_10217,N_5559,N_6843);
nand U10218 (N_10218,N_5033,N_6951);
nor U10219 (N_10219,N_9548,N_9627);
xor U10220 (N_10220,N_9570,N_6593);
and U10221 (N_10221,N_6416,N_6720);
or U10222 (N_10222,N_9591,N_9396);
nand U10223 (N_10223,N_7989,N_6732);
nand U10224 (N_10224,N_9754,N_9274);
and U10225 (N_10225,N_7534,N_6054);
nor U10226 (N_10226,N_9903,N_8164);
and U10227 (N_10227,N_7389,N_8533);
or U10228 (N_10228,N_9326,N_6069);
nor U10229 (N_10229,N_5737,N_8235);
or U10230 (N_10230,N_9783,N_5244);
nor U10231 (N_10231,N_7016,N_7516);
or U10232 (N_10232,N_8522,N_9070);
and U10233 (N_10233,N_9433,N_9693);
and U10234 (N_10234,N_8961,N_5008);
nor U10235 (N_10235,N_7674,N_9860);
or U10236 (N_10236,N_8052,N_7323);
or U10237 (N_10237,N_7691,N_7686);
nand U10238 (N_10238,N_5286,N_7730);
and U10239 (N_10239,N_8175,N_8222);
or U10240 (N_10240,N_8888,N_5872);
nor U10241 (N_10241,N_7863,N_6551);
or U10242 (N_10242,N_7785,N_9862);
and U10243 (N_10243,N_8768,N_5366);
nor U10244 (N_10244,N_7954,N_8202);
xor U10245 (N_10245,N_7009,N_7261);
or U10246 (N_10246,N_5682,N_7487);
nand U10247 (N_10247,N_8700,N_7961);
xor U10248 (N_10248,N_6644,N_9334);
or U10249 (N_10249,N_9593,N_9996);
nand U10250 (N_10250,N_9069,N_8970);
and U10251 (N_10251,N_8444,N_5253);
and U10252 (N_10252,N_7957,N_5553);
and U10253 (N_10253,N_9262,N_6417);
or U10254 (N_10254,N_6677,N_5547);
or U10255 (N_10255,N_9190,N_5332);
nand U10256 (N_10256,N_9883,N_6109);
or U10257 (N_10257,N_9247,N_7705);
nand U10258 (N_10258,N_9360,N_6785);
or U10259 (N_10259,N_8024,N_8103);
and U10260 (N_10260,N_5800,N_7846);
nor U10261 (N_10261,N_5663,N_7289);
nor U10262 (N_10262,N_9145,N_6553);
nand U10263 (N_10263,N_6782,N_6954);
or U10264 (N_10264,N_5264,N_8896);
or U10265 (N_10265,N_7575,N_9094);
or U10266 (N_10266,N_5165,N_7580);
nand U10267 (N_10267,N_8838,N_9815);
nor U10268 (N_10268,N_6764,N_9405);
and U10269 (N_10269,N_7865,N_8460);
and U10270 (N_10270,N_5922,N_5412);
or U10271 (N_10271,N_5229,N_9632);
and U10272 (N_10272,N_6751,N_5469);
nand U10273 (N_10273,N_7710,N_5078);
nand U10274 (N_10274,N_7535,N_8791);
or U10275 (N_10275,N_9061,N_6313);
or U10276 (N_10276,N_5721,N_9751);
or U10277 (N_10277,N_9611,N_9278);
xnor U10278 (N_10278,N_7975,N_9264);
or U10279 (N_10279,N_8071,N_6850);
nor U10280 (N_10280,N_7334,N_7571);
and U10281 (N_10281,N_6744,N_6647);
nor U10282 (N_10282,N_6378,N_9466);
nor U10283 (N_10283,N_9319,N_8962);
nor U10284 (N_10284,N_7542,N_9975);
xor U10285 (N_10285,N_6686,N_7394);
or U10286 (N_10286,N_6978,N_6508);
and U10287 (N_10287,N_6749,N_7031);
nor U10288 (N_10288,N_8943,N_8946);
nand U10289 (N_10289,N_9317,N_6516);
nor U10290 (N_10290,N_8056,N_7462);
nor U10291 (N_10291,N_9790,N_6917);
and U10292 (N_10292,N_8818,N_8172);
or U10293 (N_10293,N_5708,N_9567);
and U10294 (N_10294,N_6131,N_6715);
or U10295 (N_10295,N_5768,N_5820);
and U10296 (N_10296,N_8553,N_6411);
or U10297 (N_10297,N_9974,N_8387);
or U10298 (N_10298,N_7657,N_5081);
and U10299 (N_10299,N_5511,N_9807);
nor U10300 (N_10300,N_6018,N_5437);
nor U10301 (N_10301,N_8926,N_8430);
xor U10302 (N_10302,N_9121,N_9674);
nand U10303 (N_10303,N_7932,N_6351);
nand U10304 (N_10304,N_8597,N_8352);
nand U10305 (N_10305,N_9450,N_7209);
nor U10306 (N_10306,N_5191,N_6869);
nor U10307 (N_10307,N_8714,N_8992);
and U10308 (N_10308,N_5371,N_7275);
nor U10309 (N_10309,N_5401,N_8971);
xor U10310 (N_10310,N_8986,N_7613);
and U10311 (N_10311,N_5206,N_8864);
and U10312 (N_10312,N_8807,N_5961);
and U10313 (N_10313,N_9333,N_5330);
xnor U10314 (N_10314,N_7532,N_8605);
nand U10315 (N_10315,N_7798,N_5278);
xnor U10316 (N_10316,N_5851,N_5053);
xor U10317 (N_10317,N_6868,N_5064);
and U10318 (N_10318,N_9388,N_8067);
xnor U10319 (N_10319,N_5529,N_9944);
and U10320 (N_10320,N_6899,N_6483);
or U10321 (N_10321,N_5397,N_9113);
nand U10322 (N_10322,N_6297,N_9174);
nand U10323 (N_10323,N_9322,N_7378);
or U10324 (N_10324,N_8373,N_9084);
nor U10325 (N_10325,N_8027,N_6941);
and U10326 (N_10326,N_6449,N_6550);
nand U10327 (N_10327,N_6616,N_9139);
nor U10328 (N_10328,N_8206,N_5703);
and U10329 (N_10329,N_7179,N_5385);
xnor U10330 (N_10330,N_9636,N_9373);
nor U10331 (N_10331,N_6305,N_6001);
nor U10332 (N_10332,N_6910,N_6165);
nand U10333 (N_10333,N_6046,N_6095);
or U10334 (N_10334,N_7058,N_6646);
or U10335 (N_10335,N_9762,N_9128);
nor U10336 (N_10336,N_5568,N_9162);
or U10337 (N_10337,N_6522,N_9321);
or U10338 (N_10338,N_6669,N_6725);
nor U10339 (N_10339,N_8270,N_9765);
nand U10340 (N_10340,N_8908,N_8628);
nor U10341 (N_10341,N_6107,N_8025);
and U10342 (N_10342,N_7086,N_7870);
nand U10343 (N_10343,N_7225,N_6596);
and U10344 (N_10344,N_7195,N_8749);
nor U10345 (N_10345,N_7540,N_7324);
nand U10346 (N_10346,N_6286,N_6933);
and U10347 (N_10347,N_5626,N_7446);
nor U10348 (N_10348,N_7033,N_6065);
or U10349 (N_10349,N_9368,N_6307);
nand U10350 (N_10350,N_7858,N_8283);
nand U10351 (N_10351,N_8940,N_9560);
and U10352 (N_10352,N_8800,N_6671);
nor U10353 (N_10353,N_9228,N_7485);
nor U10354 (N_10354,N_6148,N_6163);
and U10355 (N_10355,N_6867,N_5557);
and U10356 (N_10356,N_9631,N_8207);
and U10357 (N_10357,N_9930,N_6160);
nand U10358 (N_10358,N_7052,N_8251);
nand U10359 (N_10359,N_7442,N_9755);
nand U10360 (N_10360,N_9572,N_9001);
nand U10361 (N_10361,N_5946,N_7513);
nand U10362 (N_10362,N_6002,N_9595);
nor U10363 (N_10363,N_7835,N_5026);
nor U10364 (N_10364,N_6479,N_9039);
or U10365 (N_10365,N_9480,N_5173);
nor U10366 (N_10366,N_6713,N_9420);
nor U10367 (N_10367,N_5112,N_8451);
nor U10368 (N_10368,N_8410,N_5569);
xor U10369 (N_10369,N_9179,N_6905);
nand U10370 (N_10370,N_9429,N_6334);
and U10371 (N_10371,N_5196,N_6623);
or U10372 (N_10372,N_7811,N_5890);
nand U10373 (N_10373,N_8137,N_9502);
or U10374 (N_10374,N_5466,N_6916);
or U10375 (N_10375,N_5502,N_9232);
and U10376 (N_10376,N_5819,N_9085);
or U10377 (N_10377,N_6090,N_5575);
or U10378 (N_10378,N_7760,N_9801);
and U10379 (N_10379,N_8059,N_6299);
and U10380 (N_10380,N_7742,N_7085);
xnor U10381 (N_10381,N_9277,N_9474);
nor U10382 (N_10382,N_8366,N_6937);
or U10383 (N_10383,N_9733,N_9779);
and U10384 (N_10384,N_9109,N_7537);
or U10385 (N_10385,N_9787,N_6562);
xnor U10386 (N_10386,N_7191,N_5793);
and U10387 (N_10387,N_7634,N_9410);
nor U10388 (N_10388,N_6173,N_6132);
and U10389 (N_10389,N_7468,N_9623);
and U10390 (N_10390,N_9081,N_9426);
nor U10391 (N_10391,N_9999,N_6841);
nor U10392 (N_10392,N_5102,N_9378);
and U10393 (N_10393,N_7278,N_8435);
xor U10394 (N_10394,N_6523,N_8901);
or U10395 (N_10395,N_8715,N_5987);
nand U10396 (N_10396,N_5434,N_9079);
and U10397 (N_10397,N_5252,N_5747);
nor U10398 (N_10398,N_8329,N_6492);
or U10399 (N_10399,N_9724,N_7396);
nor U10400 (N_10400,N_9925,N_6269);
nor U10401 (N_10401,N_6113,N_7125);
or U10402 (N_10402,N_5940,N_7357);
and U10403 (N_10403,N_5806,N_9122);
and U10404 (N_10404,N_6272,N_5828);
nand U10405 (N_10405,N_8792,N_9767);
nand U10406 (N_10406,N_8633,N_5777);
and U10407 (N_10407,N_7174,N_9600);
nand U10408 (N_10408,N_5059,N_8003);
and U10409 (N_10409,N_6093,N_7207);
nand U10410 (N_10410,N_5018,N_8519);
nor U10411 (N_10411,N_8939,N_5881);
xor U10412 (N_10412,N_8845,N_6865);
and U10413 (N_10413,N_6804,N_5322);
nor U10414 (N_10414,N_9716,N_6947);
or U10415 (N_10415,N_5859,N_8683);
nor U10416 (N_10416,N_6222,N_5296);
nand U10417 (N_10417,N_8328,N_8951);
or U10418 (N_10418,N_7823,N_6261);
or U10419 (N_10419,N_9929,N_5274);
or U10420 (N_10420,N_5647,N_8860);
nand U10421 (N_10421,N_6880,N_8324);
nor U10422 (N_10422,N_9134,N_8018);
or U10423 (N_10423,N_7818,N_5589);
nand U10424 (N_10424,N_9608,N_7567);
xor U10425 (N_10425,N_5291,N_5017);
nor U10426 (N_10426,N_6653,N_6786);
nor U10427 (N_10427,N_7899,N_5692);
nor U10428 (N_10428,N_8582,N_8799);
xor U10429 (N_10429,N_9026,N_5159);
or U10430 (N_10430,N_6747,N_7401);
nand U10431 (N_10431,N_9398,N_5615);
or U10432 (N_10432,N_8591,N_7733);
or U10433 (N_10433,N_6634,N_8100);
nor U10434 (N_10434,N_5585,N_6083);
nand U10435 (N_10435,N_9796,N_7422);
nor U10436 (N_10436,N_9092,N_5340);
nand U10437 (N_10437,N_6812,N_9272);
and U10438 (N_10438,N_8548,N_7546);
and U10439 (N_10439,N_6780,N_6673);
or U10440 (N_10440,N_8999,N_5054);
or U10441 (N_10441,N_7218,N_7797);
or U10442 (N_10442,N_5256,N_6025);
and U10443 (N_10443,N_8031,N_6008);
nor U10444 (N_10444,N_5892,N_5301);
or U10445 (N_10445,N_5298,N_7230);
nor U10446 (N_10446,N_8656,N_7912);
nor U10447 (N_10447,N_8054,N_6473);
nand U10448 (N_10448,N_8546,N_6541);
or U10449 (N_10449,N_8516,N_9886);
or U10450 (N_10450,N_9742,N_7381);
nor U10451 (N_10451,N_5262,N_5231);
nor U10452 (N_10452,N_7024,N_5959);
nor U10453 (N_10453,N_9408,N_6828);
or U10454 (N_10454,N_6276,N_7383);
and U10455 (N_10455,N_8374,N_9868);
or U10456 (N_10456,N_6121,N_6145);
or U10457 (N_10457,N_8779,N_6832);
nand U10458 (N_10458,N_9761,N_6461);
xnor U10459 (N_10459,N_8806,N_7254);
xor U10460 (N_10460,N_8390,N_9973);
nand U10461 (N_10461,N_8433,N_7761);
or U10462 (N_10462,N_7050,N_7268);
nor U10463 (N_10463,N_8486,N_6542);
or U10464 (N_10464,N_7388,N_5678);
nor U10465 (N_10465,N_9197,N_5633);
nand U10466 (N_10466,N_7145,N_7232);
and U10467 (N_10467,N_9142,N_6809);
xor U10468 (N_10468,N_6434,N_6862);
or U10469 (N_10469,N_6757,N_5227);
or U10470 (N_10470,N_8847,N_6388);
or U10471 (N_10471,N_9507,N_6601);
or U10472 (N_10472,N_9427,N_8739);
and U10473 (N_10473,N_5336,N_7198);
nand U10474 (N_10474,N_9393,N_5255);
xnor U10475 (N_10475,N_6260,N_7539);
and U10476 (N_10476,N_5534,N_9099);
nand U10477 (N_10477,N_8606,N_5025);
or U10478 (N_10478,N_8326,N_9620);
or U10479 (N_10479,N_9488,N_5832);
xor U10480 (N_10480,N_9763,N_7404);
or U10481 (N_10481,N_7724,N_5622);
nor U10482 (N_10482,N_7360,N_8890);
nand U10483 (N_10483,N_6528,N_9053);
or U10484 (N_10484,N_8977,N_8965);
nand U10485 (N_10485,N_7884,N_7978);
and U10486 (N_10486,N_8417,N_5860);
nand U10487 (N_10487,N_9810,N_6466);
nand U10488 (N_10488,N_9601,N_8017);
and U10489 (N_10489,N_6837,N_5104);
and U10490 (N_10490,N_6099,N_8191);
nand U10491 (N_10491,N_9352,N_8885);
nor U10492 (N_10492,N_9919,N_6220);
nor U10493 (N_10493,N_5488,N_7612);
nand U10494 (N_10494,N_8163,N_7092);
and U10495 (N_10495,N_7861,N_6218);
or U10496 (N_10496,N_6294,N_9708);
and U10497 (N_10497,N_7936,N_9556);
or U10498 (N_10498,N_6078,N_5480);
nand U10499 (N_10499,N_8512,N_6848);
nor U10500 (N_10500,N_6558,N_7386);
nor U10501 (N_10501,N_9731,N_7712);
xor U10502 (N_10502,N_8069,N_6377);
or U10503 (N_10503,N_5445,N_5503);
xnor U10504 (N_10504,N_9561,N_9689);
and U10505 (N_10505,N_5536,N_9106);
or U10506 (N_10506,N_7726,N_7560);
or U10507 (N_10507,N_5443,N_8935);
nor U10508 (N_10508,N_7335,N_8709);
nor U10509 (N_10509,N_9630,N_9390);
or U10510 (N_10510,N_8012,N_8747);
nor U10511 (N_10511,N_9726,N_5989);
and U10512 (N_10512,N_7151,N_6363);
and U10513 (N_10513,N_8281,N_6896);
nand U10514 (N_10514,N_7799,N_8611);
nor U10515 (N_10515,N_5399,N_9859);
nand U10516 (N_10516,N_9078,N_6203);
nand U10517 (N_10517,N_5916,N_7452);
xnor U10518 (N_10518,N_5943,N_9040);
and U10519 (N_10519,N_6795,N_8906);
nor U10520 (N_10520,N_9413,N_5007);
nor U10521 (N_10521,N_8835,N_6977);
nand U10522 (N_10522,N_6930,N_7563);
nand U10523 (N_10523,N_6717,N_7801);
or U10524 (N_10524,N_7034,N_6540);
or U10525 (N_10525,N_7193,N_8123);
and U10526 (N_10526,N_7856,N_5329);
and U10527 (N_10527,N_8049,N_5225);
and U10528 (N_10528,N_7175,N_5420);
and U10529 (N_10529,N_8592,N_9662);
nand U10530 (N_10530,N_8393,N_9432);
or U10531 (N_10531,N_9163,N_5660);
or U10532 (N_10532,N_6675,N_8731);
or U10533 (N_10533,N_8545,N_6469);
nor U10534 (N_10534,N_8996,N_8478);
nor U10535 (N_10535,N_5370,N_7987);
xnor U10536 (N_10536,N_8086,N_8034);
and U10537 (N_10537,N_5327,N_8917);
nand U10538 (N_10538,N_7548,N_9187);
nor U10539 (N_10539,N_9734,N_9415);
nand U10540 (N_10540,N_5646,N_5146);
nand U10541 (N_10541,N_7554,N_7281);
and U10542 (N_10542,N_5103,N_9180);
nor U10543 (N_10543,N_6565,N_8703);
nand U10544 (N_10544,N_8601,N_5560);
and U10545 (N_10545,N_7916,N_8445);
and U10546 (N_10546,N_5710,N_5333);
or U10547 (N_10547,N_5700,N_9969);
xnor U10548 (N_10548,N_5744,N_5694);
nand U10549 (N_10549,N_7677,N_6609);
xor U10550 (N_10550,N_7527,N_7492);
nor U10551 (N_10551,N_7124,N_5825);
and U10552 (N_10552,N_6108,N_6968);
and U10553 (N_10553,N_9802,N_5199);
and U10554 (N_10554,N_9402,N_7181);
nand U10555 (N_10555,N_7928,N_6077);
or U10556 (N_10556,N_5621,N_9425);
or U10557 (N_10557,N_7944,N_7482);
nor U10558 (N_10558,N_8617,N_7842);
and U10559 (N_10559,N_5533,N_9250);
nor U10560 (N_10560,N_7350,N_5215);
nand U10561 (N_10561,N_9245,N_8822);
or U10562 (N_10562,N_8036,N_9579);
nand U10563 (N_10563,N_7438,N_8584);
nor U10564 (N_10564,N_7326,N_7526);
nor U10565 (N_10565,N_8960,N_9819);
nor U10566 (N_10566,N_7624,N_6598);
or U10567 (N_10567,N_7087,N_7018);
and U10568 (N_10568,N_8193,N_7904);
nand U10569 (N_10569,N_6454,N_6876);
nor U10570 (N_10570,N_9112,N_5228);
nor U10571 (N_10571,N_7505,N_7509);
xor U10572 (N_10572,N_7606,N_8509);
nand U10573 (N_10573,N_7988,N_8763);
or U10574 (N_10574,N_7619,N_9265);
nand U10575 (N_10575,N_7282,N_6659);
nand U10576 (N_10576,N_5906,N_8021);
nor U10577 (N_10577,N_5882,N_6051);
and U10578 (N_10578,N_5960,N_6777);
nand U10579 (N_10579,N_8276,N_9283);
and U10580 (N_10580,N_5612,N_6074);
nand U10581 (N_10581,N_7387,N_6600);
nor U10582 (N_10582,N_7757,N_9087);
or U10583 (N_10583,N_8878,N_7149);
nor U10584 (N_10584,N_9703,N_7071);
nor U10585 (N_10585,N_7398,N_5438);
or U10586 (N_10586,N_8942,N_6386);
and U10587 (N_10587,N_5154,N_6859);
or U10588 (N_10588,N_5174,N_5857);
and U10589 (N_10589,N_5979,N_9816);
and U10590 (N_10590,N_8802,N_7493);
nand U10591 (N_10591,N_6071,N_5164);
xnor U10592 (N_10592,N_7896,N_8660);
xnor U10593 (N_10593,N_8400,N_7860);
nand U10594 (N_10594,N_9090,N_9879);
xnor U10595 (N_10595,N_8684,N_8587);
and U10596 (N_10596,N_5824,N_5599);
or U10597 (N_10597,N_9271,N_8159);
nand U10598 (N_10598,N_8242,N_7672);
nand U10599 (N_10599,N_6200,N_7019);
nand U10600 (N_10600,N_9178,N_9448);
or U10601 (N_10601,N_8277,N_5094);
nor U10602 (N_10602,N_9291,N_7678);
nand U10603 (N_10603,N_5134,N_8697);
or U10604 (N_10604,N_8169,N_7246);
xor U10605 (N_10605,N_6857,N_7333);
nand U10606 (N_10606,N_5257,N_7300);
nor U10607 (N_10607,N_6664,N_8566);
or U10608 (N_10608,N_7866,N_7640);
nand U10609 (N_10609,N_7719,N_5013);
nand U10610 (N_10610,N_8250,N_8050);
and U10611 (N_10611,N_9209,N_8981);
xnor U10612 (N_10612,N_6240,N_7110);
or U10613 (N_10613,N_9364,N_8705);
or U10614 (N_10614,N_5984,N_5745);
and U10615 (N_10615,N_8490,N_5049);
nand U10616 (N_10616,N_9945,N_7199);
or U10617 (N_10617,N_7688,N_5863);
and U10618 (N_10618,N_9843,N_8717);
nor U10619 (N_10619,N_5603,N_5994);
and U10620 (N_10620,N_9957,N_8212);
or U10621 (N_10621,N_6239,N_9865);
nor U10622 (N_10622,N_8849,N_7886);
and U10623 (N_10623,N_5226,N_9207);
nand U10624 (N_10624,N_8759,N_9628);
or U10625 (N_10625,N_8272,N_9298);
xnor U10626 (N_10626,N_7308,N_9012);
nand U10627 (N_10627,N_5346,N_7359);
and U10628 (N_10628,N_7943,N_9249);
nand U10629 (N_10629,N_7897,N_9371);
nor U10630 (N_10630,N_9728,N_6581);
or U10631 (N_10631,N_5780,N_8391);
nand U10632 (N_10632,N_5967,N_7868);
nor U10633 (N_10633,N_7395,N_5667);
nor U10634 (N_10634,N_8032,N_9997);
and U10635 (N_10635,N_8648,N_7782);
nor U10636 (N_10636,N_7481,N_8058);
xnor U10637 (N_10637,N_8581,N_9876);
nand U10638 (N_10638,N_6215,N_5381);
and U10639 (N_10639,N_9100,N_7638);
nand U10640 (N_10640,N_5235,N_8361);
and U10641 (N_10641,N_5743,N_9544);
xnor U10642 (N_10642,N_8215,N_8309);
and U10643 (N_10643,N_7557,N_8360);
and U10644 (N_10644,N_7245,N_5630);
nor U10645 (N_10645,N_5803,N_6961);
nor U10646 (N_10646,N_8974,N_8552);
and U10647 (N_10647,N_8603,N_6993);
or U10648 (N_10648,N_8803,N_9343);
or U10649 (N_10649,N_8895,N_6159);
or U10650 (N_10650,N_7711,N_8154);
nand U10651 (N_10651,N_8278,N_6919);
nand U10652 (N_10652,N_7850,N_7100);
and U10653 (N_10653,N_8448,N_6327);
nand U10654 (N_10654,N_9453,N_9266);
nor U10655 (N_10655,N_7431,N_5587);
xor U10656 (N_10656,N_8882,N_7718);
xor U10657 (N_10657,N_9829,N_5720);
and U10658 (N_10658,N_6491,N_6306);
and U10659 (N_10659,N_9893,N_8048);
and U10660 (N_10660,N_9468,N_8517);
and U10661 (N_10661,N_9050,N_6189);
or U10662 (N_10662,N_8357,N_5570);
nand U10663 (N_10663,N_8293,N_5730);
and U10664 (N_10664,N_5377,N_9086);
nand U10665 (N_10665,N_7136,N_7781);
or U10666 (N_10666,N_5883,N_9856);
nand U10667 (N_10667,N_8440,N_7942);
and U10668 (N_10668,N_6788,N_9451);
nand U10669 (N_10669,N_8394,N_8810);
and U10670 (N_10670,N_5843,N_7784);
xnor U10671 (N_10671,N_7309,N_9447);
and U10672 (N_10672,N_7032,N_9846);
or U10673 (N_10673,N_6357,N_8042);
nor U10674 (N_10674,N_5728,N_7159);
and U10675 (N_10675,N_7917,N_5738);
nor U10676 (N_10676,N_7919,N_8907);
nand U10677 (N_10677,N_8070,N_5016);
nor U10678 (N_10678,N_7443,N_7895);
xor U10679 (N_10679,N_7690,N_7558);
nand U10680 (N_10680,N_8046,N_6155);
and U10681 (N_10681,N_8784,N_7806);
and U10682 (N_10682,N_5718,N_5386);
nor U10683 (N_10683,N_5258,N_7042);
or U10684 (N_10684,N_5672,N_9155);
and U10685 (N_10685,N_9773,N_8934);
nand U10686 (N_10686,N_8734,N_7771);
nor U10687 (N_10687,N_8995,N_9290);
and U10688 (N_10688,N_6597,N_9713);
or U10689 (N_10689,N_9756,N_7337);
nand U10690 (N_10690,N_8130,N_6915);
or U10691 (N_10691,N_6519,N_8080);
nor U10692 (N_10692,N_6962,N_5373);
nor U10693 (N_10693,N_7974,N_6157);
nand U10694 (N_10694,N_7736,N_6718);
or U10695 (N_10695,N_7918,N_6017);
nand U10696 (N_10696,N_6545,N_5908);
nor U10697 (N_10697,N_8057,N_6824);
nor U10698 (N_10698,N_6587,N_9136);
and U10699 (N_10699,N_6502,N_9370);
or U10700 (N_10700,N_9744,N_6928);
and U10701 (N_10701,N_6632,N_5549);
nand U10702 (N_10702,N_8915,N_5003);
nor U10703 (N_10703,N_7594,N_5070);
and U10704 (N_10704,N_6086,N_7945);
nor U10705 (N_10705,N_6943,N_9688);
and U10706 (N_10706,N_7248,N_5283);
nor U10707 (N_10707,N_5472,N_7689);
or U10708 (N_10708,N_9214,N_7295);
nand U10709 (N_10709,N_8909,N_9284);
or U10710 (N_10710,N_6112,N_8457);
or U10711 (N_10711,N_7502,N_5209);
nand U10712 (N_10712,N_6092,N_9157);
nand U10713 (N_10713,N_9438,N_6284);
nor U10714 (N_10714,N_8183,N_7630);
nor U10715 (N_10715,N_8949,N_8736);
xnor U10716 (N_10716,N_8425,N_9532);
nor U10717 (N_10717,N_8004,N_9032);
xor U10718 (N_10718,N_8378,N_7447);
nand U10719 (N_10719,N_6343,N_5521);
or U10720 (N_10720,N_8598,N_7759);
or U10721 (N_10721,N_5831,N_9114);
nand U10722 (N_10722,N_6929,N_9093);
or U10723 (N_10723,N_7065,N_5834);
nor U10724 (N_10724,N_9914,N_8053);
or U10725 (N_10725,N_8733,N_8737);
xnor U10726 (N_10726,N_7237,N_5912);
xnor U10727 (N_10727,N_6986,N_5441);
or U10728 (N_10728,N_9854,N_7697);
or U10729 (N_10729,N_6506,N_7549);
or U10730 (N_10730,N_5523,N_6114);
and U10731 (N_10731,N_9482,N_5527);
nor U10732 (N_10732,N_9823,N_5197);
and U10733 (N_10733,N_5361,N_9234);
nand U10734 (N_10734,N_8675,N_9471);
and U10735 (N_10735,N_6965,N_8401);
and U10736 (N_10736,N_5684,N_5424);
xnor U10737 (N_10737,N_8723,N_8746);
nand U10738 (N_10738,N_7967,N_7707);
or U10739 (N_10739,N_8699,N_6105);
and U10740 (N_10740,N_8090,N_7948);
or U10741 (N_10741,N_5276,N_7969);
nand U10742 (N_10742,N_6990,N_5158);
nand U10743 (N_10743,N_6146,N_9198);
and U10744 (N_10744,N_6457,N_6726);
nand U10745 (N_10745,N_6339,N_9979);
or U10746 (N_10746,N_8881,N_5492);
nand U10747 (N_10747,N_6612,N_6818);
nand U10748 (N_10748,N_9107,N_6560);
xor U10749 (N_10749,N_7054,N_7455);
and U10750 (N_10750,N_7708,N_5545);
and U10751 (N_10751,N_5893,N_9477);
or U10752 (N_10752,N_7122,N_6622);
and U10753 (N_10753,N_9686,N_9704);
nand U10754 (N_10754,N_8081,N_9080);
nand U10755 (N_10755,N_7473,N_9347);
xor U10756 (N_10756,N_9280,N_5680);
or U10757 (N_10757,N_9148,N_6940);
xnor U10758 (N_10758,N_6452,N_7864);
nand U10759 (N_10759,N_5949,N_5794);
or U10760 (N_10760,N_6201,N_6580);
or U10761 (N_10761,N_7783,N_6216);
or U10762 (N_10762,N_8631,N_8290);
nand U10763 (N_10763,N_7459,N_9439);
nand U10764 (N_10764,N_6663,N_7569);
and U10765 (N_10765,N_6745,N_6453);
or U10766 (N_10766,N_8379,N_8542);
nand U10767 (N_10767,N_7413,N_5168);
xor U10768 (N_10768,N_7464,N_6439);
and U10769 (N_10769,N_8299,N_9225);
or U10770 (N_10770,N_5273,N_8916);
nand U10771 (N_10771,N_8184,N_7807);
and U10772 (N_10772,N_5876,N_8038);
or U10773 (N_10773,N_5931,N_9182);
nor U10774 (N_10774,N_5179,N_7568);
and U10775 (N_10775,N_6620,N_8775);
nand U10776 (N_10776,N_6115,N_9063);
nand U10777 (N_10777,N_5285,N_7940);
nor U10778 (N_10778,N_7048,N_7775);
nand U10779 (N_10779,N_9489,N_6383);
and U10780 (N_10780,N_8376,N_5066);
nand U10781 (N_10781,N_9421,N_5783);
nand U10782 (N_10782,N_5447,N_9065);
or U10783 (N_10783,N_5456,N_5929);
or U10784 (N_10784,N_6300,N_9111);
or U10785 (N_10785,N_7901,N_7094);
nor U10786 (N_10786,N_9541,N_9972);
or U10787 (N_10787,N_9023,N_6366);
or U10788 (N_10788,N_7737,N_5143);
and U10789 (N_10789,N_5713,N_5731);
or U10790 (N_10790,N_7617,N_5868);
xnor U10791 (N_10791,N_9305,N_6852);
xor U10792 (N_10792,N_5243,N_6769);
xor U10793 (N_10793,N_9146,N_6921);
nand U10794 (N_10794,N_6206,N_5021);
and U10795 (N_10795,N_5187,N_8809);
or U10796 (N_10796,N_6856,N_6110);
or U10797 (N_10797,N_5563,N_8976);
nand U10798 (N_10798,N_5249,N_6504);
nand U10799 (N_10799,N_5152,N_9690);
nor U10800 (N_10800,N_7143,N_7924);
nand U10801 (N_10801,N_8147,N_5478);
nand U10802 (N_10802,N_6731,N_7112);
or U10803 (N_10803,N_9720,N_5106);
nand U10804 (N_10804,N_8614,N_7972);
xor U10805 (N_10805,N_6643,N_8011);
or U10806 (N_10806,N_6956,N_5163);
or U10807 (N_10807,N_6624,N_8441);
nor U10808 (N_10808,N_6141,N_9839);
and U10809 (N_10809,N_6283,N_7138);
or U10810 (N_10810,N_8630,N_9075);
or U10811 (N_10811,N_9123,N_6296);
or U10812 (N_10812,N_7417,N_8596);
and U10813 (N_10813,N_6035,N_7570);
nor U10814 (N_10814,N_6242,N_7373);
or U10815 (N_10815,N_6683,N_8892);
and U10816 (N_10816,N_7553,N_5204);
nor U10817 (N_10817,N_9953,N_8349);
nor U10818 (N_10818,N_8418,N_6458);
or U10819 (N_10819,N_6496,N_7881);
nor U10820 (N_10820,N_6874,N_6384);
and U10821 (N_10821,N_6375,N_9700);
nand U10822 (N_10822,N_5221,N_7269);
xnor U10823 (N_10823,N_6872,N_7564);
nand U10824 (N_10824,N_7654,N_7150);
nor U10825 (N_10825,N_5198,N_9387);
nor U10826 (N_10826,N_9853,N_7111);
or U10827 (N_10827,N_8662,N_8990);
or U10828 (N_10828,N_6019,N_8501);
nor U10829 (N_10829,N_8900,N_8744);
xnor U10830 (N_10830,N_5328,N_6244);
or U10831 (N_10831,N_9282,N_9037);
nand U10832 (N_10832,N_6576,N_8226);
nor U10833 (N_10833,N_9991,N_7813);
xnor U10834 (N_10834,N_7292,N_5218);
and U10835 (N_10835,N_9542,N_5044);
xnor U10836 (N_10836,N_8108,N_8893);
nand U10837 (N_10837,N_8317,N_7616);
xor U10838 (N_10838,N_9663,N_6012);
nand U10839 (N_10839,N_8002,N_5352);
and U10840 (N_10840,N_6330,N_5175);
nand U10841 (N_10841,N_8858,N_9629);
nor U10842 (N_10842,N_7504,N_6654);
nor U10843 (N_10843,N_9147,N_8342);
nand U10844 (N_10844,N_7451,N_7498);
xnor U10845 (N_10845,N_8168,N_9685);
xnor U10846 (N_10846,N_6329,N_6789);
and U10847 (N_10847,N_9901,N_7667);
or U10848 (N_10848,N_8978,N_8416);
or U10849 (N_10849,N_8937,N_9933);
nor U10850 (N_10850,N_9644,N_5331);
or U10851 (N_10851,N_6518,N_8456);
nand U10852 (N_10852,N_9263,N_9792);
nor U10853 (N_10853,N_5259,N_9500);
or U10854 (N_10854,N_6342,N_5305);
nand U10855 (N_10855,N_7220,N_6234);
or U10856 (N_10856,N_6122,N_5190);
nand U10857 (N_10857,N_5150,N_9858);
and U10858 (N_10858,N_8271,N_5702);
and U10859 (N_10859,N_5607,N_8488);
and U10860 (N_10860,N_5814,N_6301);
nor U10861 (N_10861,N_5358,N_7093);
xnor U10862 (N_10862,N_5552,N_7687);
nand U10863 (N_10863,N_7930,N_8826);
nand U10864 (N_10864,N_7670,N_6588);
and U10865 (N_10865,N_5601,N_6711);
nand U10866 (N_10866,N_6311,N_7728);
nor U10867 (N_10867,N_8580,N_7922);
nor U10868 (N_10868,N_9545,N_8467);
and U10869 (N_10869,N_5795,N_9273);
nor U10870 (N_10870,N_7596,N_9652);
xnor U10871 (N_10871,N_6144,N_5411);
nor U10872 (N_10872,N_5404,N_8143);
nand U10873 (N_10873,N_7385,N_7853);
nor U10874 (N_10874,N_7890,N_5915);
nor U10875 (N_10875,N_9978,N_5476);
or U10876 (N_10876,N_6428,N_8615);
or U10877 (N_10877,N_5415,N_5457);
and U10878 (N_10878,N_5047,N_9875);
nor U10879 (N_10879,N_6413,N_8323);
or U10880 (N_10880,N_9306,N_9777);
and U10881 (N_10881,N_9725,N_8785);
or U10882 (N_10882,N_5548,N_8948);
or U10883 (N_10883,N_8029,N_8181);
nor U10884 (N_10884,N_5368,N_6511);
and U10885 (N_10885,N_8221,N_5405);
nor U10886 (N_10886,N_8616,N_9503);
nand U10887 (N_10887,N_8556,N_5334);
nor U10888 (N_10888,N_8573,N_8128);
and U10889 (N_10889,N_5676,N_9312);
or U10890 (N_10890,N_9119,N_9712);
nor U10891 (N_10891,N_7800,N_7287);
nand U10892 (N_10892,N_7913,N_7909);
nor U10893 (N_10893,N_8897,N_7288);
nor U10894 (N_10894,N_9985,N_6241);
and U10895 (N_10895,N_9452,N_5345);
and U10896 (N_10896,N_5074,N_9926);
nor U10897 (N_10897,N_8527,N_7076);
and U10898 (N_10898,N_9463,N_6101);
nor U10899 (N_10899,N_7146,N_9517);
and U10900 (N_10900,N_7082,N_6073);
nor U10901 (N_10901,N_5056,N_9173);
or U10902 (N_10902,N_9956,N_5580);
and U10903 (N_10903,N_6571,N_7131);
nand U10904 (N_10904,N_7079,N_8129);
or U10905 (N_10905,N_7310,N_8993);
nor U10906 (N_10906,N_8773,N_5619);
nor U10907 (N_10907,N_7297,N_6960);
or U10908 (N_10908,N_7351,N_7512);
xnor U10909 (N_10909,N_6679,N_7277);
or U10910 (N_10910,N_5316,N_9857);
nand U10911 (N_10911,N_8026,N_8333);
or U10912 (N_10912,N_5639,N_9506);
nor U10913 (N_10913,N_9995,N_9491);
nand U10914 (N_10914,N_7703,N_7382);
nor U10915 (N_10915,N_9131,N_5085);
nor U10916 (N_10916,N_5576,N_5661);
nor U10917 (N_10917,N_6712,N_7812);
xnor U10918 (N_10918,N_7322,N_6674);
nand U10919 (N_10919,N_6459,N_8480);
nor U10920 (N_10920,N_9607,N_9639);
and U10921 (N_10921,N_6637,N_5247);
and U10922 (N_10922,N_7479,N_6298);
and U10923 (N_10923,N_5740,N_6407);
or U10924 (N_10924,N_6337,N_6836);
nor U10925 (N_10925,N_8973,N_9314);
and U10926 (N_10926,N_6088,N_6816);
nand U10927 (N_10927,N_5784,N_7046);
xnor U10928 (N_10928,N_9992,N_6793);
and U10929 (N_10929,N_9318,N_8145);
xnor U10930 (N_10930,N_7214,N_7857);
or U10931 (N_10931,N_5130,N_6367);
nor U10932 (N_10932,N_7127,N_7577);
and U10933 (N_10933,N_8470,N_6500);
or U10934 (N_10934,N_8178,N_6405);
xnor U10935 (N_10935,N_7844,N_5119);
xor U10936 (N_10936,N_9651,N_8911);
nor U10937 (N_10937,N_8513,N_7315);
and U10938 (N_10938,N_6027,N_9133);
nand U10939 (N_10939,N_8341,N_5833);
nand U10940 (N_10940,N_5757,N_8359);
xnor U10941 (N_10941,N_7227,N_8557);
and U10942 (N_10942,N_5564,N_7979);
nand U10943 (N_10943,N_5838,N_8969);
and U10944 (N_10944,N_7397,N_6787);
nor U10945 (N_10945,N_7578,N_9464);
nand U10946 (N_10946,N_8102,N_7060);
and U10947 (N_10947,N_5635,N_9550);
and U10948 (N_10948,N_8083,N_9456);
nor U10949 (N_10949,N_9817,N_6532);
and U10950 (N_10950,N_9913,N_9916);
nor U10951 (N_10951,N_7105,N_7555);
or U10952 (N_10952,N_8098,N_8313);
xnor U10953 (N_10953,N_6752,N_9524);
and U10954 (N_10954,N_6557,N_7080);
nand U10955 (N_10955,N_9614,N_7645);
nand U10956 (N_10956,N_7375,N_8867);
nand U10957 (N_10957,N_8841,N_9863);
or U10958 (N_10958,N_7317,N_7358);
nand U10959 (N_10959,N_8404,N_6084);
nand U10960 (N_10960,N_9369,N_5037);
and U10961 (N_10961,N_6537,N_5436);
and U10962 (N_10962,N_6403,N_5812);
and U10963 (N_10963,N_7202,N_6755);
and U10964 (N_10964,N_5464,N_6976);
or U10965 (N_10965,N_5734,N_9519);
nand U10966 (N_10966,N_5941,N_5953);
nand U10967 (N_10967,N_9936,N_5864);
or U10968 (N_10968,N_6494,N_9951);
and U10969 (N_10969,N_5659,N_8913);
nand U10970 (N_10970,N_6773,N_6570);
and U10971 (N_10971,N_9495,N_7834);
nand U10972 (N_10972,N_7424,N_9215);
nand U10973 (N_10973,N_8395,N_6689);
or U10974 (N_10974,N_8358,N_8263);
xnor U10975 (N_10975,N_5042,N_8724);
nand U10976 (N_10976,N_8719,N_7740);
nand U10977 (N_10977,N_8095,N_6799);
or U10978 (N_10978,N_6164,N_7515);
xnor U10979 (N_10979,N_9775,N_9164);
or U10980 (N_10980,N_9329,N_7931);
nor U10981 (N_10981,N_7946,N_7173);
nor U10982 (N_10982,N_5889,N_6602);
nand U10983 (N_10983,N_9135,N_7190);
and U10984 (N_10984,N_6338,N_6393);
nand U10985 (N_10985,N_7774,N_8344);
or U10986 (N_10986,N_6984,N_9021);
or U10987 (N_10987,N_8726,N_5687);
nand U10988 (N_10988,N_5453,N_6087);
and U10989 (N_10989,N_5088,N_6116);
nor U10990 (N_10990,N_7015,N_9833);
nor U10991 (N_10991,N_7096,N_5981);
nor U10992 (N_10992,N_7091,N_8078);
nor U10993 (N_10993,N_9820,N_5934);
or U10994 (N_10994,N_8399,N_5491);
and U10995 (N_10995,N_7507,N_6866);
or U10996 (N_10996,N_5495,N_7073);
nor U10997 (N_10997,N_8028,N_7090);
nor U10998 (N_10998,N_9746,N_7599);
nand U10999 (N_10999,N_6372,N_7280);
xnor U11000 (N_11000,N_5609,N_5554);
nand U11001 (N_11001,N_9900,N_9336);
nor U11002 (N_11002,N_6618,N_6870);
nor U11003 (N_11003,N_9401,N_9526);
nor U11004 (N_11004,N_9154,N_6730);
and U11005 (N_11005,N_8982,N_9571);
nand U11006 (N_11006,N_5921,N_8454);
nand U11007 (N_11007,N_9323,N_7472);
nor U11008 (N_11008,N_5367,N_9308);
and U11009 (N_11009,N_7229,N_8116);
nand U11010 (N_11010,N_7029,N_8292);
or U11011 (N_11011,N_5430,N_7430);
nor U11012 (N_11012,N_9861,N_5410);
nand U11013 (N_11013,N_6985,N_5546);
or U11014 (N_11014,N_6037,N_8821);
and U11015 (N_11015,N_5423,N_5914);
nand U11016 (N_11016,N_7013,N_8832);
nand U11017 (N_11017,N_5773,N_7041);
and U11018 (N_11018,N_7374,N_6770);
and U11019 (N_11019,N_7607,N_5632);
nand U11020 (N_11020,N_9809,N_9073);
and U11021 (N_11021,N_9350,N_6263);
nand U11022 (N_11022,N_6287,N_7629);
xnor U11023 (N_11023,N_6861,N_9392);
xor U11024 (N_11024,N_9016,N_8105);
and U11025 (N_11025,N_5966,N_7905);
nand U11026 (N_11026,N_9171,N_8122);
nand U11027 (N_11027,N_9064,N_5076);
nand U11028 (N_11028,N_7631,N_6784);
and U11029 (N_11029,N_7147,N_5200);
nand U11030 (N_11030,N_8195,N_5398);
nor U11031 (N_11031,N_6688,N_6186);
nand U11032 (N_11032,N_5841,N_9719);
nor U11033 (N_11033,N_5280,N_7808);
nand U11034 (N_11034,N_7589,N_9455);
nand U11035 (N_11035,N_8602,N_6024);
xor U11036 (N_11036,N_5452,N_5815);
and U11037 (N_11037,N_6431,N_6748);
xnor U11038 (N_11038,N_6176,N_8676);
xor U11039 (N_11039,N_5470,N_8199);
nand U11040 (N_11040,N_9558,N_6783);
or U11041 (N_11041,N_8426,N_7639);
and U11042 (N_11042,N_7925,N_6354);
and U11043 (N_11043,N_8434,N_5307);
nor U11044 (N_11044,N_5666,N_8398);
or U11045 (N_11045,N_6058,N_8840);
nor U11046 (N_11046,N_8622,N_9948);
and U11047 (N_11047,N_9961,N_9747);
and U11048 (N_11048,N_9239,N_6805);
nor U11049 (N_11049,N_9669,N_9097);
or U11050 (N_11050,N_6699,N_6881);
and U11051 (N_11051,N_5939,N_9782);
or U11052 (N_11052,N_8125,N_6649);
nor U11053 (N_11053,N_9573,N_8894);
nor U11054 (N_11054,N_9736,N_9873);
nand U11055 (N_11055,N_6627,N_5281);
nor U11056 (N_11056,N_5866,N_7152);
nand U11057 (N_11057,N_7206,N_8249);
nor U11058 (N_11058,N_7313,N_5101);
nand U11059 (N_11059,N_5674,N_7256);
nand U11060 (N_11060,N_5933,N_9649);
nand U11061 (N_11061,N_9185,N_7841);
nor U11062 (N_11062,N_7832,N_5170);
nand U11063 (N_11063,N_6437,N_9457);
xnor U11064 (N_11064,N_8735,N_7602);
and U11065 (N_11065,N_7770,N_9872);
nand U11066 (N_11066,N_8008,N_7168);
nand U11067 (N_11067,N_9409,N_8674);
nand U11068 (N_11068,N_9196,N_5483);
xor U11069 (N_11069,N_6447,N_6693);
nand U11070 (N_11070,N_9619,N_5446);
nand U11071 (N_11071,N_7260,N_8197);
nand U11072 (N_11072,N_9510,N_5605);
nor U11073 (N_11073,N_5360,N_7499);
and U11074 (N_11074,N_8823,N_9301);
nand U11075 (N_11075,N_8574,N_5123);
nand U11076 (N_11076,N_8196,N_5129);
or U11077 (N_11077,N_5962,N_9960);
nor U11078 (N_11078,N_7109,N_7434);
or U11079 (N_11079,N_9005,N_8766);
nand U11080 (N_11080,N_9072,N_6471);
nand U11081 (N_11081,N_6488,N_6860);
and U11082 (N_11082,N_7040,N_8422);
or U11083 (N_11083,N_6487,N_8825);
xnor U11084 (N_11084,N_8540,N_5095);
nor U11085 (N_11085,N_5948,N_9563);
nor U11086 (N_11086,N_5402,N_5625);
nor U11087 (N_11087,N_5935,N_5867);
nand U11088 (N_11088,N_6584,N_9165);
nand U11089 (N_11089,N_6347,N_6392);
nand U11090 (N_11090,N_6489,N_5822);
and U11091 (N_11091,N_6820,N_6072);
nand U11092 (N_11092,N_8201,N_5432);
and U11093 (N_11093,N_9316,N_5433);
and U11094 (N_11094,N_6398,N_6442);
nor U11095 (N_11095,N_8866,N_5955);
xnor U11096 (N_11096,N_8837,N_5293);
or U11097 (N_11097,N_6154,N_5968);
and U11098 (N_11098,N_6882,N_9837);
nand U11099 (N_11099,N_7053,N_7005);
or U11100 (N_11100,N_7908,N_6564);
and U11101 (N_11101,N_7104,N_9348);
and U11102 (N_11102,N_5463,N_7574);
nand U11103 (N_11103,N_5485,N_9059);
nand U11104 (N_11104,N_8224,N_7900);
or U11105 (N_11105,N_9907,N_9564);
nand U11106 (N_11106,N_8006,N_6031);
and U11107 (N_11107,N_8862,N_8500);
nand U11108 (N_11108,N_5202,N_7999);
and U11109 (N_11109,N_5670,N_8583);
or U11110 (N_11110,N_9741,N_8462);
or U11111 (N_11111,N_9253,N_8431);
xor U11112 (N_11112,N_8774,N_8419);
nor U11113 (N_11113,N_8679,N_7600);
nand U11114 (N_11114,N_8180,N_9217);
nor U11115 (N_11115,N_9678,N_8409);
or U11116 (N_11116,N_8932,N_7752);
nor U11117 (N_11117,N_6578,N_5620);
nor U11118 (N_11118,N_7610,N_9418);
nor U11119 (N_11119,N_6548,N_8061);
and U11120 (N_11120,N_8253,N_5997);
nor U11121 (N_11121,N_6374,N_8740);
nor U11122 (N_11122,N_6691,N_9269);
nand U11123 (N_11123,N_9984,N_7223);
nand U11124 (N_11124,N_5723,N_9625);
or U11125 (N_11125,N_8613,N_6621);
nor U11126 (N_11126,N_5942,N_9380);
xor U11127 (N_11127,N_6125,N_9511);
nor U11128 (N_11128,N_9309,N_8585);
and U11129 (N_11129,N_7216,N_7189);
and U11130 (N_11130,N_7057,N_7448);
nor U11131 (N_11131,N_7371,N_6194);
or U11132 (N_11132,N_9403,N_7332);
nand U11133 (N_11133,N_7244,N_5741);
or U11134 (N_11134,N_7614,N_6462);
nand U11135 (N_11135,N_8682,N_9705);
nor U11136 (N_11136,N_8346,N_8427);
or U11137 (N_11137,N_7820,N_9275);
or U11138 (N_11138,N_7363,N_8941);
nand U11139 (N_11139,N_7329,N_8484);
xor U11140 (N_11140,N_6229,N_6806);
and U11141 (N_11141,N_5011,N_8502);
nand U11142 (N_11142,N_8627,N_5267);
nand U11143 (N_11143,N_9987,N_5309);
nand U11144 (N_11144,N_8353,N_8302);
and U11145 (N_11145,N_5535,N_7379);
nand U11146 (N_11146,N_8134,N_6033);
nand U11147 (N_11147,N_8788,N_6104);
nor U11148 (N_11148,N_6936,N_6486);
nand U11149 (N_11149,N_9227,N_5593);
or U11150 (N_11150,N_6332,N_5269);
or U11151 (N_11151,N_6771,N_7576);
nand U11152 (N_11152,N_8706,N_7184);
or U11153 (N_11153,N_6849,N_8577);
or U11154 (N_11154,N_6387,N_5696);
nor U11155 (N_11155,N_9462,N_6530);
and U11156 (N_11156,N_5662,N_9259);
or U11157 (N_11157,N_9004,N_9435);
nor U11158 (N_11158,N_9295,N_6433);
xor U11159 (N_11159,N_9902,N_8780);
xnor U11160 (N_11160,N_6209,N_7038);
nand U11161 (N_11161,N_7153,N_7006);
or U11162 (N_11162,N_9635,N_6640);
nor U11163 (N_11163,N_8520,N_6585);
or U11164 (N_11164,N_5005,N_8275);
nor U11165 (N_11165,N_9530,N_5726);
or U11166 (N_11166,N_7510,N_8711);
nand U11167 (N_11167,N_7274,N_5752);
and U11168 (N_11168,N_5695,N_6280);
xor U11169 (N_11169,N_5652,N_7286);
and U11170 (N_11170,N_5982,N_5624);
xor U11171 (N_11171,N_9735,N_5162);
nand U11172 (N_11172,N_6563,N_6015);
nand U11173 (N_11173,N_7968,N_5925);
nand U11174 (N_11174,N_9855,N_5875);
nand U11175 (N_11175,N_5498,N_7194);
or U11176 (N_11176,N_9424,N_6142);
xor U11177 (N_11177,N_8954,N_7906);
nor U11178 (N_11178,N_6652,N_9932);
and U11179 (N_11179,N_8991,N_6275);
or U11180 (N_11180,N_8362,N_7390);
nor U11181 (N_11181,N_8786,N_5496);
and U11182 (N_11182,N_7222,N_9950);
or U11183 (N_11183,N_6032,N_8505);
and U11184 (N_11184,N_8560,N_9200);
nand U11185 (N_11185,N_9598,N_7210);
or U11186 (N_11186,N_6168,N_9120);
xnor U11187 (N_11187,N_9565,N_9030);
and U11188 (N_11188,N_9531,N_7739);
and U11189 (N_11189,N_9102,N_9300);
or U11190 (N_11190,N_7106,N_5880);
and U11191 (N_11191,N_8839,N_9224);
xnor U11192 (N_11192,N_8696,N_5406);
or U11193 (N_11193,N_9047,N_5836);
nor U11194 (N_11194,N_8618,N_6656);
or U11195 (N_11195,N_9296,N_9981);
nand U11196 (N_11196,N_8912,N_9921);
nand U11197 (N_11197,N_7012,N_9176);
nor U11198 (N_11198,N_6059,N_9074);
and U11199 (N_11199,N_8537,N_5878);
and U11200 (N_11200,N_6219,N_6975);
nand U11201 (N_11201,N_5080,N_7741);
xor U11202 (N_11202,N_6350,N_7836);
and U11203 (N_11203,N_6359,N_6150);
nand U11204 (N_11204,N_9116,N_9941);
nor U11205 (N_11205,N_9998,N_6847);
xnor U11206 (N_11206,N_7416,N_6238);
nand U11207 (N_11207,N_6800,N_6348);
nand U11208 (N_11208,N_6346,N_7160);
nor U11209 (N_11209,N_6324,N_8343);
nor U11210 (N_11210,N_9351,N_9645);
and U11211 (N_11211,N_9118,N_7822);
nor U11212 (N_11212,N_7017,N_9289);
or U11213 (N_11213,N_7226,N_8471);
and U11214 (N_11214,N_9156,N_8685);
nor U11215 (N_11215,N_6883,N_9958);
nor U11216 (N_11216,N_6056,N_6958);
or U11217 (N_11217,N_7477,N_5132);
nand U11218 (N_11218,N_5157,N_5126);
nand U11219 (N_11219,N_6182,N_5686);
nor U11220 (N_11220,N_9208,N_9529);
and U11221 (N_11221,N_8121,N_8384);
or U11222 (N_11222,N_9129,N_6423);
and U11223 (N_11223,N_6278,N_9699);
nor U11224 (N_11224,N_9971,N_5909);
nor U11225 (N_11225,N_7533,N_8338);
and U11226 (N_11226,N_7627,N_9898);
or U11227 (N_11227,N_8139,N_8232);
nor U11228 (N_11228,N_8910,N_9753);
xnor U11229 (N_11229,N_5118,N_8868);
nor U11230 (N_11230,N_9691,N_9049);
nor U11231 (N_11231,N_6794,N_6026);
nor U11232 (N_11232,N_8564,N_5524);
or U11233 (N_11233,N_8984,N_6198);
nor U11234 (N_11234,N_9553,N_8713);
and U11235 (N_11235,N_7605,N_5897);
nor U11236 (N_11236,N_8903,N_7177);
nor U11237 (N_11237,N_7827,N_7595);
or U11238 (N_11238,N_5416,N_5214);
xnor U11239 (N_11239,N_8254,N_9575);
xnor U11240 (N_11240,N_8950,N_5359);
nor U11241 (N_11241,N_8994,N_6013);
nor U11242 (N_11242,N_6573,N_6358);
nand U11243 (N_11243,N_6885,N_7183);
or U11244 (N_11244,N_8664,N_5212);
nor U11245 (N_11245,N_9778,N_9231);
nand U11246 (N_11246,N_8072,N_6569);
or U11247 (N_11247,N_5487,N_5998);
and U11248 (N_11248,N_9009,N_8155);
and U11249 (N_11249,N_5460,N_5537);
nor U11250 (N_11250,N_6854,N_9538);
nor U11251 (N_11251,N_5421,N_6761);
or U11252 (N_11252,N_8745,N_9431);
nor U11253 (N_11253,N_8663,N_9256);
nand U11254 (N_11254,N_9483,N_9248);
xnor U11255 (N_11255,N_6741,N_5762);
or U11256 (N_11256,N_5265,N_5468);
or U11257 (N_11257,N_5320,N_6175);
xnor U11258 (N_11258,N_5138,N_7693);
or U11259 (N_11259,N_6746,N_7887);
and U11260 (N_11260,N_8141,N_5853);
nor U11261 (N_11261,N_7910,N_8795);
nor U11262 (N_11262,N_9033,N_5391);
xnor U11263 (N_11263,N_5617,N_8282);
or U11264 (N_11264,N_7211,N_5606);
nor U11265 (N_11265,N_9124,N_9311);
xnor U11266 (N_11266,N_6595,N_9555);
or U11267 (N_11267,N_9057,N_9915);
or U11268 (N_11268,N_7257,N_8808);
and U11269 (N_11269,N_6178,N_9660);
nand U11270 (N_11270,N_8953,N_7008);
nor U11271 (N_11271,N_8491,N_7064);
and U11272 (N_11272,N_8185,N_7107);
nor U11273 (N_11273,N_5232,N_9994);
or U11274 (N_11274,N_7666,N_6901);
or U11275 (N_11275,N_5396,N_5805);
nor U11276 (N_11276,N_5754,N_7077);
or U11277 (N_11277,N_7316,N_6567);
nor U11278 (N_11278,N_5354,N_6440);
or U11279 (N_11279,N_8211,N_8288);
nor U11280 (N_11280,N_7986,N_5932);
or U11281 (N_11281,N_5944,N_7480);
nand U11282 (N_11282,N_6839,N_9292);
and U11283 (N_11283,N_7120,N_8177);
nand U11284 (N_11284,N_9000,N_6039);
or U11285 (N_11285,N_6477,N_6067);
and U11286 (N_11286,N_8171,N_9490);
and U11287 (N_11287,N_9646,N_6394);
and U11288 (N_11288,N_5467,N_6169);
nor U11289 (N_11289,N_5036,N_7729);
or U11290 (N_11290,N_5392,N_9897);
or U11291 (N_11291,N_6258,N_6791);
xnor U11292 (N_11292,N_9878,N_6038);
xor U11293 (N_11293,N_8230,N_6908);
and U11294 (N_11294,N_8529,N_6753);
and U11295 (N_11295,N_7369,N_7603);
and U11296 (N_11296,N_5693,N_6291);
nand U11297 (N_11297,N_6889,N_7314);
and U11298 (N_11298,N_8957,N_6476);
and U11299 (N_11299,N_7484,N_6267);
nand U11300 (N_11300,N_7662,N_9002);
xor U11301 (N_11301,N_8023,N_8106);
nor U11302 (N_11302,N_7069,N_5571);
and U11303 (N_11303,N_6245,N_7279);
nand U11304 (N_11304,N_7349,N_5870);
nor U11305 (N_11305,N_8783,N_6817);
xor U11306 (N_11306,N_9125,N_8985);
and U11307 (N_11307,N_5725,N_9440);
and U11308 (N_11308,N_6485,N_9485);
nor U11309 (N_11309,N_7205,N_7727);
nor U11310 (N_11310,N_6172,N_5208);
nand U11311 (N_11311,N_9840,N_9622);
and U11312 (N_11312,N_5484,N_5911);
and U11313 (N_11313,N_8649,N_7847);
xor U11314 (N_11314,N_5477,N_7753);
nand U11315 (N_11315,N_7118,N_9964);
or U11316 (N_11316,N_5065,N_5844);
and U11317 (N_11317,N_6774,N_8152);
nor U11318 (N_11318,N_9258,N_6710);
or U11319 (N_11319,N_5952,N_8922);
and U11320 (N_11320,N_8653,N_5246);
xnor U11321 (N_11321,N_8824,N_5928);
or U11322 (N_11322,N_6719,N_7990);
nand U11323 (N_11323,N_9201,N_5951);
xor U11324 (N_11324,N_9596,N_8279);
nor U11325 (N_11325,N_7101,N_6735);
or U11326 (N_11326,N_9286,N_9597);
or U11327 (N_11327,N_9695,N_5827);
and U11328 (N_11328,N_7391,N_6534);
or U11329 (N_11329,N_6478,N_7503);
and U11330 (N_11330,N_6904,N_8421);
nor U11331 (N_11331,N_9082,N_5394);
and U11332 (N_11332,N_6520,N_9068);
nand U11333 (N_11333,N_8865,N_7273);
and U11334 (N_11334,N_9103,N_9534);
or U11335 (N_11335,N_7203,N_5749);
and U11336 (N_11336,N_6512,N_5032);
nor U11337 (N_11337,N_9942,N_6619);
nand U11338 (N_11338,N_5847,N_9831);
xnor U11339 (N_11339,N_6021,N_8198);
xnor U11340 (N_11340,N_7934,N_5182);
or U11341 (N_11341,N_6264,N_8524);
or U11342 (N_11342,N_8508,N_7408);
or U11343 (N_11343,N_6825,N_6266);
xor U11344 (N_11344,N_5374,N_7547);
or U11345 (N_11345,N_5898,N_7538);
and U11346 (N_11346,N_8947,N_6063);
xor U11347 (N_11347,N_9395,N_7519);
nand U11348 (N_11348,N_6391,N_7301);
nand U11349 (N_11349,N_9476,N_9687);
nor U11350 (N_11350,N_6891,N_5224);
xnor U11351 (N_11351,N_8963,N_8644);
and U11352 (N_11352,N_6098,N_5971);
or U11353 (N_11353,N_5028,N_7911);
nor U11354 (N_11354,N_6014,N_9626);
and U11355 (N_11355,N_9469,N_5057);
nor U11356 (N_11356,N_6000,N_7463);
nand U11357 (N_11357,N_8764,N_9487);
and U11358 (N_11358,N_8883,N_5518);
or U11359 (N_11359,N_8020,N_8481);
and U11360 (N_11360,N_6467,N_7636);
nand U11361 (N_11361,N_6736,N_7743);
xnor U11362 (N_11362,N_8109,N_8571);
nor U11363 (N_11363,N_8239,N_8819);
nand U11364 (N_11364,N_8590,N_6814);
and U11365 (N_11365,N_6344,N_8140);
xor U11366 (N_11366,N_9211,N_5343);
and U11367 (N_11367,N_8450,N_5976);
and U11368 (N_11368,N_5479,N_5490);
or U11369 (N_11369,N_5771,N_6167);
or U11370 (N_11370,N_7264,N_8659);
nand U11371 (N_11371,N_8161,N_8389);
or U11372 (N_11372,N_6076,N_6365);
and U11373 (N_11373,N_9797,N_6044);
nand U11374 (N_11374,N_5201,N_8624);
nor U11375 (N_11375,N_6992,N_7789);
nor U11376 (N_11376,N_5156,N_6134);
and U11377 (N_11377,N_5788,N_5513);
and U11378 (N_11378,N_7929,N_8079);
and U11379 (N_11379,N_9633,N_7241);
nand U11380 (N_11380,N_8781,N_5551);
and U11381 (N_11381,N_9568,N_6424);
or U11382 (N_11382,N_9204,N_5675);
nand U11383 (N_11383,N_7746,N_6288);
nor U11384 (N_11384,N_9965,N_9721);
or U11385 (N_11385,N_5141,N_8632);
nor U11386 (N_11386,N_6158,N_7518);
or U11387 (N_11387,N_6333,N_7128);
nand U11388 (N_11388,N_7142,N_6586);
or U11389 (N_11389,N_8712,N_9052);
nand U11390 (N_11390,N_6380,N_9218);
and U11391 (N_11391,N_7511,N_8436);
and U11392 (N_11392,N_8654,N_8610);
xor U11393 (N_11393,N_5581,N_5732);
nor U11394 (N_11394,N_8872,N_8494);
nand U11395 (N_11395,N_9847,N_5497);
or U11396 (N_11396,N_6070,N_9434);
xnor U11397 (N_11397,N_7859,N_7889);
or U11398 (N_11398,N_7721,N_6554);
nor U11399 (N_11399,N_9038,N_7514);
nor U11400 (N_11400,N_5716,N_8558);
xor U11401 (N_11401,N_7161,N_9240);
and U11402 (N_11402,N_5001,N_7787);
nor U11403 (N_11403,N_5701,N_8852);
nand U11404 (N_11404,N_7717,N_7251);
nand U11405 (N_11405,N_9814,N_9454);
nor U11406 (N_11406,N_5448,N_7845);
and U11407 (N_11407,N_9887,N_9042);
nor U11408 (N_11408,N_6758,N_6310);
or U11409 (N_11409,N_6152,N_6053);
and U11410 (N_11410,N_8828,N_8415);
xor U11411 (N_11411,N_6493,N_9341);
or U11412 (N_11412,N_6831,N_8851);
or U11413 (N_11413,N_7641,N_6151);
nand U11414 (N_11414,N_6279,N_6202);
and U11415 (N_11415,N_9653,N_5242);
nor U11416 (N_11416,N_8567,N_7788);
nor U11417 (N_11417,N_5506,N_6877);
xnor U11418 (N_11418,N_5213,N_5151);
and U11419 (N_11419,N_7551,N_9011);
xor U11420 (N_11420,N_9537,N_9605);
nor U11421 (N_11421,N_5459,N_7965);
xnor U11422 (N_11422,N_7067,N_6228);
or U11423 (N_11423,N_8729,N_7097);
xnor U11424 (N_11424,N_5679,N_5801);
and U11425 (N_11425,N_6295,N_7074);
or U11426 (N_11426,N_7347,N_7182);
and U11427 (N_11427,N_7877,N_6010);
and U11428 (N_11428,N_9397,N_5772);
or U11429 (N_11429,N_9268,N_9077);
or U11430 (N_11430,N_8043,N_8385);
and U11431 (N_11431,N_6722,N_8751);
and U11432 (N_11432,N_5640,N_5418);
or U11433 (N_11433,N_7056,N_9899);
nor U11434 (N_11434,N_9895,N_9679);
nor U11435 (N_11435,N_5069,N_9638);
or U11436 (N_11436,N_6138,N_9168);
or U11437 (N_11437,N_7664,N_5759);
nor U11438 (N_11438,N_6193,N_8370);
nor U11439 (N_11439,N_8204,N_5205);
or U11440 (N_11440,N_8902,N_7559);
nor U11441 (N_11441,N_7284,N_5840);
nand U11442 (N_11442,N_8730,N_9554);
and U11443 (N_11443,N_5699,N_6756);
nand U11444 (N_11444,N_9668,N_7247);
nand U11445 (N_11445,N_9821,N_8381);
or U11446 (N_11446,N_5389,N_7520);
nand U11447 (N_11447,N_7898,N_5178);
nand U11448 (N_11448,N_7457,N_9024);
xnor U11449 (N_11449,N_8364,N_5417);
and U11450 (N_11450,N_6608,N_6821);
and U11451 (N_11451,N_5310,N_7026);
and U11452 (N_11452,N_6991,N_5689);
nand U11453 (N_11453,N_5907,N_6429);
nand U11454 (N_11454,N_7467,N_5525);
nor U11455 (N_11455,N_6527,N_8612);
xor U11456 (N_11456,N_5735,N_5155);
nor U11457 (N_11457,N_6474,N_6135);
or U11458 (N_11458,N_6835,N_6094);
nand U11459 (N_11459,N_8308,N_8578);
and U11460 (N_11460,N_5781,N_9867);
nand U11461 (N_11461,N_5501,N_7059);
nand U11462 (N_11462,N_9297,N_8725);
or U11463 (N_11463,N_8884,N_6633);
and U11464 (N_11464,N_7469,N_5588);
and U11465 (N_11465,N_7591,N_7068);
or U11466 (N_11466,N_9365,N_5704);
and U11467 (N_11467,N_5508,N_5650);
or U11468 (N_11468,N_9151,N_6834);
nand U11469 (N_11469,N_7426,N_9533);
xnor U11470 (N_11470,N_7590,N_5767);
and U11471 (N_11471,N_9966,N_5886);
and U11472 (N_11472,N_9391,N_9242);
nor U11473 (N_11473,N_8636,N_5645);
nand U11474 (N_11474,N_7213,N_5308);
or U11475 (N_11475,N_6389,N_7490);
and U11476 (N_11476,N_9841,N_9617);
nand U11477 (N_11477,N_8551,N_8629);
nand U11478 (N_11478,N_7114,N_6430);
and U11479 (N_11479,N_7037,N_6130);
and U11480 (N_11480,N_9798,N_6988);
xor U11481 (N_11481,N_9723,N_6536);
nand U11482 (N_11482,N_8429,N_7354);
nand U11483 (N_11483,N_9055,N_8877);
nand U11484 (N_11484,N_5311,N_7586);
and U11485 (N_11485,N_7265,N_5461);
nor U11486 (N_11486,N_7021,N_7352);
or U11487 (N_11487,N_6989,N_7456);
and U11488 (N_11488,N_9967,N_8797);
and U11489 (N_11489,N_5099,N_9642);
nand U11490 (N_11490,N_7045,N_8639);
nand U11491 (N_11491,N_9813,N_5829);
or U11492 (N_11492,N_6963,N_8238);
nand U11493 (N_11493,N_6277,N_5671);
and U11494 (N_11494,N_9331,N_8704);
or U11495 (N_11495,N_7953,N_5816);
nand U11496 (N_11496,N_5673,N_8087);
or U11497 (N_11497,N_9822,N_9175);
nand U11498 (N_11498,N_8623,N_8692);
xor U11499 (N_11499,N_6322,N_8646);
nand U11500 (N_11500,N_9184,N_6082);
nor U11501 (N_11501,N_8314,N_5618);
nor U11502 (N_11502,N_9864,N_5270);
and U11503 (N_11503,N_7648,N_5629);
or U11504 (N_11504,N_7294,N_6221);
nor U11505 (N_11505,N_8925,N_6162);
nor U11506 (N_11506,N_9569,N_6660);
and U11507 (N_11507,N_8408,N_8112);
nor U11508 (N_11508,N_8424,N_8701);
and U11509 (N_11509,N_6645,N_7454);
nor U11510 (N_11510,N_9067,N_7793);
and U11511 (N_11511,N_6441,N_7497);
nand U11512 (N_11512,N_8672,N_5050);
nand U11513 (N_11513,N_8569,N_5458);
or U11514 (N_11514,N_6395,N_8013);
nand U11515 (N_11515,N_6271,N_9789);
nand U11516 (N_11516,N_6444,N_6066);
xor U11517 (N_11517,N_7355,N_5075);
or U11518 (N_11518,N_5712,N_5131);
nor U11519 (N_11519,N_8119,N_5473);
or U11520 (N_11520,N_8045,N_8170);
nand U11521 (N_11521,N_8526,N_5223);
nor U11522 (N_11522,N_7692,N_6147);
nand U11523 (N_11523,N_6262,N_8549);
xnor U11524 (N_11524,N_7892,N_7584);
nor U11525 (N_11525,N_5991,N_6185);
or U11526 (N_11526,N_6700,N_8595);
and U11527 (N_11527,N_5505,N_7882);
and U11528 (N_11528,N_6676,N_5855);
or U11529 (N_11529,N_6055,N_6995);
or U11530 (N_11530,N_5596,N_6808);
nor U11531 (N_11531,N_6192,N_9927);
and U11532 (N_11532,N_5109,N_7156);
xnor U11533 (N_11533,N_8929,N_6727);
nor U11534 (N_11534,N_8303,N_8442);
and U11535 (N_11535,N_7851,N_5985);
nand U11536 (N_11536,N_9460,N_7164);
or U11537 (N_11537,N_9095,N_8160);
nor U11538 (N_11538,N_9443,N_8075);
or U11539 (N_11539,N_7977,N_8510);
and U11540 (N_11540,N_6137,N_8966);
and U11541 (N_11541,N_6750,N_9880);
xor U11542 (N_11542,N_6970,N_5920);
or U11543 (N_11543,N_5742,N_6075);
nand U11544 (N_11544,N_8859,N_6819);
or U11545 (N_11545,N_9430,N_7722);
or U11546 (N_11546,N_6524,N_9923);
nand U11547 (N_11547,N_7002,N_7255);
xor U11548 (N_11548,N_7253,N_8312);
nand U11549 (N_11549,N_5302,N_7907);
nand U11550 (N_11550,N_9446,N_7732);
and U11551 (N_11551,N_7236,N_5039);
and U11552 (N_11552,N_8264,N_5390);
nand U11553 (N_11553,N_7491,N_8413);
and U11554 (N_11554,N_6336,N_6335);
and U11555 (N_11555,N_8014,N_7445);
and U11556 (N_11556,N_8348,N_9845);
xnor U11557 (N_11557,N_8758,N_6246);
or U11558 (N_11558,N_8099,N_9578);
or U11559 (N_11559,N_8716,N_7420);
nand U11560 (N_11560,N_9013,N_6426);
or U11561 (N_11561,N_5797,N_6971);
nand U11562 (N_11562,N_9419,N_6740);
nand U11563 (N_11563,N_6490,N_8223);
or U11564 (N_11564,N_7661,N_7824);
nor U11565 (N_11565,N_8296,N_8246);
nor U11566 (N_11566,N_9382,N_8166);
xnor U11567 (N_11567,N_8515,N_6651);
nand U11568 (N_11568,N_5765,N_5614);
or U11569 (N_11569,N_6248,N_8718);
and U11570 (N_11570,N_6034,N_6631);
nand U11571 (N_11571,N_8562,N_5375);
nand U11572 (N_11572,N_9946,N_9158);
nand U11573 (N_11573,N_9701,N_8496);
and U11574 (N_11574,N_6863,N_9098);
nor U11575 (N_11575,N_9710,N_8695);
nor U11576 (N_11576,N_7628,N_6680);
nand U11577 (N_11577,N_8886,N_7552);
nor U11578 (N_11578,N_9737,N_8816);
nand U11579 (N_11579,N_5161,N_7855);
and U11580 (N_11580,N_6591,N_7609);
xor U11581 (N_11581,N_5315,N_8115);
nand U11582 (N_11582,N_8756,N_9062);
or U11583 (N_11583,N_5097,N_7951);
nor U11584 (N_11584,N_6133,N_7172);
or U11585 (N_11585,N_8543,N_6119);
or U11586 (N_11586,N_5782,N_8138);
xnor U11587 (N_11587,N_7556,N_6801);
or U11588 (N_11588,N_8873,N_9328);
nand U11589 (N_11589,N_9357,N_5031);
and U11590 (N_11590,N_5426,N_7055);
nor U11591 (N_11591,N_9160,N_7993);
nand U11592 (N_11592,N_6503,N_5561);
nand U11593 (N_11593,N_6658,N_8208);
nand U11594 (N_11594,N_6840,N_5891);
and U11595 (N_11595,N_5356,N_7444);
nor U11596 (N_11596,N_5574,N_5758);
and U11597 (N_11597,N_7460,N_9786);
and U11598 (N_11598,N_7119,N_5148);
or U11599 (N_11599,N_9416,N_9658);
or U11600 (N_11600,N_7536,N_8593);
nor U11601 (N_11601,N_5365,N_5279);
or U11602 (N_11602,N_8748,N_6996);
or U11603 (N_11603,N_8124,N_9698);
nand U11604 (N_11604,N_8887,N_7356);
or U11605 (N_11605,N_7421,N_6464);
or U11606 (N_11606,N_8280,N_9096);
nand U11607 (N_11607,N_5555,N_7525);
nand U11608 (N_11608,N_6964,N_9805);
or U11609 (N_11609,N_7768,N_6438);
and U11610 (N_11610,N_7996,N_6707);
and U11611 (N_11611,N_5839,N_9772);
or U11612 (N_11612,N_5539,N_9917);
or U11613 (N_11613,N_5321,N_5724);
and U11614 (N_11614,N_9850,N_9648);
xor U11615 (N_11615,N_7134,N_5009);
nor U11616 (N_11616,N_8291,N_5969);
nor U11617 (N_11617,N_9144,N_5403);
nor U11618 (N_11618,N_7991,N_9400);
and U11619 (N_11619,N_6237,N_9354);
or U11620 (N_11620,N_6625,N_8643);
nor U11621 (N_11621,N_7779,N_8327);
nor U11622 (N_11622,N_8439,N_9058);
nor U11623 (N_11623,N_6521,N_5604);
nand U11624 (N_11624,N_8931,N_5861);
nor U11625 (N_11625,N_6049,N_6180);
xnor U11626 (N_11626,N_9557,N_5220);
and U11627 (N_11627,N_5045,N_6227);
xor U11628 (N_11628,N_6692,N_6894);
nand U11629 (N_11629,N_7581,N_7088);
nor U11630 (N_11630,N_7089,N_8256);
or U11631 (N_11631,N_9599,N_6212);
nand U11632 (N_11632,N_6373,N_7252);
or U11633 (N_11633,N_7366,N_6355);
and U11634 (N_11634,N_9804,N_6987);
xnor U11635 (N_11635,N_6923,N_6529);
nor U11636 (N_11636,N_6952,N_7162);
nor U11637 (N_11637,N_7885,N_5573);
and U11638 (N_11638,N_6005,N_5061);
or U11639 (N_11639,N_7025,N_5326);
or U11640 (N_11640,N_8267,N_7745);
or U11641 (N_11641,N_7751,N_6043);
or U11642 (N_11642,N_6592,N_9760);
and U11643 (N_11643,N_7365,N_6611);
nor U11644 (N_11644,N_5677,N_9132);
or U11645 (N_11645,N_9346,N_9285);
nand U11646 (N_11646,N_5147,N_8658);
nor U11647 (N_11647,N_6781,N_7367);
and U11648 (N_11648,N_8214,N_5012);
and U11649 (N_11649,N_6999,N_6370);
nand U11650 (N_11650,N_9983,N_6061);
xor U11651 (N_11651,N_9832,N_7790);
and U11652 (N_11652,N_6959,N_9676);
xor U11653 (N_11653,N_9383,N_8368);
nor U11654 (N_11654,N_9054,N_8539);
xor U11655 (N_11655,N_9244,N_8363);
nand U11656 (N_11656,N_7971,N_9656);
xor U11657 (N_11657,N_7185,N_6875);
and U11658 (N_11658,N_9752,N_6898);
and U11659 (N_11659,N_9017,N_7647);
or U11660 (N_11660,N_7764,N_5313);
and U11661 (N_11661,N_8322,N_9586);
or U11662 (N_11662,N_9784,N_7478);
nand U11663 (N_11663,N_5627,N_8114);
nor U11664 (N_11664,N_8096,N_9138);
nand U11665 (N_11665,N_7239,N_8989);
xor U11666 (N_11666,N_5387,N_9764);
nor U11667 (N_11667,N_7115,N_7419);
nand U11668 (N_11668,N_8443,N_6143);
nand U11669 (N_11669,N_5413,N_7819);
or U11670 (N_11670,N_6539,N_6325);
nand U11671 (N_11671,N_8382,N_9153);
nor U11672 (N_11672,N_7840,N_6230);
nor U11673 (N_11673,N_9041,N_7325);
and U11674 (N_11674,N_8458,N_6844);
and U11675 (N_11675,N_5811,N_5442);
and U11676 (N_11676,N_6009,N_7588);
and U11677 (N_11677,N_9481,N_9504);
xnor U11678 (N_11678,N_7839,N_8945);
nor U11679 (N_11679,N_8815,N_8833);
or U11680 (N_11680,N_8983,N_9606);
or U11681 (N_11681,N_7802,N_6945);
nand U11682 (N_11682,N_8383,N_9795);
or U11683 (N_11683,N_8572,N_6772);
xnor U11684 (N_11684,N_8016,N_6737);
xnor U11685 (N_11685,N_7345,N_7063);
and U11686 (N_11686,N_8076,N_5690);
nor U11687 (N_11687,N_5238,N_8330);
xnor U11688 (N_11688,N_6967,N_8234);
and U11689 (N_11689,N_9374,N_6052);
nor U11690 (N_11690,N_8243,N_6100);
nand U11691 (N_11691,N_8209,N_9492);
and U11692 (N_11692,N_9091,N_8265);
nor U11693 (N_11693,N_7461,N_7544);
nand U11694 (N_11694,N_9257,N_5357);
and U11695 (N_11695,N_9616,N_5818);
nor U11696 (N_11696,N_7272,N_9697);
or U11697 (N_11697,N_6446,N_6184);
or U11698 (N_11698,N_5517,N_6081);
xor U11699 (N_11699,N_5400,N_5543);
or U11700 (N_11700,N_7966,N_5936);
or U11701 (N_11701,N_7023,N_5062);
nor U11702 (N_11702,N_8933,N_9920);
nor U11703 (N_11703,N_9167,N_9338);
xor U11704 (N_11704,N_8412,N_8127);
nand U11705 (N_11705,N_6981,N_7795);
nand U11706 (N_11706,N_5510,N_7320);
or U11707 (N_11707,N_7506,N_6402);
and U11708 (N_11708,N_5567,N_6822);
or U11709 (N_11709,N_9205,N_9766);
nor U11710 (N_11710,N_5245,N_7321);
nor U11711 (N_11711,N_7318,N_9307);
nand U11712 (N_11712,N_6156,N_5739);
or U11713 (N_11713,N_5288,N_8437);
nand U11714 (N_11714,N_6903,N_6690);
or U11715 (N_11715,N_9356,N_8796);
nor U11716 (N_11716,N_8702,N_8432);
nor U11717 (N_11717,N_6900,N_7051);
xnor U11718 (N_11718,N_8638,N_5651);
or U11719 (N_11719,N_6666,N_5750);
nand U11720 (N_11720,N_9838,N_7437);
nor U11721 (N_11721,N_6191,N_6091);
or U11722 (N_11722,N_8162,N_8563);
or U11723 (N_11723,N_9757,N_6360);
nand U11724 (N_11724,N_5711,N_9869);
nand U11725 (N_11725,N_8447,N_5475);
nand U11726 (N_11726,N_9467,N_6282);
nor U11727 (N_11727,N_7659,N_8668);
xor U11728 (N_11728,N_6400,N_5705);
xnor U11729 (N_11729,N_7433,N_6102);
nand U11730 (N_11730,N_5779,N_7402);
and U11731 (N_11731,N_7530,N_5144);
xnor U11732 (N_11732,N_8146,N_8186);
nand U11733 (N_11733,N_6042,N_9349);
and U11734 (N_11734,N_9589,N_8438);
xor U11735 (N_11735,N_7488,N_7141);
nand U11736 (N_11736,N_6878,N_8149);
nor U11737 (N_11737,N_8063,N_7879);
nand U11738 (N_11738,N_5722,N_8420);
nand U11739 (N_11739,N_8830,N_7543);
nor U11740 (N_11740,N_8575,N_8182);
xnor U11741 (N_11741,N_5250,N_7956);
nand U11742 (N_11742,N_5821,N_8000);
nand U11743 (N_11743,N_7166,N_9680);
or U11744 (N_11744,N_5512,N_5289);
or U11745 (N_11745,N_6826,N_8015);
nor U11746 (N_11746,N_9889,N_7754);
nand U11747 (N_11747,N_7380,N_8216);
nand U11748 (N_11748,N_7108,N_8506);
or U11749 (N_11749,N_8151,N_7436);
nand U11750 (N_11750,N_8241,N_9372);
nand U11751 (N_11751,N_9874,N_9406);
nor U11752 (N_11752,N_9496,N_5177);
nand U11753 (N_11753,N_5210,N_9161);
nor U11754 (N_11754,N_6702,N_9003);
nand U11755 (N_11755,N_7014,N_9559);
and U11756 (N_11756,N_7838,N_6944);
nor U11757 (N_11757,N_8192,N_9367);
nand U11758 (N_11758,N_9928,N_8518);
and U11759 (N_11759,N_7319,N_7583);
xnor U11760 (N_11760,N_7231,N_6568);
nand U11761 (N_11761,N_8619,N_6939);
and U11762 (N_11762,N_6811,N_7200);
nor U11763 (N_11763,N_6139,N_9115);
nor U11764 (N_11764,N_6762,N_6323);
xnor U11765 (N_11765,N_9940,N_5462);
nand U11766 (N_11766,N_8753,N_7935);
xor U11767 (N_11767,N_6233,N_6543);
or U11768 (N_11768,N_5290,N_7955);
and U11769 (N_11769,N_9337,N_9066);
nand U11770 (N_11770,N_5299,N_5022);
and U11771 (N_11771,N_5323,N_9768);
or U11772 (N_11772,N_5251,N_8367);
or U11773 (N_11773,N_8449,N_7830);
nand U11774 (N_11774,N_8645,N_8778);
nand U11775 (N_11775,N_5122,N_6123);
xnor U11776 (N_11776,N_9884,N_5019);
and U11777 (N_11777,N_9750,N_7429);
nor U11778 (N_11778,N_8144,N_5550);
nand U11779 (N_11779,N_6935,N_5778);
or U11780 (N_11780,N_8452,N_7384);
and U11781 (N_11781,N_6927,N_6226);
or U11782 (N_11782,N_8005,N_9891);
nand U11783 (N_11783,N_8347,N_9661);
nor U11784 (N_11784,N_8955,N_8051);
nor U11785 (N_11785,N_7903,N_5715);
nor U11786 (N_11786,N_8252,N_6547);
or U11787 (N_11787,N_9407,N_5986);
nand U11788 (N_11788,N_5105,N_6668);
nor U11789 (N_11789,N_9566,N_5905);
and U11790 (N_11790,N_8547,N_6760);
nand U11791 (N_11791,N_6045,N_8728);
nor U11792 (N_11792,N_9959,N_5572);
xor U11793 (N_11793,N_5903,N_5284);
nor U11794 (N_11794,N_6409,N_9007);
nand U11795 (N_11795,N_9963,N_6510);
or U11796 (N_11796,N_8550,N_8854);
or U11797 (N_11797,N_5355,N_9577);
and U11798 (N_11798,N_9800,N_6716);
or U11799 (N_11799,N_8479,N_8874);
and U11800 (N_11800,N_5902,N_6703);
xor U11801 (N_11801,N_9461,N_6924);
nand U11802 (N_11802,N_7361,N_8743);
nor U11803 (N_11803,N_6790,N_8535);
nand U11804 (N_11804,N_5451,N_6020);
nor U11805 (N_11805,N_5856,N_6205);
and U11806 (N_11806,N_8065,N_9230);
nor U11807 (N_11807,N_9624,N_9970);
nor U11808 (N_11808,N_9740,N_5422);
and U11809 (N_11809,N_8988,N_9715);
and U11810 (N_11810,N_9389,N_8589);
and U11811 (N_11811,N_5272,N_9243);
and U11812 (N_11812,N_8188,N_8544);
nor U11813 (N_11813,N_7259,N_7123);
or U11814 (N_11814,N_7061,N_8321);
or U11815 (N_11815,N_6331,N_8650);
nand U11816 (N_11816,N_7625,N_9458);
nand U11817 (N_11817,N_6499,N_8586);
and U11818 (N_11818,N_7201,N_7875);
nand U11819 (N_11819,N_7494,N_6823);
nand U11820 (N_11820,N_7004,N_5957);
nand U11821 (N_11821,N_5746,N_7500);
and U11822 (N_11822,N_5879,N_8465);
xor U11823 (N_11823,N_7796,N_5380);
and U11824 (N_11824,N_9376,N_6111);
or U11825 (N_11825,N_6513,N_6538);
nor U11826 (N_11826,N_7671,N_7188);
nor U11827 (N_11827,N_8085,N_6140);
nand U11828 (N_11828,N_9126,N_5526);
and U11829 (N_11829,N_9183,N_8120);
and U11830 (N_11830,N_9748,N_7099);
nor U11831 (N_11831,N_6304,N_9852);
and U11832 (N_11832,N_6136,N_9799);
nor U11833 (N_11833,N_6029,N_7258);
and U11834 (N_11834,N_9666,N_7970);
or U11835 (N_11835,N_7826,N_5347);
xor U11836 (N_11836,N_9654,N_5189);
xnor U11837 (N_11837,N_6183,N_6672);
or U11838 (N_11838,N_6695,N_7927);
or U11839 (N_11839,N_9824,N_5964);
and U11840 (N_11840,N_8812,N_8247);
nor U11841 (N_11841,N_5810,N_5958);
nor U11842 (N_11842,N_8525,N_7849);
or U11843 (N_11843,N_9027,N_9199);
or U11844 (N_11844,N_5538,N_5653);
nor U11845 (N_11845,N_6270,N_7270);
or U11846 (N_11846,N_6432,N_8319);
and U11847 (N_11847,N_7007,N_6733);
and U11848 (N_11848,N_6864,N_6694);
or U11849 (N_11849,N_7192,N_5342);
nand U11850 (N_11850,N_9484,N_6858);
and U11851 (N_11851,N_6606,N_6797);
nand U11852 (N_11852,N_7915,N_9417);
and U11853 (N_11853,N_7872,N_8651);
and U11854 (N_11854,N_7137,N_7821);
nor U11855 (N_11855,N_5835,N_5349);
or U11856 (N_11856,N_5655,N_8287);
and U11857 (N_11857,N_7633,N_8834);
or U11858 (N_11858,N_5842,N_8559);
nand U11859 (N_11859,N_9219,N_6356);
and U11860 (N_11860,N_6256,N_8514);
nand U11861 (N_11861,N_8111,N_5312);
nor U11862 (N_11862,N_9220,N_6998);
and U11863 (N_11863,N_9486,N_8097);
nand U11864 (N_11864,N_8677,N_9670);
and U11865 (N_11865,N_5194,N_5027);
xor U11866 (N_11866,N_7593,N_6085);
nor U11867 (N_11867,N_8594,N_6948);
or U11868 (N_11868,N_9609,N_6641);
nand U11869 (N_11869,N_8077,N_7476);
and U11870 (N_11870,N_5786,N_6210);
and U11871 (N_11871,N_7412,N_9729);
nor U11872 (N_11872,N_9216,N_6224);
nor U11873 (N_11873,N_5996,N_9904);
nand U11874 (N_11874,N_6207,N_7980);
nor U11875 (N_11875,N_5852,N_6687);
nand U11876 (N_11876,N_7529,N_5337);
xor U11877 (N_11877,N_9584,N_5668);
nand U11878 (N_11878,N_8300,N_9381);
nor U11879 (N_11879,N_7221,N_6768);
or U11880 (N_11880,N_9527,N_5717);
or U11881 (N_11881,N_7592,N_5455);
or U11882 (N_11882,N_8055,N_7117);
nand U11883 (N_11883,N_9828,N_7276);
or U11884 (N_11884,N_6460,N_8131);
nor U11885 (N_11885,N_5092,N_8396);
or U11886 (N_11886,N_5041,N_9955);
nor U11887 (N_11887,N_5395,N_5808);
and U11888 (N_11888,N_8386,N_6404);
nor U11889 (N_11889,N_6556,N_5237);
nor U11890 (N_11890,N_8579,N_7465);
nand U11891 (N_11891,N_6455,N_5804);
or U11892 (N_11892,N_5006,N_5787);
nand U11893 (N_11893,N_9130,N_8294);
nand U11894 (N_11894,N_9325,N_7062);
nand U11895 (N_11895,N_5514,N_6738);
or U11896 (N_11896,N_9906,N_5166);
and U11897 (N_11897,N_9324,N_5924);
nor U11898 (N_11898,N_5055,N_9018);
nand U11899 (N_11899,N_5894,N_6684);
or U11900 (N_11900,N_7573,N_9019);
nor U11901 (N_11901,N_9241,N_6599);
nand U11902 (N_11902,N_5785,N_8599);
nand U11903 (N_11903,N_9189,N_7725);
and U11904 (N_11904,N_7243,N_5874);
xnor U11905 (N_11905,N_9152,N_5613);
nand U11906 (N_11906,N_5770,N_6412);
nor U11907 (N_11907,N_9896,N_6742);
nand U11908 (N_11908,N_8846,N_9363);
and U11909 (N_11909,N_8062,N_9528);
and U11910 (N_11910,N_5186,N_6040);
nand U11911 (N_11911,N_6614,N_5669);
or U11912 (N_11912,N_6312,N_8870);
nand U11913 (N_11913,N_7474,N_9871);
nor U11914 (N_11914,N_6531,N_5254);
nand U11915 (N_11915,N_5383,N_8770);
nor U11916 (N_11916,N_6408,N_7517);
nor U11917 (N_11917,N_7696,N_9657);
nand U11918 (N_11918,N_9980,N_9539);
nor U11919 (N_11919,N_7440,N_8244);
or U11920 (N_11920,N_7773,N_8641);
and U11921 (N_11921,N_5980,N_9137);
or U11922 (N_11922,N_7298,N_5598);
xnor U11923 (N_11923,N_5993,N_8455);
nand U11924 (N_11924,N_6973,N_9379);
and U11925 (N_11925,N_8179,N_5135);
and U11926 (N_11926,N_9210,N_8307);
nor U11927 (N_11927,N_8388,N_5798);
nor U11928 (N_11928,N_7428,N_7794);
nor U11929 (N_11929,N_9594,N_6685);
xor U11930 (N_11930,N_5611,N_9223);
and U11931 (N_11931,N_8405,N_7262);
nor U11932 (N_11932,N_7684,N_5823);
and U11933 (N_11933,N_7330,N_9890);
xor U11934 (N_11934,N_5324,N_8371);
or U11935 (N_11935,N_9714,N_6117);
or U11936 (N_11936,N_7923,N_8693);
or U11937 (N_11937,N_5372,N_9806);
xnor U11938 (N_11938,N_8938,N_8262);
nand U11939 (N_11939,N_6827,N_7652);
xnor U11940 (N_11940,N_7964,N_5317);
xor U11941 (N_11941,N_6629,N_9221);
and U11942 (N_11942,N_6734,N_8237);
or U11943 (N_11943,N_6997,N_8637);
xnor U11944 (N_11944,N_7714,N_9303);
nor U11945 (N_11945,N_7920,N_5282);
nand U11946 (N_11946,N_8919,N_5108);
nor U11947 (N_11947,N_7427,N_5363);
or U11948 (N_11948,N_5579,N_6231);
and U11949 (N_11949,N_5507,N_5449);
or U11950 (N_11950,N_5644,N_7327);
or U11951 (N_11951,N_8189,N_5341);
xnor U11952 (N_11952,N_6482,N_8776);
nand U11953 (N_11953,N_6435,N_8380);
and U11954 (N_11954,N_7656,N_9811);
and U11955 (N_11955,N_7758,N_8691);
or U11956 (N_11956,N_9385,N_7550);
nand U11957 (N_11957,N_5664,N_7169);
or U11958 (N_11958,N_8635,N_6181);
xnor U11959 (N_11959,N_5970,N_5145);
nand U11960 (N_11960,N_7981,N_5240);
nand U11961 (N_11961,N_5813,N_6170);
xnor U11962 (N_11962,N_7130,N_9877);
or U11963 (N_11963,N_6126,N_6723);
nor U11964 (N_11964,N_8782,N_9358);
or U11965 (N_11965,N_8721,N_9191);
nor U11966 (N_11966,N_7786,N_5769);
or U11967 (N_11967,N_7346,N_5995);
xnor U11968 (N_11968,N_5339,N_8459);
nor U11969 (N_11969,N_8690,N_7176);
nand U11970 (N_11970,N_9952,N_6247);
nand U11971 (N_11971,N_6390,N_5287);
nand U11972 (N_11972,N_6232,N_5407);
nor U11973 (N_11973,N_6704,N_5303);
or U11974 (N_11974,N_5239,N_9105);
nand U11975 (N_11975,N_5850,N_5471);
or U11976 (N_11976,N_6515,N_6481);
or U11977 (N_11977,N_6979,N_9377);
xnor U11978 (N_11978,N_8295,N_9315);
and U11979 (N_11979,N_6047,N_9681);
or U11980 (N_11980,N_7103,N_7701);
nor U11981 (N_11981,N_9501,N_9117);
and U11982 (N_11982,N_6681,N_6293);
nor U11983 (N_11983,N_6281,N_6259);
nor U11984 (N_11984,N_5610,N_7655);
xnor U11985 (N_11985,N_6648,N_7208);
or U11986 (N_11986,N_5761,N_8406);
and U11987 (N_11987,N_9672,N_5073);
or U11988 (N_11988,N_8082,N_5067);
and U11989 (N_11989,N_7399,N_6729);
nand U11990 (N_11990,N_5435,N_8316);
nor U11991 (N_11991,N_9342,N_8157);
and U11992 (N_11992,N_6525,N_5584);
nor U11993 (N_11993,N_6813,N_9281);
nor U11994 (N_11994,N_8261,N_9513);
and U11995 (N_11995,N_5207,N_5681);
and U11996 (N_11996,N_7669,N_7372);
nand U11997 (N_11997,N_8871,N_6265);
and U11998 (N_11998,N_6495,N_8001);
and U11999 (N_11999,N_5348,N_7003);
and U12000 (N_12000,N_6292,N_6526);
nand U12001 (N_12001,N_7682,N_6709);
and U12002 (N_12002,N_5090,N_9536);
nand U12003 (N_12003,N_5115,N_6815);
nor U12004 (N_12004,N_5425,N_9673);
nand U12005 (N_12005,N_5172,N_7825);
and U12006 (N_12006,N_5791,N_6533);
and U12007 (N_12007,N_6969,N_5439);
or U12008 (N_12008,N_5623,N_5052);
or U12009 (N_12009,N_6922,N_9088);
or U12010 (N_12010,N_5714,N_9924);
nor U12011 (N_12011,N_5583,N_6321);
or U12012 (N_12012,N_9020,N_8259);
or U12013 (N_12013,N_5597,N_6254);
and U12014 (N_12014,N_5918,N_8805);
or U12015 (N_12015,N_5111,N_9169);
xnor U12016 (N_12016,N_6911,N_5865);
and U12017 (N_12017,N_9718,N_7400);
and U12018 (N_12018,N_7749,N_8814);
and U12019 (N_12019,N_9375,N_9236);
and U12020 (N_12020,N_9287,N_7022);
and U12021 (N_12021,N_6096,N_7748);
or U12022 (N_12022,N_6583,N_7620);
xor U12023 (N_12023,N_8210,N_8642);
and U12024 (N_12024,N_9255,N_5641);
nor U12025 (N_12025,N_9989,N_7235);
xor U12026 (N_12026,N_6610,N_8652);
nor U12027 (N_12027,N_9497,N_6517);
nand U12028 (N_12028,N_7144,N_8093);
nand U12029 (N_12029,N_9141,N_9604);
nand U12030 (N_12030,N_6942,N_9583);
or U12031 (N_12031,N_8844,N_9613);
nand U12032 (N_12032,N_9498,N_6315);
or U12033 (N_12033,N_8009,N_7992);
nor U12034 (N_12034,N_8647,N_6318);
nand U12035 (N_12035,N_5034,N_5766);
and U12036 (N_12036,N_5072,N_7249);
and U12037 (N_12037,N_9149,N_5004);
or U12038 (N_12038,N_5431,N_7815);
nand U12039 (N_12039,N_8035,N_9170);
and U12040 (N_12040,N_7983,N_9908);
xnor U12041 (N_12041,N_6196,N_9711);
or U12042 (N_12042,N_6011,N_8231);
nor U12043 (N_12043,N_6252,N_6080);
nand U12044 (N_12044,N_5486,N_6949);
nand U12045 (N_12045,N_6062,N_7047);
nand U12046 (N_12046,N_7030,N_5450);
or U12047 (N_12047,N_9535,N_7950);
nor U12048 (N_12048,N_7078,N_8375);
nor U12049 (N_12049,N_5306,N_6199);
nand U12050 (N_12050,N_7735,N_5631);
and U12051 (N_12051,N_6873,N_6195);
nor U12052 (N_12052,N_5520,N_7803);
or U12053 (N_12053,N_9362,N_9610);
nor U12054 (N_12054,N_8528,N_9655);
and U12055 (N_12055,N_9056,N_8118);
nor U12056 (N_12056,N_8944,N_8936);
and U12057 (N_12057,N_8600,N_8968);
xnor U12058 (N_12058,N_5139,N_6480);
nand U12059 (N_12059,N_9922,N_6893);
xnor U12060 (N_12060,N_7098,N_7410);
and U12061 (N_12061,N_9521,N_5947);
nand U12062 (N_12062,N_5848,N_8772);
or U12063 (N_12063,N_6743,N_9677);
xor U12064 (N_12064,N_8228,N_8039);
and U12065 (N_12065,N_5002,N_9882);
nand U12066 (N_12066,N_7541,N_8495);
and U12067 (N_12067,N_7998,N_7618);
and U12068 (N_12068,N_6635,N_8921);
or U12069 (N_12069,N_7715,N_9618);
nor U12070 (N_12070,N_7139,N_9675);
nor U12071 (N_12071,N_8019,N_5388);
xnor U12072 (N_12072,N_8842,N_6505);
nand U12073 (N_12073,N_7675,N_7704);
xor U12074 (N_12074,N_6124,N_5910);
nor U12075 (N_12075,N_9621,N_6235);
and U12076 (N_12076,N_7075,N_7364);
xor U12077 (N_12077,N_6022,N_6399);
xnor U12078 (N_12078,N_7694,N_5084);
and U12079 (N_12079,N_5862,N_7044);
or U12080 (N_12080,N_7043,N_5160);
or U12081 (N_12081,N_5972,N_8485);
nor U12082 (N_12082,N_7810,N_7305);
nor U12083 (N_12083,N_8670,N_7939);
nor U12084 (N_12084,N_8972,N_7495);
and U12085 (N_12085,N_9423,N_5988);
nand U12086 (N_12086,N_7995,N_6759);
nor U12087 (N_12087,N_9574,N_8355);
and U12088 (N_12088,N_6484,N_8831);
nand U12089 (N_12089,N_5755,N_9194);
nor U12090 (N_12090,N_5393,N_9758);
or U12091 (N_12091,N_7393,N_8377);
and U12092 (N_12092,N_5493,N_7224);
nor U12093 (N_12093,N_9665,N_9842);
nand U12094 (N_12094,N_9083,N_5978);
nor U12095 (N_12095,N_6931,N_9254);
or U12096 (N_12096,N_5376,N_6385);
or U12097 (N_12097,N_8461,N_9931);
xnor U12098 (N_12098,N_6914,N_8588);
or U12099 (N_12099,N_8066,N_5351);
or U12100 (N_12100,N_8269,N_5294);
nor U12101 (N_12101,N_7947,N_5707);
and U12102 (N_12102,N_8720,N_8203);
nand U12103 (N_12103,N_9585,N_8068);
nand U12104 (N_12104,N_5051,N_9634);
nor U12105 (N_12105,N_5884,N_9785);
or U12106 (N_12106,N_9937,N_9386);
and U12107 (N_12107,N_8007,N_8033);
or U12108 (N_12108,N_7196,N_8334);
xnor U12109 (N_12109,N_8089,N_7158);
nand U12110 (N_12110,N_9706,N_5124);
nor U12111 (N_12111,N_5142,N_9043);
or U12112 (N_12112,N_8372,N_9246);
or U12113 (N_12113,N_8523,N_8790);
nand U12114 (N_12114,N_7328,N_9912);
or U12115 (N_12115,N_6211,N_9010);
nand U12116 (N_12116,N_6667,N_5304);
or U12117 (N_12117,N_8041,N_8318);
and U12118 (N_12118,N_5895,N_7852);
nand U12119 (N_12119,N_6268,N_8769);
and U12120 (N_12120,N_7644,N_5060);
nor U12121 (N_12121,N_8793,N_9602);
or U12122 (N_12122,N_8657,N_7713);
or U12123 (N_12123,N_5950,N_8956);
and U12124 (N_12124,N_7960,N_6983);
nor U12125 (N_12125,N_8414,N_6353);
nand U12126 (N_12126,N_5727,N_9442);
or U12127 (N_12127,N_5973,N_5086);
or U12128 (N_12128,N_7888,N_7341);
and U12129 (N_12129,N_6980,N_9918);
nor U12130 (N_12130,N_5656,N_8354);
and U12131 (N_12131,N_9547,N_6974);
nand U12132 (N_12132,N_7914,N_5901);
nand U12133 (N_12133,N_5125,N_7303);
nor U12134 (N_12134,N_8680,N_8997);
nand U12135 (N_12135,N_5350,N_7336);
and U12136 (N_12136,N_7049,N_6617);
nor U12137 (N_12137,N_6546,N_9771);
nor U12138 (N_12138,N_7604,N_5698);
or U12139 (N_12139,N_5133,N_9581);
and U12140 (N_12140,N_8044,N_8092);
and U12141 (N_12141,N_7976,N_6120);
nand U12142 (N_12142,N_7804,N_7376);
xnor U12143 (N_12143,N_9939,N_9444);
xor U12144 (N_12144,N_8843,N_8407);
and U12145 (N_12145,N_5058,N_8853);
nor U12146 (N_12146,N_9071,N_5127);
nor U12147 (N_12147,N_7072,N_5595);
or U12148 (N_12148,N_6705,N_9399);
or U12149 (N_12149,N_6888,N_5499);
xnor U12150 (N_12150,N_8255,N_8037);
or U12151 (N_12151,N_7921,N_9110);
nor U12152 (N_12152,N_5082,N_7197);
nor U12153 (N_12153,N_7285,N_5079);
or U12154 (N_12154,N_6895,N_5826);
nand U12155 (N_12155,N_5649,N_6352);
or U12156 (N_12156,N_8794,N_7651);
nand U12157 (N_12157,N_7668,N_5858);
nor U12158 (N_12158,N_8920,N_9836);
and U12159 (N_12159,N_6406,N_7228);
or U12160 (N_12160,N_6422,N_6048);
xnor U12161 (N_12161,N_9683,N_6662);
and U12162 (N_12162,N_5763,N_9791);
or U12163 (N_12163,N_6950,N_5594);
nand U12164 (N_12164,N_9045,N_9516);
nor U12165 (N_12165,N_9422,N_9441);
or U12166 (N_12166,N_8666,N_5113);
nand U12167 (N_12167,N_7716,N_9770);
and U12168 (N_12168,N_6451,N_8561);
and U12169 (N_12169,N_5719,N_5419);
nor U12170 (N_12170,N_9894,N_9404);
or U12171 (N_12171,N_5817,N_8742);
and U12172 (N_12172,N_7731,N_9650);
or U12173 (N_12173,N_5494,N_9345);
or U12174 (N_12174,N_7407,N_5087);
nand U12175 (N_12175,N_8655,N_7873);
nand U12176 (N_12176,N_7763,N_8980);
nor U12177 (N_12177,N_6934,N_7475);
or U12178 (N_12178,N_7623,N_5733);
nor U12179 (N_12179,N_7418,N_9702);
xor U12180 (N_12180,N_5236,N_6425);
nand U12181 (N_12181,N_6468,N_5481);
nor U12182 (N_12182,N_8576,N_8392);
nand U12183 (N_12183,N_6630,N_9590);
and U12184 (N_12184,N_7403,N_7458);
nand U12185 (N_12185,N_9793,N_8176);
or U12186 (N_12186,N_9962,N_5192);
or U12187 (N_12187,N_6603,N_8771);
nand U12188 (N_12188,N_5558,N_9905);
or U12189 (N_12189,N_6913,N_8472);
and U12190 (N_12190,N_6920,N_6636);
xnor U12191 (N_12191,N_5751,N_8787);
or U12192 (N_12192,N_7267,N_9177);
or U12193 (N_12193,N_6149,N_9159);
and U12194 (N_12194,N_6361,N_6214);
and U12195 (N_12195,N_7135,N_7891);
or U12196 (N_12196,N_5937,N_6579);
nand U12197 (N_12197,N_5544,N_8727);
nor U12198 (N_12198,N_6443,N_9993);
or U12199 (N_12199,N_5683,N_9514);
nand U12200 (N_12200,N_6129,N_6982);
or U12201 (N_12201,N_6274,N_6303);
and U12202 (N_12202,N_5219,N_6549);
nand U12203 (N_12203,N_8469,N_8667);
and U12204 (N_12204,N_7902,N_5530);
nand U12205 (N_12205,N_8689,N_7304);
nor U12206 (N_12206,N_5149,N_6853);
or U12207 (N_12207,N_7148,N_8694);
nand U12208 (N_12208,N_6128,N_5577);
nand U12209 (N_12209,N_5409,N_5233);
nand U12210 (N_12210,N_7871,N_8710);
or U12211 (N_12211,N_6401,N_8958);
nand U12212 (N_12212,N_8904,N_7679);
or U12213 (N_12213,N_8315,N_8489);
nor U12214 (N_12214,N_8755,N_6845);
nor U12215 (N_12215,N_6721,N_6846);
and U12216 (N_12216,N_6179,N_6057);
nor U12217 (N_12217,N_6465,N_9612);
nand U12218 (N_12218,N_7848,N_6507);
nand U12219 (N_12219,N_8365,N_9525);
nand U12220 (N_12220,N_6023,N_7791);
or U12221 (N_12221,N_5344,N_6225);
xor U12222 (N_12222,N_9493,N_7266);
nor U12223 (N_12223,N_9304,N_7963);
nor U12224 (N_12224,N_6257,N_5181);
nor U12225 (N_12225,N_5176,N_8487);
nand U12226 (N_12226,N_8930,N_5709);
or U12227 (N_12227,N_7414,N_5098);
xor U12228 (N_12228,N_5120,N_8604);
nand U12229 (N_12229,N_5216,N_8918);
and U12230 (N_12230,N_8707,N_7985);
or U12231 (N_12231,N_7299,N_6792);
and U12232 (N_12232,N_9659,N_8475);
and U12233 (N_12233,N_5314,N_5277);
or U12234 (N_12234,N_5556,N_8351);
or U12235 (N_12235,N_7632,N_6590);
nand U12236 (N_12236,N_9717,N_6957);
nor U12237 (N_12237,N_6436,N_8350);
and U12238 (N_12238,N_6559,N_5888);
nand U12239 (N_12239,N_8088,N_9251);
nand U12240 (N_12240,N_9803,N_6362);
xor U12241 (N_12241,N_7561,N_5871);
nor U12242 (N_12242,N_9730,N_6906);
nor U12243 (N_12243,N_6701,N_8928);
and U12244 (N_12244,N_5068,N_8340);
xor U12245 (N_12245,N_8634,N_6103);
and U12246 (N_12246,N_8428,N_8132);
and U12247 (N_12247,N_6739,N_6382);
or U12248 (N_12248,N_9935,N_8091);
nor U12249 (N_12249,N_7973,N_9769);
xor U12250 (N_12250,N_5775,N_9844);
nor U12251 (N_12251,N_9976,N_9212);
and U12252 (N_12252,N_5030,N_9947);
or U12253 (N_12253,N_7409,N_5428);
nand U12254 (N_12254,N_5697,N_7095);
nor U12255 (N_12255,N_5930,N_8369);
nand U12256 (N_12256,N_6670,N_8345);
and U12257 (N_12257,N_5999,N_8220);
nand U12258 (N_12258,N_5110,N_5602);
xnor U12259 (N_12259,N_9885,N_6068);
or U12260 (N_12260,N_8565,N_8325);
or U12261 (N_12261,N_5634,N_6594);
nand U12262 (N_12262,N_7545,N_7709);
and U12263 (N_12263,N_7126,N_9603);
or U12264 (N_12264,N_8765,N_6004);
or U12265 (N_12265,N_6030,N_9339);
xor U12266 (N_12266,N_6041,N_9108);
nand U12267 (N_12267,N_6714,N_5096);
nor U12268 (N_12268,N_6097,N_9826);
and U12269 (N_12269,N_9192,N_5089);
or U12270 (N_12270,N_6902,N_6767);
nand U12271 (N_12271,N_8905,N_5230);
and U12272 (N_12272,N_9202,N_5956);
xor U12273 (N_12273,N_5854,N_6376);
nor U12274 (N_12274,N_5519,N_5474);
nor U12275 (N_12275,N_5900,N_7734);
or U12276 (N_12276,N_5789,N_7598);
or U12277 (N_12277,N_6953,N_6064);
nor U12278 (N_12278,N_8889,N_5136);
or U12279 (N_12279,N_7883,N_5515);
nor U12280 (N_12280,N_8466,N_5516);
nand U12281 (N_12281,N_6309,N_9031);
nor U12282 (N_12282,N_7772,N_7611);
nor U12283 (N_12283,N_8722,N_7001);
or U12284 (N_12284,N_7876,N_8503);
xnor U12285 (N_12285,N_8274,N_9788);
nor U12286 (N_12286,N_8101,N_7528);
nor U12287 (N_12287,N_7020,N_5540);
and U12288 (N_12288,N_5790,N_9051);
nand U12289 (N_12289,N_7486,N_7121);
and U12290 (N_12290,N_5020,N_9193);
and U12291 (N_12291,N_7621,N_9692);
xnor U12292 (N_12292,N_9237,N_8752);
nor U12293 (N_12293,N_6514,N_8924);
and U12294 (N_12294,N_5100,N_5362);
and U12295 (N_12295,N_5542,N_7406);
nand U12296 (N_12296,N_5107,N_7163);
nand U12297 (N_12297,N_9696,N_8698);
or U12298 (N_12298,N_8273,N_9834);
or U12299 (N_12299,N_8010,N_5364);
and U12300 (N_12300,N_6912,N_7155);
nor U12301 (N_12301,N_5877,N_9739);
or U12302 (N_12302,N_7432,N_5222);
nand U12303 (N_12303,N_8482,N_7937);
xor U12304 (N_12304,N_7343,N_7862);
nand U12305 (N_12305,N_6188,N_5185);
nor U12306 (N_12306,N_8801,N_7723);
xnor U12307 (N_12307,N_6341,N_8568);
nand U12308 (N_12308,N_8848,N_7765);
and U12309 (N_12309,N_5706,N_5117);
or U12310 (N_12310,N_8094,N_8190);
nand U12311 (N_12311,N_5248,N_8245);
nor U12312 (N_12312,N_6118,N_9549);
nand U12313 (N_12313,N_5379,N_6475);
nor U12314 (N_12314,N_6926,N_7531);
xnor U12315 (N_12315,N_8899,N_7081);
xor U12316 (N_12316,N_6887,N_5318);
nand U12317 (N_12317,N_7339,N_5378);
and U12318 (N_12318,N_5642,N_9830);
nand U12319 (N_12319,N_5046,N_8861);
nor U12320 (N_12320,N_8074,N_6036);
xnor U12321 (N_12321,N_9166,N_7816);
and U12322 (N_12322,N_8150,N_6830);
nor U12323 (N_12323,N_7649,N_5992);
nor U12324 (N_12324,N_6197,N_5444);
or U12325 (N_12325,N_7762,N_6089);
nor U12326 (N_12326,N_8927,N_5748);
and U12327 (N_12327,N_5268,N_5658);
or U12328 (N_12328,N_6605,N_7646);
nor U12329 (N_12329,N_8117,N_7240);
and U12330 (N_12330,N_6364,N_7700);
and U12331 (N_12331,N_7362,N_8305);
nand U12332 (N_12332,N_6223,N_6607);
or U12333 (N_12333,N_8483,N_5873);
and U12334 (N_12334,N_7958,N_5846);
nor U12335 (N_12335,N_9359,N_7982);
and U12336 (N_12336,N_8687,N_5919);
or U12337 (N_12337,N_8541,N_7312);
nand U12338 (N_12338,N_5369,N_6994);
and U12339 (N_12339,N_9104,N_9587);
and U12340 (N_12340,N_7242,N_9934);
nand U12341 (N_12341,N_6217,N_8258);
xor U12342 (N_12342,N_5760,N_7411);
nor U12343 (N_12343,N_9213,N_6316);
nor U12344 (N_12344,N_5600,N_6535);
nand U12345 (N_12345,N_9034,N_9938);
nor U12346 (N_12346,N_9794,N_6638);
and U12347 (N_12347,N_8301,N_5974);
or U12348 (N_12348,N_8158,N_9330);
and U12349 (N_12349,N_8213,N_5522);
and U12350 (N_12350,N_7894,N_7489);
nand U12351 (N_12351,N_6448,N_9682);
nand U12352 (N_12352,N_8304,N_8022);
and U12353 (N_12353,N_6589,N_5063);
or U12354 (N_12354,N_7952,N_5509);
nor U12355 (N_12355,N_6938,N_5799);
or U12356 (N_12356,N_5353,N_6174);
and U12357 (N_12357,N_6897,N_7302);
and U12358 (N_12358,N_9186,N_7831);
or U12359 (N_12359,N_9172,N_6396);
nand U12360 (N_12360,N_8555,N_9848);
or U12361 (N_12361,N_7984,N_8476);
nand U12362 (N_12362,N_7776,N_8298);
nor U12363 (N_12363,N_7180,N_6803);
xor U12364 (N_12364,N_6615,N_5500);
nor U12365 (N_12365,N_6445,N_5038);
or U12366 (N_12366,N_8310,N_6456);
nand U12367 (N_12367,N_7941,N_7587);
or U12368 (N_12368,N_8285,N_5565);
nor U12369 (N_12369,N_7997,N_8879);
or U12370 (N_12370,N_9745,N_7466);
nand U12371 (N_12371,N_9776,N_8173);
nor U12372 (N_12372,N_6697,N_8863);
and U12373 (N_12373,N_8998,N_8492);
and U12374 (N_12374,N_7441,N_8474);
nand U12375 (N_12375,N_6253,N_9022);
nor U12376 (N_12376,N_6678,N_6966);
or U12377 (N_12377,N_9006,N_9982);
nand U12378 (N_12378,N_5756,N_9977);
nand U12379 (N_12379,N_6320,N_7665);
and U12380 (N_12380,N_8297,N_9036);
or U12381 (N_12381,N_6410,N_6907);
nand U12382 (N_12382,N_9195,N_7926);
nand U12383 (N_12383,N_5688,N_9029);
or U12384 (N_12384,N_5657,N_5083);
and U12385 (N_12385,N_9781,N_9818);
and U12386 (N_12386,N_6613,N_6497);
nor U12387 (N_12387,N_5983,N_5531);
and U12388 (N_12388,N_6340,N_8165);
and U12389 (N_12389,N_9494,N_7706);
nand U12390 (N_12390,N_9667,N_9643);
or U12391 (N_12391,N_8857,N_8538);
and U12392 (N_12392,N_9509,N_9637);
nor U12393 (N_12393,N_9684,N_9988);
or U12394 (N_12394,N_7263,N_6776);
nand U12395 (N_12395,N_5184,N_8804);
or U12396 (N_12396,N_6833,N_7658);
nand U12397 (N_12397,N_9647,N_9238);
or U12398 (N_12398,N_6190,N_5845);
nor U12399 (N_12399,N_7521,N_5963);
or U12400 (N_12400,N_9866,N_7234);
or U12401 (N_12401,N_9943,N_8511);
nand U12402 (N_12402,N_9437,N_6273);
nand U12403 (N_12403,N_9881,N_8813);
nor U12404 (N_12404,N_8609,N_5636);
nand U12405 (N_12405,N_9512,N_5807);
or U12406 (N_12406,N_7187,N_9580);
or U12407 (N_12407,N_5887,N_7792);
xor U12408 (N_12408,N_9270,N_9888);
and U12409 (N_12409,N_5764,N_5586);
or U12410 (N_12410,N_5913,N_6932);
nor U12411 (N_12411,N_8669,N_7769);
or U12412 (N_12412,N_5169,N_8320);
xor U12413 (N_12413,N_8829,N_9101);
xor U12414 (N_12414,N_8987,N_8665);
nor U12415 (N_12415,N_7660,N_5093);
nand U12416 (N_12416,N_7994,N_5562);
or U12417 (N_12417,N_8498,N_8754);
or U12418 (N_12418,N_9143,N_7450);
and U12419 (N_12419,N_8532,N_6604);
and U12420 (N_12420,N_6285,N_9986);
xnor U12421 (N_12421,N_7778,N_5643);
or U12422 (N_12422,N_6802,N_6763);
nor U12423 (N_12423,N_9588,N_7837);
and U12424 (N_12424,N_7501,N_8477);
and U12425 (N_12425,N_7470,N_9293);
or U12426 (N_12426,N_5091,N_7171);
and U12427 (N_12427,N_8536,N_7219);
nand U12428 (N_12428,N_9709,N_8142);
xnor U12429 (N_12429,N_7829,N_8620);
nor U12430 (N_12430,N_9459,N_6972);
nand U12431 (N_12431,N_6415,N_9465);
nand U12432 (N_12432,N_7562,N_9150);
xnor U12433 (N_12433,N_6050,N_6106);
and U12434 (N_12434,N_8236,N_6450);
nor U12435 (N_12435,N_6498,N_6778);
and U12436 (N_12436,N_6775,N_5776);
nor U12437 (N_12437,N_9025,N_9911);
nor U12438 (N_12438,N_9344,N_8678);
and U12439 (N_12439,N_9470,N_6842);
nor U12440 (N_12440,N_9181,N_9732);
nand U12441 (N_12441,N_9235,N_8738);
and U12442 (N_12442,N_5193,N_5638);
and U12443 (N_12443,N_7415,N_7653);
and U12444 (N_12444,N_7291,N_5465);
xnor U12445 (N_12445,N_5608,N_6575);
nor U12446 (N_12446,N_9505,N_5024);
or U12447 (N_12447,N_8507,N_9229);
nor U12448 (N_12448,N_6006,N_9412);
or U12449 (N_12449,N_6855,N_7744);
nand U12450 (N_12450,N_6544,N_5325);
and U12451 (N_12451,N_5408,N_9641);
nor U12452 (N_12452,N_6328,N_9414);
or U12453 (N_12453,N_6572,N_9576);
nand U12454 (N_12454,N_7116,N_7738);
nor U12455 (N_12455,N_9849,N_9127);
or U12456 (N_12456,N_9518,N_5180);
nand U12457 (N_12457,N_9320,N_5592);
nand U12458 (N_12458,N_8811,N_6829);
or U12459 (N_12459,N_7698,N_6871);
xnor U12460 (N_12460,N_5382,N_9949);
or U12461 (N_12461,N_7685,N_5260);
nor U12462 (N_12462,N_9267,N_9015);
nand U12463 (N_12463,N_8260,N_7608);
nor U12464 (N_12464,N_6345,N_6472);
and U12465 (N_12465,N_9910,N_8227);
nand U12466 (N_12466,N_7140,N_9353);
or U12467 (N_12467,N_6326,N_5338);
or U12468 (N_12468,N_9089,N_8741);
and U12469 (N_12469,N_9540,N_7392);
or U12470 (N_12470,N_9222,N_5429);
nor U12471 (N_12471,N_9428,N_9473);
and U12472 (N_12472,N_7353,N_9436);
nand U12473 (N_12473,N_7178,N_7027);
or U12474 (N_12474,N_9140,N_6884);
nand U12475 (N_12475,N_8453,N_5489);
nor U12476 (N_12476,N_7011,N_6886);
nor U12477 (N_12477,N_8073,N_6249);
nor U12478 (N_12478,N_6250,N_5899);
or U12479 (N_12479,N_9327,N_6308);
and U12480 (N_12480,N_9035,N_7000);
or U12481 (N_12481,N_6650,N_5975);
nand U12482 (N_12482,N_6255,N_8060);
nand U12483 (N_12483,N_7695,N_5319);
and U12484 (N_12484,N_8850,N_5591);
or U12485 (N_12485,N_9445,N_5965);
nor U12486 (N_12486,N_9499,N_7579);
nand U12487 (N_12487,N_7039,N_8499);
or U12488 (N_12488,N_8493,N_6724);
or U12489 (N_12489,N_5927,N_6879);
nand U12490 (N_12490,N_7597,N_9808);
nor U12491 (N_12491,N_9552,N_8673);
nand U12492 (N_12492,N_7217,N_9472);
and U12493 (N_12493,N_5029,N_8289);
and U12494 (N_12494,N_6414,N_8403);
nand U12495 (N_12495,N_6208,N_5736);
nand U12496 (N_12496,N_7307,N_9774);
xnor U12497 (N_12497,N_8686,N_8979);
nor U12498 (N_12498,N_6810,N_5628);
nand U12499 (N_12499,N_9479,N_8240);
xnor U12500 (N_12500,N_8008,N_9654);
and U12501 (N_12501,N_8412,N_9220);
nand U12502 (N_12502,N_5940,N_9404);
nand U12503 (N_12503,N_6982,N_9557);
or U12504 (N_12504,N_5462,N_6385);
nor U12505 (N_12505,N_5189,N_5638);
nor U12506 (N_12506,N_7078,N_7146);
nor U12507 (N_12507,N_6123,N_7211);
nor U12508 (N_12508,N_6022,N_8262);
nor U12509 (N_12509,N_8164,N_8788);
nor U12510 (N_12510,N_7529,N_9149);
or U12511 (N_12511,N_8250,N_7489);
and U12512 (N_12512,N_9661,N_7911);
and U12513 (N_12513,N_7583,N_8794);
nor U12514 (N_12514,N_9815,N_6563);
xnor U12515 (N_12515,N_5173,N_8392);
nand U12516 (N_12516,N_6652,N_7302);
nand U12517 (N_12517,N_5072,N_6791);
and U12518 (N_12518,N_6646,N_6579);
nand U12519 (N_12519,N_9379,N_7259);
nand U12520 (N_12520,N_6044,N_7560);
or U12521 (N_12521,N_8915,N_7147);
nand U12522 (N_12522,N_6642,N_8096);
or U12523 (N_12523,N_5797,N_8382);
xor U12524 (N_12524,N_6086,N_5154);
nand U12525 (N_12525,N_6726,N_8673);
nand U12526 (N_12526,N_9898,N_7223);
or U12527 (N_12527,N_5751,N_9136);
and U12528 (N_12528,N_7976,N_5501);
nor U12529 (N_12529,N_8937,N_7960);
nor U12530 (N_12530,N_8532,N_5342);
or U12531 (N_12531,N_7408,N_7343);
nand U12532 (N_12532,N_8308,N_6585);
nor U12533 (N_12533,N_8496,N_6488);
nand U12534 (N_12534,N_5394,N_9423);
or U12535 (N_12535,N_5820,N_9574);
nand U12536 (N_12536,N_6100,N_7926);
nand U12537 (N_12537,N_5422,N_6366);
or U12538 (N_12538,N_5776,N_5445);
nor U12539 (N_12539,N_5099,N_9518);
nand U12540 (N_12540,N_7338,N_7263);
and U12541 (N_12541,N_9900,N_5237);
nor U12542 (N_12542,N_9207,N_8057);
nand U12543 (N_12543,N_5089,N_9024);
xnor U12544 (N_12544,N_7410,N_7824);
nor U12545 (N_12545,N_9931,N_5908);
and U12546 (N_12546,N_5939,N_5914);
nor U12547 (N_12547,N_7258,N_6772);
or U12548 (N_12548,N_7541,N_9135);
or U12549 (N_12549,N_7542,N_9901);
xnor U12550 (N_12550,N_8272,N_5881);
and U12551 (N_12551,N_5444,N_5050);
nand U12552 (N_12552,N_9634,N_8181);
or U12553 (N_12553,N_5654,N_9637);
nor U12554 (N_12554,N_9028,N_9971);
and U12555 (N_12555,N_9712,N_8022);
nand U12556 (N_12556,N_9472,N_8187);
and U12557 (N_12557,N_9117,N_5017);
nor U12558 (N_12558,N_6207,N_6571);
xnor U12559 (N_12559,N_6041,N_9181);
nor U12560 (N_12560,N_9023,N_7808);
xor U12561 (N_12561,N_5356,N_7357);
and U12562 (N_12562,N_7915,N_5763);
nor U12563 (N_12563,N_7307,N_6119);
nand U12564 (N_12564,N_5897,N_7163);
and U12565 (N_12565,N_8374,N_9473);
and U12566 (N_12566,N_5059,N_5378);
or U12567 (N_12567,N_7309,N_9946);
nand U12568 (N_12568,N_8874,N_5079);
nand U12569 (N_12569,N_5619,N_8058);
or U12570 (N_12570,N_5064,N_7030);
nor U12571 (N_12571,N_7331,N_9677);
nor U12572 (N_12572,N_7502,N_7515);
nor U12573 (N_12573,N_8124,N_6743);
nand U12574 (N_12574,N_7425,N_8725);
or U12575 (N_12575,N_5198,N_5313);
nor U12576 (N_12576,N_7718,N_6399);
xnor U12577 (N_12577,N_8049,N_9043);
nand U12578 (N_12578,N_5105,N_5136);
and U12579 (N_12579,N_6824,N_7724);
nand U12580 (N_12580,N_6858,N_8149);
xnor U12581 (N_12581,N_5009,N_7743);
nor U12582 (N_12582,N_5706,N_6177);
and U12583 (N_12583,N_9078,N_8787);
nand U12584 (N_12584,N_6207,N_8400);
and U12585 (N_12585,N_8432,N_8729);
or U12586 (N_12586,N_7638,N_5976);
or U12587 (N_12587,N_5426,N_7275);
or U12588 (N_12588,N_8262,N_8956);
or U12589 (N_12589,N_8231,N_8455);
nand U12590 (N_12590,N_9362,N_5767);
nor U12591 (N_12591,N_7437,N_8039);
nor U12592 (N_12592,N_8322,N_7335);
or U12593 (N_12593,N_8651,N_5111);
and U12594 (N_12594,N_7814,N_9373);
nand U12595 (N_12595,N_6035,N_7081);
nand U12596 (N_12596,N_7541,N_5556);
or U12597 (N_12597,N_6023,N_7191);
xnor U12598 (N_12598,N_9293,N_5093);
and U12599 (N_12599,N_7338,N_6414);
nand U12600 (N_12600,N_5283,N_9288);
and U12601 (N_12601,N_6151,N_8853);
nand U12602 (N_12602,N_6298,N_6651);
nand U12603 (N_12603,N_5763,N_8780);
nor U12604 (N_12604,N_9584,N_5143);
nand U12605 (N_12605,N_7919,N_8169);
and U12606 (N_12606,N_8845,N_9222);
xor U12607 (N_12607,N_5767,N_8421);
nor U12608 (N_12608,N_9802,N_7444);
and U12609 (N_12609,N_7027,N_9634);
nor U12610 (N_12610,N_6181,N_7691);
nand U12611 (N_12611,N_5853,N_5401);
and U12612 (N_12612,N_5047,N_8732);
nor U12613 (N_12613,N_5218,N_8979);
or U12614 (N_12614,N_6313,N_9859);
and U12615 (N_12615,N_5241,N_9416);
nor U12616 (N_12616,N_8704,N_5635);
nor U12617 (N_12617,N_7910,N_7791);
nor U12618 (N_12618,N_5792,N_8412);
nand U12619 (N_12619,N_8053,N_8616);
or U12620 (N_12620,N_6329,N_6926);
nand U12621 (N_12621,N_5517,N_9330);
xnor U12622 (N_12622,N_9788,N_9697);
xor U12623 (N_12623,N_8200,N_9064);
nand U12624 (N_12624,N_6127,N_7414);
nand U12625 (N_12625,N_9944,N_9521);
xor U12626 (N_12626,N_6771,N_8613);
and U12627 (N_12627,N_5816,N_8068);
or U12628 (N_12628,N_8732,N_9729);
or U12629 (N_12629,N_7846,N_8012);
nand U12630 (N_12630,N_8634,N_6208);
nor U12631 (N_12631,N_5808,N_9047);
xor U12632 (N_12632,N_7048,N_5583);
or U12633 (N_12633,N_5310,N_8464);
nand U12634 (N_12634,N_9637,N_7590);
or U12635 (N_12635,N_8103,N_8087);
or U12636 (N_12636,N_7209,N_6206);
nand U12637 (N_12637,N_8118,N_6825);
and U12638 (N_12638,N_6479,N_6641);
or U12639 (N_12639,N_9688,N_5036);
nor U12640 (N_12640,N_7938,N_7105);
and U12641 (N_12641,N_9728,N_8834);
or U12642 (N_12642,N_7643,N_8179);
and U12643 (N_12643,N_8064,N_5234);
nand U12644 (N_12644,N_5394,N_5424);
xor U12645 (N_12645,N_9816,N_8209);
or U12646 (N_12646,N_6208,N_5157);
nand U12647 (N_12647,N_9808,N_7890);
xor U12648 (N_12648,N_5058,N_6188);
nor U12649 (N_12649,N_7120,N_7844);
nand U12650 (N_12650,N_8987,N_8005);
nor U12651 (N_12651,N_5389,N_9149);
nor U12652 (N_12652,N_8379,N_8005);
and U12653 (N_12653,N_5602,N_9972);
nand U12654 (N_12654,N_6201,N_5727);
or U12655 (N_12655,N_7853,N_8286);
nand U12656 (N_12656,N_9306,N_5705);
or U12657 (N_12657,N_5123,N_6277);
nand U12658 (N_12658,N_6157,N_7564);
nor U12659 (N_12659,N_7305,N_9632);
or U12660 (N_12660,N_5314,N_9118);
or U12661 (N_12661,N_5902,N_7495);
nor U12662 (N_12662,N_9195,N_9092);
nor U12663 (N_12663,N_5043,N_6211);
and U12664 (N_12664,N_7794,N_9020);
nor U12665 (N_12665,N_7599,N_9391);
nor U12666 (N_12666,N_5035,N_7896);
nand U12667 (N_12667,N_6370,N_5013);
or U12668 (N_12668,N_7069,N_5243);
nand U12669 (N_12669,N_7312,N_6147);
or U12670 (N_12670,N_8099,N_9643);
or U12671 (N_12671,N_5878,N_5665);
or U12672 (N_12672,N_7384,N_8117);
nand U12673 (N_12673,N_9898,N_8175);
xnor U12674 (N_12674,N_8654,N_6554);
and U12675 (N_12675,N_6257,N_9314);
or U12676 (N_12676,N_6032,N_7932);
nand U12677 (N_12677,N_7497,N_5775);
and U12678 (N_12678,N_7962,N_5525);
and U12679 (N_12679,N_5524,N_5425);
nor U12680 (N_12680,N_5393,N_5282);
and U12681 (N_12681,N_7689,N_9565);
or U12682 (N_12682,N_8111,N_5397);
nand U12683 (N_12683,N_9153,N_6565);
or U12684 (N_12684,N_5941,N_7411);
xnor U12685 (N_12685,N_7664,N_7371);
nor U12686 (N_12686,N_7572,N_6053);
or U12687 (N_12687,N_9814,N_7227);
and U12688 (N_12688,N_6991,N_5559);
or U12689 (N_12689,N_8261,N_9023);
nand U12690 (N_12690,N_7753,N_8780);
or U12691 (N_12691,N_9566,N_6751);
nand U12692 (N_12692,N_9011,N_9074);
nand U12693 (N_12693,N_7405,N_8175);
nor U12694 (N_12694,N_5232,N_5977);
or U12695 (N_12695,N_5526,N_7501);
nand U12696 (N_12696,N_7324,N_9591);
nand U12697 (N_12697,N_6863,N_5398);
or U12698 (N_12698,N_8813,N_5619);
or U12699 (N_12699,N_8207,N_8451);
nand U12700 (N_12700,N_7427,N_9301);
nand U12701 (N_12701,N_9066,N_9839);
or U12702 (N_12702,N_6251,N_8357);
and U12703 (N_12703,N_5373,N_8102);
nand U12704 (N_12704,N_6804,N_8491);
nor U12705 (N_12705,N_7813,N_9477);
or U12706 (N_12706,N_5406,N_7294);
and U12707 (N_12707,N_5375,N_8959);
or U12708 (N_12708,N_6700,N_8088);
or U12709 (N_12709,N_7508,N_5102);
nor U12710 (N_12710,N_9533,N_7807);
and U12711 (N_12711,N_8374,N_9312);
nor U12712 (N_12712,N_6027,N_6581);
nor U12713 (N_12713,N_5567,N_9193);
or U12714 (N_12714,N_8050,N_9481);
or U12715 (N_12715,N_5240,N_6795);
or U12716 (N_12716,N_5947,N_8847);
or U12717 (N_12717,N_5268,N_8134);
nand U12718 (N_12718,N_9386,N_8351);
xnor U12719 (N_12719,N_6290,N_9776);
nor U12720 (N_12720,N_9619,N_8613);
or U12721 (N_12721,N_6750,N_7321);
or U12722 (N_12722,N_5973,N_8789);
xnor U12723 (N_12723,N_5650,N_9950);
and U12724 (N_12724,N_9216,N_8067);
nor U12725 (N_12725,N_7843,N_5727);
nor U12726 (N_12726,N_6202,N_5130);
and U12727 (N_12727,N_5879,N_9419);
nand U12728 (N_12728,N_9215,N_7038);
and U12729 (N_12729,N_5193,N_8530);
or U12730 (N_12730,N_5487,N_6323);
and U12731 (N_12731,N_7500,N_7906);
or U12732 (N_12732,N_5973,N_9309);
nand U12733 (N_12733,N_9550,N_6776);
nand U12734 (N_12734,N_6125,N_7629);
nor U12735 (N_12735,N_5874,N_6844);
nor U12736 (N_12736,N_9938,N_7676);
xnor U12737 (N_12737,N_9881,N_7758);
nand U12738 (N_12738,N_9223,N_8228);
nor U12739 (N_12739,N_6744,N_7597);
or U12740 (N_12740,N_9071,N_5345);
and U12741 (N_12741,N_7633,N_6712);
nand U12742 (N_12742,N_5919,N_5336);
or U12743 (N_12743,N_5878,N_6522);
nand U12744 (N_12744,N_8374,N_6764);
nor U12745 (N_12745,N_6344,N_5501);
nor U12746 (N_12746,N_7397,N_5086);
or U12747 (N_12747,N_6733,N_5239);
nand U12748 (N_12748,N_9113,N_9294);
and U12749 (N_12749,N_8499,N_6862);
nand U12750 (N_12750,N_7199,N_6214);
or U12751 (N_12751,N_9492,N_5253);
or U12752 (N_12752,N_7241,N_7712);
xor U12753 (N_12753,N_5783,N_9830);
nor U12754 (N_12754,N_6849,N_5301);
nand U12755 (N_12755,N_7575,N_5391);
nor U12756 (N_12756,N_9517,N_9901);
nand U12757 (N_12757,N_5662,N_7198);
and U12758 (N_12758,N_7508,N_9872);
and U12759 (N_12759,N_6103,N_7515);
nor U12760 (N_12760,N_6653,N_5096);
nor U12761 (N_12761,N_8301,N_7277);
nand U12762 (N_12762,N_7654,N_8963);
and U12763 (N_12763,N_5541,N_8377);
xor U12764 (N_12764,N_6165,N_5815);
and U12765 (N_12765,N_5260,N_7274);
nand U12766 (N_12766,N_9584,N_6516);
and U12767 (N_12767,N_7091,N_6789);
or U12768 (N_12768,N_9499,N_5199);
xnor U12769 (N_12769,N_5315,N_9562);
nor U12770 (N_12770,N_9719,N_5370);
nor U12771 (N_12771,N_8113,N_6614);
nor U12772 (N_12772,N_9947,N_5326);
nor U12773 (N_12773,N_6253,N_6521);
xnor U12774 (N_12774,N_9249,N_7652);
xnor U12775 (N_12775,N_6390,N_8411);
or U12776 (N_12776,N_6611,N_9853);
or U12777 (N_12777,N_5893,N_8527);
xnor U12778 (N_12778,N_8351,N_5069);
and U12779 (N_12779,N_9661,N_6584);
nor U12780 (N_12780,N_9486,N_6962);
or U12781 (N_12781,N_7944,N_8808);
nor U12782 (N_12782,N_5437,N_8808);
and U12783 (N_12783,N_5669,N_9733);
nor U12784 (N_12784,N_5074,N_6375);
or U12785 (N_12785,N_7140,N_7229);
nand U12786 (N_12786,N_7277,N_7041);
nand U12787 (N_12787,N_8282,N_8902);
nand U12788 (N_12788,N_8600,N_7547);
xnor U12789 (N_12789,N_5524,N_9012);
or U12790 (N_12790,N_8614,N_5423);
nand U12791 (N_12791,N_6120,N_7823);
xnor U12792 (N_12792,N_6192,N_5106);
nor U12793 (N_12793,N_5896,N_6489);
xnor U12794 (N_12794,N_9264,N_9683);
or U12795 (N_12795,N_6893,N_6567);
nor U12796 (N_12796,N_8372,N_9107);
xnor U12797 (N_12797,N_9603,N_7935);
xnor U12798 (N_12798,N_6747,N_8745);
or U12799 (N_12799,N_8910,N_6726);
nor U12800 (N_12800,N_7172,N_8413);
nor U12801 (N_12801,N_8234,N_7457);
nor U12802 (N_12802,N_7575,N_5623);
or U12803 (N_12803,N_5076,N_8908);
and U12804 (N_12804,N_8656,N_6885);
nor U12805 (N_12805,N_9543,N_9038);
and U12806 (N_12806,N_6996,N_5951);
nor U12807 (N_12807,N_7344,N_9872);
and U12808 (N_12808,N_6863,N_5055);
nand U12809 (N_12809,N_5587,N_5802);
nor U12810 (N_12810,N_8211,N_8892);
nor U12811 (N_12811,N_5822,N_9277);
and U12812 (N_12812,N_9706,N_7492);
xnor U12813 (N_12813,N_5777,N_8159);
and U12814 (N_12814,N_7956,N_5878);
and U12815 (N_12815,N_5089,N_9157);
and U12816 (N_12816,N_6652,N_7091);
xor U12817 (N_12817,N_6022,N_7798);
nand U12818 (N_12818,N_6755,N_8647);
and U12819 (N_12819,N_8998,N_8709);
or U12820 (N_12820,N_6617,N_7408);
and U12821 (N_12821,N_5299,N_6393);
and U12822 (N_12822,N_6540,N_8129);
nor U12823 (N_12823,N_7777,N_8008);
nand U12824 (N_12824,N_5559,N_5523);
nor U12825 (N_12825,N_9101,N_8866);
and U12826 (N_12826,N_6933,N_9856);
nand U12827 (N_12827,N_7765,N_7904);
or U12828 (N_12828,N_9537,N_9148);
and U12829 (N_12829,N_6141,N_6140);
and U12830 (N_12830,N_9556,N_5576);
nand U12831 (N_12831,N_5693,N_5154);
or U12832 (N_12832,N_5485,N_9432);
and U12833 (N_12833,N_6811,N_6855);
nor U12834 (N_12834,N_8821,N_6161);
or U12835 (N_12835,N_6665,N_5744);
or U12836 (N_12836,N_9380,N_8398);
and U12837 (N_12837,N_5305,N_9308);
nand U12838 (N_12838,N_5375,N_8988);
nand U12839 (N_12839,N_7489,N_5020);
nand U12840 (N_12840,N_9898,N_9506);
xnor U12841 (N_12841,N_5442,N_7147);
nand U12842 (N_12842,N_6638,N_7584);
or U12843 (N_12843,N_9974,N_6485);
and U12844 (N_12844,N_8522,N_8912);
or U12845 (N_12845,N_6930,N_5383);
and U12846 (N_12846,N_6271,N_8094);
or U12847 (N_12847,N_5970,N_8497);
nand U12848 (N_12848,N_8580,N_5210);
nor U12849 (N_12849,N_5509,N_8163);
or U12850 (N_12850,N_8748,N_6200);
or U12851 (N_12851,N_9401,N_6175);
or U12852 (N_12852,N_6278,N_5803);
nand U12853 (N_12853,N_9734,N_6332);
or U12854 (N_12854,N_9132,N_6499);
nor U12855 (N_12855,N_5149,N_7886);
nand U12856 (N_12856,N_8688,N_5212);
nand U12857 (N_12857,N_8527,N_6136);
nor U12858 (N_12858,N_6514,N_8501);
nor U12859 (N_12859,N_7399,N_5860);
nor U12860 (N_12860,N_5265,N_6168);
nand U12861 (N_12861,N_7829,N_5020);
nand U12862 (N_12862,N_6222,N_9195);
or U12863 (N_12863,N_7520,N_9820);
or U12864 (N_12864,N_8428,N_7707);
nand U12865 (N_12865,N_8728,N_9942);
nor U12866 (N_12866,N_9944,N_5498);
and U12867 (N_12867,N_9815,N_7075);
or U12868 (N_12868,N_9736,N_9108);
nand U12869 (N_12869,N_7565,N_8281);
and U12870 (N_12870,N_5649,N_5901);
nand U12871 (N_12871,N_9784,N_7424);
nor U12872 (N_12872,N_8744,N_8755);
nand U12873 (N_12873,N_7204,N_9994);
or U12874 (N_12874,N_8967,N_8056);
and U12875 (N_12875,N_6396,N_8837);
nor U12876 (N_12876,N_8739,N_9501);
or U12877 (N_12877,N_9301,N_6787);
nand U12878 (N_12878,N_8755,N_7338);
or U12879 (N_12879,N_8581,N_9805);
nor U12880 (N_12880,N_6235,N_8513);
nor U12881 (N_12881,N_7442,N_9244);
and U12882 (N_12882,N_5882,N_7895);
nor U12883 (N_12883,N_7631,N_7605);
nand U12884 (N_12884,N_5218,N_7939);
nor U12885 (N_12885,N_5816,N_5885);
nand U12886 (N_12886,N_6139,N_9171);
or U12887 (N_12887,N_6390,N_9205);
nor U12888 (N_12888,N_6575,N_5578);
nor U12889 (N_12889,N_8775,N_9271);
or U12890 (N_12890,N_8660,N_5354);
nor U12891 (N_12891,N_7284,N_5098);
or U12892 (N_12892,N_7019,N_6872);
and U12893 (N_12893,N_5985,N_6042);
and U12894 (N_12894,N_6542,N_6175);
nand U12895 (N_12895,N_7975,N_5171);
nand U12896 (N_12896,N_6062,N_5741);
or U12897 (N_12897,N_5381,N_9011);
and U12898 (N_12898,N_7736,N_5929);
nor U12899 (N_12899,N_7960,N_7183);
nor U12900 (N_12900,N_9700,N_8550);
or U12901 (N_12901,N_6635,N_5539);
nand U12902 (N_12902,N_7734,N_5311);
nor U12903 (N_12903,N_7740,N_8655);
or U12904 (N_12904,N_6563,N_6815);
nand U12905 (N_12905,N_5403,N_9452);
nor U12906 (N_12906,N_9854,N_7591);
and U12907 (N_12907,N_6127,N_9746);
or U12908 (N_12908,N_8581,N_9100);
nand U12909 (N_12909,N_8494,N_8350);
nand U12910 (N_12910,N_7459,N_6297);
nor U12911 (N_12911,N_9582,N_7637);
or U12912 (N_12912,N_7118,N_5771);
or U12913 (N_12913,N_7735,N_7097);
and U12914 (N_12914,N_6373,N_5022);
or U12915 (N_12915,N_8467,N_9768);
and U12916 (N_12916,N_6780,N_5743);
or U12917 (N_12917,N_9338,N_7033);
nor U12918 (N_12918,N_5550,N_9179);
nor U12919 (N_12919,N_7610,N_7007);
or U12920 (N_12920,N_7033,N_9511);
or U12921 (N_12921,N_7267,N_9803);
nand U12922 (N_12922,N_6256,N_7410);
or U12923 (N_12923,N_6413,N_7891);
and U12924 (N_12924,N_9416,N_6882);
xor U12925 (N_12925,N_8249,N_5825);
or U12926 (N_12926,N_8277,N_8903);
or U12927 (N_12927,N_9177,N_5087);
nand U12928 (N_12928,N_7686,N_8851);
or U12929 (N_12929,N_9130,N_7675);
or U12930 (N_12930,N_6182,N_8871);
or U12931 (N_12931,N_8985,N_6605);
and U12932 (N_12932,N_7063,N_7603);
and U12933 (N_12933,N_6339,N_5293);
and U12934 (N_12934,N_6445,N_5072);
or U12935 (N_12935,N_6536,N_7215);
nor U12936 (N_12936,N_9872,N_9341);
nor U12937 (N_12937,N_8262,N_8546);
and U12938 (N_12938,N_8337,N_8583);
or U12939 (N_12939,N_7946,N_5704);
or U12940 (N_12940,N_9684,N_8824);
xor U12941 (N_12941,N_8268,N_9937);
nor U12942 (N_12942,N_7385,N_9627);
nor U12943 (N_12943,N_7170,N_8800);
xor U12944 (N_12944,N_8155,N_6341);
or U12945 (N_12945,N_5588,N_5362);
nor U12946 (N_12946,N_9206,N_9455);
or U12947 (N_12947,N_7370,N_7781);
or U12948 (N_12948,N_7214,N_5052);
and U12949 (N_12949,N_9853,N_8874);
nand U12950 (N_12950,N_9231,N_8282);
nand U12951 (N_12951,N_6656,N_7961);
or U12952 (N_12952,N_5530,N_7478);
nand U12953 (N_12953,N_8663,N_7992);
xnor U12954 (N_12954,N_8249,N_8162);
nand U12955 (N_12955,N_8797,N_8742);
or U12956 (N_12956,N_8680,N_5567);
or U12957 (N_12957,N_6109,N_7790);
and U12958 (N_12958,N_7641,N_9677);
and U12959 (N_12959,N_6133,N_8614);
nor U12960 (N_12960,N_5988,N_9989);
nand U12961 (N_12961,N_5567,N_6403);
nor U12962 (N_12962,N_7666,N_5616);
nand U12963 (N_12963,N_8916,N_5800);
nand U12964 (N_12964,N_6511,N_9921);
xor U12965 (N_12965,N_7827,N_7844);
or U12966 (N_12966,N_5803,N_8627);
nand U12967 (N_12967,N_5952,N_8110);
nand U12968 (N_12968,N_5676,N_6299);
and U12969 (N_12969,N_6987,N_8699);
and U12970 (N_12970,N_7041,N_7128);
and U12971 (N_12971,N_6651,N_8741);
nand U12972 (N_12972,N_9814,N_8103);
and U12973 (N_12973,N_9014,N_7409);
and U12974 (N_12974,N_6913,N_7400);
xnor U12975 (N_12975,N_7530,N_8213);
xnor U12976 (N_12976,N_8152,N_7794);
nand U12977 (N_12977,N_5046,N_9307);
nor U12978 (N_12978,N_6639,N_8379);
nor U12979 (N_12979,N_6367,N_9650);
nor U12980 (N_12980,N_6170,N_9751);
and U12981 (N_12981,N_6208,N_6560);
nand U12982 (N_12982,N_6663,N_6458);
and U12983 (N_12983,N_9184,N_8721);
nor U12984 (N_12984,N_9427,N_9271);
nand U12985 (N_12985,N_9171,N_6945);
nor U12986 (N_12986,N_7672,N_9990);
nand U12987 (N_12987,N_7915,N_5799);
and U12988 (N_12988,N_6399,N_9851);
or U12989 (N_12989,N_6563,N_6115);
and U12990 (N_12990,N_7679,N_6714);
and U12991 (N_12991,N_7557,N_5245);
xnor U12992 (N_12992,N_7414,N_9720);
or U12993 (N_12993,N_8020,N_6419);
nand U12994 (N_12994,N_5103,N_9853);
nor U12995 (N_12995,N_8943,N_6752);
or U12996 (N_12996,N_6965,N_6913);
nor U12997 (N_12997,N_5481,N_7344);
nand U12998 (N_12998,N_9862,N_9384);
and U12999 (N_12999,N_9957,N_9048);
nor U13000 (N_13000,N_6930,N_6737);
nor U13001 (N_13001,N_7352,N_9904);
or U13002 (N_13002,N_6136,N_5285);
or U13003 (N_13003,N_6138,N_8185);
xnor U13004 (N_13004,N_6840,N_5204);
and U13005 (N_13005,N_6024,N_7052);
nor U13006 (N_13006,N_6583,N_5341);
or U13007 (N_13007,N_5686,N_5448);
and U13008 (N_13008,N_8281,N_8242);
or U13009 (N_13009,N_9961,N_6565);
or U13010 (N_13010,N_8018,N_7296);
nor U13011 (N_13011,N_7779,N_9445);
nor U13012 (N_13012,N_6574,N_9696);
or U13013 (N_13013,N_5123,N_7728);
and U13014 (N_13014,N_8118,N_7943);
or U13015 (N_13015,N_7084,N_9954);
or U13016 (N_13016,N_9024,N_5868);
or U13017 (N_13017,N_9035,N_8651);
nand U13018 (N_13018,N_5874,N_8710);
nor U13019 (N_13019,N_9173,N_9956);
nor U13020 (N_13020,N_9705,N_6308);
or U13021 (N_13021,N_7935,N_7285);
nand U13022 (N_13022,N_7164,N_6775);
nor U13023 (N_13023,N_6877,N_9443);
nor U13024 (N_13024,N_9669,N_8112);
nor U13025 (N_13025,N_9575,N_7714);
nand U13026 (N_13026,N_6960,N_9110);
nand U13027 (N_13027,N_9864,N_7494);
and U13028 (N_13028,N_5778,N_5219);
and U13029 (N_13029,N_7068,N_9941);
nand U13030 (N_13030,N_7131,N_9937);
and U13031 (N_13031,N_8089,N_6939);
xnor U13032 (N_13032,N_7383,N_6110);
nor U13033 (N_13033,N_8379,N_9370);
nand U13034 (N_13034,N_6695,N_5340);
nor U13035 (N_13035,N_6482,N_8231);
and U13036 (N_13036,N_7580,N_8498);
nand U13037 (N_13037,N_7327,N_8137);
or U13038 (N_13038,N_5669,N_7176);
nand U13039 (N_13039,N_9222,N_7263);
nor U13040 (N_13040,N_9820,N_5544);
nor U13041 (N_13041,N_8086,N_7267);
and U13042 (N_13042,N_8887,N_9749);
nor U13043 (N_13043,N_7524,N_9519);
xnor U13044 (N_13044,N_7442,N_7038);
nand U13045 (N_13045,N_7211,N_9721);
and U13046 (N_13046,N_6260,N_7763);
nor U13047 (N_13047,N_8067,N_6700);
nor U13048 (N_13048,N_6596,N_8235);
or U13049 (N_13049,N_7854,N_7305);
and U13050 (N_13050,N_6528,N_5816);
and U13051 (N_13051,N_8748,N_7231);
and U13052 (N_13052,N_7335,N_5176);
or U13053 (N_13053,N_6355,N_9125);
xnor U13054 (N_13054,N_8319,N_8705);
and U13055 (N_13055,N_8874,N_5728);
and U13056 (N_13056,N_8482,N_6858);
nor U13057 (N_13057,N_6147,N_5325);
or U13058 (N_13058,N_6404,N_5225);
xnor U13059 (N_13059,N_9365,N_8490);
xnor U13060 (N_13060,N_9448,N_5207);
nand U13061 (N_13061,N_6276,N_7970);
or U13062 (N_13062,N_5798,N_6962);
or U13063 (N_13063,N_5350,N_7243);
nor U13064 (N_13064,N_8579,N_8770);
nand U13065 (N_13065,N_7067,N_9179);
xor U13066 (N_13066,N_9236,N_5123);
and U13067 (N_13067,N_7677,N_8869);
nand U13068 (N_13068,N_8128,N_6376);
and U13069 (N_13069,N_7870,N_6025);
or U13070 (N_13070,N_5877,N_8480);
xor U13071 (N_13071,N_7815,N_7909);
and U13072 (N_13072,N_7496,N_8164);
nor U13073 (N_13073,N_8558,N_8417);
or U13074 (N_13074,N_7746,N_9282);
nand U13075 (N_13075,N_6980,N_7205);
and U13076 (N_13076,N_6935,N_9926);
nand U13077 (N_13077,N_7188,N_5954);
or U13078 (N_13078,N_7151,N_6787);
nand U13079 (N_13079,N_8516,N_5331);
and U13080 (N_13080,N_8119,N_5120);
nand U13081 (N_13081,N_5938,N_7153);
or U13082 (N_13082,N_9528,N_5959);
and U13083 (N_13083,N_8601,N_7644);
nand U13084 (N_13084,N_7685,N_7569);
nand U13085 (N_13085,N_6221,N_5442);
and U13086 (N_13086,N_7817,N_9435);
nor U13087 (N_13087,N_9949,N_6336);
and U13088 (N_13088,N_8712,N_9640);
nand U13089 (N_13089,N_6563,N_8653);
nand U13090 (N_13090,N_9269,N_8433);
and U13091 (N_13091,N_8793,N_8668);
or U13092 (N_13092,N_7997,N_7056);
and U13093 (N_13093,N_7782,N_5433);
and U13094 (N_13094,N_8240,N_5596);
or U13095 (N_13095,N_5356,N_8701);
and U13096 (N_13096,N_5812,N_5193);
nand U13097 (N_13097,N_5327,N_5555);
and U13098 (N_13098,N_9123,N_8543);
or U13099 (N_13099,N_5808,N_6682);
nor U13100 (N_13100,N_6114,N_5962);
or U13101 (N_13101,N_8988,N_9573);
or U13102 (N_13102,N_5082,N_8645);
and U13103 (N_13103,N_7387,N_8574);
and U13104 (N_13104,N_5933,N_6183);
nor U13105 (N_13105,N_5100,N_6046);
nand U13106 (N_13106,N_9851,N_6236);
nor U13107 (N_13107,N_9041,N_7919);
or U13108 (N_13108,N_5234,N_9982);
or U13109 (N_13109,N_5266,N_9022);
nand U13110 (N_13110,N_5863,N_8265);
nand U13111 (N_13111,N_7173,N_6283);
and U13112 (N_13112,N_8039,N_7639);
or U13113 (N_13113,N_7541,N_7936);
nor U13114 (N_13114,N_6916,N_7269);
nor U13115 (N_13115,N_9323,N_6764);
nand U13116 (N_13116,N_9765,N_6032);
nor U13117 (N_13117,N_9849,N_6259);
or U13118 (N_13118,N_9039,N_5115);
nor U13119 (N_13119,N_9930,N_5581);
nor U13120 (N_13120,N_8005,N_7704);
or U13121 (N_13121,N_7310,N_5735);
and U13122 (N_13122,N_7682,N_7047);
nand U13123 (N_13123,N_6951,N_8198);
and U13124 (N_13124,N_8782,N_5515);
nor U13125 (N_13125,N_5406,N_8910);
nand U13126 (N_13126,N_8363,N_6335);
or U13127 (N_13127,N_7679,N_5303);
nor U13128 (N_13128,N_5381,N_5230);
and U13129 (N_13129,N_9946,N_5419);
and U13130 (N_13130,N_8956,N_7077);
and U13131 (N_13131,N_8685,N_5318);
nand U13132 (N_13132,N_7851,N_7281);
nor U13133 (N_13133,N_7891,N_6193);
xor U13134 (N_13134,N_9233,N_8143);
and U13135 (N_13135,N_7990,N_5974);
nand U13136 (N_13136,N_7623,N_5115);
nand U13137 (N_13137,N_6230,N_8909);
nand U13138 (N_13138,N_5505,N_7844);
nand U13139 (N_13139,N_9485,N_6066);
or U13140 (N_13140,N_8588,N_7618);
nor U13141 (N_13141,N_5901,N_7252);
and U13142 (N_13142,N_6784,N_7957);
or U13143 (N_13143,N_8602,N_7020);
and U13144 (N_13144,N_5733,N_8713);
nand U13145 (N_13145,N_9661,N_7457);
or U13146 (N_13146,N_6716,N_6906);
and U13147 (N_13147,N_8390,N_8488);
or U13148 (N_13148,N_8272,N_7794);
and U13149 (N_13149,N_7080,N_8911);
and U13150 (N_13150,N_8150,N_8626);
nor U13151 (N_13151,N_9375,N_7943);
nand U13152 (N_13152,N_7202,N_8695);
nor U13153 (N_13153,N_6158,N_5142);
or U13154 (N_13154,N_5506,N_9867);
and U13155 (N_13155,N_6773,N_8787);
nand U13156 (N_13156,N_8842,N_6957);
or U13157 (N_13157,N_8744,N_9891);
nand U13158 (N_13158,N_6440,N_5516);
nand U13159 (N_13159,N_8258,N_6821);
nand U13160 (N_13160,N_9490,N_9949);
nor U13161 (N_13161,N_5159,N_5606);
nand U13162 (N_13162,N_7245,N_8117);
nor U13163 (N_13163,N_7938,N_7578);
nor U13164 (N_13164,N_5847,N_6328);
or U13165 (N_13165,N_8112,N_8951);
nor U13166 (N_13166,N_9531,N_8049);
nand U13167 (N_13167,N_5775,N_9123);
or U13168 (N_13168,N_9915,N_5809);
nor U13169 (N_13169,N_5355,N_8617);
xnor U13170 (N_13170,N_8727,N_6854);
or U13171 (N_13171,N_8398,N_8264);
nor U13172 (N_13172,N_6244,N_9135);
or U13173 (N_13173,N_7344,N_9674);
and U13174 (N_13174,N_8541,N_7834);
or U13175 (N_13175,N_6199,N_5160);
nor U13176 (N_13176,N_7328,N_8072);
and U13177 (N_13177,N_8439,N_9275);
and U13178 (N_13178,N_5372,N_7688);
or U13179 (N_13179,N_7596,N_8700);
nor U13180 (N_13180,N_6033,N_6589);
nand U13181 (N_13181,N_6579,N_6436);
nand U13182 (N_13182,N_8848,N_6648);
and U13183 (N_13183,N_7356,N_8537);
nand U13184 (N_13184,N_8158,N_6455);
and U13185 (N_13185,N_9057,N_9330);
nor U13186 (N_13186,N_5135,N_6680);
and U13187 (N_13187,N_6180,N_5118);
or U13188 (N_13188,N_9722,N_8314);
nor U13189 (N_13189,N_9172,N_8251);
or U13190 (N_13190,N_9032,N_5423);
or U13191 (N_13191,N_5093,N_7465);
nor U13192 (N_13192,N_5184,N_6751);
nor U13193 (N_13193,N_5918,N_6896);
xor U13194 (N_13194,N_7087,N_9519);
and U13195 (N_13195,N_8315,N_5447);
or U13196 (N_13196,N_8944,N_7552);
nor U13197 (N_13197,N_5152,N_6576);
xor U13198 (N_13198,N_8294,N_5496);
nand U13199 (N_13199,N_6139,N_8316);
nand U13200 (N_13200,N_9389,N_5269);
nand U13201 (N_13201,N_7565,N_9064);
nor U13202 (N_13202,N_9072,N_5628);
xnor U13203 (N_13203,N_5486,N_8171);
nor U13204 (N_13204,N_9051,N_9860);
xnor U13205 (N_13205,N_5468,N_9480);
or U13206 (N_13206,N_5705,N_9082);
nor U13207 (N_13207,N_7640,N_5985);
or U13208 (N_13208,N_8579,N_9068);
and U13209 (N_13209,N_8690,N_5000);
nand U13210 (N_13210,N_6614,N_5120);
nor U13211 (N_13211,N_6748,N_6205);
nand U13212 (N_13212,N_5173,N_8357);
nor U13213 (N_13213,N_9942,N_8999);
nor U13214 (N_13214,N_5582,N_5277);
and U13215 (N_13215,N_5086,N_6991);
nand U13216 (N_13216,N_6863,N_5659);
nor U13217 (N_13217,N_6519,N_7928);
and U13218 (N_13218,N_7394,N_5269);
or U13219 (N_13219,N_8365,N_6929);
or U13220 (N_13220,N_7093,N_6174);
and U13221 (N_13221,N_9872,N_8137);
nor U13222 (N_13222,N_9933,N_6617);
nor U13223 (N_13223,N_7135,N_5433);
nor U13224 (N_13224,N_8480,N_9178);
nand U13225 (N_13225,N_6336,N_6080);
nand U13226 (N_13226,N_6820,N_5178);
nand U13227 (N_13227,N_9507,N_9960);
or U13228 (N_13228,N_5549,N_8637);
nand U13229 (N_13229,N_7136,N_5305);
and U13230 (N_13230,N_7766,N_5557);
nand U13231 (N_13231,N_6082,N_6262);
nand U13232 (N_13232,N_6420,N_8036);
nor U13233 (N_13233,N_9519,N_7810);
or U13234 (N_13234,N_5399,N_9390);
nand U13235 (N_13235,N_8624,N_7204);
or U13236 (N_13236,N_7275,N_9594);
or U13237 (N_13237,N_8854,N_8992);
nand U13238 (N_13238,N_8781,N_6954);
nand U13239 (N_13239,N_6712,N_7767);
and U13240 (N_13240,N_6109,N_9701);
nor U13241 (N_13241,N_9764,N_9115);
nor U13242 (N_13242,N_9133,N_6991);
nand U13243 (N_13243,N_7078,N_7244);
xnor U13244 (N_13244,N_7120,N_5421);
nor U13245 (N_13245,N_8867,N_7241);
and U13246 (N_13246,N_5485,N_5111);
nor U13247 (N_13247,N_8362,N_7306);
nand U13248 (N_13248,N_7098,N_6826);
nor U13249 (N_13249,N_5525,N_7596);
or U13250 (N_13250,N_9038,N_7730);
nand U13251 (N_13251,N_9807,N_8605);
and U13252 (N_13252,N_8299,N_7764);
nand U13253 (N_13253,N_6791,N_5463);
nand U13254 (N_13254,N_7175,N_7901);
nor U13255 (N_13255,N_7330,N_8108);
nor U13256 (N_13256,N_7205,N_5302);
nand U13257 (N_13257,N_9971,N_7072);
nand U13258 (N_13258,N_8338,N_6399);
or U13259 (N_13259,N_7216,N_7618);
or U13260 (N_13260,N_9285,N_9376);
nor U13261 (N_13261,N_8848,N_7648);
nor U13262 (N_13262,N_8329,N_7483);
or U13263 (N_13263,N_9553,N_5526);
xnor U13264 (N_13264,N_9206,N_6315);
nand U13265 (N_13265,N_8372,N_9275);
nor U13266 (N_13266,N_8430,N_6149);
or U13267 (N_13267,N_6098,N_7134);
and U13268 (N_13268,N_7374,N_8090);
and U13269 (N_13269,N_6228,N_6691);
or U13270 (N_13270,N_9355,N_6518);
nor U13271 (N_13271,N_9791,N_8397);
xnor U13272 (N_13272,N_7652,N_9876);
or U13273 (N_13273,N_8889,N_6422);
nand U13274 (N_13274,N_8301,N_7459);
nor U13275 (N_13275,N_7938,N_8564);
nor U13276 (N_13276,N_6920,N_5203);
or U13277 (N_13277,N_9736,N_7389);
and U13278 (N_13278,N_8647,N_8916);
nand U13279 (N_13279,N_8391,N_7862);
xnor U13280 (N_13280,N_6312,N_9867);
and U13281 (N_13281,N_8276,N_8234);
nand U13282 (N_13282,N_5877,N_7725);
nor U13283 (N_13283,N_9304,N_7044);
nor U13284 (N_13284,N_6318,N_7013);
nand U13285 (N_13285,N_6339,N_5916);
nor U13286 (N_13286,N_9967,N_6581);
or U13287 (N_13287,N_8829,N_5780);
xor U13288 (N_13288,N_6080,N_7191);
and U13289 (N_13289,N_5308,N_8022);
xnor U13290 (N_13290,N_6452,N_5913);
nand U13291 (N_13291,N_9809,N_9357);
nor U13292 (N_13292,N_5250,N_5143);
and U13293 (N_13293,N_5211,N_8317);
nand U13294 (N_13294,N_6919,N_6563);
and U13295 (N_13295,N_6474,N_8278);
and U13296 (N_13296,N_7978,N_9683);
nand U13297 (N_13297,N_8441,N_7678);
and U13298 (N_13298,N_6644,N_8501);
nand U13299 (N_13299,N_5707,N_8760);
or U13300 (N_13300,N_5000,N_7217);
and U13301 (N_13301,N_7840,N_5588);
nor U13302 (N_13302,N_8602,N_9505);
xor U13303 (N_13303,N_6599,N_6243);
and U13304 (N_13304,N_5617,N_9436);
or U13305 (N_13305,N_6402,N_7040);
nor U13306 (N_13306,N_9533,N_7993);
nor U13307 (N_13307,N_5517,N_6238);
nor U13308 (N_13308,N_5023,N_9211);
and U13309 (N_13309,N_6078,N_5039);
and U13310 (N_13310,N_8896,N_7212);
and U13311 (N_13311,N_5138,N_7453);
nand U13312 (N_13312,N_8641,N_5946);
xnor U13313 (N_13313,N_6924,N_5617);
nand U13314 (N_13314,N_6191,N_6562);
or U13315 (N_13315,N_9177,N_5063);
or U13316 (N_13316,N_6899,N_9695);
nand U13317 (N_13317,N_8355,N_7054);
nand U13318 (N_13318,N_7647,N_5219);
or U13319 (N_13319,N_7739,N_5916);
or U13320 (N_13320,N_8404,N_6602);
nand U13321 (N_13321,N_8706,N_5217);
nand U13322 (N_13322,N_7861,N_6231);
or U13323 (N_13323,N_8275,N_7384);
nand U13324 (N_13324,N_7650,N_6075);
nor U13325 (N_13325,N_9224,N_7439);
or U13326 (N_13326,N_8674,N_9657);
or U13327 (N_13327,N_9809,N_7296);
nor U13328 (N_13328,N_7404,N_5563);
or U13329 (N_13329,N_7525,N_8661);
or U13330 (N_13330,N_7259,N_5033);
or U13331 (N_13331,N_9722,N_7667);
nand U13332 (N_13332,N_9460,N_5708);
or U13333 (N_13333,N_9393,N_9956);
nor U13334 (N_13334,N_5759,N_8106);
or U13335 (N_13335,N_7148,N_5687);
or U13336 (N_13336,N_9568,N_6310);
nor U13337 (N_13337,N_5544,N_7379);
or U13338 (N_13338,N_9423,N_7097);
nor U13339 (N_13339,N_7640,N_7371);
and U13340 (N_13340,N_9071,N_9050);
or U13341 (N_13341,N_8291,N_5998);
or U13342 (N_13342,N_6824,N_6715);
nand U13343 (N_13343,N_6042,N_5578);
and U13344 (N_13344,N_5700,N_5077);
nor U13345 (N_13345,N_5834,N_5145);
or U13346 (N_13346,N_8487,N_6386);
or U13347 (N_13347,N_7118,N_5661);
and U13348 (N_13348,N_7335,N_8593);
xor U13349 (N_13349,N_5332,N_5233);
nand U13350 (N_13350,N_5165,N_5033);
and U13351 (N_13351,N_7416,N_7902);
and U13352 (N_13352,N_9664,N_8372);
or U13353 (N_13353,N_9358,N_8004);
nor U13354 (N_13354,N_8491,N_7490);
nand U13355 (N_13355,N_5224,N_9264);
and U13356 (N_13356,N_5825,N_8435);
or U13357 (N_13357,N_5198,N_9415);
nor U13358 (N_13358,N_7638,N_8574);
xor U13359 (N_13359,N_5429,N_5281);
nor U13360 (N_13360,N_6776,N_9622);
and U13361 (N_13361,N_8355,N_6631);
xor U13362 (N_13362,N_6025,N_8346);
nand U13363 (N_13363,N_8229,N_9376);
nor U13364 (N_13364,N_6050,N_8664);
or U13365 (N_13365,N_9084,N_8121);
and U13366 (N_13366,N_6511,N_7775);
nand U13367 (N_13367,N_9284,N_7652);
nand U13368 (N_13368,N_9557,N_8917);
nor U13369 (N_13369,N_6876,N_6404);
and U13370 (N_13370,N_8002,N_5954);
nor U13371 (N_13371,N_5697,N_5314);
or U13372 (N_13372,N_7320,N_8633);
and U13373 (N_13373,N_7534,N_9594);
nor U13374 (N_13374,N_7639,N_9859);
nor U13375 (N_13375,N_5151,N_5164);
nand U13376 (N_13376,N_5734,N_7830);
and U13377 (N_13377,N_8274,N_7193);
nor U13378 (N_13378,N_5222,N_8168);
xor U13379 (N_13379,N_7208,N_9117);
or U13380 (N_13380,N_5590,N_6078);
or U13381 (N_13381,N_6043,N_9980);
or U13382 (N_13382,N_9390,N_9131);
xnor U13383 (N_13383,N_5429,N_5235);
nor U13384 (N_13384,N_8988,N_8027);
nor U13385 (N_13385,N_6763,N_6813);
nand U13386 (N_13386,N_8144,N_9431);
nor U13387 (N_13387,N_9321,N_5563);
or U13388 (N_13388,N_7757,N_7930);
or U13389 (N_13389,N_6518,N_5117);
and U13390 (N_13390,N_6199,N_8756);
xnor U13391 (N_13391,N_5196,N_9925);
or U13392 (N_13392,N_6779,N_7430);
or U13393 (N_13393,N_9971,N_5598);
and U13394 (N_13394,N_7296,N_5198);
xor U13395 (N_13395,N_9764,N_7851);
or U13396 (N_13396,N_7391,N_8976);
nand U13397 (N_13397,N_9401,N_9172);
nand U13398 (N_13398,N_6217,N_8232);
xor U13399 (N_13399,N_5734,N_6405);
nor U13400 (N_13400,N_6937,N_8923);
nand U13401 (N_13401,N_5965,N_7504);
nor U13402 (N_13402,N_7807,N_6072);
xnor U13403 (N_13403,N_5383,N_5275);
and U13404 (N_13404,N_8712,N_8547);
nor U13405 (N_13405,N_8763,N_8592);
nand U13406 (N_13406,N_6652,N_6351);
and U13407 (N_13407,N_6032,N_6927);
and U13408 (N_13408,N_7251,N_8490);
nand U13409 (N_13409,N_9353,N_9889);
nor U13410 (N_13410,N_7651,N_6470);
or U13411 (N_13411,N_8541,N_7793);
nand U13412 (N_13412,N_9157,N_5921);
and U13413 (N_13413,N_5700,N_8051);
nor U13414 (N_13414,N_9125,N_8597);
nand U13415 (N_13415,N_5722,N_7764);
and U13416 (N_13416,N_8430,N_8786);
and U13417 (N_13417,N_7767,N_6760);
nor U13418 (N_13418,N_7371,N_5885);
nor U13419 (N_13419,N_9460,N_7327);
or U13420 (N_13420,N_6697,N_9198);
and U13421 (N_13421,N_5611,N_9822);
and U13422 (N_13422,N_9732,N_6166);
xor U13423 (N_13423,N_9931,N_5671);
nor U13424 (N_13424,N_8705,N_9571);
xnor U13425 (N_13425,N_9739,N_6024);
or U13426 (N_13426,N_9938,N_7620);
nand U13427 (N_13427,N_8651,N_6230);
or U13428 (N_13428,N_5145,N_7801);
nor U13429 (N_13429,N_6114,N_8809);
or U13430 (N_13430,N_7170,N_5654);
nor U13431 (N_13431,N_9354,N_7842);
xnor U13432 (N_13432,N_8891,N_7562);
nand U13433 (N_13433,N_6732,N_7589);
and U13434 (N_13434,N_6844,N_7391);
nor U13435 (N_13435,N_7046,N_7761);
nand U13436 (N_13436,N_9342,N_7700);
nand U13437 (N_13437,N_9977,N_6520);
nand U13438 (N_13438,N_7222,N_6011);
and U13439 (N_13439,N_8862,N_8160);
and U13440 (N_13440,N_9017,N_7025);
nor U13441 (N_13441,N_7961,N_6194);
nand U13442 (N_13442,N_8999,N_7400);
nor U13443 (N_13443,N_5311,N_5247);
and U13444 (N_13444,N_9490,N_6210);
or U13445 (N_13445,N_7947,N_6010);
nand U13446 (N_13446,N_5064,N_5799);
or U13447 (N_13447,N_6847,N_8851);
xnor U13448 (N_13448,N_5881,N_9032);
nand U13449 (N_13449,N_7659,N_8323);
nor U13450 (N_13450,N_8207,N_7675);
nand U13451 (N_13451,N_8715,N_6600);
or U13452 (N_13452,N_6506,N_5518);
nand U13453 (N_13453,N_9512,N_7393);
nor U13454 (N_13454,N_7690,N_7839);
nand U13455 (N_13455,N_9755,N_5267);
or U13456 (N_13456,N_8958,N_8027);
nand U13457 (N_13457,N_6837,N_6001);
or U13458 (N_13458,N_5349,N_9494);
and U13459 (N_13459,N_7722,N_7301);
or U13460 (N_13460,N_8378,N_6739);
and U13461 (N_13461,N_7272,N_5461);
and U13462 (N_13462,N_9170,N_7308);
or U13463 (N_13463,N_9317,N_6807);
and U13464 (N_13464,N_7980,N_9392);
and U13465 (N_13465,N_5514,N_9434);
or U13466 (N_13466,N_7082,N_6950);
nand U13467 (N_13467,N_8287,N_7452);
nand U13468 (N_13468,N_6147,N_6295);
and U13469 (N_13469,N_5639,N_7256);
xor U13470 (N_13470,N_5676,N_5107);
nand U13471 (N_13471,N_7739,N_9136);
or U13472 (N_13472,N_8127,N_7678);
or U13473 (N_13473,N_6730,N_8837);
nand U13474 (N_13474,N_6036,N_6353);
nor U13475 (N_13475,N_7888,N_6870);
or U13476 (N_13476,N_9382,N_9181);
nor U13477 (N_13477,N_9963,N_7264);
nor U13478 (N_13478,N_5790,N_8309);
xor U13479 (N_13479,N_8517,N_8349);
nor U13480 (N_13480,N_8512,N_8241);
nor U13481 (N_13481,N_5343,N_8778);
nor U13482 (N_13482,N_7232,N_8717);
nand U13483 (N_13483,N_9856,N_5680);
nand U13484 (N_13484,N_7016,N_7838);
and U13485 (N_13485,N_7101,N_7601);
and U13486 (N_13486,N_6673,N_5264);
nand U13487 (N_13487,N_6063,N_7041);
and U13488 (N_13488,N_7286,N_5840);
nand U13489 (N_13489,N_7671,N_7928);
nor U13490 (N_13490,N_6887,N_8044);
nand U13491 (N_13491,N_9343,N_9078);
and U13492 (N_13492,N_5884,N_5523);
nor U13493 (N_13493,N_7835,N_7135);
or U13494 (N_13494,N_7631,N_5448);
nand U13495 (N_13495,N_7096,N_5676);
nor U13496 (N_13496,N_8504,N_8930);
or U13497 (N_13497,N_6851,N_6653);
nor U13498 (N_13498,N_7845,N_6107);
or U13499 (N_13499,N_6530,N_9143);
nor U13500 (N_13500,N_7275,N_5983);
and U13501 (N_13501,N_7321,N_9594);
and U13502 (N_13502,N_8206,N_9625);
nand U13503 (N_13503,N_8056,N_6202);
nand U13504 (N_13504,N_9603,N_8876);
nand U13505 (N_13505,N_6648,N_8465);
and U13506 (N_13506,N_8340,N_8237);
and U13507 (N_13507,N_8180,N_8382);
nor U13508 (N_13508,N_7191,N_8497);
nor U13509 (N_13509,N_5857,N_6537);
nand U13510 (N_13510,N_7549,N_9232);
or U13511 (N_13511,N_7611,N_5721);
and U13512 (N_13512,N_9354,N_9843);
or U13513 (N_13513,N_9152,N_7376);
nand U13514 (N_13514,N_7937,N_8739);
or U13515 (N_13515,N_9552,N_7346);
xor U13516 (N_13516,N_5988,N_7365);
or U13517 (N_13517,N_9093,N_5176);
and U13518 (N_13518,N_9802,N_5459);
nor U13519 (N_13519,N_5270,N_7908);
and U13520 (N_13520,N_9099,N_7184);
nand U13521 (N_13521,N_9936,N_8848);
and U13522 (N_13522,N_8638,N_7906);
and U13523 (N_13523,N_5246,N_9931);
or U13524 (N_13524,N_8434,N_5962);
nor U13525 (N_13525,N_5264,N_8559);
or U13526 (N_13526,N_6685,N_7385);
or U13527 (N_13527,N_5815,N_6918);
nand U13528 (N_13528,N_7675,N_6479);
nand U13529 (N_13529,N_6319,N_9350);
or U13530 (N_13530,N_7996,N_7432);
xor U13531 (N_13531,N_8079,N_7219);
and U13532 (N_13532,N_7392,N_9459);
and U13533 (N_13533,N_9275,N_8852);
nand U13534 (N_13534,N_8338,N_7982);
nor U13535 (N_13535,N_9555,N_6271);
or U13536 (N_13536,N_7477,N_7210);
nor U13537 (N_13537,N_7832,N_9999);
or U13538 (N_13538,N_9457,N_7895);
nor U13539 (N_13539,N_9888,N_7928);
nand U13540 (N_13540,N_5273,N_9326);
or U13541 (N_13541,N_6028,N_8480);
and U13542 (N_13542,N_9409,N_9843);
nor U13543 (N_13543,N_7188,N_6297);
nand U13544 (N_13544,N_5222,N_6280);
nor U13545 (N_13545,N_7329,N_8596);
and U13546 (N_13546,N_8961,N_5488);
nor U13547 (N_13547,N_8632,N_6483);
and U13548 (N_13548,N_9498,N_9536);
nand U13549 (N_13549,N_6075,N_9850);
or U13550 (N_13550,N_6137,N_9515);
nand U13551 (N_13551,N_9163,N_6641);
and U13552 (N_13552,N_5530,N_5570);
and U13553 (N_13553,N_7909,N_6282);
and U13554 (N_13554,N_5141,N_9550);
or U13555 (N_13555,N_9177,N_7600);
nor U13556 (N_13556,N_9058,N_7469);
nor U13557 (N_13557,N_7994,N_9114);
or U13558 (N_13558,N_5849,N_9849);
xnor U13559 (N_13559,N_7052,N_6506);
nand U13560 (N_13560,N_5821,N_5049);
and U13561 (N_13561,N_7842,N_9789);
nand U13562 (N_13562,N_6251,N_5993);
or U13563 (N_13563,N_8722,N_7474);
and U13564 (N_13564,N_5844,N_5127);
nand U13565 (N_13565,N_8373,N_5900);
nand U13566 (N_13566,N_5180,N_9861);
nor U13567 (N_13567,N_9399,N_7171);
nor U13568 (N_13568,N_5137,N_9377);
and U13569 (N_13569,N_7354,N_5310);
nor U13570 (N_13570,N_9103,N_9675);
nor U13571 (N_13571,N_9565,N_8873);
nor U13572 (N_13572,N_7899,N_7503);
or U13573 (N_13573,N_5070,N_8885);
nand U13574 (N_13574,N_9882,N_6567);
or U13575 (N_13575,N_8833,N_5514);
or U13576 (N_13576,N_8936,N_9547);
and U13577 (N_13577,N_6411,N_8396);
xor U13578 (N_13578,N_7517,N_9956);
nand U13579 (N_13579,N_9508,N_5337);
nand U13580 (N_13580,N_6676,N_9133);
or U13581 (N_13581,N_9921,N_6634);
nor U13582 (N_13582,N_8185,N_9369);
nand U13583 (N_13583,N_9297,N_8334);
nor U13584 (N_13584,N_7353,N_7401);
nand U13585 (N_13585,N_5533,N_9608);
and U13586 (N_13586,N_8329,N_6620);
xnor U13587 (N_13587,N_6130,N_6338);
or U13588 (N_13588,N_9521,N_7927);
nor U13589 (N_13589,N_8557,N_5906);
and U13590 (N_13590,N_6586,N_6116);
xor U13591 (N_13591,N_5721,N_7719);
and U13592 (N_13592,N_5400,N_9511);
nand U13593 (N_13593,N_9257,N_6788);
xnor U13594 (N_13594,N_6911,N_7850);
xor U13595 (N_13595,N_5110,N_5895);
or U13596 (N_13596,N_7860,N_9053);
nand U13597 (N_13597,N_5471,N_9492);
and U13598 (N_13598,N_8107,N_5500);
or U13599 (N_13599,N_6003,N_6840);
nor U13600 (N_13600,N_7170,N_5926);
nand U13601 (N_13601,N_9691,N_5876);
nor U13602 (N_13602,N_8947,N_5083);
nand U13603 (N_13603,N_9098,N_9822);
or U13604 (N_13604,N_5252,N_5273);
nor U13605 (N_13605,N_8500,N_7258);
xnor U13606 (N_13606,N_7586,N_7423);
nand U13607 (N_13607,N_6010,N_6962);
nor U13608 (N_13608,N_9301,N_8788);
nand U13609 (N_13609,N_9422,N_9858);
xnor U13610 (N_13610,N_7753,N_7140);
nand U13611 (N_13611,N_9584,N_6955);
or U13612 (N_13612,N_8399,N_6029);
and U13613 (N_13613,N_7670,N_9433);
nor U13614 (N_13614,N_8034,N_7274);
and U13615 (N_13615,N_9152,N_5325);
nand U13616 (N_13616,N_9245,N_8505);
and U13617 (N_13617,N_8851,N_5669);
or U13618 (N_13618,N_9226,N_7750);
nand U13619 (N_13619,N_9256,N_7776);
xnor U13620 (N_13620,N_7425,N_9404);
and U13621 (N_13621,N_6960,N_8917);
and U13622 (N_13622,N_6619,N_5712);
or U13623 (N_13623,N_8795,N_9803);
and U13624 (N_13624,N_5499,N_8240);
nor U13625 (N_13625,N_6063,N_8093);
nor U13626 (N_13626,N_7313,N_6116);
nand U13627 (N_13627,N_5476,N_8723);
nor U13628 (N_13628,N_8280,N_9186);
or U13629 (N_13629,N_8236,N_6295);
xnor U13630 (N_13630,N_6892,N_7640);
xor U13631 (N_13631,N_7084,N_7163);
nand U13632 (N_13632,N_9775,N_7160);
and U13633 (N_13633,N_9313,N_7084);
nand U13634 (N_13634,N_5867,N_5401);
nor U13635 (N_13635,N_5913,N_6059);
nor U13636 (N_13636,N_9657,N_7294);
nor U13637 (N_13637,N_6184,N_7720);
or U13638 (N_13638,N_9004,N_5819);
nand U13639 (N_13639,N_6921,N_5926);
and U13640 (N_13640,N_9053,N_9168);
nand U13641 (N_13641,N_8831,N_9907);
and U13642 (N_13642,N_8980,N_8329);
nand U13643 (N_13643,N_6832,N_9019);
or U13644 (N_13644,N_8744,N_8053);
nor U13645 (N_13645,N_8115,N_5432);
nand U13646 (N_13646,N_6918,N_5410);
and U13647 (N_13647,N_8172,N_6260);
and U13648 (N_13648,N_5328,N_7066);
nand U13649 (N_13649,N_8130,N_9636);
nand U13650 (N_13650,N_7058,N_5507);
nand U13651 (N_13651,N_5581,N_8906);
xnor U13652 (N_13652,N_8788,N_9116);
and U13653 (N_13653,N_7805,N_9111);
and U13654 (N_13654,N_5574,N_9813);
or U13655 (N_13655,N_8280,N_7341);
or U13656 (N_13656,N_6701,N_9931);
or U13657 (N_13657,N_5439,N_8344);
nand U13658 (N_13658,N_5178,N_5923);
nor U13659 (N_13659,N_5615,N_8962);
and U13660 (N_13660,N_6622,N_5044);
or U13661 (N_13661,N_5160,N_7025);
or U13662 (N_13662,N_6743,N_9857);
or U13663 (N_13663,N_8644,N_9648);
nor U13664 (N_13664,N_6763,N_7462);
or U13665 (N_13665,N_9450,N_8922);
nor U13666 (N_13666,N_8165,N_6283);
or U13667 (N_13667,N_6237,N_9079);
or U13668 (N_13668,N_5825,N_8336);
and U13669 (N_13669,N_6733,N_9671);
nand U13670 (N_13670,N_9167,N_9658);
and U13671 (N_13671,N_5667,N_6469);
nor U13672 (N_13672,N_6803,N_5925);
and U13673 (N_13673,N_8349,N_7355);
nor U13674 (N_13674,N_5788,N_7988);
or U13675 (N_13675,N_9797,N_6431);
and U13676 (N_13676,N_7488,N_5797);
and U13677 (N_13677,N_7925,N_6350);
nor U13678 (N_13678,N_8403,N_9007);
nor U13679 (N_13679,N_7450,N_5714);
and U13680 (N_13680,N_6208,N_5209);
nor U13681 (N_13681,N_8432,N_6626);
and U13682 (N_13682,N_6947,N_9446);
and U13683 (N_13683,N_7259,N_8006);
xnor U13684 (N_13684,N_7840,N_9128);
and U13685 (N_13685,N_7240,N_6154);
and U13686 (N_13686,N_5685,N_9631);
or U13687 (N_13687,N_7013,N_7288);
or U13688 (N_13688,N_6594,N_9661);
xnor U13689 (N_13689,N_5167,N_5653);
nor U13690 (N_13690,N_8659,N_7782);
nand U13691 (N_13691,N_7587,N_8663);
or U13692 (N_13692,N_9183,N_8634);
nand U13693 (N_13693,N_9830,N_5418);
or U13694 (N_13694,N_8697,N_5474);
xor U13695 (N_13695,N_5587,N_9998);
xnor U13696 (N_13696,N_7007,N_9794);
or U13697 (N_13697,N_6832,N_5432);
xor U13698 (N_13698,N_7408,N_6117);
or U13699 (N_13699,N_5685,N_6641);
nand U13700 (N_13700,N_6379,N_6727);
nand U13701 (N_13701,N_6965,N_6589);
nand U13702 (N_13702,N_5610,N_9402);
or U13703 (N_13703,N_5849,N_8946);
xnor U13704 (N_13704,N_6815,N_5839);
and U13705 (N_13705,N_6132,N_6608);
nor U13706 (N_13706,N_9697,N_5680);
and U13707 (N_13707,N_6917,N_8749);
nand U13708 (N_13708,N_9715,N_8239);
and U13709 (N_13709,N_5034,N_5435);
or U13710 (N_13710,N_7268,N_8304);
and U13711 (N_13711,N_5314,N_8266);
nor U13712 (N_13712,N_9699,N_8625);
nand U13713 (N_13713,N_6390,N_6401);
nand U13714 (N_13714,N_8990,N_9019);
or U13715 (N_13715,N_9523,N_8354);
nand U13716 (N_13716,N_8783,N_8509);
nand U13717 (N_13717,N_8281,N_7071);
or U13718 (N_13718,N_9556,N_5427);
or U13719 (N_13719,N_7793,N_9188);
or U13720 (N_13720,N_6942,N_8536);
or U13721 (N_13721,N_8823,N_7551);
nand U13722 (N_13722,N_8738,N_7565);
and U13723 (N_13723,N_8613,N_7438);
or U13724 (N_13724,N_7061,N_7506);
or U13725 (N_13725,N_6564,N_9893);
xor U13726 (N_13726,N_8535,N_8594);
or U13727 (N_13727,N_8066,N_6206);
nand U13728 (N_13728,N_8246,N_8890);
xnor U13729 (N_13729,N_7326,N_9074);
and U13730 (N_13730,N_6367,N_8194);
nand U13731 (N_13731,N_6669,N_6833);
nand U13732 (N_13732,N_8574,N_5611);
nor U13733 (N_13733,N_8499,N_7320);
nand U13734 (N_13734,N_6502,N_8181);
or U13735 (N_13735,N_8979,N_8180);
nor U13736 (N_13736,N_9739,N_8160);
xnor U13737 (N_13737,N_7145,N_5497);
xnor U13738 (N_13738,N_9318,N_7554);
and U13739 (N_13739,N_8444,N_7880);
nand U13740 (N_13740,N_9752,N_6721);
nor U13741 (N_13741,N_5705,N_9798);
nand U13742 (N_13742,N_6749,N_9457);
xnor U13743 (N_13743,N_7277,N_9300);
nand U13744 (N_13744,N_7142,N_6021);
and U13745 (N_13745,N_6996,N_6072);
nand U13746 (N_13746,N_6413,N_9823);
nand U13747 (N_13747,N_5814,N_9518);
and U13748 (N_13748,N_6103,N_9274);
and U13749 (N_13749,N_8698,N_7972);
nor U13750 (N_13750,N_7539,N_6974);
nor U13751 (N_13751,N_6900,N_5530);
nor U13752 (N_13752,N_9277,N_8737);
nor U13753 (N_13753,N_8249,N_8246);
and U13754 (N_13754,N_9111,N_6611);
or U13755 (N_13755,N_7703,N_5364);
and U13756 (N_13756,N_5893,N_5587);
nor U13757 (N_13757,N_7826,N_5049);
or U13758 (N_13758,N_9959,N_9224);
nand U13759 (N_13759,N_8882,N_5764);
or U13760 (N_13760,N_7825,N_8599);
nand U13761 (N_13761,N_6507,N_8293);
nor U13762 (N_13762,N_6294,N_7056);
and U13763 (N_13763,N_8588,N_5387);
or U13764 (N_13764,N_8823,N_9796);
nand U13765 (N_13765,N_7578,N_5599);
and U13766 (N_13766,N_9377,N_5704);
xnor U13767 (N_13767,N_9658,N_8057);
nor U13768 (N_13768,N_7270,N_9343);
nand U13769 (N_13769,N_6748,N_8490);
nor U13770 (N_13770,N_7832,N_8117);
and U13771 (N_13771,N_9408,N_8166);
and U13772 (N_13772,N_7646,N_5054);
or U13773 (N_13773,N_8607,N_7854);
nor U13774 (N_13774,N_5373,N_7167);
and U13775 (N_13775,N_6020,N_8888);
and U13776 (N_13776,N_9511,N_8784);
nor U13777 (N_13777,N_6646,N_9199);
or U13778 (N_13778,N_9319,N_7759);
and U13779 (N_13779,N_7998,N_7679);
or U13780 (N_13780,N_7833,N_9944);
nor U13781 (N_13781,N_6737,N_5913);
or U13782 (N_13782,N_7992,N_5254);
or U13783 (N_13783,N_8303,N_5083);
xnor U13784 (N_13784,N_7389,N_6805);
or U13785 (N_13785,N_6515,N_9041);
and U13786 (N_13786,N_8641,N_6709);
nor U13787 (N_13787,N_8513,N_8208);
nor U13788 (N_13788,N_9465,N_5462);
or U13789 (N_13789,N_8314,N_6299);
or U13790 (N_13790,N_6672,N_7874);
nand U13791 (N_13791,N_7146,N_9885);
and U13792 (N_13792,N_8726,N_9887);
nand U13793 (N_13793,N_9167,N_5723);
nor U13794 (N_13794,N_8726,N_8222);
and U13795 (N_13795,N_6477,N_8619);
and U13796 (N_13796,N_6192,N_5010);
nor U13797 (N_13797,N_8817,N_7807);
nand U13798 (N_13798,N_7799,N_7145);
and U13799 (N_13799,N_6560,N_7043);
nor U13800 (N_13800,N_7414,N_6201);
nand U13801 (N_13801,N_9505,N_8286);
nand U13802 (N_13802,N_9907,N_9865);
nor U13803 (N_13803,N_9523,N_7210);
and U13804 (N_13804,N_8361,N_9641);
nor U13805 (N_13805,N_8332,N_7755);
nor U13806 (N_13806,N_9765,N_7989);
nand U13807 (N_13807,N_8660,N_6750);
xnor U13808 (N_13808,N_9183,N_6072);
nor U13809 (N_13809,N_5520,N_8572);
nand U13810 (N_13810,N_9579,N_7852);
or U13811 (N_13811,N_8053,N_5693);
nand U13812 (N_13812,N_7673,N_5992);
nand U13813 (N_13813,N_7861,N_7930);
or U13814 (N_13814,N_8144,N_6454);
or U13815 (N_13815,N_7741,N_9979);
and U13816 (N_13816,N_9771,N_9308);
and U13817 (N_13817,N_9901,N_7107);
or U13818 (N_13818,N_6293,N_5838);
nand U13819 (N_13819,N_7537,N_5286);
xor U13820 (N_13820,N_6065,N_5789);
nand U13821 (N_13821,N_9143,N_5123);
nor U13822 (N_13822,N_9004,N_7359);
nand U13823 (N_13823,N_9551,N_9621);
or U13824 (N_13824,N_5788,N_7246);
nand U13825 (N_13825,N_7689,N_9512);
nor U13826 (N_13826,N_9380,N_9718);
and U13827 (N_13827,N_8854,N_9294);
nor U13828 (N_13828,N_8713,N_7846);
nor U13829 (N_13829,N_7277,N_6193);
and U13830 (N_13830,N_5210,N_6591);
or U13831 (N_13831,N_6894,N_9504);
or U13832 (N_13832,N_9605,N_8329);
nand U13833 (N_13833,N_9996,N_7150);
nand U13834 (N_13834,N_8626,N_7101);
xnor U13835 (N_13835,N_5401,N_7544);
nor U13836 (N_13836,N_9037,N_5223);
nor U13837 (N_13837,N_8473,N_6923);
and U13838 (N_13838,N_8937,N_9697);
or U13839 (N_13839,N_6871,N_5653);
and U13840 (N_13840,N_7286,N_7021);
nor U13841 (N_13841,N_8113,N_9671);
nand U13842 (N_13842,N_7769,N_7224);
nor U13843 (N_13843,N_9593,N_7596);
nor U13844 (N_13844,N_7529,N_6276);
or U13845 (N_13845,N_7948,N_7238);
and U13846 (N_13846,N_6281,N_8768);
or U13847 (N_13847,N_7988,N_5115);
nor U13848 (N_13848,N_5021,N_7884);
and U13849 (N_13849,N_6872,N_6347);
nand U13850 (N_13850,N_9807,N_9639);
or U13851 (N_13851,N_6716,N_5832);
nor U13852 (N_13852,N_6965,N_8888);
and U13853 (N_13853,N_5039,N_5863);
or U13854 (N_13854,N_6392,N_7452);
and U13855 (N_13855,N_9715,N_5772);
nor U13856 (N_13856,N_8931,N_8373);
nand U13857 (N_13857,N_5552,N_6561);
and U13858 (N_13858,N_8719,N_9178);
or U13859 (N_13859,N_5849,N_5465);
nand U13860 (N_13860,N_6335,N_6468);
nor U13861 (N_13861,N_5245,N_9846);
nor U13862 (N_13862,N_9699,N_8465);
or U13863 (N_13863,N_7969,N_5412);
and U13864 (N_13864,N_7277,N_8417);
or U13865 (N_13865,N_7262,N_9438);
or U13866 (N_13866,N_6152,N_7016);
nand U13867 (N_13867,N_6916,N_6774);
nor U13868 (N_13868,N_9728,N_9178);
nand U13869 (N_13869,N_8239,N_7743);
or U13870 (N_13870,N_8856,N_6835);
and U13871 (N_13871,N_5228,N_6542);
nor U13872 (N_13872,N_5911,N_9451);
nand U13873 (N_13873,N_8284,N_5169);
nand U13874 (N_13874,N_6708,N_7842);
nand U13875 (N_13875,N_9013,N_5488);
nand U13876 (N_13876,N_6243,N_8198);
nand U13877 (N_13877,N_8952,N_7098);
and U13878 (N_13878,N_7271,N_6167);
and U13879 (N_13879,N_6139,N_8540);
or U13880 (N_13880,N_5751,N_7857);
or U13881 (N_13881,N_6041,N_9198);
or U13882 (N_13882,N_6213,N_5509);
xnor U13883 (N_13883,N_6858,N_5905);
and U13884 (N_13884,N_6783,N_7341);
or U13885 (N_13885,N_7259,N_9727);
nand U13886 (N_13886,N_8090,N_6419);
nand U13887 (N_13887,N_6082,N_7107);
nor U13888 (N_13888,N_6795,N_7479);
xor U13889 (N_13889,N_9140,N_6168);
or U13890 (N_13890,N_5246,N_5644);
and U13891 (N_13891,N_5464,N_7383);
and U13892 (N_13892,N_7892,N_8114);
nor U13893 (N_13893,N_7822,N_6461);
and U13894 (N_13894,N_5225,N_7704);
nand U13895 (N_13895,N_7876,N_8611);
and U13896 (N_13896,N_5516,N_8023);
nand U13897 (N_13897,N_7971,N_6216);
nor U13898 (N_13898,N_5197,N_5241);
or U13899 (N_13899,N_5720,N_6166);
nor U13900 (N_13900,N_7576,N_8298);
nand U13901 (N_13901,N_7230,N_6418);
and U13902 (N_13902,N_7675,N_7235);
nor U13903 (N_13903,N_7902,N_5528);
and U13904 (N_13904,N_5627,N_9764);
nor U13905 (N_13905,N_6698,N_5459);
and U13906 (N_13906,N_9930,N_5849);
nand U13907 (N_13907,N_8113,N_7844);
nand U13908 (N_13908,N_7070,N_5666);
nor U13909 (N_13909,N_9224,N_8554);
or U13910 (N_13910,N_8009,N_9521);
nor U13911 (N_13911,N_7476,N_6012);
nor U13912 (N_13912,N_9253,N_7854);
nand U13913 (N_13913,N_6334,N_7182);
nor U13914 (N_13914,N_7587,N_6959);
or U13915 (N_13915,N_9524,N_6143);
and U13916 (N_13916,N_5188,N_6811);
or U13917 (N_13917,N_9269,N_7585);
or U13918 (N_13918,N_7571,N_9385);
and U13919 (N_13919,N_7087,N_8807);
nand U13920 (N_13920,N_7649,N_8550);
or U13921 (N_13921,N_7593,N_6410);
nand U13922 (N_13922,N_5079,N_8841);
or U13923 (N_13923,N_8792,N_9930);
xor U13924 (N_13924,N_9336,N_9660);
and U13925 (N_13925,N_5727,N_5375);
nor U13926 (N_13926,N_9597,N_8519);
xor U13927 (N_13927,N_9072,N_7407);
xnor U13928 (N_13928,N_7119,N_6690);
xor U13929 (N_13929,N_9023,N_9618);
nor U13930 (N_13930,N_9357,N_9382);
and U13931 (N_13931,N_5584,N_8732);
and U13932 (N_13932,N_6217,N_6495);
and U13933 (N_13933,N_8962,N_6929);
nand U13934 (N_13934,N_5926,N_6165);
nor U13935 (N_13935,N_7672,N_8362);
nand U13936 (N_13936,N_6935,N_9889);
nor U13937 (N_13937,N_7450,N_8684);
nor U13938 (N_13938,N_9061,N_6496);
and U13939 (N_13939,N_9686,N_6560);
and U13940 (N_13940,N_6688,N_5322);
and U13941 (N_13941,N_7716,N_6357);
nor U13942 (N_13942,N_9728,N_9003);
nor U13943 (N_13943,N_6305,N_7627);
or U13944 (N_13944,N_5384,N_9975);
nor U13945 (N_13945,N_5713,N_7888);
and U13946 (N_13946,N_8779,N_6330);
nand U13947 (N_13947,N_5039,N_9859);
nand U13948 (N_13948,N_8435,N_7505);
xor U13949 (N_13949,N_6350,N_6626);
nand U13950 (N_13950,N_6125,N_8494);
and U13951 (N_13951,N_6048,N_8959);
nor U13952 (N_13952,N_9867,N_9018);
xor U13953 (N_13953,N_8012,N_8231);
nor U13954 (N_13954,N_9454,N_5707);
or U13955 (N_13955,N_8800,N_5405);
nand U13956 (N_13956,N_7815,N_7771);
or U13957 (N_13957,N_9452,N_9068);
and U13958 (N_13958,N_8155,N_8867);
nor U13959 (N_13959,N_6120,N_7521);
or U13960 (N_13960,N_9751,N_8334);
or U13961 (N_13961,N_5444,N_9857);
nor U13962 (N_13962,N_5084,N_7972);
xnor U13963 (N_13963,N_5460,N_6311);
nand U13964 (N_13964,N_9248,N_8090);
nor U13965 (N_13965,N_6882,N_6619);
or U13966 (N_13966,N_8904,N_6788);
and U13967 (N_13967,N_5152,N_5772);
nor U13968 (N_13968,N_8173,N_7293);
nor U13969 (N_13969,N_7240,N_7335);
and U13970 (N_13970,N_5598,N_9826);
or U13971 (N_13971,N_7936,N_8874);
nand U13972 (N_13972,N_9616,N_7000);
nor U13973 (N_13973,N_5723,N_7172);
nor U13974 (N_13974,N_6246,N_5126);
nand U13975 (N_13975,N_5576,N_9047);
and U13976 (N_13976,N_6909,N_9817);
nand U13977 (N_13977,N_7435,N_6434);
nor U13978 (N_13978,N_6750,N_9630);
xor U13979 (N_13979,N_9283,N_7593);
xnor U13980 (N_13980,N_5315,N_9423);
or U13981 (N_13981,N_8706,N_9851);
and U13982 (N_13982,N_9003,N_9806);
nor U13983 (N_13983,N_9187,N_8350);
nand U13984 (N_13984,N_9144,N_9191);
nor U13985 (N_13985,N_9546,N_6110);
nand U13986 (N_13986,N_7804,N_8465);
nor U13987 (N_13987,N_7711,N_6995);
and U13988 (N_13988,N_6625,N_6163);
xnor U13989 (N_13989,N_7447,N_5684);
nand U13990 (N_13990,N_5386,N_7623);
and U13991 (N_13991,N_6593,N_5005);
and U13992 (N_13992,N_5702,N_6710);
xnor U13993 (N_13993,N_6074,N_8419);
nor U13994 (N_13994,N_7087,N_7620);
and U13995 (N_13995,N_9469,N_6076);
and U13996 (N_13996,N_8260,N_8244);
and U13997 (N_13997,N_8311,N_5281);
and U13998 (N_13998,N_7539,N_5062);
nand U13999 (N_13999,N_7454,N_7832);
or U14000 (N_14000,N_7380,N_9062);
nor U14001 (N_14001,N_7035,N_6028);
or U14002 (N_14002,N_9069,N_7357);
nor U14003 (N_14003,N_9520,N_9678);
and U14004 (N_14004,N_5694,N_8694);
xnor U14005 (N_14005,N_5067,N_7253);
nand U14006 (N_14006,N_5529,N_5975);
and U14007 (N_14007,N_6986,N_8554);
nor U14008 (N_14008,N_6368,N_8838);
or U14009 (N_14009,N_9750,N_9612);
and U14010 (N_14010,N_9306,N_7913);
nand U14011 (N_14011,N_7240,N_6557);
nand U14012 (N_14012,N_9563,N_6606);
xnor U14013 (N_14013,N_8491,N_8193);
and U14014 (N_14014,N_8563,N_5927);
nand U14015 (N_14015,N_9590,N_8004);
and U14016 (N_14016,N_5587,N_9513);
nand U14017 (N_14017,N_5673,N_6288);
or U14018 (N_14018,N_8373,N_8579);
or U14019 (N_14019,N_8977,N_6142);
xnor U14020 (N_14020,N_8051,N_9644);
and U14021 (N_14021,N_8347,N_8021);
xor U14022 (N_14022,N_8659,N_8825);
nor U14023 (N_14023,N_6167,N_7373);
xnor U14024 (N_14024,N_9392,N_9710);
nand U14025 (N_14025,N_5128,N_8970);
or U14026 (N_14026,N_8479,N_5543);
nand U14027 (N_14027,N_9788,N_7016);
or U14028 (N_14028,N_7598,N_9088);
xor U14029 (N_14029,N_9374,N_5994);
and U14030 (N_14030,N_8750,N_5632);
nand U14031 (N_14031,N_8253,N_7458);
xnor U14032 (N_14032,N_6225,N_6300);
nor U14033 (N_14033,N_5470,N_6548);
nand U14034 (N_14034,N_6744,N_9106);
nand U14035 (N_14035,N_7938,N_9770);
nor U14036 (N_14036,N_7702,N_6206);
or U14037 (N_14037,N_7834,N_9576);
nand U14038 (N_14038,N_6523,N_9267);
nand U14039 (N_14039,N_9724,N_5367);
and U14040 (N_14040,N_6647,N_7427);
and U14041 (N_14041,N_5744,N_5673);
nor U14042 (N_14042,N_9830,N_5677);
xor U14043 (N_14043,N_7884,N_5738);
nand U14044 (N_14044,N_5721,N_8115);
and U14045 (N_14045,N_5472,N_7586);
nand U14046 (N_14046,N_9576,N_6425);
nand U14047 (N_14047,N_8570,N_6135);
xor U14048 (N_14048,N_8546,N_8896);
and U14049 (N_14049,N_6976,N_9091);
nand U14050 (N_14050,N_5096,N_7430);
nand U14051 (N_14051,N_5623,N_8036);
nor U14052 (N_14052,N_9977,N_9128);
or U14053 (N_14053,N_8678,N_9481);
nand U14054 (N_14054,N_8049,N_7194);
nand U14055 (N_14055,N_7996,N_6212);
nor U14056 (N_14056,N_9179,N_6559);
nand U14057 (N_14057,N_6765,N_8336);
and U14058 (N_14058,N_7083,N_8458);
nand U14059 (N_14059,N_5496,N_6591);
xor U14060 (N_14060,N_8059,N_7465);
nand U14061 (N_14061,N_6200,N_6073);
nor U14062 (N_14062,N_8025,N_9250);
or U14063 (N_14063,N_9999,N_9910);
and U14064 (N_14064,N_6457,N_8306);
nand U14065 (N_14065,N_5116,N_8133);
nand U14066 (N_14066,N_7108,N_5104);
and U14067 (N_14067,N_7771,N_6772);
nand U14068 (N_14068,N_6903,N_8989);
or U14069 (N_14069,N_7175,N_8711);
nor U14070 (N_14070,N_7107,N_6645);
and U14071 (N_14071,N_7730,N_8339);
nand U14072 (N_14072,N_8466,N_6430);
and U14073 (N_14073,N_5708,N_6584);
or U14074 (N_14074,N_6218,N_9273);
nor U14075 (N_14075,N_6850,N_9269);
xnor U14076 (N_14076,N_6132,N_7492);
nand U14077 (N_14077,N_8765,N_7335);
or U14078 (N_14078,N_7215,N_8303);
or U14079 (N_14079,N_9455,N_9747);
nand U14080 (N_14080,N_8495,N_6362);
and U14081 (N_14081,N_8289,N_8187);
nor U14082 (N_14082,N_5907,N_6401);
xnor U14083 (N_14083,N_7505,N_5007);
and U14084 (N_14084,N_7875,N_7450);
nand U14085 (N_14085,N_8114,N_8452);
and U14086 (N_14086,N_6351,N_6085);
nor U14087 (N_14087,N_9621,N_5333);
nor U14088 (N_14088,N_7495,N_5124);
or U14089 (N_14089,N_7449,N_9839);
or U14090 (N_14090,N_7829,N_9136);
nor U14091 (N_14091,N_7252,N_5088);
or U14092 (N_14092,N_8166,N_8719);
nand U14093 (N_14093,N_9117,N_5068);
or U14094 (N_14094,N_6283,N_5912);
nand U14095 (N_14095,N_5901,N_5987);
nand U14096 (N_14096,N_8685,N_9158);
or U14097 (N_14097,N_6342,N_6582);
nand U14098 (N_14098,N_9413,N_6653);
and U14099 (N_14099,N_6085,N_7895);
or U14100 (N_14100,N_8530,N_7328);
nand U14101 (N_14101,N_6523,N_9196);
or U14102 (N_14102,N_6220,N_7934);
and U14103 (N_14103,N_9671,N_6368);
nand U14104 (N_14104,N_5692,N_9433);
and U14105 (N_14105,N_6400,N_7264);
nand U14106 (N_14106,N_6117,N_5318);
nor U14107 (N_14107,N_8735,N_6437);
nor U14108 (N_14108,N_7735,N_7723);
and U14109 (N_14109,N_6800,N_8414);
or U14110 (N_14110,N_6863,N_9915);
xor U14111 (N_14111,N_7645,N_5615);
and U14112 (N_14112,N_9482,N_7799);
or U14113 (N_14113,N_8851,N_9474);
nor U14114 (N_14114,N_7816,N_5781);
or U14115 (N_14115,N_5825,N_8973);
nand U14116 (N_14116,N_9243,N_6063);
or U14117 (N_14117,N_7645,N_5618);
and U14118 (N_14118,N_6817,N_7625);
nor U14119 (N_14119,N_7952,N_6784);
and U14120 (N_14120,N_8658,N_8094);
and U14121 (N_14121,N_9503,N_8405);
and U14122 (N_14122,N_6134,N_5426);
nor U14123 (N_14123,N_9952,N_6062);
or U14124 (N_14124,N_5264,N_6696);
nor U14125 (N_14125,N_5514,N_8154);
and U14126 (N_14126,N_9912,N_9507);
or U14127 (N_14127,N_9586,N_9198);
or U14128 (N_14128,N_6028,N_6714);
and U14129 (N_14129,N_5576,N_5716);
nand U14130 (N_14130,N_7937,N_9221);
nor U14131 (N_14131,N_6238,N_7728);
or U14132 (N_14132,N_6775,N_8249);
and U14133 (N_14133,N_7597,N_8421);
xor U14134 (N_14134,N_8747,N_6522);
nor U14135 (N_14135,N_8534,N_8237);
xor U14136 (N_14136,N_8269,N_5029);
xnor U14137 (N_14137,N_8390,N_6538);
and U14138 (N_14138,N_6837,N_7991);
or U14139 (N_14139,N_9376,N_6717);
nor U14140 (N_14140,N_9542,N_5420);
or U14141 (N_14141,N_6633,N_9458);
or U14142 (N_14142,N_7141,N_6401);
nor U14143 (N_14143,N_9378,N_5825);
or U14144 (N_14144,N_9554,N_7180);
and U14145 (N_14145,N_7093,N_7318);
and U14146 (N_14146,N_8230,N_8406);
nand U14147 (N_14147,N_5532,N_7355);
xnor U14148 (N_14148,N_7269,N_5059);
and U14149 (N_14149,N_5185,N_8443);
nor U14150 (N_14150,N_9384,N_7524);
or U14151 (N_14151,N_6152,N_6458);
nor U14152 (N_14152,N_9371,N_8789);
and U14153 (N_14153,N_9450,N_8752);
or U14154 (N_14154,N_7230,N_6944);
nand U14155 (N_14155,N_6056,N_7055);
and U14156 (N_14156,N_7383,N_9621);
xnor U14157 (N_14157,N_5032,N_6651);
or U14158 (N_14158,N_9562,N_8608);
nor U14159 (N_14159,N_9308,N_7329);
nor U14160 (N_14160,N_5862,N_9095);
nand U14161 (N_14161,N_5124,N_7869);
and U14162 (N_14162,N_8462,N_7149);
and U14163 (N_14163,N_8680,N_5279);
nor U14164 (N_14164,N_5678,N_9069);
xnor U14165 (N_14165,N_7159,N_9400);
nor U14166 (N_14166,N_7567,N_9835);
or U14167 (N_14167,N_8759,N_8903);
and U14168 (N_14168,N_8387,N_7933);
or U14169 (N_14169,N_7839,N_9785);
or U14170 (N_14170,N_5967,N_5893);
nand U14171 (N_14171,N_6055,N_9969);
nor U14172 (N_14172,N_6540,N_6708);
or U14173 (N_14173,N_9977,N_7576);
nand U14174 (N_14174,N_9767,N_8910);
or U14175 (N_14175,N_8306,N_5098);
and U14176 (N_14176,N_5228,N_7378);
or U14177 (N_14177,N_6672,N_9121);
nor U14178 (N_14178,N_8789,N_7108);
or U14179 (N_14179,N_5396,N_9309);
nand U14180 (N_14180,N_6651,N_5162);
and U14181 (N_14181,N_8954,N_9585);
or U14182 (N_14182,N_9353,N_6809);
nor U14183 (N_14183,N_9609,N_9117);
nand U14184 (N_14184,N_7925,N_9878);
nor U14185 (N_14185,N_5028,N_8948);
xor U14186 (N_14186,N_8593,N_8886);
xnor U14187 (N_14187,N_5095,N_6862);
nand U14188 (N_14188,N_7732,N_8261);
or U14189 (N_14189,N_9975,N_8499);
nor U14190 (N_14190,N_6859,N_7220);
and U14191 (N_14191,N_5421,N_9494);
or U14192 (N_14192,N_5207,N_9159);
nor U14193 (N_14193,N_9103,N_8781);
nand U14194 (N_14194,N_8195,N_5694);
nand U14195 (N_14195,N_7309,N_7130);
or U14196 (N_14196,N_8280,N_6926);
nor U14197 (N_14197,N_5940,N_5736);
nand U14198 (N_14198,N_9982,N_6893);
and U14199 (N_14199,N_8263,N_8343);
or U14200 (N_14200,N_7863,N_7210);
and U14201 (N_14201,N_8002,N_6364);
or U14202 (N_14202,N_6228,N_7673);
nand U14203 (N_14203,N_8835,N_7665);
or U14204 (N_14204,N_8934,N_5883);
and U14205 (N_14205,N_8877,N_9086);
and U14206 (N_14206,N_7833,N_5896);
nor U14207 (N_14207,N_9644,N_9151);
xnor U14208 (N_14208,N_7977,N_9498);
or U14209 (N_14209,N_7556,N_8177);
nor U14210 (N_14210,N_8886,N_9896);
nand U14211 (N_14211,N_6093,N_6969);
nor U14212 (N_14212,N_6386,N_8749);
and U14213 (N_14213,N_7194,N_7421);
nand U14214 (N_14214,N_5686,N_8496);
nor U14215 (N_14215,N_7503,N_7934);
xor U14216 (N_14216,N_7451,N_9547);
or U14217 (N_14217,N_8503,N_6955);
or U14218 (N_14218,N_6009,N_8478);
nor U14219 (N_14219,N_8177,N_8901);
xor U14220 (N_14220,N_9644,N_5102);
and U14221 (N_14221,N_6863,N_8310);
or U14222 (N_14222,N_6040,N_9878);
xor U14223 (N_14223,N_8342,N_8796);
and U14224 (N_14224,N_8691,N_7799);
or U14225 (N_14225,N_5221,N_9596);
or U14226 (N_14226,N_5116,N_9266);
and U14227 (N_14227,N_8422,N_6548);
xor U14228 (N_14228,N_7358,N_8454);
nor U14229 (N_14229,N_7011,N_7909);
or U14230 (N_14230,N_9993,N_5499);
or U14231 (N_14231,N_9563,N_6251);
or U14232 (N_14232,N_5714,N_7562);
xor U14233 (N_14233,N_5708,N_6051);
nand U14234 (N_14234,N_9333,N_8546);
or U14235 (N_14235,N_6901,N_8033);
and U14236 (N_14236,N_9572,N_9457);
or U14237 (N_14237,N_8102,N_7017);
and U14238 (N_14238,N_7377,N_9143);
and U14239 (N_14239,N_5319,N_5617);
nand U14240 (N_14240,N_5376,N_5469);
xor U14241 (N_14241,N_8887,N_7548);
and U14242 (N_14242,N_5200,N_6930);
and U14243 (N_14243,N_8047,N_5314);
xnor U14244 (N_14244,N_7688,N_9976);
or U14245 (N_14245,N_7767,N_9535);
xor U14246 (N_14246,N_9008,N_7863);
nor U14247 (N_14247,N_5481,N_6219);
or U14248 (N_14248,N_7424,N_7549);
nand U14249 (N_14249,N_9163,N_7300);
and U14250 (N_14250,N_7708,N_9494);
nand U14251 (N_14251,N_7090,N_6732);
nor U14252 (N_14252,N_6201,N_9619);
nor U14253 (N_14253,N_6871,N_9880);
or U14254 (N_14254,N_5502,N_9393);
and U14255 (N_14255,N_8164,N_8291);
nor U14256 (N_14256,N_6309,N_5894);
or U14257 (N_14257,N_9410,N_5958);
or U14258 (N_14258,N_9202,N_7029);
or U14259 (N_14259,N_6758,N_5648);
or U14260 (N_14260,N_5926,N_7230);
or U14261 (N_14261,N_8491,N_7581);
or U14262 (N_14262,N_8568,N_8432);
and U14263 (N_14263,N_5625,N_7037);
or U14264 (N_14264,N_5624,N_9920);
nor U14265 (N_14265,N_5855,N_6411);
nor U14266 (N_14266,N_5629,N_8111);
and U14267 (N_14267,N_9477,N_8579);
nor U14268 (N_14268,N_5078,N_5081);
and U14269 (N_14269,N_5109,N_5659);
nand U14270 (N_14270,N_6540,N_5820);
nand U14271 (N_14271,N_6949,N_7800);
nor U14272 (N_14272,N_8624,N_8735);
or U14273 (N_14273,N_8056,N_7717);
nor U14274 (N_14274,N_6386,N_5239);
nor U14275 (N_14275,N_7239,N_8651);
and U14276 (N_14276,N_7032,N_9900);
nand U14277 (N_14277,N_9951,N_6428);
nand U14278 (N_14278,N_5879,N_8943);
or U14279 (N_14279,N_9297,N_9056);
nand U14280 (N_14280,N_7335,N_6357);
nor U14281 (N_14281,N_7165,N_6766);
and U14282 (N_14282,N_6139,N_8511);
nor U14283 (N_14283,N_8049,N_9727);
or U14284 (N_14284,N_6655,N_6358);
or U14285 (N_14285,N_8022,N_5080);
and U14286 (N_14286,N_6163,N_6037);
or U14287 (N_14287,N_9029,N_7477);
nand U14288 (N_14288,N_6716,N_9116);
or U14289 (N_14289,N_8985,N_8589);
nor U14290 (N_14290,N_9630,N_6186);
or U14291 (N_14291,N_6611,N_9173);
and U14292 (N_14292,N_9263,N_5491);
and U14293 (N_14293,N_6483,N_7222);
xor U14294 (N_14294,N_9559,N_8138);
or U14295 (N_14295,N_7263,N_7530);
or U14296 (N_14296,N_5262,N_5167);
nor U14297 (N_14297,N_7507,N_8319);
and U14298 (N_14298,N_5665,N_6285);
or U14299 (N_14299,N_7605,N_8106);
and U14300 (N_14300,N_8113,N_6017);
or U14301 (N_14301,N_7043,N_9742);
xor U14302 (N_14302,N_9839,N_5106);
nand U14303 (N_14303,N_9732,N_7514);
nor U14304 (N_14304,N_6765,N_9901);
and U14305 (N_14305,N_5198,N_8242);
nand U14306 (N_14306,N_6400,N_9945);
or U14307 (N_14307,N_8960,N_5330);
nor U14308 (N_14308,N_9749,N_6763);
nor U14309 (N_14309,N_6064,N_7993);
nor U14310 (N_14310,N_6419,N_9851);
nor U14311 (N_14311,N_9526,N_5650);
nor U14312 (N_14312,N_7221,N_8230);
nor U14313 (N_14313,N_9557,N_7528);
nand U14314 (N_14314,N_6446,N_5542);
nor U14315 (N_14315,N_7790,N_8208);
nand U14316 (N_14316,N_5684,N_5343);
nand U14317 (N_14317,N_6238,N_8843);
nand U14318 (N_14318,N_5854,N_9879);
nand U14319 (N_14319,N_9197,N_7386);
or U14320 (N_14320,N_5632,N_7987);
or U14321 (N_14321,N_6090,N_8479);
nand U14322 (N_14322,N_5223,N_9186);
xnor U14323 (N_14323,N_5225,N_7680);
xnor U14324 (N_14324,N_8009,N_5819);
nor U14325 (N_14325,N_5905,N_8890);
or U14326 (N_14326,N_8061,N_5957);
or U14327 (N_14327,N_9630,N_7886);
nor U14328 (N_14328,N_9459,N_5782);
nor U14329 (N_14329,N_6379,N_8641);
nand U14330 (N_14330,N_9810,N_9868);
nand U14331 (N_14331,N_6275,N_9950);
nand U14332 (N_14332,N_6578,N_8444);
and U14333 (N_14333,N_7466,N_6041);
xor U14334 (N_14334,N_8322,N_7101);
and U14335 (N_14335,N_6836,N_5159);
or U14336 (N_14336,N_9333,N_9428);
nand U14337 (N_14337,N_9060,N_8285);
nor U14338 (N_14338,N_7708,N_6403);
and U14339 (N_14339,N_8444,N_7344);
nor U14340 (N_14340,N_9245,N_5885);
nand U14341 (N_14341,N_7510,N_9904);
and U14342 (N_14342,N_5938,N_5063);
xor U14343 (N_14343,N_9707,N_5133);
and U14344 (N_14344,N_8598,N_8167);
or U14345 (N_14345,N_8616,N_8146);
and U14346 (N_14346,N_5838,N_9581);
nor U14347 (N_14347,N_5749,N_8839);
xor U14348 (N_14348,N_7620,N_5167);
nand U14349 (N_14349,N_9561,N_5022);
or U14350 (N_14350,N_8083,N_9578);
nor U14351 (N_14351,N_8023,N_5386);
nand U14352 (N_14352,N_9908,N_8674);
nand U14353 (N_14353,N_8557,N_9723);
nand U14354 (N_14354,N_7987,N_7753);
or U14355 (N_14355,N_5904,N_8619);
or U14356 (N_14356,N_9665,N_5840);
or U14357 (N_14357,N_5852,N_7779);
and U14358 (N_14358,N_5638,N_7031);
or U14359 (N_14359,N_6689,N_8668);
and U14360 (N_14360,N_7030,N_7878);
nand U14361 (N_14361,N_7681,N_6833);
and U14362 (N_14362,N_8396,N_5667);
nand U14363 (N_14363,N_5790,N_6236);
nand U14364 (N_14364,N_7640,N_8624);
nor U14365 (N_14365,N_8476,N_6145);
and U14366 (N_14366,N_9648,N_8648);
nand U14367 (N_14367,N_5563,N_7295);
nand U14368 (N_14368,N_5625,N_6219);
or U14369 (N_14369,N_7421,N_5931);
nand U14370 (N_14370,N_6405,N_8127);
nand U14371 (N_14371,N_5761,N_7088);
and U14372 (N_14372,N_6300,N_6186);
and U14373 (N_14373,N_8848,N_7989);
xnor U14374 (N_14374,N_6610,N_7945);
and U14375 (N_14375,N_7033,N_7552);
nand U14376 (N_14376,N_7729,N_6805);
nor U14377 (N_14377,N_5422,N_6470);
xor U14378 (N_14378,N_7974,N_8401);
nand U14379 (N_14379,N_5436,N_6856);
nand U14380 (N_14380,N_7478,N_6554);
and U14381 (N_14381,N_8849,N_5569);
and U14382 (N_14382,N_7108,N_5853);
nand U14383 (N_14383,N_8052,N_9819);
or U14384 (N_14384,N_9157,N_9084);
or U14385 (N_14385,N_8195,N_7048);
nor U14386 (N_14386,N_7324,N_6698);
and U14387 (N_14387,N_5508,N_5256);
and U14388 (N_14388,N_6803,N_7425);
nor U14389 (N_14389,N_5577,N_8932);
nand U14390 (N_14390,N_6917,N_9444);
nand U14391 (N_14391,N_8216,N_5194);
or U14392 (N_14392,N_5423,N_9615);
nand U14393 (N_14393,N_9002,N_8263);
nand U14394 (N_14394,N_6611,N_9845);
and U14395 (N_14395,N_5354,N_9824);
or U14396 (N_14396,N_9268,N_5730);
and U14397 (N_14397,N_6490,N_7122);
nor U14398 (N_14398,N_7241,N_6536);
nor U14399 (N_14399,N_8521,N_7171);
nand U14400 (N_14400,N_9965,N_8544);
nor U14401 (N_14401,N_5429,N_9607);
or U14402 (N_14402,N_9625,N_8697);
xnor U14403 (N_14403,N_7973,N_8384);
nor U14404 (N_14404,N_8626,N_6668);
nand U14405 (N_14405,N_7879,N_7542);
nor U14406 (N_14406,N_9097,N_8002);
or U14407 (N_14407,N_7939,N_5012);
nor U14408 (N_14408,N_7491,N_9483);
nor U14409 (N_14409,N_9624,N_7300);
nand U14410 (N_14410,N_9482,N_8864);
nand U14411 (N_14411,N_5833,N_7869);
and U14412 (N_14412,N_8095,N_8104);
or U14413 (N_14413,N_9353,N_9555);
or U14414 (N_14414,N_8282,N_6771);
and U14415 (N_14415,N_9140,N_9258);
nor U14416 (N_14416,N_7418,N_7394);
and U14417 (N_14417,N_5258,N_5420);
xnor U14418 (N_14418,N_5290,N_8095);
xnor U14419 (N_14419,N_5955,N_7729);
nand U14420 (N_14420,N_6141,N_7189);
nand U14421 (N_14421,N_9971,N_7442);
nand U14422 (N_14422,N_9937,N_8535);
and U14423 (N_14423,N_7323,N_5282);
nand U14424 (N_14424,N_8655,N_9595);
nor U14425 (N_14425,N_8245,N_6262);
nand U14426 (N_14426,N_7206,N_7122);
or U14427 (N_14427,N_9020,N_5828);
or U14428 (N_14428,N_5890,N_5790);
xor U14429 (N_14429,N_6255,N_9997);
or U14430 (N_14430,N_5782,N_5744);
or U14431 (N_14431,N_5597,N_9355);
and U14432 (N_14432,N_9757,N_5618);
nor U14433 (N_14433,N_8794,N_5640);
and U14434 (N_14434,N_6905,N_6315);
nand U14435 (N_14435,N_6794,N_7330);
nand U14436 (N_14436,N_5631,N_6116);
nor U14437 (N_14437,N_5475,N_6775);
nor U14438 (N_14438,N_9265,N_9922);
and U14439 (N_14439,N_8132,N_9376);
or U14440 (N_14440,N_7384,N_6678);
nand U14441 (N_14441,N_8709,N_9769);
and U14442 (N_14442,N_5478,N_8855);
nand U14443 (N_14443,N_6203,N_5204);
nor U14444 (N_14444,N_8464,N_5137);
or U14445 (N_14445,N_5849,N_6810);
or U14446 (N_14446,N_5440,N_7130);
and U14447 (N_14447,N_5702,N_8759);
nand U14448 (N_14448,N_7249,N_5630);
or U14449 (N_14449,N_5603,N_6300);
nor U14450 (N_14450,N_5136,N_5152);
nor U14451 (N_14451,N_7305,N_9698);
nand U14452 (N_14452,N_8323,N_6433);
and U14453 (N_14453,N_8862,N_7636);
and U14454 (N_14454,N_8405,N_6290);
nand U14455 (N_14455,N_6505,N_8461);
or U14456 (N_14456,N_7170,N_7914);
xnor U14457 (N_14457,N_9559,N_7427);
or U14458 (N_14458,N_6085,N_5644);
or U14459 (N_14459,N_9136,N_6165);
or U14460 (N_14460,N_9759,N_8956);
nor U14461 (N_14461,N_6587,N_5409);
nand U14462 (N_14462,N_7501,N_5667);
or U14463 (N_14463,N_8061,N_7547);
or U14464 (N_14464,N_6172,N_7498);
nand U14465 (N_14465,N_9335,N_6997);
or U14466 (N_14466,N_6356,N_9770);
nand U14467 (N_14467,N_7918,N_5254);
or U14468 (N_14468,N_5063,N_6158);
nand U14469 (N_14469,N_6607,N_8896);
nor U14470 (N_14470,N_8464,N_8091);
and U14471 (N_14471,N_8797,N_8259);
nor U14472 (N_14472,N_7994,N_9951);
and U14473 (N_14473,N_6029,N_8927);
and U14474 (N_14474,N_5362,N_7847);
nor U14475 (N_14475,N_6204,N_6798);
nor U14476 (N_14476,N_9533,N_9527);
xnor U14477 (N_14477,N_8451,N_7853);
xnor U14478 (N_14478,N_8375,N_7917);
and U14479 (N_14479,N_9974,N_9930);
nor U14480 (N_14480,N_5314,N_8954);
and U14481 (N_14481,N_5751,N_8891);
xor U14482 (N_14482,N_8444,N_9775);
nor U14483 (N_14483,N_7106,N_5724);
nor U14484 (N_14484,N_7774,N_9449);
nor U14485 (N_14485,N_5655,N_5352);
xnor U14486 (N_14486,N_7188,N_7080);
nor U14487 (N_14487,N_9985,N_5205);
and U14488 (N_14488,N_8887,N_5898);
or U14489 (N_14489,N_9481,N_9693);
or U14490 (N_14490,N_8367,N_5216);
nand U14491 (N_14491,N_6344,N_5089);
nand U14492 (N_14492,N_8842,N_6007);
or U14493 (N_14493,N_8898,N_7823);
or U14494 (N_14494,N_7605,N_5425);
and U14495 (N_14495,N_9157,N_7947);
nand U14496 (N_14496,N_9581,N_9127);
nor U14497 (N_14497,N_6391,N_6510);
or U14498 (N_14498,N_7037,N_9881);
and U14499 (N_14499,N_5496,N_8656);
nor U14500 (N_14500,N_5221,N_9278);
nand U14501 (N_14501,N_8960,N_7721);
nor U14502 (N_14502,N_6632,N_7701);
nand U14503 (N_14503,N_5208,N_7951);
nand U14504 (N_14504,N_7954,N_7903);
nor U14505 (N_14505,N_5774,N_7840);
xor U14506 (N_14506,N_9241,N_7784);
or U14507 (N_14507,N_5110,N_7927);
nand U14508 (N_14508,N_7897,N_9454);
nor U14509 (N_14509,N_8423,N_6229);
and U14510 (N_14510,N_8969,N_8665);
and U14511 (N_14511,N_7217,N_9669);
xnor U14512 (N_14512,N_7208,N_7822);
nand U14513 (N_14513,N_8275,N_9173);
nand U14514 (N_14514,N_5484,N_7231);
or U14515 (N_14515,N_8876,N_6503);
and U14516 (N_14516,N_9788,N_7182);
nor U14517 (N_14517,N_8410,N_5683);
nand U14518 (N_14518,N_6883,N_8168);
or U14519 (N_14519,N_6686,N_7552);
xor U14520 (N_14520,N_9949,N_8744);
nand U14521 (N_14521,N_6280,N_9899);
xor U14522 (N_14522,N_6160,N_7952);
nor U14523 (N_14523,N_7073,N_5809);
and U14524 (N_14524,N_7451,N_6174);
nor U14525 (N_14525,N_7010,N_9560);
xnor U14526 (N_14526,N_9821,N_9406);
and U14527 (N_14527,N_8194,N_9105);
nand U14528 (N_14528,N_5298,N_9151);
and U14529 (N_14529,N_8865,N_8987);
nand U14530 (N_14530,N_7011,N_7638);
nor U14531 (N_14531,N_5137,N_6154);
or U14532 (N_14532,N_8417,N_6432);
and U14533 (N_14533,N_8200,N_8217);
or U14534 (N_14534,N_5437,N_6924);
nor U14535 (N_14535,N_9692,N_5756);
and U14536 (N_14536,N_5880,N_7851);
nor U14537 (N_14537,N_8473,N_9188);
or U14538 (N_14538,N_6713,N_7451);
nor U14539 (N_14539,N_7374,N_5014);
nand U14540 (N_14540,N_8857,N_9081);
nand U14541 (N_14541,N_7388,N_7161);
nor U14542 (N_14542,N_7716,N_9900);
and U14543 (N_14543,N_5413,N_8465);
xnor U14544 (N_14544,N_6035,N_6283);
nand U14545 (N_14545,N_9078,N_5756);
nand U14546 (N_14546,N_7780,N_7853);
nand U14547 (N_14547,N_5846,N_8546);
nor U14548 (N_14548,N_7792,N_7884);
or U14549 (N_14549,N_7665,N_8812);
or U14550 (N_14550,N_6363,N_6602);
or U14551 (N_14551,N_7843,N_5515);
and U14552 (N_14552,N_6949,N_5076);
nor U14553 (N_14553,N_5543,N_8744);
nor U14554 (N_14554,N_8456,N_7870);
or U14555 (N_14555,N_8839,N_5499);
or U14556 (N_14556,N_8156,N_9390);
and U14557 (N_14557,N_8384,N_5538);
xnor U14558 (N_14558,N_9994,N_9047);
or U14559 (N_14559,N_7630,N_7756);
and U14560 (N_14560,N_9502,N_9451);
nand U14561 (N_14561,N_7900,N_6875);
nor U14562 (N_14562,N_9877,N_7761);
nor U14563 (N_14563,N_5999,N_9301);
nor U14564 (N_14564,N_7327,N_6599);
and U14565 (N_14565,N_8437,N_6458);
and U14566 (N_14566,N_8297,N_6665);
nand U14567 (N_14567,N_7684,N_6926);
xor U14568 (N_14568,N_7987,N_9675);
and U14569 (N_14569,N_6502,N_8930);
and U14570 (N_14570,N_5868,N_9737);
nand U14571 (N_14571,N_9552,N_5590);
and U14572 (N_14572,N_8595,N_9248);
nand U14573 (N_14573,N_7485,N_7495);
nor U14574 (N_14574,N_8185,N_7633);
xor U14575 (N_14575,N_6442,N_8987);
or U14576 (N_14576,N_5956,N_6903);
nor U14577 (N_14577,N_7201,N_8617);
nand U14578 (N_14578,N_9408,N_5862);
nand U14579 (N_14579,N_8079,N_9267);
nand U14580 (N_14580,N_6748,N_5696);
xor U14581 (N_14581,N_6988,N_7466);
nand U14582 (N_14582,N_7169,N_8740);
nor U14583 (N_14583,N_6072,N_6628);
or U14584 (N_14584,N_5114,N_5862);
xnor U14585 (N_14585,N_7057,N_9973);
nor U14586 (N_14586,N_9876,N_6826);
nand U14587 (N_14587,N_9881,N_7103);
and U14588 (N_14588,N_5104,N_9992);
nor U14589 (N_14589,N_8427,N_5249);
and U14590 (N_14590,N_7661,N_9511);
nor U14591 (N_14591,N_9614,N_7482);
or U14592 (N_14592,N_8362,N_5190);
nand U14593 (N_14593,N_9551,N_5587);
nor U14594 (N_14594,N_9671,N_7244);
nor U14595 (N_14595,N_7689,N_7565);
nand U14596 (N_14596,N_7471,N_9676);
nand U14597 (N_14597,N_5184,N_6685);
xnor U14598 (N_14598,N_9243,N_5781);
and U14599 (N_14599,N_8677,N_9950);
and U14600 (N_14600,N_5641,N_5284);
nor U14601 (N_14601,N_7731,N_7010);
xor U14602 (N_14602,N_6217,N_5512);
nor U14603 (N_14603,N_9007,N_9682);
and U14604 (N_14604,N_5085,N_6705);
and U14605 (N_14605,N_5599,N_9992);
xor U14606 (N_14606,N_7007,N_6241);
nand U14607 (N_14607,N_6101,N_7723);
or U14608 (N_14608,N_9953,N_5608);
nand U14609 (N_14609,N_6443,N_5202);
xnor U14610 (N_14610,N_7199,N_7575);
nand U14611 (N_14611,N_8177,N_9870);
and U14612 (N_14612,N_8422,N_6415);
nor U14613 (N_14613,N_5123,N_6128);
or U14614 (N_14614,N_5105,N_5986);
or U14615 (N_14615,N_8186,N_8529);
nand U14616 (N_14616,N_8255,N_5094);
nand U14617 (N_14617,N_9476,N_6724);
and U14618 (N_14618,N_9260,N_6399);
xnor U14619 (N_14619,N_9495,N_5117);
nand U14620 (N_14620,N_9655,N_5460);
nor U14621 (N_14621,N_9461,N_6314);
and U14622 (N_14622,N_5673,N_8755);
and U14623 (N_14623,N_7124,N_8915);
xnor U14624 (N_14624,N_7424,N_7936);
and U14625 (N_14625,N_8351,N_5986);
xnor U14626 (N_14626,N_5997,N_5647);
and U14627 (N_14627,N_8819,N_6732);
and U14628 (N_14628,N_6441,N_7337);
or U14629 (N_14629,N_8547,N_8718);
and U14630 (N_14630,N_6627,N_5310);
nand U14631 (N_14631,N_7545,N_9642);
xor U14632 (N_14632,N_6281,N_6859);
or U14633 (N_14633,N_7083,N_6782);
and U14634 (N_14634,N_7216,N_9861);
nor U14635 (N_14635,N_6714,N_6419);
and U14636 (N_14636,N_7585,N_9126);
nor U14637 (N_14637,N_5873,N_9617);
xnor U14638 (N_14638,N_5007,N_5811);
xor U14639 (N_14639,N_8222,N_7706);
and U14640 (N_14640,N_6840,N_9352);
or U14641 (N_14641,N_8792,N_5553);
and U14642 (N_14642,N_9122,N_6185);
or U14643 (N_14643,N_7524,N_5465);
xnor U14644 (N_14644,N_9810,N_8585);
nand U14645 (N_14645,N_5778,N_6046);
nand U14646 (N_14646,N_6252,N_6166);
and U14647 (N_14647,N_8912,N_6176);
nand U14648 (N_14648,N_8310,N_7718);
nor U14649 (N_14649,N_7964,N_9232);
nor U14650 (N_14650,N_9689,N_6963);
nand U14651 (N_14651,N_7080,N_9815);
nand U14652 (N_14652,N_8949,N_6361);
or U14653 (N_14653,N_8116,N_5201);
or U14654 (N_14654,N_6753,N_6304);
nand U14655 (N_14655,N_9551,N_9229);
nand U14656 (N_14656,N_8286,N_5995);
nand U14657 (N_14657,N_8030,N_7806);
nand U14658 (N_14658,N_6924,N_7784);
or U14659 (N_14659,N_7349,N_9175);
nor U14660 (N_14660,N_5377,N_7737);
nor U14661 (N_14661,N_6214,N_7714);
nor U14662 (N_14662,N_9158,N_5039);
nor U14663 (N_14663,N_6502,N_9547);
xor U14664 (N_14664,N_6094,N_9039);
or U14665 (N_14665,N_7617,N_5277);
nand U14666 (N_14666,N_5661,N_7441);
and U14667 (N_14667,N_9465,N_7947);
nor U14668 (N_14668,N_5231,N_9406);
or U14669 (N_14669,N_6481,N_8122);
or U14670 (N_14670,N_5215,N_5983);
nand U14671 (N_14671,N_6335,N_9890);
nor U14672 (N_14672,N_9678,N_5257);
nand U14673 (N_14673,N_7019,N_8370);
nor U14674 (N_14674,N_8066,N_5309);
nand U14675 (N_14675,N_5532,N_8292);
nor U14676 (N_14676,N_7493,N_9060);
nand U14677 (N_14677,N_6908,N_5201);
or U14678 (N_14678,N_7386,N_8066);
or U14679 (N_14679,N_6786,N_5131);
or U14680 (N_14680,N_7642,N_6768);
nor U14681 (N_14681,N_9764,N_9015);
xnor U14682 (N_14682,N_7339,N_8752);
and U14683 (N_14683,N_9183,N_8181);
nor U14684 (N_14684,N_7645,N_7224);
nand U14685 (N_14685,N_8292,N_8744);
or U14686 (N_14686,N_8076,N_9461);
nor U14687 (N_14687,N_7464,N_5973);
nor U14688 (N_14688,N_8224,N_8092);
nand U14689 (N_14689,N_9769,N_7466);
xor U14690 (N_14690,N_6174,N_8011);
or U14691 (N_14691,N_5528,N_6796);
nand U14692 (N_14692,N_5554,N_9811);
nor U14693 (N_14693,N_7751,N_5831);
nor U14694 (N_14694,N_6913,N_9044);
and U14695 (N_14695,N_6095,N_8297);
nor U14696 (N_14696,N_6101,N_7755);
nand U14697 (N_14697,N_8298,N_8498);
nand U14698 (N_14698,N_5286,N_9965);
nand U14699 (N_14699,N_8763,N_8224);
or U14700 (N_14700,N_9496,N_8105);
or U14701 (N_14701,N_6549,N_8191);
xnor U14702 (N_14702,N_8987,N_6641);
nor U14703 (N_14703,N_7429,N_7528);
or U14704 (N_14704,N_5772,N_7259);
nand U14705 (N_14705,N_8854,N_9256);
and U14706 (N_14706,N_6956,N_6347);
or U14707 (N_14707,N_9711,N_6748);
nor U14708 (N_14708,N_7199,N_6079);
or U14709 (N_14709,N_7738,N_9781);
and U14710 (N_14710,N_7551,N_9979);
xnor U14711 (N_14711,N_5648,N_9516);
nor U14712 (N_14712,N_7859,N_6231);
nor U14713 (N_14713,N_9897,N_5762);
and U14714 (N_14714,N_9044,N_9709);
nand U14715 (N_14715,N_8516,N_6654);
and U14716 (N_14716,N_7170,N_5847);
and U14717 (N_14717,N_8483,N_5492);
or U14718 (N_14718,N_9675,N_8959);
nor U14719 (N_14719,N_8497,N_9218);
nand U14720 (N_14720,N_7470,N_8368);
nor U14721 (N_14721,N_6242,N_5693);
and U14722 (N_14722,N_5131,N_5219);
nor U14723 (N_14723,N_6409,N_8420);
and U14724 (N_14724,N_9908,N_7276);
and U14725 (N_14725,N_9494,N_7262);
or U14726 (N_14726,N_9445,N_8968);
and U14727 (N_14727,N_7495,N_6125);
and U14728 (N_14728,N_9530,N_9994);
and U14729 (N_14729,N_6939,N_6575);
xor U14730 (N_14730,N_9530,N_6808);
or U14731 (N_14731,N_9089,N_8631);
nand U14732 (N_14732,N_9060,N_6201);
or U14733 (N_14733,N_6620,N_9703);
or U14734 (N_14734,N_6249,N_9236);
nand U14735 (N_14735,N_5467,N_9917);
or U14736 (N_14736,N_6203,N_5809);
xnor U14737 (N_14737,N_5112,N_8958);
or U14738 (N_14738,N_9753,N_5774);
and U14739 (N_14739,N_8962,N_6135);
nand U14740 (N_14740,N_5157,N_6786);
nor U14741 (N_14741,N_9633,N_8780);
or U14742 (N_14742,N_9455,N_5446);
and U14743 (N_14743,N_8618,N_8482);
or U14744 (N_14744,N_6049,N_6252);
nor U14745 (N_14745,N_5213,N_6795);
and U14746 (N_14746,N_9045,N_6523);
nor U14747 (N_14747,N_8720,N_9554);
or U14748 (N_14748,N_5708,N_5493);
and U14749 (N_14749,N_5620,N_6962);
or U14750 (N_14750,N_7768,N_9127);
nor U14751 (N_14751,N_9017,N_8568);
and U14752 (N_14752,N_5944,N_9017);
and U14753 (N_14753,N_9467,N_9356);
and U14754 (N_14754,N_7570,N_5744);
and U14755 (N_14755,N_8437,N_7392);
nand U14756 (N_14756,N_7319,N_5535);
or U14757 (N_14757,N_8389,N_6352);
nand U14758 (N_14758,N_5545,N_7572);
or U14759 (N_14759,N_8999,N_9540);
and U14760 (N_14760,N_5530,N_6135);
nor U14761 (N_14761,N_9618,N_9904);
nand U14762 (N_14762,N_6146,N_7431);
xor U14763 (N_14763,N_5672,N_7573);
or U14764 (N_14764,N_6246,N_9102);
nor U14765 (N_14765,N_8198,N_5474);
or U14766 (N_14766,N_7049,N_6736);
xnor U14767 (N_14767,N_7128,N_9285);
nand U14768 (N_14768,N_7670,N_6357);
and U14769 (N_14769,N_6256,N_5843);
or U14770 (N_14770,N_9158,N_9292);
xnor U14771 (N_14771,N_9270,N_5300);
nand U14772 (N_14772,N_7130,N_9703);
and U14773 (N_14773,N_7500,N_8594);
xor U14774 (N_14774,N_5359,N_9504);
or U14775 (N_14775,N_8865,N_7732);
and U14776 (N_14776,N_7775,N_6604);
and U14777 (N_14777,N_5128,N_6433);
nor U14778 (N_14778,N_7462,N_6481);
and U14779 (N_14779,N_8723,N_9987);
or U14780 (N_14780,N_7954,N_5455);
and U14781 (N_14781,N_7002,N_9078);
and U14782 (N_14782,N_9167,N_8470);
nand U14783 (N_14783,N_8066,N_9589);
nor U14784 (N_14784,N_8434,N_9419);
nor U14785 (N_14785,N_9275,N_7192);
and U14786 (N_14786,N_6212,N_5703);
nand U14787 (N_14787,N_8396,N_7253);
nor U14788 (N_14788,N_5586,N_9611);
xnor U14789 (N_14789,N_8325,N_6137);
nand U14790 (N_14790,N_9563,N_8354);
xor U14791 (N_14791,N_9762,N_9511);
nand U14792 (N_14792,N_8254,N_8120);
or U14793 (N_14793,N_7521,N_7851);
and U14794 (N_14794,N_7285,N_8009);
and U14795 (N_14795,N_5316,N_8331);
nor U14796 (N_14796,N_5117,N_6845);
nor U14797 (N_14797,N_7470,N_7721);
or U14798 (N_14798,N_8369,N_7303);
nor U14799 (N_14799,N_8828,N_6499);
and U14800 (N_14800,N_9467,N_9669);
xnor U14801 (N_14801,N_5511,N_6011);
nor U14802 (N_14802,N_9059,N_8263);
or U14803 (N_14803,N_9959,N_9560);
or U14804 (N_14804,N_8265,N_5231);
nand U14805 (N_14805,N_8632,N_6366);
or U14806 (N_14806,N_5227,N_5840);
and U14807 (N_14807,N_9070,N_5771);
nor U14808 (N_14808,N_9957,N_7548);
and U14809 (N_14809,N_7733,N_5405);
or U14810 (N_14810,N_9987,N_7680);
nor U14811 (N_14811,N_6027,N_8841);
and U14812 (N_14812,N_8339,N_9370);
nor U14813 (N_14813,N_7363,N_6275);
or U14814 (N_14814,N_8693,N_6632);
or U14815 (N_14815,N_7121,N_8979);
and U14816 (N_14816,N_8819,N_6340);
or U14817 (N_14817,N_8975,N_7545);
nor U14818 (N_14818,N_8268,N_7993);
xor U14819 (N_14819,N_5261,N_5884);
nand U14820 (N_14820,N_7386,N_8070);
nor U14821 (N_14821,N_7820,N_7547);
nor U14822 (N_14822,N_7848,N_8883);
or U14823 (N_14823,N_7877,N_6755);
nor U14824 (N_14824,N_5241,N_5560);
or U14825 (N_14825,N_8838,N_6730);
and U14826 (N_14826,N_9980,N_9571);
nand U14827 (N_14827,N_5470,N_6730);
nand U14828 (N_14828,N_5629,N_5334);
nand U14829 (N_14829,N_9715,N_5587);
nor U14830 (N_14830,N_5804,N_6390);
and U14831 (N_14831,N_7094,N_9827);
nand U14832 (N_14832,N_7538,N_9500);
nand U14833 (N_14833,N_7689,N_7739);
or U14834 (N_14834,N_8668,N_9559);
nor U14835 (N_14835,N_5137,N_9667);
nor U14836 (N_14836,N_9142,N_9357);
nand U14837 (N_14837,N_6129,N_6336);
or U14838 (N_14838,N_5968,N_5719);
and U14839 (N_14839,N_8306,N_6452);
or U14840 (N_14840,N_6322,N_7668);
xnor U14841 (N_14841,N_5799,N_5897);
and U14842 (N_14842,N_7556,N_8699);
or U14843 (N_14843,N_8355,N_5686);
nand U14844 (N_14844,N_5381,N_5089);
xnor U14845 (N_14845,N_7378,N_8318);
and U14846 (N_14846,N_5694,N_8576);
nand U14847 (N_14847,N_7584,N_7313);
or U14848 (N_14848,N_9643,N_9414);
nand U14849 (N_14849,N_9493,N_5082);
or U14850 (N_14850,N_6908,N_6007);
or U14851 (N_14851,N_9019,N_7615);
nor U14852 (N_14852,N_9606,N_7723);
nand U14853 (N_14853,N_7961,N_6529);
or U14854 (N_14854,N_8672,N_7449);
xnor U14855 (N_14855,N_7281,N_5627);
nor U14856 (N_14856,N_6616,N_7589);
xor U14857 (N_14857,N_9476,N_9927);
xnor U14858 (N_14858,N_5255,N_8647);
nor U14859 (N_14859,N_9316,N_6685);
or U14860 (N_14860,N_5004,N_7287);
or U14861 (N_14861,N_7425,N_7535);
nand U14862 (N_14862,N_8915,N_6192);
and U14863 (N_14863,N_8623,N_8631);
or U14864 (N_14864,N_8659,N_9991);
and U14865 (N_14865,N_8894,N_5822);
or U14866 (N_14866,N_8949,N_7010);
or U14867 (N_14867,N_6912,N_6832);
nand U14868 (N_14868,N_6150,N_8669);
or U14869 (N_14869,N_5905,N_5153);
or U14870 (N_14870,N_9360,N_6141);
nor U14871 (N_14871,N_7379,N_9633);
or U14872 (N_14872,N_9349,N_7633);
nand U14873 (N_14873,N_8175,N_7846);
nor U14874 (N_14874,N_6509,N_6494);
and U14875 (N_14875,N_8246,N_8716);
nor U14876 (N_14876,N_9905,N_6059);
or U14877 (N_14877,N_6314,N_8647);
xnor U14878 (N_14878,N_8412,N_8542);
or U14879 (N_14879,N_7157,N_6612);
nand U14880 (N_14880,N_6549,N_7585);
and U14881 (N_14881,N_9938,N_6988);
or U14882 (N_14882,N_8251,N_5261);
nand U14883 (N_14883,N_5858,N_7594);
or U14884 (N_14884,N_7386,N_7047);
or U14885 (N_14885,N_6579,N_8426);
or U14886 (N_14886,N_7604,N_5894);
nand U14887 (N_14887,N_7953,N_9289);
xnor U14888 (N_14888,N_5703,N_5586);
xor U14889 (N_14889,N_8896,N_9010);
or U14890 (N_14890,N_9546,N_5681);
and U14891 (N_14891,N_5751,N_9929);
or U14892 (N_14892,N_6243,N_6545);
and U14893 (N_14893,N_5298,N_5641);
xnor U14894 (N_14894,N_8326,N_8512);
nor U14895 (N_14895,N_6807,N_7269);
nand U14896 (N_14896,N_6837,N_6971);
nor U14897 (N_14897,N_7779,N_5109);
nand U14898 (N_14898,N_6290,N_5727);
nor U14899 (N_14899,N_9056,N_8627);
and U14900 (N_14900,N_7322,N_6927);
nor U14901 (N_14901,N_6003,N_5966);
nand U14902 (N_14902,N_7823,N_5760);
nor U14903 (N_14903,N_7568,N_9815);
nand U14904 (N_14904,N_8253,N_6067);
nor U14905 (N_14905,N_8359,N_9208);
nand U14906 (N_14906,N_7522,N_5903);
xor U14907 (N_14907,N_8781,N_8118);
or U14908 (N_14908,N_9570,N_8901);
or U14909 (N_14909,N_7629,N_9795);
and U14910 (N_14910,N_5317,N_5581);
nand U14911 (N_14911,N_7774,N_9441);
or U14912 (N_14912,N_5767,N_6395);
xnor U14913 (N_14913,N_7231,N_7448);
or U14914 (N_14914,N_8730,N_6689);
nor U14915 (N_14915,N_8682,N_5604);
nand U14916 (N_14916,N_5273,N_7553);
or U14917 (N_14917,N_7151,N_8042);
or U14918 (N_14918,N_7274,N_8345);
xor U14919 (N_14919,N_6125,N_8282);
and U14920 (N_14920,N_8869,N_6953);
nor U14921 (N_14921,N_5214,N_9786);
and U14922 (N_14922,N_5319,N_9818);
xor U14923 (N_14923,N_9319,N_5191);
or U14924 (N_14924,N_7669,N_5519);
and U14925 (N_14925,N_7734,N_7182);
or U14926 (N_14926,N_8188,N_7012);
nand U14927 (N_14927,N_6299,N_9345);
and U14928 (N_14928,N_5287,N_9217);
nor U14929 (N_14929,N_6219,N_9598);
nand U14930 (N_14930,N_9008,N_6253);
or U14931 (N_14931,N_8884,N_6682);
nor U14932 (N_14932,N_8495,N_5488);
xnor U14933 (N_14933,N_5670,N_9912);
nand U14934 (N_14934,N_7438,N_8101);
and U14935 (N_14935,N_9608,N_7532);
nor U14936 (N_14936,N_7543,N_7576);
nor U14937 (N_14937,N_6047,N_6444);
and U14938 (N_14938,N_5477,N_5320);
and U14939 (N_14939,N_8254,N_6774);
nand U14940 (N_14940,N_7627,N_7962);
nand U14941 (N_14941,N_8304,N_6204);
xor U14942 (N_14942,N_7885,N_8295);
nor U14943 (N_14943,N_9864,N_6692);
nand U14944 (N_14944,N_9038,N_5075);
or U14945 (N_14945,N_5359,N_9177);
nand U14946 (N_14946,N_6576,N_7382);
or U14947 (N_14947,N_9436,N_9332);
nand U14948 (N_14948,N_5454,N_9319);
nand U14949 (N_14949,N_6776,N_5863);
xor U14950 (N_14950,N_6184,N_8723);
nor U14951 (N_14951,N_5054,N_9683);
or U14952 (N_14952,N_8590,N_6245);
and U14953 (N_14953,N_9792,N_5927);
and U14954 (N_14954,N_7772,N_6414);
or U14955 (N_14955,N_9266,N_7284);
nor U14956 (N_14956,N_7181,N_7329);
and U14957 (N_14957,N_9840,N_8156);
and U14958 (N_14958,N_6689,N_9891);
and U14959 (N_14959,N_8572,N_7287);
or U14960 (N_14960,N_9251,N_8277);
nor U14961 (N_14961,N_5586,N_9850);
xnor U14962 (N_14962,N_8756,N_9495);
or U14963 (N_14963,N_8287,N_9152);
nand U14964 (N_14964,N_7028,N_8141);
nor U14965 (N_14965,N_5110,N_8210);
or U14966 (N_14966,N_7436,N_7805);
nand U14967 (N_14967,N_6039,N_7618);
or U14968 (N_14968,N_8063,N_6962);
nor U14969 (N_14969,N_9507,N_8537);
nor U14970 (N_14970,N_6487,N_5722);
nand U14971 (N_14971,N_6465,N_7348);
or U14972 (N_14972,N_5204,N_6694);
or U14973 (N_14973,N_6919,N_6978);
nand U14974 (N_14974,N_6628,N_7880);
nand U14975 (N_14975,N_5225,N_8703);
nor U14976 (N_14976,N_9809,N_9811);
nand U14977 (N_14977,N_5405,N_8054);
nor U14978 (N_14978,N_6975,N_7466);
nand U14979 (N_14979,N_8016,N_9276);
nor U14980 (N_14980,N_8570,N_7999);
nor U14981 (N_14981,N_6477,N_8173);
nand U14982 (N_14982,N_9214,N_9250);
nand U14983 (N_14983,N_8555,N_7721);
nand U14984 (N_14984,N_5535,N_5473);
nand U14985 (N_14985,N_8516,N_6714);
nor U14986 (N_14986,N_9430,N_8155);
nand U14987 (N_14987,N_7614,N_9844);
nand U14988 (N_14988,N_5948,N_8090);
xor U14989 (N_14989,N_6606,N_5317);
nand U14990 (N_14990,N_5253,N_6949);
and U14991 (N_14991,N_9860,N_8351);
or U14992 (N_14992,N_9405,N_9236);
nor U14993 (N_14993,N_7125,N_8633);
xor U14994 (N_14994,N_5759,N_5024);
or U14995 (N_14995,N_6249,N_5816);
or U14996 (N_14996,N_9581,N_9070);
nand U14997 (N_14997,N_5248,N_7308);
and U14998 (N_14998,N_9404,N_6777);
and U14999 (N_14999,N_5058,N_6378);
nor U15000 (N_15000,N_14473,N_14561);
nand U15001 (N_15001,N_11648,N_11878);
or U15002 (N_15002,N_13035,N_13236);
and U15003 (N_15003,N_11346,N_10224);
nand U15004 (N_15004,N_14775,N_13162);
nand U15005 (N_15005,N_13893,N_14957);
or U15006 (N_15006,N_14964,N_12245);
nand U15007 (N_15007,N_12834,N_10936);
nand U15008 (N_15008,N_10497,N_10937);
nand U15009 (N_15009,N_12380,N_12450);
or U15010 (N_15010,N_10354,N_13498);
or U15011 (N_15011,N_10459,N_13001);
nor U15012 (N_15012,N_10480,N_14532);
or U15013 (N_15013,N_14710,N_12371);
nor U15014 (N_15014,N_11125,N_13937);
or U15015 (N_15015,N_11457,N_10609);
nand U15016 (N_15016,N_14848,N_11991);
xor U15017 (N_15017,N_13476,N_13770);
nand U15018 (N_15018,N_12694,N_14625);
and U15019 (N_15019,N_13972,N_11859);
and U15020 (N_15020,N_10218,N_14427);
and U15021 (N_15021,N_10665,N_13737);
or U15022 (N_15022,N_13612,N_11203);
nand U15023 (N_15023,N_13724,N_11679);
nor U15024 (N_15024,N_12099,N_10831);
nor U15025 (N_15025,N_11479,N_10106);
xnor U15026 (N_15026,N_11711,N_13928);
nor U15027 (N_15027,N_11004,N_10349);
and U15028 (N_15028,N_11860,N_14339);
or U15029 (N_15029,N_11423,N_11867);
nand U15030 (N_15030,N_13089,N_14713);
or U15031 (N_15031,N_14833,N_12370);
and U15032 (N_15032,N_12187,N_11396);
and U15033 (N_15033,N_12131,N_11613);
and U15034 (N_15034,N_10985,N_14590);
or U15035 (N_15035,N_11987,N_12574);
nand U15036 (N_15036,N_13884,N_13273);
xnor U15037 (N_15037,N_11221,N_10439);
nand U15038 (N_15038,N_10689,N_13073);
nor U15039 (N_15039,N_12066,N_14390);
and U15040 (N_15040,N_14988,N_13912);
or U15041 (N_15041,N_11535,N_10920);
or U15042 (N_15042,N_12218,N_14409);
xor U15043 (N_15043,N_13016,N_12394);
nor U15044 (N_15044,N_14628,N_13753);
nand U15045 (N_15045,N_11704,N_11851);
nand U15046 (N_15046,N_14684,N_14800);
and U15047 (N_15047,N_13627,N_13916);
nand U15048 (N_15048,N_12193,N_11803);
nand U15049 (N_15049,N_10592,N_10591);
nand U15050 (N_15050,N_10488,N_12182);
and U15051 (N_15051,N_13167,N_11124);
nand U15052 (N_15052,N_10393,N_10377);
or U15053 (N_15053,N_14661,N_10191);
or U15054 (N_15054,N_13925,N_10658);
nand U15055 (N_15055,N_12138,N_11498);
and U15056 (N_15056,N_13606,N_13015);
nand U15057 (N_15057,N_11507,N_12952);
nand U15058 (N_15058,N_13397,N_13227);
or U15059 (N_15059,N_10722,N_10257);
or U15060 (N_15060,N_14444,N_14969);
and U15061 (N_15061,N_12803,N_11841);
nor U15062 (N_15062,N_12223,N_12310);
nor U15063 (N_15063,N_12510,N_14051);
xnor U15064 (N_15064,N_12012,N_12351);
or U15065 (N_15065,N_10775,N_10928);
or U15066 (N_15066,N_11487,N_13908);
and U15067 (N_15067,N_12392,N_14048);
or U15068 (N_15068,N_12408,N_14574);
or U15069 (N_15069,N_14616,N_14973);
nor U15070 (N_15070,N_12515,N_11254);
xor U15071 (N_15071,N_14242,N_14451);
and U15072 (N_15072,N_10790,N_10039);
nor U15073 (N_15073,N_12585,N_11961);
nor U15074 (N_15074,N_12856,N_13889);
nor U15075 (N_15075,N_12070,N_13607);
nor U15076 (N_15076,N_14088,N_10863);
and U15077 (N_15077,N_10995,N_13269);
nor U15078 (N_15078,N_13096,N_13598);
and U15079 (N_15079,N_11119,N_14068);
or U15080 (N_15080,N_14058,N_11585);
or U15081 (N_15081,N_11531,N_10067);
nor U15082 (N_15082,N_13404,N_12091);
and U15083 (N_15083,N_14569,N_13883);
and U15084 (N_15084,N_11989,N_11559);
nand U15085 (N_15085,N_11111,N_11511);
xor U15086 (N_15086,N_10312,N_10091);
and U15087 (N_15087,N_13938,N_12242);
xor U15088 (N_15088,N_12640,N_11085);
or U15089 (N_15089,N_11975,N_10172);
and U15090 (N_15090,N_10291,N_11243);
nand U15091 (N_15091,N_13689,N_12887);
or U15092 (N_15092,N_12477,N_11730);
and U15093 (N_15093,N_10421,N_12651);
or U15094 (N_15094,N_12650,N_12054);
and U15095 (N_15095,N_14116,N_11709);
nand U15096 (N_15096,N_14660,N_11224);
xnor U15097 (N_15097,N_10960,N_14239);
or U15098 (N_15098,N_14344,N_13617);
nor U15099 (N_15099,N_11637,N_11425);
and U15100 (N_15100,N_11015,N_10918);
or U15101 (N_15101,N_12215,N_13481);
or U15102 (N_15102,N_14378,N_11642);
nand U15103 (N_15103,N_10938,N_14172);
or U15104 (N_15104,N_13773,N_10803);
or U15105 (N_15105,N_14460,N_11395);
or U15106 (N_15106,N_12334,N_13847);
nor U15107 (N_15107,N_13364,N_10254);
nand U15108 (N_15108,N_11029,N_10650);
nand U15109 (N_15109,N_11121,N_11104);
nand U15110 (N_15110,N_11355,N_10616);
nand U15111 (N_15111,N_10269,N_10746);
or U15112 (N_15112,N_13163,N_14562);
nor U15113 (N_15113,N_13699,N_14555);
nor U15114 (N_15114,N_13479,N_11021);
and U15115 (N_15115,N_12830,N_11343);
or U15116 (N_15116,N_12583,N_11393);
or U15117 (N_15117,N_13741,N_12202);
and U15118 (N_15118,N_13160,N_10756);
or U15119 (N_15119,N_14915,N_11264);
and U15120 (N_15120,N_13556,N_14137);
nand U15121 (N_15121,N_10783,N_11633);
nor U15122 (N_15122,N_14948,N_14982);
nor U15123 (N_15123,N_11672,N_13246);
or U15124 (N_15124,N_10453,N_11326);
xnor U15125 (N_15125,N_11097,N_10483);
nor U15126 (N_15126,N_12929,N_10390);
or U15127 (N_15127,N_11936,N_14691);
nand U15128 (N_15128,N_10123,N_10478);
and U15129 (N_15129,N_14272,N_12098);
and U15130 (N_15130,N_11918,N_11078);
and U15131 (N_15131,N_14154,N_14284);
nand U15132 (N_15132,N_14762,N_14405);
xor U15133 (N_15133,N_11509,N_11342);
nand U15134 (N_15134,N_13866,N_13906);
and U15135 (N_15135,N_10119,N_11474);
nor U15136 (N_15136,N_11536,N_13903);
or U15137 (N_15137,N_10024,N_13164);
or U15138 (N_15138,N_13472,N_10889);
nor U15139 (N_15139,N_10629,N_14345);
nand U15140 (N_15140,N_14872,N_13718);
or U15141 (N_15141,N_12199,N_10214);
or U15142 (N_15142,N_14765,N_12917);
xor U15143 (N_15143,N_13102,N_12417);
and U15144 (N_15144,N_12431,N_12002);
and U15145 (N_15145,N_14977,N_13584);
nor U15146 (N_15146,N_12522,N_12372);
and U15147 (N_15147,N_13858,N_11280);
and U15148 (N_15148,N_12220,N_12543);
nand U15149 (N_15149,N_10401,N_12879);
or U15150 (N_15150,N_10990,N_10595);
nand U15151 (N_15151,N_14208,N_10880);
or U15152 (N_15152,N_11900,N_11998);
nand U15153 (N_15153,N_12764,N_13203);
or U15154 (N_15154,N_11994,N_11389);
or U15155 (N_15155,N_14004,N_14580);
and U15156 (N_15156,N_12566,N_13595);
nand U15157 (N_15157,N_11093,N_11786);
xor U15158 (N_15158,N_10799,N_12126);
nand U15159 (N_15159,N_14269,N_11504);
or U15160 (N_15160,N_11107,N_13253);
nand U15161 (N_15161,N_14479,N_13958);
nor U15162 (N_15162,N_13511,N_10289);
and U15163 (N_15163,N_13275,N_14793);
nor U15164 (N_15164,N_12827,N_14712);
nor U15165 (N_15165,N_12071,N_10597);
nand U15166 (N_15166,N_14032,N_11359);
and U15167 (N_15167,N_11740,N_10249);
and U15168 (N_15168,N_10639,N_12303);
or U15169 (N_15169,N_13949,N_14146);
xor U15170 (N_15170,N_14448,N_10034);
and U15171 (N_15171,N_11824,N_12934);
or U15172 (N_15172,N_12143,N_14653);
or U15173 (N_15173,N_14624,N_11741);
and U15174 (N_15174,N_14276,N_13134);
xnor U15175 (N_15175,N_14851,N_10409);
or U15176 (N_15176,N_10149,N_14753);
nand U15177 (N_15177,N_10809,N_12254);
xnor U15178 (N_15178,N_10352,N_11083);
nand U15179 (N_15179,N_13545,N_14862);
xor U15180 (N_15180,N_14059,N_14501);
nand U15181 (N_15181,N_13447,N_13790);
nor U15182 (N_15182,N_14845,N_11174);
or U15183 (N_15183,N_12086,N_12068);
and U15184 (N_15184,N_12795,N_12038);
nor U15185 (N_15185,N_12471,N_13927);
and U15186 (N_15186,N_10202,N_13169);
or U15187 (N_15187,N_11007,N_11819);
and U15188 (N_15188,N_10178,N_11069);
xor U15189 (N_15189,N_14490,N_14241);
or U15190 (N_15190,N_14159,N_13292);
and U15191 (N_15191,N_10819,N_14464);
or U15192 (N_15192,N_14296,N_10963);
nand U15193 (N_15193,N_14924,N_11297);
or U15194 (N_15194,N_14268,N_11022);
nor U15195 (N_15195,N_13546,N_11896);
and U15196 (N_15196,N_13457,N_14402);
and U15197 (N_15197,N_14736,N_14437);
and U15198 (N_15198,N_12339,N_12556);
or U15199 (N_15199,N_14544,N_11148);
and U15200 (N_15200,N_13146,N_12229);
nand U15201 (N_15201,N_11318,N_11311);
and U15202 (N_15202,N_11818,N_14425);
xor U15203 (N_15203,N_10387,N_13775);
and U15204 (N_15204,N_13542,N_11590);
and U15205 (N_15205,N_13856,N_13824);
and U15206 (N_15206,N_14905,N_11300);
nor U15207 (N_15207,N_14138,N_13034);
nor U15208 (N_15208,N_11696,N_11041);
xor U15209 (N_15209,N_12781,N_10222);
nor U15210 (N_15210,N_11322,N_13522);
nor U15211 (N_15211,N_14792,N_13738);
nor U15212 (N_15212,N_12172,N_10988);
nand U15213 (N_15213,N_13781,N_14103);
nand U15214 (N_15214,N_10824,N_14538);
nand U15215 (N_15215,N_10890,N_14306);
nor U15216 (N_15216,N_11495,N_14618);
nor U15217 (N_15217,N_10089,N_13212);
nand U15218 (N_15218,N_12999,N_12540);
xnor U15219 (N_15219,N_14282,N_12949);
or U15220 (N_15220,N_13168,N_14166);
nor U15221 (N_15221,N_11059,N_10014);
nand U15222 (N_15222,N_12058,N_10964);
or U15223 (N_15223,N_12107,N_14070);
and U15224 (N_15224,N_13643,N_14334);
nor U15225 (N_15225,N_10281,N_12634);
nor U15226 (N_15226,N_13580,N_14553);
nand U15227 (N_15227,N_14916,N_10523);
xor U15228 (N_15228,N_10558,N_12652);
or U15229 (N_15229,N_14175,N_14831);
nor U15230 (N_15230,N_11833,N_11910);
or U15231 (N_15231,N_12684,N_14978);
xnor U15232 (N_15232,N_14387,N_10822);
nand U15233 (N_15233,N_14584,N_14453);
nor U15234 (N_15234,N_10734,N_12327);
and U15235 (N_15235,N_10036,N_13859);
nor U15236 (N_15236,N_13571,N_12366);
or U15237 (N_15237,N_10848,N_13049);
or U15238 (N_15238,N_12889,N_14413);
or U15239 (N_15239,N_12397,N_14097);
and U15240 (N_15240,N_10777,N_14098);
nor U15241 (N_15241,N_14745,N_11647);
xnor U15242 (N_15242,N_14568,N_10400);
or U15243 (N_15243,N_12293,N_11189);
nor U15244 (N_15244,N_14057,N_10787);
or U15245 (N_15245,N_10651,N_11766);
nor U15246 (N_15246,N_14811,N_13503);
and U15247 (N_15247,N_14535,N_11050);
and U15248 (N_15248,N_10926,N_14053);
xnor U15249 (N_15249,N_11809,N_10223);
and U15250 (N_15250,N_14498,N_11312);
nor U15251 (N_15251,N_14355,N_11657);
nor U15252 (N_15252,N_11887,N_11133);
nor U15253 (N_15253,N_13304,N_14906);
and U15254 (N_15254,N_13195,N_14335);
and U15255 (N_15255,N_13998,N_12864);
nor U15256 (N_15256,N_14860,N_13252);
nor U15257 (N_15257,N_11876,N_14152);
nand U15258 (N_15258,N_12641,N_14621);
or U15259 (N_15259,N_13974,N_11475);
nand U15260 (N_15260,N_12601,N_10950);
nor U15261 (N_15261,N_11829,N_13105);
nor U15262 (N_15262,N_12336,N_11020);
and U15263 (N_15263,N_12527,N_12564);
or U15264 (N_15264,N_11090,N_12860);
nor U15265 (N_15265,N_14417,N_10786);
or U15266 (N_15266,N_10753,N_14856);
xnor U15267 (N_15267,N_14258,N_13529);
nand U15268 (N_15268,N_14773,N_11413);
or U15269 (N_15269,N_14442,N_10837);
and U15270 (N_15270,N_14510,N_12854);
or U15271 (N_15271,N_10700,N_10672);
and U15272 (N_15272,N_13002,N_11634);
and U15273 (N_15273,N_12765,N_11886);
nor U15274 (N_15274,N_13356,N_10046);
and U15275 (N_15275,N_13576,N_13991);
nand U15276 (N_15276,N_11156,N_10571);
and U15277 (N_15277,N_10104,N_12315);
or U15278 (N_15278,N_10452,N_13551);
nand U15279 (N_15279,N_13415,N_11151);
or U15280 (N_15280,N_12643,N_14828);
nor U15281 (N_15281,N_14690,N_10945);
or U15282 (N_15282,N_11478,N_11820);
and U15283 (N_15283,N_14126,N_14746);
nand U15284 (N_15284,N_14377,N_10431);
and U15285 (N_15285,N_10503,N_10278);
and U15286 (N_15286,N_11565,N_13181);
nand U15287 (N_15287,N_12951,N_13459);
nor U15288 (N_15288,N_11489,N_14252);
nor U15289 (N_15289,N_14733,N_11341);
and U15290 (N_15290,N_10198,N_12969);
nor U15291 (N_15291,N_10195,N_10953);
and U15292 (N_15292,N_12981,N_10369);
nand U15293 (N_15293,N_14943,N_14468);
nor U15294 (N_15294,N_10060,N_14664);
or U15295 (N_15295,N_10263,N_12359);
or U15296 (N_15296,N_12939,N_11211);
and U15297 (N_15297,N_12841,N_10697);
nand U15298 (N_15298,N_10931,N_11967);
nor U15299 (N_15299,N_14730,N_11246);
nand U15300 (N_15300,N_10048,N_10433);
or U15301 (N_15301,N_13501,N_13987);
and U15302 (N_15302,N_11248,N_14100);
nor U15303 (N_15303,N_14229,N_14682);
nor U15304 (N_15304,N_11282,N_10517);
nor U15305 (N_15305,N_13967,N_10314);
nor U15306 (N_15306,N_13418,N_14187);
nor U15307 (N_15307,N_11979,N_13319);
xor U15308 (N_15308,N_10838,N_12845);
and U15309 (N_15309,N_10407,N_14844);
and U15310 (N_15310,N_11617,N_14949);
or U15311 (N_15311,N_14549,N_12148);
xnor U15312 (N_15312,N_12790,N_13044);
nor U15313 (N_15313,N_14686,N_11601);
or U15314 (N_15314,N_12383,N_12579);
nand U15315 (N_15315,N_12966,N_13180);
and U15316 (N_15316,N_11421,N_14260);
nor U15317 (N_15317,N_13301,N_13762);
or U15318 (N_15318,N_11473,N_13682);
nand U15319 (N_15319,N_12913,N_12858);
and U15320 (N_15320,N_14285,N_10136);
nand U15321 (N_15321,N_11168,N_12532);
or U15322 (N_15322,N_14917,N_10562);
nor U15323 (N_15323,N_13450,N_13358);
or U15324 (N_15324,N_12658,N_10417);
xor U15325 (N_15325,N_14692,N_13182);
nor U15326 (N_15326,N_11849,N_14842);
xnor U15327 (N_15327,N_11361,N_12051);
and U15328 (N_15328,N_14958,N_14997);
and U15329 (N_15329,N_13478,N_14696);
xnor U15330 (N_15330,N_13351,N_11921);
nor U15331 (N_15331,N_12046,N_14374);
and U15332 (N_15332,N_14771,N_10414);
nand U15333 (N_15333,N_13314,N_10551);
or U15334 (N_15334,N_11924,N_14222);
nor U15335 (N_15335,N_10978,N_12622);
and U15336 (N_15336,N_12816,N_10299);
and U15337 (N_15337,N_12575,N_12873);
and U15338 (N_15338,N_14799,N_12196);
nor U15339 (N_15339,N_11321,N_12709);
and U15340 (N_15340,N_14271,N_14830);
nor U15341 (N_15341,N_10802,N_10573);
and U15342 (N_15342,N_12171,N_11414);
nand U15343 (N_15343,N_13065,N_11606);
or U15344 (N_15344,N_10501,N_12089);
and U15345 (N_15345,N_10887,N_10647);
nand U15346 (N_15346,N_11232,N_12619);
nor U15347 (N_15347,N_13072,N_10923);
nand U15348 (N_15348,N_10396,N_14368);
and U15349 (N_15349,N_12629,N_13067);
nor U15350 (N_15350,N_13873,N_14962);
xnor U15351 (N_15351,N_10556,N_13367);
xnor U15352 (N_15352,N_10723,N_10232);
nor U15353 (N_15353,N_11079,N_12778);
nand U15354 (N_15354,N_10676,N_14247);
or U15355 (N_15355,N_10972,N_13448);
and U15356 (N_15356,N_10662,N_10916);
xnor U15357 (N_15357,N_10096,N_14434);
or U15358 (N_15358,N_10944,N_11238);
nor U15359 (N_15359,N_13821,N_13804);
or U15360 (N_15360,N_10427,N_12998);
nand U15361 (N_15361,N_12085,N_13649);
nand U15362 (N_15362,N_14256,N_10835);
nand U15363 (N_15363,N_10652,N_13727);
nand U15364 (N_15364,N_11893,N_10548);
nand U15365 (N_15365,N_10628,N_13539);
or U15366 (N_15366,N_11800,N_12094);
xor U15367 (N_15367,N_14323,N_11703);
or U15368 (N_15368,N_11656,N_14316);
and U15369 (N_15369,N_13726,N_12598);
nor U15370 (N_15370,N_12783,N_12480);
nor U15371 (N_15371,N_14201,N_11720);
xnor U15372 (N_15372,N_12298,N_13149);
nor U15373 (N_15373,N_12004,N_10490);
nand U15374 (N_15374,N_11619,N_14760);
xor U15375 (N_15375,N_13553,N_14465);
xnor U15376 (N_15376,N_12558,N_10436);
and U15377 (N_15377,N_11728,N_11775);
and U15378 (N_15378,N_12679,N_11623);
or U15379 (N_15379,N_14114,N_12479);
nor U15380 (N_15380,N_11659,N_12978);
or U15381 (N_15381,N_13083,N_11873);
or U15382 (N_15382,N_14497,N_13868);
and U15383 (N_15383,N_12063,N_10348);
or U15384 (N_15384,N_10566,N_13919);
nand U15385 (N_15385,N_14592,N_14700);
nor U15386 (N_15386,N_10482,N_14426);
and U15387 (N_15387,N_10408,N_11816);
nand U15388 (N_15388,N_12580,N_11171);
nand U15389 (N_15389,N_14517,N_14396);
nand U15390 (N_15390,N_12707,N_14761);
nor U15391 (N_15391,N_11747,N_11195);
xnor U15392 (N_15392,N_12531,N_14983);
and U15393 (N_15393,N_12914,N_14363);
nand U15394 (N_15394,N_14240,N_11739);
nor U15395 (N_15395,N_13780,N_11530);
nor U15396 (N_15396,N_10134,N_13975);
or U15397 (N_15397,N_10472,N_13765);
xnor U15398 (N_15398,N_11713,N_10213);
nor U15399 (N_15399,N_12693,N_10321);
xor U15400 (N_15400,N_14708,N_14614);
nor U15401 (N_15401,N_13876,N_12446);
or U15402 (N_15402,N_11862,N_13907);
or U15403 (N_15403,N_10773,N_13784);
and U15404 (N_15404,N_13909,N_10242);
nand U15405 (N_15405,N_12428,N_11272);
or U15406 (N_15406,N_14440,N_12581);
nand U15407 (N_15407,N_11985,N_13281);
nor U15408 (N_15408,N_13347,N_13887);
xnor U15409 (N_15409,N_13944,N_14836);
or U15410 (N_15410,N_12142,N_10004);
nand U15411 (N_15411,N_11988,N_13139);
and U15412 (N_15412,N_11661,N_13854);
or U15413 (N_15413,N_11751,N_12040);
nand U15414 (N_15414,N_10815,N_13899);
nor U15415 (N_15415,N_10617,N_12452);
xnor U15416 (N_15416,N_10817,N_12839);
nor U15417 (N_15417,N_11087,N_10107);
nand U15418 (N_15418,N_14195,N_13288);
nand U15419 (N_15419,N_11769,N_12101);
or U15420 (N_15420,N_11467,N_13039);
and U15421 (N_15421,N_12065,N_14896);
and U15422 (N_15422,N_12015,N_10788);
or U15423 (N_15423,N_13911,N_10821);
and U15424 (N_15424,N_12685,N_13045);
and U15425 (N_15425,N_11388,N_13350);
nor U15426 (N_15426,N_12608,N_13636);
xor U15427 (N_15427,N_12307,N_10906);
nor U15428 (N_15428,N_10250,N_11000);
xnor U15429 (N_15429,N_10533,N_13036);
or U15430 (N_15430,N_12319,N_12927);
nand U15431 (N_15431,N_14236,N_10580);
nand U15432 (N_15432,N_10295,N_13814);
or U15433 (N_15433,N_14122,N_11266);
nor U15434 (N_15434,N_13059,N_10555);
or U15435 (N_15435,N_14227,N_10686);
or U15436 (N_15436,N_13337,N_12796);
nor U15437 (N_15437,N_14864,N_14940);
nor U15438 (N_15438,N_11969,N_13735);
xor U15439 (N_15439,N_10507,N_11700);
or U15440 (N_15440,N_12486,N_10322);
or U15441 (N_15441,N_10684,N_10845);
nor U15442 (N_15442,N_11347,N_10765);
or U15443 (N_15443,N_14496,N_13694);
or U15444 (N_15444,N_13370,N_13956);
nand U15445 (N_15445,N_14613,N_10582);
and U15446 (N_15446,N_11150,N_12160);
nor U15447 (N_15447,N_11438,N_13708);
and U15448 (N_15448,N_13813,N_11812);
xnor U15449 (N_15449,N_12149,N_11813);
or U15450 (N_15450,N_14920,N_12430);
xor U15451 (N_15451,N_12669,N_10008);
nor U15452 (N_15452,N_14814,N_13009);
nor U15453 (N_15453,N_13455,N_10443);
or U15454 (N_15454,N_10781,N_12635);
or U15455 (N_15455,N_11673,N_11611);
or U15456 (N_15456,N_14859,N_14125);
xnor U15457 (N_15457,N_11576,N_12758);
or U15458 (N_15458,N_11398,N_14687);
or U15459 (N_15459,N_10428,N_12426);
or U15460 (N_15460,N_12509,N_12767);
nor U15461 (N_15461,N_10994,N_11428);
and U15462 (N_15462,N_10277,N_14475);
or U15463 (N_15463,N_13074,N_13965);
or U15464 (N_15464,N_11579,N_10664);
nor U15465 (N_15465,N_10830,N_11954);
nor U15466 (N_15466,N_11014,N_10381);
xnor U15467 (N_15467,N_10741,N_12258);
and U15468 (N_15468,N_10457,N_13834);
or U15469 (N_15469,N_11060,N_14231);
nor U15470 (N_15470,N_13714,N_14646);
nand U15471 (N_15471,N_11476,N_14416);
xor U15472 (N_15472,N_12291,N_12292);
and U15473 (N_15473,N_12717,N_14834);
nor U15474 (N_15474,N_12209,N_11554);
nand U15475 (N_15475,N_10818,N_13808);
nor U15476 (N_15476,N_14140,N_13559);
nand U15477 (N_15477,N_13177,N_13355);
nand U15478 (N_15478,N_14533,N_10557);
and U15479 (N_15479,N_13691,N_11970);
or U15480 (N_15480,N_14027,N_11830);
or U15481 (N_15481,N_14902,N_13698);
or U15482 (N_15482,N_10274,N_12485);
nand U15483 (N_15483,N_14560,N_13502);
nand U15484 (N_15484,N_12542,N_10353);
and U15485 (N_15485,N_14403,N_10740);
or U15486 (N_15486,N_11027,N_11333);
and U15487 (N_15487,N_14254,N_13122);
and U15488 (N_15488,N_12139,N_12920);
nand U15489 (N_15489,N_14343,N_10405);
nor U15490 (N_15490,N_10430,N_11144);
xor U15491 (N_15491,N_12059,N_12401);
or U15492 (N_15492,N_12869,N_10154);
nand U15493 (N_15493,N_10898,N_12469);
and U15494 (N_15494,N_12241,N_13508);
nor U15495 (N_15495,N_10640,N_11604);
nor U15496 (N_15496,N_14234,N_13100);
nand U15497 (N_15497,N_14457,N_12434);
nand U15498 (N_15498,N_10133,N_14850);
and U15499 (N_15499,N_12751,N_11332);
nor U15500 (N_15500,N_10709,N_14565);
or U15501 (N_15501,N_12769,N_13175);
nand U15502 (N_15502,N_10999,N_14155);
nor U15503 (N_15503,N_11768,N_12541);
xnor U15504 (N_15504,N_12926,N_11194);
nor U15505 (N_15505,N_11615,N_10760);
or U15506 (N_15506,N_13760,N_12244);
nor U15507 (N_15507,N_13148,N_11750);
nor U15508 (N_15508,N_11653,N_12667);
and U15509 (N_15509,N_14499,N_10248);
xnor U15510 (N_15510,N_13525,N_14768);
xnor U15511 (N_15511,N_10294,N_13131);
xor U15512 (N_15512,N_12356,N_12627);
nor U15513 (N_15513,N_10304,N_12174);
xor U15514 (N_15514,N_13756,N_12178);
and U15515 (N_15515,N_10878,N_13189);
nand U15516 (N_15516,N_14168,N_10090);
nor U15517 (N_15517,N_14295,N_14891);
or U15518 (N_15518,N_12724,N_14963);
or U15519 (N_15519,N_11483,N_14536);
nor U15520 (N_15520,N_14463,N_14291);
nand U15521 (N_15521,N_11826,N_12195);
and U15522 (N_15522,N_11912,N_11685);
or U15523 (N_15523,N_13043,N_12922);
and U15524 (N_15524,N_11652,N_13801);
or U15525 (N_15525,N_10454,N_12021);
and U15526 (N_15526,N_13565,N_10696);
or U15527 (N_15527,N_10323,N_13900);
nand U15528 (N_15528,N_14723,N_13621);
nor U15529 (N_15529,N_10121,N_14852);
nor U15530 (N_15530,N_12523,N_14832);
and U15531 (N_15531,N_10093,N_14633);
nor U15532 (N_15532,N_10515,N_13817);
or U15533 (N_15533,N_14790,N_13506);
and U15534 (N_15534,N_10521,N_11444);
nor U15535 (N_15535,N_13210,N_10441);
nand U15536 (N_15536,N_13379,N_10082);
nor U15537 (N_15537,N_14865,N_11367);
nor U15538 (N_15538,N_13357,N_11005);
nand U15539 (N_15539,N_13994,N_14216);
xor U15540 (N_15540,N_14423,N_11274);
and U15541 (N_15541,N_10940,N_12146);
nand U15542 (N_15542,N_13431,N_10206);
nor U15543 (N_15543,N_10416,N_13218);
and U15544 (N_15544,N_14035,N_13445);
nand U15545 (N_15545,N_12849,N_11785);
nor U15546 (N_15546,N_13130,N_12508);
or U15547 (N_15547,N_13297,N_14446);
xor U15548 (N_15548,N_13101,N_12982);
or U15549 (N_15549,N_12593,N_11360);
nand U15550 (N_15550,N_12487,N_11746);
nor U15551 (N_15551,N_14304,N_12276);
and U15552 (N_15552,N_12453,N_14975);
or U15553 (N_15553,N_11067,N_10240);
nand U15554 (N_15554,N_12726,N_11181);
or U15555 (N_15555,N_11888,N_11607);
xnor U15556 (N_15556,N_13620,N_12036);
or U15557 (N_15557,N_14545,N_14482);
nand U15558 (N_15558,N_14644,N_11911);
xor U15559 (N_15559,N_12774,N_10601);
or U15560 (N_15560,N_13376,N_12072);
nor U15561 (N_15561,N_12017,N_12528);
nor U15562 (N_15562,N_10162,N_10981);
or U15563 (N_15563,N_10952,N_11305);
nand U15564 (N_15564,N_12167,N_14557);
or U15565 (N_15565,N_12547,N_11870);
or U15566 (N_15566,N_12819,N_14670);
nand U15567 (N_15567,N_13754,N_14807);
or U15568 (N_15568,N_10019,N_10255);
nor U15569 (N_15569,N_12777,N_14677);
or U15570 (N_15570,N_10267,N_13192);
and U15571 (N_15571,N_13420,N_14581);
nor U15572 (N_15572,N_12637,N_14351);
or U15573 (N_15573,N_13660,N_12490);
nor U15574 (N_15574,N_11049,N_12409);
or U15575 (N_15575,N_12552,N_12899);
and U15576 (N_15576,N_14798,N_12782);
and U15577 (N_15577,N_11780,N_12088);
nor U15578 (N_15578,N_14158,N_10007);
nand U15579 (N_15579,N_14090,N_10770);
nor U15580 (N_15580,N_11907,N_12151);
and U15581 (N_15581,N_12559,N_11285);
or U15582 (N_15582,N_10315,N_13852);
nor U15583 (N_15583,N_13572,N_13451);
nor U15584 (N_15584,N_12944,N_11117);
nor U15585 (N_15585,N_13326,N_13678);
nor U15586 (N_15586,N_12711,N_12141);
nor U15587 (N_15587,N_12355,N_12248);
or U15588 (N_15588,N_10066,N_11167);
or U15589 (N_15589,N_10153,N_11089);
nor U15590 (N_15590,N_13853,N_10053);
nand U15591 (N_15591,N_14747,N_10867);
and U15592 (N_15592,N_10166,N_11184);
xnor U15593 (N_15593,N_11273,N_14766);
nand U15594 (N_15594,N_14612,N_14109);
or U15595 (N_15595,N_12586,N_11153);
and U15596 (N_15596,N_11006,N_13230);
or U15597 (N_15597,N_11584,N_12247);
nor U15598 (N_15598,N_14589,N_13964);
or U15599 (N_15599,N_11971,N_14266);
nand U15600 (N_15600,N_12030,N_12925);
nor U15601 (N_15601,N_12780,N_10143);
and U15602 (N_15602,N_12217,N_12263);
nor U15603 (N_15603,N_12984,N_12988);
nor U15604 (N_15604,N_10059,N_13792);
nor U15605 (N_15605,N_13797,N_13260);
and U15606 (N_15606,N_14481,N_14563);
nor U15607 (N_15607,N_11242,N_10701);
nand U15608 (N_15608,N_13352,N_12230);
nor U15609 (N_15609,N_10759,N_10702);
or U15610 (N_15610,N_11159,N_14056);
xnor U15611 (N_15611,N_10332,N_13135);
nor U15612 (N_15612,N_14876,N_12096);
and U15613 (N_15613,N_13681,N_13206);
xnor U15614 (N_15614,N_13618,N_10745);
or U15615 (N_15615,N_13709,N_12108);
and U15616 (N_15616,N_14907,N_13662);
or U15617 (N_15617,N_10212,N_12013);
xor U15618 (N_15618,N_12587,N_14748);
nor U15619 (N_15619,N_14701,N_14827);
nand U15620 (N_15620,N_13703,N_12124);
nand U15621 (N_15621,N_14754,N_12549);
nor U15622 (N_15622,N_10545,N_13342);
nor U15623 (N_15623,N_10270,N_14751);
and U15624 (N_15624,N_10128,N_12871);
nand U15625 (N_15625,N_12620,N_13561);
and U15626 (N_15626,N_10273,N_14996);
or U15627 (N_15627,N_13411,N_13022);
nand U15628 (N_15628,N_13778,N_13097);
nand U15629 (N_15629,N_14893,N_11122);
nand U15630 (N_15630,N_14724,N_12388);
nor U15631 (N_15631,N_13645,N_13133);
or U15632 (N_15632,N_14318,N_11736);
nor U15633 (N_15633,N_12538,N_11905);
nand U15634 (N_15634,N_14952,N_12970);
nor U15635 (N_15635,N_13632,N_14188);
nand U15636 (N_15636,N_10144,N_10194);
nand U15637 (N_15637,N_13611,N_13902);
nand U15638 (N_15638,N_12642,N_10968);
nand U15639 (N_15639,N_11324,N_10516);
nand U15640 (N_15640,N_13500,N_10912);
nor U15641 (N_15641,N_12743,N_13187);
or U15642 (N_15642,N_12533,N_12440);
and U15643 (N_15643,N_12023,N_11735);
and U15644 (N_15644,N_13848,N_14076);
nand U15645 (N_15645,N_10719,N_14685);
xor U15646 (N_15646,N_11126,N_10469);
or U15647 (N_15647,N_10301,N_12470);
and U15648 (N_15648,N_10670,N_11056);
nand U15649 (N_15649,N_13391,N_12491);
xor U15650 (N_15650,N_11278,N_12340);
nand U15651 (N_15651,N_14846,N_10750);
nor U15652 (N_15652,N_13138,N_10247);
or U15653 (N_15653,N_11368,N_11108);
or U15654 (N_15654,N_12266,N_14530);
and U15655 (N_15655,N_14688,N_13461);
or U15656 (N_15656,N_10886,N_12662);
nor U15657 (N_15657,N_10462,N_11962);
or U15658 (N_15658,N_12432,N_12915);
or U15659 (N_15659,N_13194,N_13228);
nand U15660 (N_15660,N_14812,N_12916);
xnor U15661 (N_15661,N_14855,N_14518);
nor U15662 (N_15662,N_12865,N_10204);
and U15663 (N_15663,N_12407,N_13136);
nand U15664 (N_15664,N_14777,N_12514);
nand U15665 (N_15665,N_11538,N_11625);
or U15666 (N_15666,N_13264,N_10833);
nand U15667 (N_15667,N_12398,N_12053);
nor U15668 (N_15668,N_10547,N_11110);
nand U15669 (N_15669,N_13557,N_11302);
nor U15670 (N_15670,N_14130,N_10241);
nand U15671 (N_15671,N_11697,N_11017);
nor U15672 (N_15672,N_12192,N_11922);
nand U15673 (N_15673,N_14414,N_11743);
or U15674 (N_15674,N_11338,N_10644);
and U15675 (N_15675,N_13533,N_10768);
xnor U15676 (N_15676,N_12333,N_10245);
nand U15677 (N_15677,N_11034,N_14976);
xor U15678 (N_15678,N_11291,N_12648);
or U15679 (N_15679,N_10069,N_11410);
nor U15680 (N_15680,N_12727,N_10575);
or U15681 (N_15681,N_12048,N_11100);
and U15682 (N_15682,N_11185,N_10411);
nand U15683 (N_15683,N_10905,N_10692);
nand U15684 (N_15684,N_12275,N_13635);
nor U15685 (N_15685,N_10581,N_13318);
nor U15686 (N_15686,N_10437,N_13021);
nor U15687 (N_15687,N_11680,N_11146);
or U15688 (N_15688,N_12368,N_12255);
nand U15689 (N_15689,N_14406,N_13262);
and U15690 (N_15690,N_10116,N_11649);
and U15691 (N_15691,N_13805,N_13591);
nand U15692 (N_15692,N_14105,N_13989);
or U15693 (N_15693,N_12181,N_10203);
and U15694 (N_15694,N_14181,N_11761);
nand U15695 (N_15695,N_14503,N_11503);
nor U15696 (N_15696,N_13282,N_13099);
or U15697 (N_15697,N_10861,N_12921);
and U15698 (N_15698,N_11676,N_13159);
or U15699 (N_15699,N_12381,N_10329);
nor U15700 (N_15700,N_11113,N_14650);
or U15701 (N_15701,N_10062,N_13063);
and U15702 (N_15702,N_10820,N_14466);
nor U15703 (N_15703,N_14881,N_10659);
or U15704 (N_15704,N_13720,N_14106);
nor U15705 (N_15705,N_11094,N_11433);
or U15706 (N_15706,N_13107,N_12569);
nand U15707 (N_15707,N_12930,N_13575);
xor U15708 (N_15708,N_13343,N_14895);
nand U15709 (N_15709,N_10225,N_13910);
and U15710 (N_15710,N_14418,N_13622);
nor U15711 (N_15711,N_10005,N_11702);
nor U15712 (N_15712,N_11596,N_12001);
nor U15713 (N_15713,N_13939,N_11430);
and U15714 (N_15714,N_11043,N_12859);
or U15715 (N_15715,N_12797,N_13658);
or U15716 (N_15716,N_10577,N_10654);
nand U15717 (N_15717,N_13396,N_11491);
or U15718 (N_15718,N_14186,N_12467);
and U15719 (N_15719,N_14635,N_12349);
or U15720 (N_15720,N_13142,N_11293);
and U15721 (N_15721,N_13843,N_10574);
nand U15722 (N_15722,N_14302,N_13215);
xnor U15723 (N_15723,N_14139,N_11790);
or U15724 (N_15724,N_14731,N_14037);
nor U15725 (N_15725,N_12779,N_12557);
nor U15726 (N_15726,N_10292,N_13441);
or U15727 (N_15727,N_11627,N_11035);
nand U15728 (N_15728,N_10869,N_11283);
nor U15729 (N_15729,N_14348,N_12855);
nor U15730 (N_15730,N_12596,N_14566);
or U15731 (N_15731,N_13878,N_10406);
or U15732 (N_15732,N_14489,N_10092);
xor U15733 (N_15733,N_10442,N_13941);
and U15734 (N_15734,N_14632,N_14824);
xnor U15735 (N_15735,N_13986,N_14627);
nand U15736 (N_15736,N_12260,N_11624);
nor U15737 (N_15737,N_12867,N_12135);
and U15738 (N_15738,N_13038,N_10418);
nor U15739 (N_15739,N_13454,N_12844);
nor U15740 (N_15740,N_12618,N_12868);
nand U15741 (N_15741,N_10588,N_12611);
nand U15742 (N_15742,N_13325,N_11805);
nand U15743 (N_15743,N_10174,N_14816);
or U15744 (N_15744,N_11881,N_13332);
xor U15745 (N_15745,N_13983,N_10509);
and U15746 (N_15746,N_14120,N_13128);
or U15747 (N_15747,N_14511,N_13597);
and U15748 (N_15748,N_13000,N_11539);
nand U15749 (N_15749,N_12129,N_14235);
or U15750 (N_15750,N_13121,N_14995);
nand U15751 (N_15751,N_12813,N_14069);
or U15752 (N_15752,N_12968,N_14022);
or U15753 (N_15753,N_11582,N_10856);
or U15754 (N_15754,N_13763,N_11493);
nor U15755 (N_15755,N_10021,N_13010);
or U15756 (N_15756,N_13600,N_12236);
and U15757 (N_15757,N_12332,N_14806);
nor U15758 (N_15758,N_11468,N_12657);
or U15759 (N_15759,N_12425,N_13151);
nor U15760 (N_15760,N_14698,N_12517);
or U15761 (N_15761,N_11265,N_11136);
nor U15762 (N_15762,N_11386,N_10615);
and U15763 (N_15763,N_12696,N_14034);
or U15764 (N_15764,N_10572,N_10852);
or U15765 (N_15765,N_11852,N_13064);
or U15766 (N_15766,N_11522,N_11047);
and U15767 (N_15767,N_11417,N_11434);
or U15768 (N_15768,N_11024,N_14955);
or U15769 (N_15769,N_10440,N_12102);
nand U15770 (N_15770,N_13085,N_10506);
or U15771 (N_15771,N_12318,N_11884);
xor U15772 (N_15772,N_12708,N_14430);
or U15773 (N_15773,N_13922,N_12603);
nand U15774 (N_15774,N_12518,N_13145);
nand U15775 (N_15775,N_14010,N_13715);
nor U15776 (N_15776,N_11256,N_13232);
or U15777 (N_15777,N_14605,N_11892);
xor U15778 (N_15778,N_12621,N_12663);
nand U15779 (N_15779,N_14767,N_13186);
and U15780 (N_15780,N_13031,N_10237);
and U15781 (N_15781,N_11044,N_13581);
nor U15782 (N_15782,N_10170,N_11456);
or U15783 (N_15783,N_10882,N_14994);
nor U15784 (N_15784,N_10010,N_11875);
or U15785 (N_15785,N_14221,N_12103);
or U15786 (N_15786,N_13521,N_14220);
xor U15787 (N_15787,N_12449,N_11667);
nand U15788 (N_15788,N_12200,N_13693);
or U15789 (N_15789,N_12512,N_11038);
nor U15790 (N_15790,N_13103,N_13920);
nor U15791 (N_15791,N_10584,N_13725);
and U15792 (N_15792,N_13412,N_11400);
nor U15793 (N_15793,N_10398,N_12308);
or U15794 (N_15794,N_14123,N_11866);
nor U15795 (N_15795,N_13165,N_13857);
and U15796 (N_15796,N_14358,N_10355);
xnor U15797 (N_15797,N_14791,N_14892);
and U15798 (N_15798,N_12787,N_13458);
nand U15799 (N_15799,N_13125,N_10780);
nand U15800 (N_15800,N_14238,N_13340);
and U15801 (N_15801,N_12385,N_13748);
xor U15802 (N_15802,N_10043,N_12847);
and U15803 (N_15803,N_12870,N_14450);
or U15804 (N_15804,N_11187,N_12137);
nand U15805 (N_15805,N_11102,N_14823);
and U15806 (N_15806,N_10447,N_13183);
and U15807 (N_15807,N_13048,N_14937);
nand U15808 (N_15808,N_12008,N_13582);
or U15809 (N_15809,N_12752,N_10504);
nor U15810 (N_15810,N_13882,N_12670);
nand U15811 (N_15811,N_11407,N_14206);
nor U15812 (N_15812,N_11934,N_12261);
nand U15813 (N_15813,N_14121,N_13905);
nand U15814 (N_15814,N_12285,N_12660);
and U15815 (N_15815,N_11532,N_13213);
nor U15816 (N_15816,N_12773,N_12599);
nand U15817 (N_15817,N_11929,N_12617);
nor U15818 (N_15818,N_13872,N_10751);
or U15819 (N_15819,N_14429,N_10251);
and U15820 (N_15820,N_13605,N_12173);
and U15821 (N_15821,N_10632,N_11252);
or U15822 (N_15822,N_14929,N_11313);
and U15823 (N_15823,N_12721,N_10736);
nor U15824 (N_15824,N_14672,N_11628);
nor U15825 (N_15825,N_14398,N_13783);
nor U15826 (N_15826,N_10302,N_12447);
or U15827 (N_15827,N_11635,N_10610);
xor U15828 (N_15828,N_10265,N_13639);
nand U15829 (N_15829,N_11555,N_12763);
nor U15830 (N_15830,N_10841,N_11654);
or U15831 (N_15831,N_10720,N_11115);
or U15832 (N_15832,N_11502,N_10140);
and U15833 (N_15833,N_14129,N_10167);
nand U15834 (N_15834,N_13274,N_14092);
nor U15835 (N_15835,N_11180,N_13901);
and U15836 (N_15836,N_11040,N_11621);
xnor U15837 (N_15837,N_10681,N_11556);
nor U15838 (N_15838,N_12936,N_10563);
nor U15839 (N_15839,N_11973,N_10487);
or U15840 (N_15840,N_10177,N_13219);
and U15841 (N_15841,N_12731,N_10682);
and U15842 (N_15842,N_14491,N_13025);
nand U15843 (N_15843,N_14023,N_14619);
nand U15844 (N_15844,N_12155,N_12924);
and U15845 (N_15845,N_10456,N_10145);
xor U15846 (N_15846,N_11880,N_11542);
nand U15847 (N_15847,N_11758,N_11540);
nand U15848 (N_15848,N_12127,N_11401);
and U15849 (N_15849,N_13436,N_10816);
nand U15850 (N_15850,N_12850,N_14087);
and U15851 (N_15851,N_14781,N_11898);
nand U15852 (N_15852,N_10598,N_11753);
or U15853 (N_15853,N_14312,N_10413);
and U15854 (N_15854,N_12365,N_11854);
and U15855 (N_15855,N_14528,N_12950);
nand U15856 (N_15856,N_11525,N_12358);
and U15857 (N_15857,N_11890,N_13731);
nand U15858 (N_15858,N_11404,N_12279);
and U15859 (N_15859,N_13403,N_13517);
nor U15860 (N_15860,N_14292,N_13665);
and U15861 (N_15861,N_14091,N_14327);
and U15862 (N_15862,N_12852,N_10135);
nand U15863 (N_15863,N_13943,N_11533);
xnor U15864 (N_15864,N_11052,N_10993);
nor U15865 (N_15865,N_14061,N_12043);
and U15866 (N_15866,N_10137,N_12405);
nor U15867 (N_15867,N_13463,N_13241);
nand U15868 (N_15868,N_11142,N_12186);
nand U15869 (N_15869,N_14575,N_12818);
nand U15870 (N_15870,N_12184,N_13120);
and U15871 (N_15871,N_12794,N_12537);
or U15872 (N_15872,N_14849,N_10989);
nand U15873 (N_15873,N_14847,N_14540);
nand U15874 (N_15874,N_12006,N_10002);
nand U15875 (N_15875,N_13839,N_11213);
and U15876 (N_15876,N_11843,N_11670);
and U15877 (N_15877,N_12227,N_10947);
or U15878 (N_15878,N_12749,N_11128);
or U15879 (N_15879,N_14819,N_13093);
nor U15880 (N_15880,N_11217,N_10675);
or U15881 (N_15881,N_10371,N_14868);
xor U15882 (N_15882,N_14990,N_11289);
xor U15883 (N_15883,N_12993,N_14835);
nand U15884 (N_15884,N_14054,N_13810);
nor U15885 (N_15885,N_13936,N_13524);
nand U15886 (N_15886,N_11446,N_12702);
nor U15887 (N_15887,N_10283,N_10744);
or U15888 (N_15888,N_10395,N_12373);
xnor U15889 (N_15889,N_14298,N_10375);
or U15890 (N_15890,N_14267,N_11692);
or U15891 (N_15891,N_11992,N_10018);
nor U15892 (N_15892,N_14273,N_12503);
nand U15893 (N_15893,N_11950,N_12115);
or U15894 (N_15894,N_10896,N_10666);
and U15895 (N_15895,N_14301,N_13242);
nand U15896 (N_15896,N_12418,N_11942);
and U15897 (N_15897,N_10331,N_12840);
nand U15898 (N_15898,N_13117,N_11996);
nand U15899 (N_15899,N_10738,N_10849);
nand U15900 (N_15900,N_12744,N_14822);
nor U15901 (N_15901,N_11080,N_11724);
and U15902 (N_15902,N_12766,N_14289);
nor U15903 (N_15903,N_12314,N_10489);
or U15904 (N_15904,N_14210,N_13327);
or U15905 (N_15905,N_14841,N_11399);
and U15906 (N_15906,N_14991,N_10813);
and U15907 (N_15907,N_12214,N_13400);
nor U15908 (N_15908,N_11470,N_10226);
xnor U15909 (N_15909,N_10392,N_11465);
xnor U15910 (N_15910,N_13568,N_11737);
and U15911 (N_15911,N_11963,N_14945);
and U15912 (N_15912,N_12616,N_13362);
nand U15913 (N_15913,N_14861,N_13394);
and U15914 (N_15914,N_10704,N_10097);
and U15915 (N_15915,N_10677,N_10310);
or U15916 (N_15916,N_10948,N_11143);
or U15917 (N_15917,N_14340,N_13329);
or U15918 (N_15918,N_11380,N_11299);
nor U15919 (N_15919,N_13578,N_11390);
nand U15920 (N_15920,N_14428,N_12825);
or U15921 (N_15921,N_14780,N_13076);
nand U15922 (N_15922,N_13812,N_12990);
or U15923 (N_15923,N_10866,N_11682);
nor U15924 (N_15924,N_10868,N_13050);
or U15925 (N_15925,N_11101,N_11206);
nand U15926 (N_15926,N_11548,N_13336);
nor U15927 (N_15927,N_10725,N_14484);
nor U15928 (N_15928,N_11891,N_11009);
and U15929 (N_15929,N_14265,N_12891);
or U15930 (N_15930,N_14537,N_11091);
nand U15931 (N_15931,N_14815,N_10190);
and U15932 (N_15932,N_10410,N_11323);
or U15933 (N_15933,N_13896,N_13029);
and U15934 (N_15934,N_12460,N_14840);
xnor U15935 (N_15935,N_14215,N_12029);
nand U15936 (N_15936,N_10827,N_11325);
nor U15937 (N_15937,N_11541,N_12695);
nor U15938 (N_15938,N_11258,N_14593);
nor U15939 (N_15939,N_11365,N_11908);
or U15940 (N_15940,N_14472,N_11214);
or U15941 (N_15941,N_10716,N_14826);
xor U15942 (N_15942,N_13971,N_11534);
and U15943 (N_15943,N_11344,N_14000);
nor U15944 (N_15944,N_13798,N_10244);
and U15945 (N_15945,N_10187,N_12835);
nor U15946 (N_15946,N_12806,N_14099);
nor U15947 (N_15947,N_13483,N_12277);
or U15948 (N_15948,N_12312,N_12747);
and U15949 (N_15949,N_14877,N_10337);
xnor U15950 (N_15950,N_11953,N_12252);
and U15951 (N_15951,N_14055,N_12690);
or U15952 (N_15952,N_10631,N_10297);
and U15953 (N_15953,N_11406,N_14884);
nor U15954 (N_15954,N_13642,N_11403);
nand U15955 (N_15955,N_12228,N_13012);
and U15956 (N_15956,N_11230,N_13863);
nor U15957 (N_15957,N_13528,N_10621);
and U15958 (N_15958,N_14030,N_13293);
nor U15959 (N_15959,N_13886,N_13446);
nor U15960 (N_15960,N_14548,N_12578);
or U15961 (N_15961,N_14725,N_14506);
nor U15962 (N_15962,N_13933,N_11543);
and U15963 (N_15963,N_14029,N_14987);
nand U15964 (N_15964,N_11130,N_11372);
nor U15965 (N_15965,N_13184,N_13062);
nand U15966 (N_15966,N_12226,N_13384);
or U15967 (N_15967,N_13716,N_13239);
or U15968 (N_15968,N_11183,N_11269);
or U15969 (N_15969,N_11053,N_11757);
and U15970 (N_15970,N_13650,N_10823);
xor U15971 (N_15971,N_10510,N_14384);
nor U15972 (N_15972,N_10636,N_13794);
nand U15973 (N_15973,N_14454,N_13205);
nand U15974 (N_15974,N_10648,N_10959);
and U15975 (N_15975,N_12203,N_14364);
nor U15976 (N_15976,N_13712,N_14369);
and U15977 (N_15977,N_12492,N_12386);
and U15978 (N_15978,N_13221,N_12000);
or U15979 (N_15979,N_12957,N_10227);
or U15980 (N_15980,N_11927,N_12977);
nand U15981 (N_15981,N_14050,N_13697);
nor U15982 (N_15982,N_11591,N_10596);
or U15983 (N_15983,N_13722,N_12093);
xnor U15984 (N_15984,N_10669,N_11701);
nand U15985 (N_15985,N_12893,N_11861);
nor U15986 (N_15986,N_10217,N_13652);
or U15987 (N_15987,N_12798,N_14461);
and U15988 (N_15988,N_11058,N_12083);
or U15989 (N_15989,N_10854,N_11949);
nor U15990 (N_15990,N_13657,N_11557);
or U15991 (N_15991,N_12659,N_14346);
nor U15992 (N_15992,N_14763,N_10769);
nand U15993 (N_15993,N_11384,N_13027);
or U15994 (N_15994,N_12412,N_12473);
or U15995 (N_15995,N_11842,N_14117);
and U15996 (N_15996,N_13894,N_13387);
or U15997 (N_15997,N_13862,N_14066);
or U15998 (N_15998,N_10015,N_14714);
or U15999 (N_15999,N_13676,N_11139);
or U16000 (N_16000,N_14576,N_11527);
and U16001 (N_16001,N_11909,N_10455);
xnor U16002 (N_16002,N_14253,N_10607);
nand U16003 (N_16003,N_12791,N_12438);
or U16004 (N_16004,N_12876,N_11135);
or U16005 (N_16005,N_13985,N_13330);
nor U16006 (N_16006,N_11846,N_14667);
nor U16007 (N_16007,N_13978,N_13942);
and U16008 (N_16008,N_10844,N_13263);
nor U16009 (N_16009,N_10911,N_10946);
nand U16010 (N_16010,N_12716,N_12996);
nor U16011 (N_16011,N_13249,N_10793);
or U16012 (N_16012,N_10151,N_11772);
nand U16013 (N_16013,N_14542,N_11340);
nor U16014 (N_16014,N_12423,N_13833);
or U16015 (N_16015,N_13018,N_13088);
nor U16016 (N_16016,N_10451,N_11378);
and U16017 (N_16017,N_10749,N_10518);
and U16018 (N_16018,N_13444,N_12706);
nor U16019 (N_16019,N_13348,N_13881);
or U16020 (N_16020,N_14707,N_11481);
xnor U16021 (N_16021,N_14397,N_13926);
nand U16022 (N_16022,N_14717,N_13023);
nand U16023 (N_16023,N_11199,N_12555);
or U16024 (N_16024,N_10138,N_10054);
and U16025 (N_16025,N_12390,N_11817);
and U16026 (N_16026,N_10642,N_14083);
or U16027 (N_16027,N_11436,N_14421);
xor U16028 (N_16028,N_10674,N_11202);
nor U16029 (N_16029,N_13816,N_11166);
xor U16030 (N_16030,N_10434,N_14729);
nor U16031 (N_16031,N_10003,N_10929);
and U16032 (N_16032,N_10368,N_14697);
nand U16033 (N_16033,N_14458,N_13871);
nor U16034 (N_16034,N_11245,N_14774);
xor U16035 (N_16035,N_12673,N_10376);
or U16036 (N_16036,N_11705,N_12760);
nand U16037 (N_16037,N_10977,N_10874);
and U16038 (N_16038,N_12728,N_12396);
or U16039 (N_16039,N_14934,N_13729);
and U16040 (N_16040,N_10967,N_14173);
or U16041 (N_16041,N_11141,N_13217);
nand U16042 (N_16042,N_14399,N_10626);
and U16043 (N_16043,N_14889,N_10895);
nand U16044 (N_16044,N_14758,N_12983);
and U16045 (N_16045,N_13771,N_10864);
and U16046 (N_16046,N_14319,N_12570);
nand U16047 (N_16047,N_12842,N_13574);
nand U16048 (N_16048,N_11286,N_12521);
nand U16049 (N_16049,N_11749,N_14594);
and U16050 (N_16050,N_10256,N_14922);
or U16051 (N_16051,N_10179,N_14809);
and U16052 (N_16052,N_14492,N_11952);
xor U16053 (N_16053,N_11959,N_12588);
and U16054 (N_16054,N_11965,N_14786);
or U16055 (N_16055,N_13058,N_13838);
xnor U16056 (N_16056,N_10220,N_13374);
and U16057 (N_16057,N_11831,N_12125);
xor U16058 (N_16058,N_10544,N_14110);
and U16059 (N_16059,N_13789,N_13924);
and U16060 (N_16060,N_13037,N_11082);
and U16061 (N_16061,N_11799,N_14392);
or U16062 (N_16062,N_10448,N_14541);
nor U16063 (N_16063,N_13491,N_12128);
nor U16064 (N_16064,N_13091,N_13291);
or U16065 (N_16065,N_12748,N_10234);
and U16066 (N_16066,N_11447,N_13480);
and U16067 (N_16067,N_10280,N_11574);
and U16068 (N_16068,N_10789,N_13294);
nand U16069 (N_16069,N_13124,N_10385);
or U16070 (N_16070,N_10806,N_10496);
nor U16071 (N_16071,N_14744,N_12745);
xnor U16072 (N_16072,N_13226,N_11415);
nor U16073 (N_16073,N_14246,N_14615);
nand U16074 (N_16074,N_13671,N_13518);
nand U16075 (N_16075,N_10884,N_11003);
and U16076 (N_16076,N_11485,N_14160);
nand U16077 (N_16077,N_11220,N_10111);
and U16078 (N_16078,N_11620,N_13057);
and U16079 (N_16079,N_13406,N_13423);
nor U16080 (N_16080,N_12116,N_14966);
or U16081 (N_16081,N_12573,N_12087);
or U16082 (N_16082,N_14551,N_13669);
nand U16083 (N_16083,N_10735,N_13141);
nand U16084 (N_16084,N_11666,N_10991);
nor U16085 (N_16085,N_13054,N_11899);
nor U16086 (N_16086,N_11550,N_12507);
or U16087 (N_16087,N_10894,N_10942);
nor U16088 (N_16088,N_14796,N_12057);
nor U16089 (N_16089,N_14757,N_12338);
xor U16090 (N_16090,N_11699,N_11715);
or U16091 (N_16091,N_14443,N_14556);
or U16092 (N_16092,N_12804,N_14134);
xnor U16093 (N_16093,N_10871,N_14586);
or U16094 (N_16094,N_11508,N_10085);
nand U16095 (N_16095,N_14903,N_12233);
and U16096 (N_16096,N_13870,N_12212);
or U16097 (N_16097,N_11872,N_13945);
and U16098 (N_16098,N_13467,N_12833);
nand U16099 (N_16099,N_14951,N_14078);
nor U16100 (N_16100,N_13537,N_10892);
or U16101 (N_16101,N_11716,N_14180);
nor U16102 (N_16102,N_14329,N_14193);
and U16103 (N_16103,N_13979,N_12019);
or U16104 (N_16104,N_11320,N_13877);
nand U16105 (N_16105,N_11863,N_10877);
nor U16106 (N_16106,N_12264,N_12897);
or U16107 (N_16107,N_12361,N_12746);
xnor U16108 (N_16108,N_13328,N_10951);
and U16109 (N_16109,N_12799,N_11366);
nor U16110 (N_16110,N_12378,N_10484);
and U16111 (N_16111,N_12565,N_10721);
or U16112 (N_16112,N_10156,N_13526);
and U16113 (N_16113,N_13822,N_11284);
and U16114 (N_16114,N_13654,N_14342);
nor U16115 (N_16115,N_11773,N_10543);
or U16116 (N_16116,N_10146,N_10101);
nand U16117 (N_16117,N_14894,N_10049);
or U16118 (N_16118,N_10083,N_11466);
xor U16119 (N_16119,N_12630,N_14162);
nor U16120 (N_16120,N_10035,N_13875);
xor U16121 (N_16121,N_13823,N_13492);
nand U16122 (N_16122,N_12232,N_12052);
and U16123 (N_16123,N_14115,N_12723);
nand U16124 (N_16124,N_12654,N_12462);
nor U16125 (N_16125,N_10712,N_12197);
nor U16126 (N_16126,N_11048,N_14354);
and U16127 (N_16127,N_10714,N_10604);
nand U16128 (N_16128,N_12632,N_10657);
nand U16129 (N_16129,N_13413,N_12069);
nand U16130 (N_16130,N_11581,N_12545);
nor U16131 (N_16131,N_11426,N_14887);
nor U16132 (N_16132,N_10290,N_10673);
nand U16133 (N_16133,N_13477,N_12831);
and U16134 (N_16134,N_12156,N_13590);
xnor U16135 (N_16135,N_11229,N_13898);
xor U16136 (N_16136,N_14634,N_13512);
nand U16137 (N_16137,N_13723,N_10071);
nor U16138 (N_16138,N_14918,N_11336);
nand U16139 (N_16139,N_10973,N_13443);
or U16140 (N_16140,N_12363,N_14972);
and U16141 (N_16141,N_12826,N_10383);
or U16142 (N_16142,N_12326,N_14651);
or U16143 (N_16143,N_10074,N_10678);
nor U16144 (N_16144,N_14743,N_12710);
nand U16145 (N_16145,N_12287,N_11416);
or U16146 (N_16146,N_14347,N_12493);
nand U16147 (N_16147,N_13265,N_13730);
and U16148 (N_16148,N_12584,N_10924);
or U16149 (N_16149,N_14064,N_14866);
nand U16150 (N_16150,N_11545,N_13111);
or U16151 (N_16151,N_13849,N_14243);
and U16152 (N_16152,N_11754,N_13030);
and U16153 (N_16153,N_10955,N_14147);
xor U16154 (N_16154,N_11065,N_11132);
nor U16155 (N_16155,N_11351,N_11553);
or U16156 (N_16156,N_10238,N_10727);
xor U16157 (N_16157,N_14526,N_13686);
nand U16158 (N_16158,N_12862,N_14196);
xor U16159 (N_16159,N_14500,N_12645);
or U16160 (N_16160,N_11490,N_14337);
and U16161 (N_16161,N_13828,N_14182);
nand U16162 (N_16162,N_14470,N_10679);
nand U16163 (N_16163,N_10061,N_14512);
nand U16164 (N_16164,N_11155,N_12896);
nand U16165 (N_16165,N_14950,N_14145);
nor U16166 (N_16166,N_13519,N_11147);
xnor U16167 (N_16167,N_14879,N_14944);
nor U16168 (N_16168,N_14602,N_11571);
nand U16169 (N_16169,N_10468,N_10330);
and U16170 (N_16170,N_13353,N_11810);
xnor U16171 (N_16171,N_12025,N_13835);
nand U16172 (N_16172,N_13800,N_10196);
or U16173 (N_16173,N_10603,N_14954);
or U16174 (N_16174,N_13630,N_13383);
or U16175 (N_16175,N_12185,N_12007);
nor U16176 (N_16176,N_10360,N_10933);
nand U16177 (N_16177,N_13462,N_12457);
nor U16178 (N_16178,N_10380,N_13250);
nand U16179 (N_16179,N_13201,N_11823);
and U16180 (N_16180,N_10761,N_12832);
nand U16181 (N_16181,N_13255,N_10549);
nand U16182 (N_16182,N_13471,N_13047);
or U16183 (N_16183,N_14853,N_10498);
and U16184 (N_16184,N_12625,N_14164);
nand U16185 (N_16185,N_13317,N_14366);
nand U16186 (N_16186,N_12810,N_10029);
and U16187 (N_16187,N_13324,N_11231);
or U16188 (N_16188,N_11660,N_12987);
or U16189 (N_16189,N_10209,N_11678);
nor U16190 (N_16190,N_14654,N_13497);
or U16191 (N_16191,N_14169,N_11412);
and U16192 (N_16192,N_11387,N_10637);
nand U16193 (N_16193,N_11062,N_11477);
and U16194 (N_16194,N_10914,N_11317);
and U16195 (N_16195,N_10219,N_14689);
nor U16196 (N_16196,N_14939,N_14564);
xnor U16197 (N_16197,N_13710,N_11742);
and U16198 (N_16198,N_10359,N_14156);
xnor U16199 (N_16199,N_13626,N_13119);
nor U16200 (N_16200,N_11877,N_13934);
nand U16201 (N_16201,N_12931,N_14674);
xor U16202 (N_16202,N_12940,N_12973);
nor U16203 (N_16203,N_11092,N_13155);
nand U16204 (N_16204,N_12606,N_10285);
and U16205 (N_16205,N_14520,N_12656);
nor U16206 (N_16206,N_14082,N_12009);
xor U16207 (N_16207,N_12631,N_10103);
nor U16208 (N_16208,N_13410,N_10528);
and U16209 (N_16209,N_12189,N_10041);
nand U16210 (N_16210,N_11602,N_12304);
or U16211 (N_16211,N_10127,N_14559);
nand U16212 (N_16212,N_10646,N_14232);
or U16213 (N_16213,N_14938,N_14360);
and U16214 (N_16214,N_10272,N_12316);
nand U16215 (N_16215,N_11529,N_13433);
nor U16216 (N_16216,N_12504,N_12050);
and U16217 (N_16217,N_12400,N_11725);
nor U16218 (N_16218,N_13046,N_12649);
nand U16219 (N_16219,N_14449,N_13127);
and U16220 (N_16220,N_13191,N_11776);
nand U16221 (N_16221,N_11638,N_14142);
and U16222 (N_16222,N_12055,N_11759);
nand U16223 (N_16223,N_13256,N_13108);
xor U16224 (N_16224,N_13302,N_12097);
xor U16225 (N_16225,N_11718,N_11207);
or U16226 (N_16226,N_13019,N_10389);
and U16227 (N_16227,N_14656,N_13851);
nor U16228 (N_16228,N_12890,N_13706);
nand U16229 (N_16229,N_11774,N_12162);
and U16230 (N_16230,N_10108,N_10531);
nor U16231 (N_16231,N_12811,N_12207);
and U16232 (N_16232,N_12222,N_13229);
and U16233 (N_16233,N_13690,N_14300);
nor U16234 (N_16234,N_11131,N_13081);
and U16235 (N_16235,N_13592,N_14133);
xor U16236 (N_16236,N_12971,N_13266);
nor U16237 (N_16237,N_12208,N_12877);
nand U16238 (N_16238,N_11904,N_13960);
and U16239 (N_16239,N_11304,N_11631);
nand U16240 (N_16240,N_12597,N_12678);
xor U16241 (N_16241,N_12330,N_14308);
and U16242 (N_16242,N_13401,N_13452);
nor U16243 (N_16243,N_13644,N_10423);
nand U16244 (N_16244,N_10513,N_11589);
xnor U16245 (N_16245,N_14325,N_12109);
nor U16246 (N_16246,N_11145,N_13389);
nor U16247 (N_16247,N_11182,N_14299);
and U16248 (N_16248,N_13335,N_13567);
xor U16249 (N_16249,N_13114,N_11453);
and U16250 (N_16250,N_14522,N_14509);
nor U16251 (N_16251,N_14046,N_12965);
nor U16252 (N_16252,N_14531,N_10086);
nor U16253 (N_16253,N_12754,N_14550);
or U16254 (N_16254,N_10313,N_10339);
and U16255 (N_16255,N_14328,N_10065);
xor U16256 (N_16256,N_14165,N_10717);
nand U16257 (N_16257,N_14184,N_11832);
and U16258 (N_16258,N_11018,N_13113);
or U16259 (N_16259,N_10192,N_10229);
nand U16260 (N_16260,N_13947,N_13071);
and U16261 (N_16261,N_14028,N_12904);
and U16262 (N_16262,N_10435,N_10534);
xor U16263 (N_16263,N_14788,N_13806);
or U16264 (N_16264,N_10667,N_11316);
and U16265 (N_16265,N_14356,N_13077);
nand U16266 (N_16266,N_12535,N_12455);
nor U16267 (N_16267,N_11240,N_10718);
nand U16268 (N_16268,N_14759,N_10559);
nor U16269 (N_16269,N_12551,N_14107);
nor U16270 (N_16270,N_13825,N_14259);
nor U16271 (N_16271,N_14467,N_12676);
nand U16272 (N_16272,N_10426,N_12892);
nand U16273 (N_16273,N_12403,N_14926);
and U16274 (N_16274,N_14407,N_10899);
nand U16275 (N_16275,N_14679,N_14021);
and U16276 (N_16276,N_12820,N_10356);
nor U16277 (N_16277,N_13981,N_10197);
xor U16278 (N_16278,N_13564,N_13717);
nor U16279 (N_16279,N_12439,N_13493);
nand U16280 (N_16280,N_12342,N_11191);
nor U16281 (N_16281,N_12299,N_14740);
nand U16282 (N_16282,N_12190,N_12980);
xor U16283 (N_16283,N_13196,N_12100);
xor U16284 (N_16284,N_14669,N_11636);
nor U16285 (N_16285,N_10463,N_12610);
and U16286 (N_16286,N_12823,N_12848);
or U16287 (N_16287,N_14810,N_14089);
or U16288 (N_16288,N_11309,N_13439);
nor U16289 (N_16289,N_12577,N_11193);
and U16290 (N_16290,N_14127,N_11855);
and U16291 (N_16291,N_11566,N_13315);
nor U16292 (N_16292,N_11218,N_13380);
nand U16293 (N_16293,N_13534,N_12060);
and U16294 (N_16294,N_12562,N_11460);
nand U16295 (N_16295,N_14719,N_14171);
xor U16296 (N_16296,N_12005,N_12201);
or U16297 (N_16297,N_10997,N_10467);
or U16298 (N_16298,N_10785,N_12605);
nand U16299 (N_16299,N_13473,N_12908);
nand U16300 (N_16300,N_10782,N_12044);
xor U16301 (N_16301,N_12822,N_12636);
or U16302 (N_16302,N_11723,N_11138);
xor U16303 (N_16303,N_14483,N_14959);
xnor U16304 (N_16304,N_12268,N_10965);
nor U16305 (N_16305,N_10708,N_11165);
and U16306 (N_16306,N_10623,N_13957);
or U16307 (N_16307,N_12807,N_14608);
nand U16308 (N_16308,N_14113,N_13566);
nor U16309 (N_16309,N_13587,N_12379);
or U16310 (N_16310,N_13306,N_11528);
nor U16311 (N_16311,N_13268,N_14071);
nand U16312 (N_16312,N_12111,N_13005);
and U16313 (N_16313,N_10471,N_13704);
or U16314 (N_16314,N_12288,N_11719);
and U16315 (N_16315,N_14203,N_11913);
or U16316 (N_16316,N_11161,N_14970);
or U16317 (N_16317,N_12120,N_14519);
nand U16318 (N_16318,N_14931,N_13675);
nand U16319 (N_16319,N_12489,N_14317);
nor U16320 (N_16320,N_11710,N_10527);
nor U16321 (N_16321,N_11629,N_11437);
or U16322 (N_16322,N_14303,N_12677);
and U16323 (N_16323,N_10715,N_10279);
nand U16324 (N_16324,N_10693,N_10031);
nor U16325 (N_16325,N_14436,N_11216);
and U16326 (N_16326,N_13855,N_12302);
xnor U16327 (N_16327,N_12866,N_12836);
nor U16328 (N_16328,N_12666,N_14967);
and U16329 (N_16329,N_14513,N_12235);
xor U16330 (N_16330,N_12134,N_14419);
xor U16331 (N_16331,N_11928,N_11463);
and U16332 (N_16332,N_14357,N_11668);
xor U16333 (N_16333,N_13588,N_12175);
and U16334 (N_16334,N_11681,N_11834);
or U16335 (N_16335,N_13802,N_10525);
and U16336 (N_16336,N_10124,N_13244);
nor U16337 (N_16337,N_10420,N_12478);
or U16338 (N_16338,N_14578,N_13390);
or U16339 (N_16339,N_13914,N_10009);
nand U16340 (N_16340,N_12880,N_13233);
nand U16341 (N_16341,N_12122,N_10728);
nor U16342 (N_16342,N_10150,N_10378);
nand U16343 (N_16343,N_12688,N_12883);
nor U16344 (N_16344,N_11825,N_12967);
xnor U16345 (N_16345,N_11612,N_13673);
and U16346 (N_16346,N_10794,N_10879);
nor U16347 (N_16347,N_11518,N_11262);
xnor U16348 (N_16348,N_11588,N_11114);
nor U16349 (N_16349,N_12159,N_11640);
nor U16350 (N_16350,N_14603,N_14185);
nand U16351 (N_16351,N_13634,N_11459);
nand U16352 (N_16352,N_14486,N_10971);
and U16353 (N_16353,N_13369,N_10475);
and U16354 (N_16354,N_14529,N_10748);
and U16355 (N_16355,N_12296,N_14198);
or U16356 (N_16356,N_13280,N_12461);
or U16357 (N_16357,N_14878,N_11349);
nor U16358 (N_16358,N_14947,N_11974);
xor U16359 (N_16359,N_11903,N_11448);
or U16360 (N_16360,N_10893,N_10183);
and U16361 (N_16361,N_11960,N_10842);
nand U16362 (N_16362,N_14207,N_14077);
nand U16363 (N_16363,N_12933,N_11074);
nor U16364 (N_16364,N_10535,N_13004);
nor U16365 (N_16365,N_11170,N_12323);
nor U16366 (N_16366,N_13633,N_13311);
nand U16367 (N_16367,N_11946,N_11951);
and U16368 (N_16368,N_13982,N_13570);
or U16369 (N_16369,N_10834,N_11392);
and U16370 (N_16370,N_11310,N_14795);
or U16371 (N_16371,N_14488,N_12771);
and U16372 (N_16372,N_11916,N_10068);
xnor U16373 (N_16373,N_11564,N_10047);
nand U16374 (N_16374,N_11505,N_10846);
and U16375 (N_16375,N_14248,N_10579);
nand U16376 (N_16376,N_14205,N_14394);
nor U16377 (N_16377,N_10585,N_14543);
nand U16378 (N_16378,N_10661,N_12901);
or U16379 (N_16379,N_10077,N_14270);
xor U16380 (N_16380,N_12433,N_14311);
nor U16381 (N_16381,N_13486,N_13796);
xor U16382 (N_16382,N_14081,N_10752);
or U16383 (N_16383,N_12964,N_14359);
nand U16384 (N_16384,N_13285,N_10771);
nor U16385 (N_16385,N_11307,N_10625);
nand U16386 (N_16386,N_14485,N_13954);
nor U16387 (N_16387,N_13740,N_10287);
and U16388 (N_16388,N_13751,N_14752);
and U16389 (N_16389,N_10215,N_14885);
nand U16390 (N_16390,N_10446,N_11198);
nand U16391 (N_16391,N_10807,N_14001);
nor U16392 (N_16392,N_12145,N_12337);
nand U16393 (N_16393,N_11734,N_11271);
nor U16394 (N_16394,N_10633,N_10094);
nor U16395 (N_16395,N_13864,N_10318);
or U16396 (N_16396,N_13589,N_13787);
nand U16397 (N_16397,N_12759,N_10465);
nor U16398 (N_16398,N_11496,N_14843);
nand U16399 (N_16399,N_11013,N_12309);
nand U16400 (N_16400,N_14673,N_13033);
nand U16401 (N_16401,N_10493,N_11691);
nand U16402 (N_16402,N_11451,N_13466);
nand U16403 (N_16403,N_13276,N_11783);
xnor U16404 (N_16404,N_13300,N_11608);
or U16405 (N_16405,N_10169,N_12720);
nand U16406 (N_16406,N_14539,N_10055);
or U16407 (N_16407,N_13656,N_11294);
nor U16408 (N_16408,N_12402,N_10638);
or U16409 (N_16409,N_11149,N_11001);
nor U16410 (N_16410,N_10466,N_12801);
nand U16411 (N_16411,N_11733,N_10904);
and U16412 (N_16412,N_12335,N_11990);
nand U16413 (N_16413,N_13153,N_11938);
or U16414 (N_16414,N_14607,N_14264);
or U16415 (N_16415,N_13623,N_11237);
xnor U16416 (N_16416,N_12775,N_13267);
or U16417 (N_16417,N_11836,N_13995);
and U16418 (N_16418,N_13548,N_10537);
or U16419 (N_16419,N_14583,N_11594);
nor U16420 (N_16420,N_14974,N_14036);
or U16421 (N_16421,N_14965,N_11275);
nor U16422 (N_16422,N_12152,N_12738);
nor U16423 (N_16423,N_12881,N_12576);
nor U16424 (N_16424,N_14389,N_14157);
or U16425 (N_16425,N_10115,N_13247);
nor U16426 (N_16426,N_14829,N_10184);
and U16427 (N_16427,N_12113,N_12935);
or U16428 (N_16428,N_11169,N_12919);
nand U16429 (N_16429,N_11577,N_13610);
nor U16430 (N_16430,N_13583,N_14722);
or U16431 (N_16431,N_10757,N_13961);
nand U16432 (N_16432,N_14217,N_12144);
nand U16433 (N_16433,N_14307,N_12413);
xnor U16434 (N_16434,N_14388,N_10624);
nor U16435 (N_16435,N_14445,N_13428);
nor U16436 (N_16436,N_10165,N_11381);
nand U16437 (N_16437,N_10182,N_12410);
or U16438 (N_16438,N_13349,N_11292);
and U16439 (N_16439,N_12391,N_14230);
and U16440 (N_16440,N_13156,N_10843);
nand U16441 (N_16441,N_12639,N_13307);
and U16442 (N_16442,N_14998,N_13485);
xor U16443 (N_16443,N_12198,N_10266);
nor U16444 (N_16444,N_14025,N_14018);
or U16445 (N_16445,N_13918,N_13437);
nor U16446 (N_16446,N_12354,N_12526);
xor U16447 (N_16447,N_10199,N_13550);
nor U16448 (N_16448,N_11901,N_12444);
nor U16449 (N_16449,N_11839,N_12382);
nor U16450 (N_16450,N_11419,N_10552);
nor U16451 (N_16451,N_12062,N_11134);
and U16452 (N_16452,N_10026,N_13070);
xor U16453 (N_16453,N_10120,N_10839);
nor U16454 (N_16454,N_11244,N_11233);
nand U16455 (N_16455,N_13495,N_14349);
and U16456 (N_16456,N_13254,N_11597);
or U16457 (N_16457,N_12034,N_13295);
nand U16458 (N_16458,N_13504,N_12166);
or U16459 (N_16459,N_14639,N_11046);
xnor U16460 (N_16460,N_14704,N_10155);
nor U16461 (N_16461,N_13090,N_13154);
nor U16462 (N_16462,N_14718,N_11609);
nor U16463 (N_16463,N_13638,N_12084);
nand U16464 (N_16464,N_14447,N_12468);
or U16465 (N_16465,N_14570,N_13007);
nor U16466 (N_16466,N_11259,N_10541);
or U16467 (N_16467,N_14393,N_13432);
nor U16468 (N_16468,N_10363,N_13963);
xnor U16469 (N_16469,N_11337,N_14721);
and U16470 (N_16470,N_10286,N_14153);
and U16471 (N_16471,N_14128,N_12714);
nand U16472 (N_16472,N_12411,N_14953);
xnor U16473 (N_16473,N_12348,N_12092);
nor U16474 (N_16474,N_12080,N_14093);
or U16475 (N_16475,N_13303,N_13593);
xor U16476 (N_16476,N_14880,N_14874);
nand U16477 (N_16477,N_11449,N_13666);
nand U16478 (N_16478,N_13625,N_13456);
and U16479 (N_16479,N_13631,N_11717);
or U16480 (N_16480,N_14794,N_10589);
nor U16481 (N_16481,N_12163,N_14060);
nand U16482 (N_16482,N_10460,N_10023);
nand U16483 (N_16483,N_14631,N_12003);
nor U16484 (N_16484,N_13766,N_11055);
or U16485 (N_16485,N_11537,N_13869);
and U16486 (N_16486,N_11972,N_12519);
and U16487 (N_16487,N_13684,N_10683);
or U16488 (N_16488,N_14890,N_11940);
nand U16489 (N_16489,N_11154,N_13728);
xor U16490 (N_16490,N_14214,N_13440);
or U16491 (N_16491,N_12594,N_12907);
nor U16492 (N_16492,N_10373,N_11917);
nand U16493 (N_16493,N_14380,N_10713);
and U16494 (N_16494,N_12843,N_13331);
nor U16495 (N_16495,N_12353,N_12018);
or U16496 (N_16496,N_11815,N_11677);
and U16497 (N_16497,N_12683,N_11845);
nor U16498 (N_16498,N_10284,N_14245);
nand U16499 (N_16499,N_12238,N_14376);
nand U16500 (N_16500,N_14476,N_12560);
xnor U16501 (N_16501,N_10954,N_12325);
nand U16502 (N_16502,N_11603,N_14321);
nor U16503 (N_16503,N_14711,N_11002);
and U16504 (N_16504,N_14297,N_11674);
or U16505 (N_16505,N_11228,N_10763);
nor U16506 (N_16506,N_10317,N_14011);
and U16507 (N_16507,N_13106,N_12032);
xnor U16508 (N_16508,N_13837,N_14999);
nand U16509 (N_16509,N_12733,N_11042);
and U16510 (N_16510,N_11084,N_12289);
nand U16511 (N_16511,N_14779,N_12414);
or U16512 (N_16512,N_10976,N_11068);
nor U16513 (N_16513,N_12437,N_11643);
and U16514 (N_16514,N_12536,N_12665);
nor U16515 (N_16515,N_10221,N_12406);
xor U16516 (N_16516,N_13895,N_12300);
or U16517 (N_16517,N_14275,N_11106);
nor U16518 (N_16518,N_11512,N_10934);
or U16519 (N_16519,N_12320,N_11031);
nor U16520 (N_16520,N_12341,N_12219);
or U16521 (N_16521,N_12563,N_10152);
nor U16522 (N_16522,N_10316,N_14283);
nor U16523 (N_16523,N_10532,N_11201);
and U16524 (N_16524,N_10118,N_12077);
or U16525 (N_16525,N_10444,N_13946);
nor U16526 (N_16526,N_12991,N_14211);
nor U16527 (N_16527,N_14993,N_13430);
and U16528 (N_16528,N_11335,N_10876);
and U16529 (N_16529,N_11209,N_10252);
or U16530 (N_16530,N_13768,N_11651);
or U16531 (N_16531,N_10909,N_12466);
and U16532 (N_16532,N_14194,N_11793);
nand U16533 (N_16533,N_11744,N_11290);
or U16534 (N_16534,N_14867,N_13655);
and U16535 (N_16535,N_14502,N_11563);
and U16536 (N_16536,N_10050,N_10445);
and U16537 (N_16537,N_12249,N_12882);
nor U16538 (N_16538,N_12857,N_11919);
nor U16539 (N_16539,N_12064,N_10685);
nand U16540 (N_16540,N_12352,N_12305);
or U16541 (N_16541,N_10275,N_12736);
nor U16542 (N_16542,N_10519,N_12592);
xor U16543 (N_16543,N_13056,N_13157);
nor U16544 (N_16544,N_13664,N_12306);
or U16545 (N_16545,N_14985,N_12026);
nor U16546 (N_16546,N_10282,N_11472);
or U16547 (N_16547,N_14315,N_10309);
nand U16548 (N_16548,N_11329,N_14370);
and U16549 (N_16549,N_14992,N_13344);
or U16550 (N_16550,N_10347,N_10038);
and U16551 (N_16551,N_13211,N_11241);
nand U16552 (N_16552,N_13743,N_11729);
and U16553 (N_16553,N_13779,N_10764);
and U16554 (N_16554,N_14379,N_14960);
xnor U16555 (N_16555,N_14224,N_14063);
or U16556 (N_16556,N_10690,N_13032);
and U16557 (N_16557,N_14119,N_12851);
nand U16558 (N_16558,N_13759,N_14237);
or U16559 (N_16559,N_10594,N_13087);
nor U16560 (N_16560,N_14040,N_10479);
nand U16561 (N_16561,N_12838,N_12516);
nand U16562 (N_16562,N_12812,N_10526);
nand U16563 (N_16563,N_13615,N_10168);
and U16564 (N_16564,N_11694,N_13333);
nand U16565 (N_16565,N_10645,N_14582);
or U16566 (N_16566,N_10058,N_12808);
or U16567 (N_16567,N_11560,N_14433);
and U16568 (N_16568,N_12768,N_10865);
or U16569 (N_16569,N_14202,N_11432);
nor U16570 (N_16570,N_10186,N_12123);
and U16571 (N_16571,N_12750,N_11319);
and U16572 (N_16572,N_10346,N_10643);
nand U16573 (N_16573,N_12589,N_12623);
and U16574 (N_16574,N_12756,N_10766);
or U16575 (N_16575,N_11944,N_10826);
and U16576 (N_16576,N_12705,N_11781);
or U16577 (N_16577,N_13399,N_12436);
nand U16578 (N_16578,N_10730,N_14263);
and U16579 (N_16579,N_14942,N_11391);
or U16580 (N_16580,N_12267,N_11469);
xnor U16581 (N_16581,N_12730,N_10932);
and U16582 (N_16582,N_10141,N_11858);
nand U16583 (N_16583,N_12164,N_11175);
nand U16584 (N_16584,N_10606,N_13237);
nor U16585 (N_16585,N_11738,N_13609);
nor U16586 (N_16586,N_11036,N_12056);
xnor U16587 (N_16587,N_14455,N_12454);
nor U16588 (N_16588,N_10342,N_10795);
and U16589 (N_16589,N_14326,N_13060);
and U16590 (N_16590,N_14658,N_14287);
or U16591 (N_16591,N_12037,N_11353);
or U16592 (N_16592,N_13640,N_10193);
or U16593 (N_16593,N_13809,N_12561);
nor U16594 (N_16594,N_13118,N_14324);
nand U16595 (N_16595,N_14524,N_12994);
nand U16596 (N_16596,N_14008,N_13313);
nor U16597 (N_16597,N_14212,N_11731);
nand U16598 (N_16598,N_12262,N_11763);
or U16599 (N_16599,N_10388,N_13272);
nor U16600 (N_16600,N_12329,N_10176);
nor U16601 (N_16601,N_13601,N_13951);
or U16602 (N_16602,N_13360,N_11868);
xor U16603 (N_16603,N_10798,N_12112);
nor U16604 (N_16604,N_11263,N_13261);
nor U16605 (N_16605,N_12010,N_12387);
or U16606 (N_16606,N_10975,N_12350);
nor U16607 (N_16607,N_13788,N_12664);
and U16608 (N_16608,N_12761,N_13243);
xnor U16609 (N_16609,N_13190,N_10707);
or U16610 (N_16610,N_13305,N_10792);
xor U16611 (N_16611,N_14805,N_12886);
nor U16612 (N_16612,N_11840,N_11443);
and U16613 (N_16613,N_12211,N_11937);
or U16614 (N_16614,N_13646,N_12472);
xor U16615 (N_16615,N_13826,N_13392);
nor U16616 (N_16616,N_14638,N_11105);
and U16617 (N_16617,N_11771,N_12231);
xor U16618 (N_16618,N_14043,N_10012);
and U16619 (N_16619,N_10958,N_10211);
nand U16620 (N_16620,N_11255,N_14320);
nand U16621 (N_16621,N_12317,N_13041);
nor U16622 (N_16622,N_12903,N_12377);
nor U16623 (N_16623,N_13323,N_14280);
and U16624 (N_16624,N_12272,N_14250);
and U16625 (N_16625,N_12484,N_11665);
and U16626 (N_16626,N_14072,N_14641);
nor U16627 (N_16627,N_12256,N_13560);
nand U16628 (N_16628,N_13540,N_12740);
and U16629 (N_16629,N_11808,N_10160);
or U16630 (N_16630,N_10635,N_13312);
or U16631 (N_16631,N_11418,N_14412);
nor U16632 (N_16632,N_14310,N_11357);
nand U16633 (N_16633,N_12567,N_14177);
nand U16634 (N_16634,N_10370,N_14226);
or U16635 (N_16635,N_10320,N_13346);
nand U16636 (N_16636,N_14435,N_10477);
or U16637 (N_16637,N_10334,N_11352);
xor U16638 (N_16638,N_11356,N_11501);
or U16639 (N_16639,N_11054,N_10605);
nor U16640 (N_16640,N_12894,N_10508);
nor U16641 (N_16641,N_13969,N_13782);
nor U16642 (N_16642,N_10350,N_13750);
or U16643 (N_16643,N_13322,N_11129);
nand U16644 (N_16644,N_14322,N_13586);
and U16645 (N_16645,N_10611,N_12074);
nor U16646 (N_16646,N_12443,N_12347);
and U16647 (N_16647,N_12602,N_10164);
xnor U16648 (N_16648,N_10260,N_13791);
nor U16649 (N_16649,N_13984,N_11086);
nand U16650 (N_16650,N_11767,N_14642);
and U16651 (N_16651,N_11348,N_12529);
and U16652 (N_16652,N_13116,N_11061);
and U16653 (N_16653,N_10470,N_10362);
nor U16654 (N_16654,N_11023,N_13702);
nor U16655 (N_16655,N_12739,N_12961);
nand U16656 (N_16656,N_10619,N_14769);
and U16657 (N_16657,N_13172,N_11558);
xnor U16658 (N_16658,N_12130,N_14898);
xnor U16659 (N_16659,N_13366,N_13171);
nor U16660 (N_16660,N_13487,N_10268);
and U16661 (N_16661,N_14585,N_13465);
and U16662 (N_16662,N_13104,N_14980);
nor U16663 (N_16663,N_11012,N_14170);
xor U16664 (N_16664,N_14424,N_11422);
nor U16665 (N_16665,N_11778,N_12785);
nor U16666 (N_16666,N_11978,N_12674);
nor U16667 (N_16667,N_12875,N_13082);
and U16668 (N_16668,N_12614,N_13238);
nor U16669 (N_16669,N_12735,N_12090);
or U16670 (N_16670,N_13200,N_10485);
and U16671 (N_16671,N_12902,N_13980);
or U16672 (N_16672,N_14727,N_14655);
nor U16673 (N_16673,N_12301,N_11788);
xnor U16674 (N_16674,N_11510,N_14755);
xor U16675 (N_16675,N_14567,N_13345);
and U16676 (N_16676,N_14462,N_14386);
nor U16677 (N_16677,N_11614,N_13860);
nand U16678 (N_16678,N_10524,N_14932);
nand U16679 (N_16679,N_10438,N_13661);
nor U16680 (N_16680,N_14314,N_10495);
nand U16681 (N_16681,N_10296,N_10512);
and U16682 (N_16682,N_10030,N_14257);
nor U16683 (N_16683,N_11308,N_13585);
nand U16684 (N_16684,N_10351,N_11983);
nand U16685 (N_16685,N_10814,N_10602);
xnor U16686 (N_16686,N_14012,N_14016);
nand U16687 (N_16687,N_10811,N_14671);
xor U16688 (N_16688,N_12421,N_14219);
or U16689 (N_16689,N_10481,N_10327);
and U16690 (N_16690,N_14143,N_14770);
or U16691 (N_16691,N_14802,N_11573);
and U16692 (N_16692,N_14124,N_13628);
or U16693 (N_16693,N_14546,N_13199);
nor U16694 (N_16694,N_12888,N_13003);
or U16695 (N_16695,N_13523,N_11755);
xor U16696 (N_16696,N_10870,N_13532);
xor U16697 (N_16697,N_14927,N_11095);
nor U16698 (N_16698,N_12225,N_10855);
and U16699 (N_16699,N_12502,N_14213);
or U16700 (N_16700,N_11526,N_14441);
and U16701 (N_16701,N_13080,N_11445);
xor U16702 (N_16702,N_12011,N_10052);
nand U16703 (N_16703,N_13904,N_11157);
nor U16704 (N_16704,N_10979,N_12638);
nor U16705 (N_16705,N_13417,N_12633);
nor U16706 (N_16706,N_11669,N_14367);
nor U16707 (N_16707,N_13040,N_10476);
or U16708 (N_16708,N_14649,N_10538);
and U16709 (N_16709,N_11770,N_12906);
xnor U16710 (N_16710,N_14118,N_14901);
nor U16711 (N_16711,N_11137,N_10126);
nand U16712 (N_16712,N_11405,N_14610);
or U16713 (N_16713,N_11618,N_14277);
nor U16714 (N_16714,N_10564,N_12158);
nand U16715 (N_16715,N_11798,N_13464);
nand U16716 (N_16716,N_13677,N_14131);
xnor U16717 (N_16717,N_12539,N_11427);
nand U16718 (N_16718,N_13402,N_10367);
nand U16719 (N_16719,N_10907,N_10857);
or U16720 (N_16720,N_10159,N_10982);
nor U16721 (N_16721,N_12805,N_12224);
nor U16722 (N_16722,N_10500,N_11190);
xor U16723 (N_16723,N_11315,N_12898);
and U16724 (N_16724,N_10671,N_10100);
nor U16725 (N_16725,N_12259,N_14591);
nor U16726 (N_16726,N_13844,N_11077);
or U16727 (N_16727,N_13321,N_14643);
nand U16728 (N_16728,N_11688,N_10883);
or U16729 (N_16729,N_13398,N_12095);
or U16730 (N_16730,N_14020,N_14601);
or U16731 (N_16731,N_12495,N_10569);
nand U16732 (N_16732,N_14961,N_14797);
or U16733 (N_16733,N_14936,N_11707);
or U16734 (N_16734,N_11764,N_14385);
or U16735 (N_16735,N_12114,N_10365);
and U16736 (N_16736,N_14471,N_10560);
or U16737 (N_16737,N_11777,N_11377);
or U16738 (N_16738,N_11641,N_12177);
or U16739 (N_16739,N_13891,N_11958);
and U16740 (N_16740,N_13515,N_10984);
nand U16741 (N_16741,N_10189,N_10344);
nand U16742 (N_16742,N_11499,N_10694);
or U16743 (N_16743,N_10117,N_11486);
nand U16744 (N_16744,N_11794,N_12976);
xor U16745 (N_16745,N_13287,N_11804);
nand U16746 (N_16746,N_10051,N_10655);
xor U16747 (N_16747,N_10474,N_12802);
nand U16748 (N_16748,N_12367,N_13084);
nor U16749 (N_16749,N_14331,N_12821);
nor U16750 (N_16750,N_10306,N_13278);
nor U16751 (N_16751,N_13395,N_14897);
or U16752 (N_16752,N_14288,N_12941);
or U16753 (N_16753,N_10382,N_12985);
or U16754 (N_16754,N_13393,N_10630);
nor U16755 (N_16755,N_14968,N_14946);
and U16756 (N_16756,N_13377,N_11616);
and U16757 (N_16757,N_10105,N_10529);
and U16758 (N_16758,N_14353,N_14863);
xor U16759 (N_16759,N_13732,N_13222);
nand U16760 (N_16760,N_14913,N_10705);
and U16761 (N_16761,N_13739,N_12544);
or U16762 (N_16762,N_14882,N_10881);
or U16763 (N_16763,N_14261,N_13674);
and U16764 (N_16764,N_14044,N_11520);
nor U16765 (N_16765,N_10461,N_11383);
xnor U16766 (N_16766,N_14233,N_14045);
nand U16767 (N_16767,N_13259,N_10338);
and U16768 (N_16768,N_11251,N_12374);
nor U16769 (N_16769,N_12456,N_14620);
or U16770 (N_16770,N_13755,N_10522);
nor U16771 (N_16771,N_11976,N_11632);
nand U16772 (N_16772,N_14647,N_14629);
nand U16773 (N_16773,N_14680,N_14666);
and U16774 (N_16774,N_10885,N_13799);
nand U16775 (N_16775,N_11037,N_13310);
nand U16776 (N_16776,N_12294,N_10372);
nor U16777 (N_16777,N_10022,N_12568);
and U16778 (N_16778,N_13094,N_10587);
and U16779 (N_16779,N_12772,N_13109);
or U16780 (N_16780,N_11488,N_13688);
or U16781 (N_16781,N_13614,N_10796);
and U16782 (N_16782,N_11906,N_11658);
nand U16783 (N_16783,N_13558,N_10825);
xor U16784 (N_16784,N_14163,N_14652);
nor U16785 (N_16785,N_11452,N_13897);
or U16786 (N_16786,N_13308,N_14693);
nor U16787 (N_16787,N_13198,N_11523);
and U16788 (N_16788,N_10897,N_14534);
xnor U16789 (N_16789,N_13161,N_14204);
and U16790 (N_16790,N_11440,N_11897);
or U16791 (N_16791,N_14925,N_12800);
nor U16792 (N_16792,N_14784,N_11663);
nor U16793 (N_16793,N_12448,N_14478);
xnor U16794 (N_16794,N_14108,N_14274);
xor U16795 (N_16795,N_10087,N_14933);
or U16796 (N_16796,N_14006,N_14333);
nor U16797 (N_16797,N_13251,N_12364);
nor U16798 (N_16798,N_10590,N_13747);
and U16799 (N_16799,N_11215,N_12014);
and U16800 (N_16800,N_11098,N_13513);
nand U16801 (N_16801,N_10962,N_13341);
nand U16802 (N_16802,N_11689,N_12494);
or U16803 (N_16803,N_13147,N_13752);
nor U16804 (N_16804,N_11915,N_14648);
and U16805 (N_16805,N_14726,N_11208);
and U16806 (N_16806,N_13867,N_13736);
nand U16807 (N_16807,N_14604,N_12715);
nor U16808 (N_16808,N_12250,N_13494);
xor U16809 (N_16809,N_13619,N_14135);
nand U16810 (N_16810,N_14383,N_11420);
or U16811 (N_16811,N_11032,N_11298);
or U16812 (N_16812,N_11385,N_11708);
or U16813 (N_16813,N_10424,N_12809);
nor U16814 (N_16814,N_14571,N_13368);
nand U16815 (N_16815,N_10230,N_11301);
and U16816 (N_16816,N_10311,N_12554);
nand U16817 (N_16817,N_12946,N_12497);
or U16818 (N_16818,N_10875,N_14341);
and U16819 (N_16819,N_10536,N_10253);
nor U16820 (N_16820,N_12445,N_13885);
and U16821 (N_16821,N_11821,N_13334);
xnor U16822 (N_16822,N_10634,N_12376);
nor U16823 (N_16823,N_12872,N_14038);
or U16824 (N_16824,N_14005,N_14785);
or U16825 (N_16825,N_13685,N_13613);
nor U16826 (N_16826,N_11706,N_14873);
nand U16827 (N_16827,N_12958,N_12923);
nand U16828 (N_16828,N_10450,N_12082);
nand U16829 (N_16829,N_11411,N_14899);
or U16830 (N_16830,N_13637,N_11109);
nand U16831 (N_16831,N_12168,N_14657);
nor U16832 (N_16832,N_12240,N_12604);
and U16833 (N_16833,N_12686,N_14244);
nor U16834 (N_16834,N_11966,N_13749);
or U16835 (N_16835,N_10663,N_12615);
nor U16836 (N_16836,N_12725,N_14183);
nand U16837 (N_16837,N_12701,N_13453);
xnor U16838 (N_16838,N_13123,N_14789);
or U16839 (N_16839,N_11484,N_10969);
and U16840 (N_16840,N_11045,N_10620);
xor U16841 (N_16841,N_13996,N_10110);
nor U16842 (N_16842,N_12506,N_10016);
nor U16843 (N_16843,N_14956,N_11461);
nand U16844 (N_16844,N_12188,N_14587);
or U16845 (N_16845,N_10737,N_10568);
or U16846 (N_16846,N_13764,N_10987);
nor U16847 (N_16847,N_10612,N_13831);
nand U16848 (N_16848,N_13086,N_13772);
nand U16849 (N_16849,N_11072,N_10328);
or U16850 (N_16850,N_12524,N_11424);
or U16851 (N_16851,N_11334,N_10711);
xnor U16852 (N_16852,N_10175,N_12176);
nor U16853 (N_16853,N_12786,N_11394);
nor U16854 (N_16854,N_11152,N_13541);
xnor U16855 (N_16855,N_13490,N_10554);
xnor U16856 (N_16856,N_14439,N_14372);
nand U16857 (N_16857,N_12719,N_12499);
xor U16858 (N_16858,N_11570,N_12476);
or U16859 (N_16859,N_13668,N_10570);
or U16860 (N_16860,N_11995,N_14622);
nor U16861 (N_16861,N_13776,N_13815);
nor U16862 (N_16862,N_12828,N_11455);
nand U16863 (N_16863,N_13705,N_12590);
or U16864 (N_16864,N_13769,N_14255);
or U16865 (N_16865,N_14923,N_14675);
or U16866 (N_16866,N_13425,N_14778);
nand U16867 (N_16867,N_13803,N_14715);
nand U16868 (N_16868,N_10853,N_13940);
or U16869 (N_16869,N_14678,N_10872);
nand U16870 (N_16870,N_11645,N_10915);
nand U16871 (N_16871,N_11955,N_14085);
nor U16872 (N_16872,N_13687,N_14408);
nor U16873 (N_16873,N_14228,N_13679);
or U16874 (N_16874,N_11583,N_11328);
or U16875 (N_16875,N_14225,N_13520);
nand U16876 (N_16876,N_11162,N_12295);
or U16877 (N_16877,N_13530,N_13197);
and U16878 (N_16878,N_11303,N_11575);
or U16879 (N_16879,N_11330,N_10561);
nand U16880 (N_16880,N_13257,N_10706);
or U16881 (N_16881,N_11889,N_10276);
and U16882 (N_16882,N_10384,N_12273);
and U16883 (N_16883,N_12937,N_11277);
nand U16884 (N_16884,N_12609,N_14609);
nor U16885 (N_16885,N_12505,N_12463);
or U16886 (N_16886,N_13745,N_12481);
and U16887 (N_16887,N_13932,N_11865);
nor U16888 (N_16888,N_10040,N_11572);
nand U16889 (N_16889,N_14420,N_14776);
nand U16890 (N_16890,N_14305,N_14552);
and U16891 (N_16891,N_13535,N_11856);
nand U16892 (N_16892,N_11932,N_12253);
or U16893 (N_16893,N_14474,N_12932);
nand U16894 (N_16894,N_10919,N_14096);
or U16895 (N_16895,N_12427,N_11026);
and U16896 (N_16896,N_11225,N_11064);
and U16897 (N_16897,N_13320,N_13573);
xnor U16898 (N_16898,N_10860,N_13966);
and U16899 (N_16899,N_11568,N_13993);
or U16900 (N_16900,N_12424,N_14787);
nand U16901 (N_16901,N_11103,N_14167);
nand U16902 (N_16902,N_12713,N_10397);
or U16903 (N_16903,N_14981,N_11172);
xnor U16904 (N_16904,N_10000,N_10262);
and U16905 (N_16905,N_14141,N_13132);
nor U16906 (N_16906,N_12345,N_12647);
and U16907 (N_16907,N_14452,N_13277);
nor U16908 (N_16908,N_14742,N_10691);
nor U16909 (N_16909,N_13144,N_11857);
nor U16910 (N_16910,N_10943,N_10966);
nand U16911 (N_16911,N_10680,N_11516);
xor U16912 (N_16912,N_14577,N_13193);
and U16913 (N_16913,N_10599,N_14516);
and U16914 (N_16914,N_13599,N_13427);
and U16915 (N_16915,N_13129,N_13235);
or U16916 (N_16916,N_11176,N_14415);
nand U16917 (N_16917,N_11025,N_13700);
and U16918 (N_16918,N_11787,N_14401);
nand U16919 (N_16919,N_14411,N_14636);
and U16920 (N_16920,N_13861,N_14668);
nand U16921 (N_16921,N_12697,N_13746);
and U16922 (N_16922,N_13785,N_14391);
or U16923 (N_16923,N_10361,N_13240);
nor U16924 (N_16924,N_10079,N_14818);
nor U16925 (N_16925,N_14251,N_12104);
nor U16926 (N_16926,N_11279,N_13407);
nand U16927 (N_16927,N_14373,N_10425);
nor U16928 (N_16928,N_11977,N_11930);
and U16929 (N_16929,N_13733,N_14505);
xnor U16930 (N_16930,N_13429,N_10084);
nor U16931 (N_16931,N_10037,N_14681);
and U16932 (N_16932,N_12963,N_11695);
nor U16933 (N_16933,N_14870,N_10687);
nor U16934 (N_16934,N_14914,N_11008);
nand U16935 (N_16935,N_14007,N_14031);
or U16936 (N_16936,N_13489,N_10913);
and U16937 (N_16937,N_10862,N_10941);
nand U16938 (N_16938,N_11982,N_10996);
nand U16939 (N_16939,N_14508,N_10305);
xor U16940 (N_16940,N_12429,N_13248);
nor U16941 (N_16941,N_12237,N_13850);
and U16942 (N_16942,N_13549,N_10163);
and U16943 (N_16943,N_10064,N_10261);
or U16944 (N_16944,N_14111,N_12117);
or U16945 (N_16945,N_12079,N_12691);
and U16946 (N_16946,N_10171,N_14024);
nor U16947 (N_16947,N_13174,N_14013);
and U16948 (N_16948,N_13527,N_10271);
xnor U16949 (N_16949,N_12118,N_13378);
or U16950 (N_16950,N_10335,N_12500);
nand U16951 (N_16951,N_13110,N_14223);
xor U16952 (N_16952,N_13220,N_10158);
nand U16953 (N_16953,N_11276,N_10733);
and U16954 (N_16954,N_13793,N_11605);
and U16955 (N_16955,N_11806,N_12698);
nor U16956 (N_16956,N_13185,N_13962);
or U16957 (N_16957,N_10762,N_11257);
or U16958 (N_16958,N_13419,N_14663);
nor U16959 (N_16959,N_14716,N_12910);
nor U16960 (N_16960,N_13915,N_10502);
or U16961 (N_16961,N_11011,N_13408);
or U16962 (N_16962,N_14209,N_10258);
or U16963 (N_16963,N_13052,N_14480);
and U16964 (N_16964,N_11267,N_13758);
nor U16965 (N_16965,N_12027,N_12073);
nor U16966 (N_16966,N_13594,N_14854);
nand U16967 (N_16967,N_13381,N_11376);
nor U16968 (N_16968,N_13976,N_11562);
nor U16969 (N_16969,N_11039,N_13719);
nand U16970 (N_16970,N_10812,N_11578);
or U16971 (N_16971,N_14174,N_10147);
or U16972 (N_16972,N_12283,N_11339);
nor U16973 (N_16973,N_10974,N_12321);
or U16974 (N_16974,N_10980,N_13997);
xor U16975 (N_16975,N_13053,N_13475);
or U16976 (N_16976,N_12671,N_12274);
nand U16977 (N_16977,N_11827,N_10805);
xor U16978 (N_16978,N_11140,N_12076);
nor U16979 (N_16979,N_14728,N_11789);
and U16980 (N_16980,N_10505,N_14148);
nor U16981 (N_16981,N_11370,N_10797);
and U16982 (N_16982,N_11760,N_10228);
and U16983 (N_16983,N_10033,N_12297);
nor U16984 (N_16984,N_11296,N_13990);
nor U16985 (N_16985,N_10205,N_11837);
xor U16986 (N_16986,N_10754,N_11853);
nand U16987 (N_16987,N_13840,N_11450);
or U16988 (N_16988,N_13422,N_10326);
nand U16989 (N_16989,N_13140,N_10900);
nand U16990 (N_16990,N_11943,N_10888);
nor U16991 (N_16991,N_12313,N_12420);
or U16992 (N_16992,N_10858,N_13562);
nor U16993 (N_16993,N_13061,N_14309);
or U16994 (N_16994,N_12995,N_14003);
nor U16995 (N_16995,N_13024,N_12360);
nand U16996 (N_16996,N_11902,N_14732);
or U16997 (N_16997,N_14709,N_11599);
xor U16998 (N_16998,N_10772,N_13604);
nor U16999 (N_16999,N_14971,N_11327);
or U17000 (N_17000,N_12045,N_12884);
or U17001 (N_17001,N_10970,N_10726);
nand U17002 (N_17002,N_12550,N_11948);
or U17003 (N_17003,N_10336,N_14290);
nor U17004 (N_17004,N_14477,N_11587);
nor U17005 (N_17005,N_11883,N_14676);
or U17006 (N_17006,N_13216,N_10001);
or U17007 (N_17007,N_12375,N_11204);
xnor U17008 (N_17008,N_11885,N_14262);
or U17009 (N_17009,N_10288,N_14869);
nor U17010 (N_17010,N_12311,N_14313);
nor U17011 (N_17011,N_13774,N_11028);
nor U17012 (N_17012,N_11547,N_11722);
nand U17013 (N_17013,N_10057,N_14504);
nor U17014 (N_17014,N_12075,N_11524);
nor U17015 (N_17015,N_14249,N_10829);
or U17016 (N_17016,N_14825,N_10325);
nand U17017 (N_17017,N_14739,N_13214);
nand U17018 (N_17018,N_10530,N_10925);
nor U17019 (N_17019,N_10340,N_12482);
or U17020 (N_17020,N_12395,N_11253);
or U17021 (N_17021,N_10236,N_13178);
and U17022 (N_17022,N_13536,N_10961);
nand U17023 (N_17023,N_14911,N_11160);
or U17024 (N_17024,N_10366,N_12704);
xnor U17025 (N_17025,N_12033,N_14662);
nor U17026 (N_17026,N_12369,N_10847);
nor U17027 (N_17027,N_10747,N_10930);
nor U17028 (N_17028,N_10758,N_10063);
or U17029 (N_17029,N_11287,N_11431);
nand U17030 (N_17030,N_10243,N_10767);
nor U17031 (N_17031,N_13299,N_13388);
nand U17032 (N_17032,N_14352,N_13298);
and U17033 (N_17033,N_11382,N_13603);
nor U17034 (N_17034,N_13069,N_14371);
nor U17035 (N_17035,N_10161,N_13006);
and U17036 (N_17036,N_13930,N_13316);
nand U17037 (N_17037,N_12204,N_10622);
or U17038 (N_17038,N_13173,N_11514);
or U17039 (N_17039,N_10142,N_11580);
nor U17040 (N_17040,N_11073,N_10078);
or U17041 (N_17041,N_14074,N_13468);
nor U17042 (N_17042,N_11686,N_14190);
nand U17043 (N_17043,N_12675,N_10027);
nand U17044 (N_17044,N_12911,N_11693);
nor U17045 (N_17045,N_13414,N_10494);
nand U17046 (N_17046,N_14112,N_12331);
nor U17047 (N_17047,N_13469,N_12732);
xor U17048 (N_17048,N_14073,N_14041);
and U17049 (N_17049,N_11784,N_11373);
nor U17050 (N_17050,N_11698,N_11822);
or U17051 (N_17051,N_11592,N_14857);
and U17052 (N_17052,N_10044,N_11748);
nor U17053 (N_17053,N_10774,N_10072);
nand U17054 (N_17054,N_13373,N_10076);
and U17055 (N_17055,N_12234,N_13284);
or U17056 (N_17056,N_11250,N_14132);
and U17057 (N_17057,N_10703,N_13832);
nand U17058 (N_17058,N_13095,N_14588);
or U17059 (N_17059,N_14151,N_11497);
xnor U17060 (N_17060,N_13929,N_13409);
and U17061 (N_17061,N_14456,N_12280);
nand U17062 (N_17062,N_14820,N_13442);
nand U17063 (N_17063,N_13968,N_11517);
and U17064 (N_17064,N_13680,N_11752);
and U17065 (N_17065,N_10828,N_10180);
xor U17066 (N_17066,N_14102,N_14640);
and U17067 (N_17067,N_10081,N_13482);
nor U17068 (N_17068,N_10308,N_13245);
nand U17069 (N_17069,N_10921,N_10114);
xnor U17070 (N_17070,N_11223,N_10080);
nand U17071 (N_17071,N_10859,N_11732);
and U17072 (N_17072,N_13055,N_14361);
and U17073 (N_17073,N_14150,N_12612);
or U17074 (N_17074,N_11163,N_12817);
or U17075 (N_17075,N_14595,N_12885);
nor U17076 (N_17076,N_12278,N_11684);
and U17077 (N_17077,N_12753,N_11675);
nor U17078 (N_17078,N_11726,N_11935);
nor U17079 (N_17079,N_12419,N_11178);
and U17080 (N_17080,N_11569,N_11435);
xor U17081 (N_17081,N_12251,N_13158);
or U17082 (N_17082,N_13066,N_10668);
nor U17083 (N_17083,N_12863,N_14919);
nand U17084 (N_17084,N_12997,N_10201);
or U17085 (N_17085,N_12655,N_12464);
or U17086 (N_17086,N_12136,N_12362);
and U17087 (N_17087,N_13296,N_14375);
or U17088 (N_17088,N_10804,N_10358);
or U17089 (N_17089,N_10319,N_11561);
and U17090 (N_17090,N_10600,N_10303);
nor U17091 (N_17091,N_11506,N_10902);
or U17092 (N_17092,N_14197,N_14189);
nor U17093 (N_17093,N_14278,N_11081);
and U17094 (N_17094,N_11549,N_10851);
nor U17095 (N_17095,N_10404,N_12938);
nand U17096 (N_17096,N_11226,N_14052);
nor U17097 (N_17097,N_11261,N_14192);
and U17098 (N_17098,N_11622,N_10873);
and U17099 (N_17099,N_14062,N_11358);
or U17100 (N_17100,N_11186,N_10473);
xnor U17101 (N_17101,N_12729,N_10492);
nor U17102 (N_17102,N_12206,N_13713);
nand U17103 (N_17103,N_10743,N_14136);
nor U17104 (N_17104,N_12755,N_13279);
or U17105 (N_17105,N_11811,N_13474);
and U17106 (N_17106,N_11941,N_12281);
nor U17107 (N_17107,N_10688,N_10429);
and U17108 (N_17108,N_11212,N_11546);
and U17109 (N_17109,N_13449,N_14554);
nand U17110 (N_17110,N_13544,N_11227);
nand U17111 (N_17111,N_13385,N_10020);
or U17112 (N_17112,N_10013,N_10698);
or U17113 (N_17113,N_12183,N_12905);
and U17114 (N_17114,N_13078,N_12422);
nand U17115 (N_17115,N_14547,N_11712);
xnor U17116 (N_17116,N_12959,N_10565);
or U17117 (N_17117,N_14527,N_11980);
nand U17118 (N_17118,N_13554,N_14598);
and U17119 (N_17119,N_10957,N_14941);
and U17120 (N_17120,N_12943,N_14912);
xor U17121 (N_17121,N_12689,N_11828);
and U17122 (N_17122,N_11593,N_14782);
nand U17123 (N_17123,N_10935,N_13988);
and U17124 (N_17124,N_14908,N_10386);
nor U17125 (N_17125,N_10017,N_10208);
nor U17126 (N_17126,N_13416,N_11791);
nand U17127 (N_17127,N_13711,N_13359);
nand U17128 (N_17128,N_12955,N_14703);
nor U17129 (N_17129,N_14979,N_11120);
or U17130 (N_17130,N_13829,N_14803);
nor U17131 (N_17131,N_14738,N_12824);
or U17132 (N_17132,N_14989,N_11464);
and U17133 (N_17133,N_13484,N_12290);
xor U17134 (N_17134,N_10540,N_11598);
nand U17135 (N_17135,N_12624,N_10200);
or U17136 (N_17136,N_14706,N_13651);
nand U17137 (N_17137,N_10641,N_13372);
nand U17138 (N_17138,N_14900,N_10032);
and U17139 (N_17139,N_12661,N_13179);
and U17140 (N_17140,N_14514,N_13354);
nand U17141 (N_17141,N_10586,N_10724);
nand U17142 (N_17142,N_12221,N_10235);
and U17143 (N_17143,N_12792,N_11158);
or U17144 (N_17144,N_12956,N_11551);
nor U17145 (N_17145,N_11480,N_14065);
nand U17146 (N_17146,N_14886,N_14218);
nor U17147 (N_17147,N_11864,N_13338);
and U17148 (N_17148,N_11947,N_13223);
and U17149 (N_17149,N_11626,N_14596);
nor U17150 (N_17150,N_14084,N_12945);
and U17151 (N_17151,N_14813,N_10300);
nand U17152 (N_17152,N_10415,N_10514);
nand U17153 (N_17153,N_10157,N_12458);
or U17154 (N_17154,N_10028,N_12180);
nor U17155 (N_17155,N_11882,N_12132);
and U17156 (N_17156,N_10231,N_13999);
and U17157 (N_17157,N_12737,N_13008);
nand U17158 (N_17158,N_11369,N_11762);
or U17159 (N_17159,N_14930,N_11844);
or U17160 (N_17160,N_12024,N_11205);
or U17161 (N_17161,N_13892,N_11515);
nor U17162 (N_17162,N_14178,N_11968);
or U17163 (N_17163,N_13846,N_14459);
nor U17164 (N_17164,N_11112,N_12757);
and U17165 (N_17165,N_10025,N_11118);
xor U17166 (N_17166,N_12814,N_12699);
nand U17167 (N_17167,N_10399,N_13150);
nand U17168 (N_17168,N_14875,N_11838);
xor U17169 (N_17169,N_11782,N_10113);
nand U17170 (N_17170,N_10917,N_13973);
nand U17171 (N_17171,N_10891,N_12105);
nor U17172 (N_17172,N_10432,N_13207);
or U17173 (N_17173,N_14431,N_11188);
xnor U17174 (N_17174,N_12909,N_10122);
nor U17175 (N_17175,N_11920,N_10109);
or U17176 (N_17176,N_13202,N_11792);
nor U17177 (N_17177,N_10618,N_14986);
nor U17178 (N_17178,N_11364,N_11964);
or U17179 (N_17179,N_12829,N_12776);
and U17180 (N_17180,N_13283,N_13435);
or U17181 (N_17181,N_14579,N_14804);
xor U17182 (N_17182,N_14049,N_11016);
xnor U17183 (N_17183,N_12947,N_11295);
and U17184 (N_17184,N_10379,N_13955);
nand U17185 (N_17185,N_12133,N_11690);
or U17186 (N_17186,N_12646,N_13865);
nor U17187 (N_17187,N_14645,N_14720);
and U17188 (N_17188,N_10656,N_14438);
xnor U17189 (N_17189,N_12918,N_11454);
nand U17190 (N_17190,N_10298,N_10784);
nand U17191 (N_17191,N_10927,N_10710);
or U17192 (N_17192,N_14033,N_13270);
nand U17193 (N_17193,N_12147,N_13786);
and U17194 (N_17194,N_11462,N_13258);
nor U17195 (N_17195,N_10412,N_11247);
and U17196 (N_17196,N_12861,N_13092);
or U17197 (N_17197,N_12488,N_11727);
nor U17198 (N_17198,N_14101,N_14095);
nand U17199 (N_17199,N_12213,N_14200);
or U17200 (N_17200,N_13020,N_10129);
or U17201 (N_17201,N_10653,N_13761);
or U17202 (N_17202,N_12078,N_13225);
nor U17203 (N_17203,N_14665,N_13516);
and U17204 (N_17204,N_10998,N_11931);
nand U17205 (N_17205,N_13507,N_11923);
and U17206 (N_17206,N_10419,N_10422);
and U17207 (N_17207,N_14294,N_13514);
nand U17208 (N_17208,N_11402,N_14350);
or U17209 (N_17209,N_12324,N_10608);
and U17210 (N_17210,N_13579,N_11179);
xnor U17211 (N_17211,N_13143,N_14015);
nor U17212 (N_17212,N_11177,N_13842);
nand U17213 (N_17213,N_11057,N_13879);
and U17214 (N_17214,N_11552,N_14161);
nor U17215 (N_17215,N_12815,N_14808);
nor U17216 (N_17216,N_14702,N_13051);
nor U17217 (N_17217,N_14191,N_10239);
nand U17218 (N_17218,N_11458,N_11925);
xnor U17219 (N_17219,N_12081,N_11033);
nand U17220 (N_17220,N_12243,N_10808);
or U17221 (N_17221,N_14338,N_13209);
xor U17222 (N_17222,N_10264,N_14017);
and U17223 (N_17223,N_13170,N_10185);
or U17224 (N_17224,N_11196,N_10374);
nor U17225 (N_17225,N_12269,N_10173);
or U17226 (N_17226,N_12284,N_11847);
nand U17227 (N_17227,N_11331,N_11521);
nor U17228 (N_17228,N_14928,N_10778);
nor U17229 (N_17229,N_12742,N_12553);
nor U17230 (N_17230,N_13880,N_13672);
or U17231 (N_17231,N_12989,N_12191);
and U17232 (N_17232,N_12257,N_10992);
xnor U17233 (N_17233,N_13653,N_12404);
nor U17234 (N_17234,N_11088,N_10832);
and U17235 (N_17235,N_11070,N_10394);
and U17236 (N_17236,N_12682,N_11721);
and U17237 (N_17237,N_10695,N_12520);
nand U17238 (N_17238,N_13707,N_12979);
nor U17239 (N_17239,N_11268,N_14756);
or U17240 (N_17240,N_14699,N_12942);
and U17241 (N_17241,N_14494,N_11071);
nor U17242 (N_17242,N_13382,N_11939);
or U17243 (N_17243,N_11374,N_13629);
nor U17244 (N_17244,N_10546,N_14149);
and U17245 (N_17245,N_11362,N_14293);
and U17246 (N_17246,N_10403,N_10593);
nand U17247 (N_17247,N_11802,N_11835);
nor U17248 (N_17248,N_12607,N_14883);
and U17249 (N_17249,N_10939,N_10486);
or U17250 (N_17250,N_12416,N_13670);
xnor U17251 (N_17251,N_11471,N_12591);
nand U17252 (N_17252,N_11595,N_10011);
nor U17253 (N_17253,N_13424,N_11895);
or U17254 (N_17254,N_12770,N_14821);
or U17255 (N_17255,N_14381,N_14838);
nand U17256 (N_17256,N_13505,N_14199);
or U17257 (N_17257,N_11981,N_12530);
nand U17258 (N_17258,N_10731,N_12953);
nand U17259 (N_17259,N_14026,N_14469);
xor U17260 (N_17260,N_12498,N_11051);
and U17261 (N_17261,N_11796,N_11848);
or U17262 (N_17262,N_10307,N_14695);
and U17263 (N_17263,N_11249,N_10578);
nor U17264 (N_17264,N_12501,N_13935);
and U17265 (N_17265,N_13647,N_12644);
nand U17266 (N_17266,N_13641,N_13659);
and U17267 (N_17267,N_10542,N_13309);
and U17268 (N_17268,N_14079,N_14839);
or U17269 (N_17269,N_14623,N_14523);
nor U17270 (N_17270,N_13807,N_14525);
or U17271 (N_17271,N_14858,N_11914);
or U17272 (N_17272,N_12672,N_10345);
xor U17273 (N_17273,N_11600,N_12712);
nor U17274 (N_17274,N_14179,N_10073);
or U17275 (N_17275,N_10139,N_11683);
nor U17276 (N_17276,N_11544,N_12975);
nor U17277 (N_17277,N_14521,N_10491);
and U17278 (N_17278,N_13375,N_13079);
or U17279 (N_17279,N_10099,N_11192);
and U17280 (N_17280,N_13531,N_13721);
and U17281 (N_17281,N_11630,N_12415);
nor U17282 (N_17282,N_14422,N_13224);
nor U17283 (N_17283,N_14935,N_14626);
and U17284 (N_17284,N_13496,N_12784);
or U17285 (N_17285,N_10216,N_10755);
or U17286 (N_17286,N_11482,N_13438);
nand U17287 (N_17287,N_10576,N_13959);
nor U17288 (N_17288,N_13470,N_12626);
nand U17289 (N_17289,N_11513,N_10791);
or U17290 (N_17290,N_12465,N_14104);
or U17291 (N_17291,N_14772,N_13112);
or U17292 (N_17292,N_10956,N_13992);
or U17293 (N_17293,N_10259,N_14336);
nor U17294 (N_17294,N_10801,N_11644);
and U17295 (N_17295,N_11010,N_14741);
xnor U17296 (N_17296,N_10583,N_14694);
nor U17297 (N_17297,N_14558,N_10910);
nor U17298 (N_17298,N_13948,N_14330);
xor U17299 (N_17299,N_12600,N_11687);
nand U17300 (N_17300,N_13098,N_12282);
and U17301 (N_17301,N_14404,N_14487);
nand U17302 (N_17302,N_13913,N_13115);
nor U17303 (N_17303,N_12441,N_10098);
nand U17304 (N_17304,N_13421,N_11639);
or U17305 (N_17305,N_11306,N_10511);
or U17306 (N_17306,N_13757,N_10742);
nand U17307 (N_17307,N_11795,N_13075);
or U17308 (N_17308,N_11127,N_11671);
nand U17309 (N_17309,N_10729,N_14410);
nand U17310 (N_17310,N_14279,N_10627);
and U17311 (N_17311,N_14495,N_12680);
and U17312 (N_17312,N_12992,N_13577);
and U17313 (N_17313,N_12205,N_12047);
nor U17314 (N_17314,N_13499,N_13510);
or U17315 (N_17315,N_14750,N_10095);
and U17316 (N_17316,N_12322,N_10739);
or U17317 (N_17317,N_13011,N_13602);
xnor U17318 (N_17318,N_13126,N_10056);
or U17319 (N_17319,N_12239,N_11379);
or U17320 (N_17320,N_12572,N_13509);
and U17321 (N_17321,N_11314,N_12121);
or U17322 (N_17322,N_11288,N_12049);
and U17323 (N_17323,N_14067,N_14286);
and U17324 (N_17324,N_11281,N_14572);
nand U17325 (N_17325,N_14888,N_11019);
nand U17326 (N_17326,N_13696,N_10357);
xor U17327 (N_17327,N_10908,N_11745);
or U17328 (N_17328,N_12474,N_12571);
nor U17329 (N_17329,N_12119,N_11075);
nor U17330 (N_17330,N_13950,N_12022);
nor U17331 (N_17331,N_10075,N_13742);
or U17332 (N_17332,N_14611,N_11662);
and U17333 (N_17333,N_10567,N_14047);
nand U17334 (N_17334,N_13836,N_13204);
and U17335 (N_17335,N_14705,N_12442);
or U17336 (N_17336,N_12962,N_14737);
and U17337 (N_17337,N_14039,N_11408);
or U17338 (N_17338,N_11076,N_11850);
and U17339 (N_17339,N_13569,N_10210);
nor U17340 (N_17340,N_10660,N_13777);
or U17341 (N_17341,N_11219,N_10614);
or U17342 (N_17342,N_13361,N_11096);
and U17343 (N_17343,N_11197,N_13701);
and U17344 (N_17344,N_11030,N_11371);
xor U17345 (N_17345,N_13552,N_12246);
nand U17346 (N_17346,N_13977,N_10132);
nand U17347 (N_17347,N_11409,N_12061);
nand U17348 (N_17348,N_12613,N_12986);
or U17349 (N_17349,N_14659,N_10800);
nor U17350 (N_17350,N_12020,N_12343);
or U17351 (N_17351,N_10130,N_11492);
nand U17352 (N_17352,N_13608,N_14362);
nor U17353 (N_17353,N_12106,N_13188);
or U17354 (N_17354,N_11871,N_12216);
and U17355 (N_17355,N_11610,N_14002);
nor U17356 (N_17356,N_13460,N_10699);
or U17357 (N_17357,N_12110,N_12161);
and U17358 (N_17358,N_11354,N_10402);
or U17359 (N_17359,N_12384,N_13013);
or U17360 (N_17360,N_12346,N_13152);
and U17361 (N_17361,N_11984,N_11957);
or U17362 (N_17362,N_10131,N_10045);
or U17363 (N_17363,N_12668,N_13692);
xor U17364 (N_17364,N_14080,N_12628);
and U17365 (N_17365,N_12150,N_12513);
xnor U17366 (N_17366,N_14801,N_12140);
nor U17367 (N_17367,N_10810,N_12874);
or U17368 (N_17368,N_12451,N_14600);
and U17369 (N_17369,N_12960,N_13767);
and U17370 (N_17370,N_12435,N_11164);
xor U17371 (N_17371,N_13208,N_10449);
nor U17372 (N_17372,N_14783,N_13563);
nor U17373 (N_17373,N_13426,N_14683);
nor U17374 (N_17374,N_10364,N_13616);
and U17375 (N_17375,N_10148,N_10006);
and U17376 (N_17376,N_10520,N_11063);
nor U17377 (N_17377,N_10779,N_12948);
nand U17378 (N_17378,N_14630,N_12028);
or U17379 (N_17379,N_12389,N_13166);
xor U17380 (N_17380,N_13017,N_11270);
xor U17381 (N_17381,N_11123,N_11797);
nor U17382 (N_17382,N_12157,N_11200);
nor U17383 (N_17383,N_14871,N_12681);
nor U17384 (N_17384,N_14597,N_12393);
or U17385 (N_17385,N_13820,N_12210);
and U17386 (N_17386,N_10986,N_12687);
or U17387 (N_17387,N_12928,N_14493);
or U17388 (N_17388,N_14817,N_10343);
xnor U17389 (N_17389,N_12595,N_14400);
xnor U17390 (N_17390,N_14365,N_12154);
and U17391 (N_17391,N_10207,N_11586);
and U17392 (N_17392,N_13543,N_11066);
nand U17393 (N_17393,N_13405,N_12846);
nor U17394 (N_17394,N_10333,N_11993);
and U17395 (N_17395,N_14984,N_13818);
nor U17396 (N_17396,N_12016,N_14910);
and U17397 (N_17397,N_12357,N_14176);
nand U17398 (N_17398,N_12788,N_13538);
xor U17399 (N_17399,N_11350,N_13683);
nand U17400 (N_17400,N_13819,N_13744);
and U17401 (N_17401,N_12344,N_10102);
or U17402 (N_17402,N_12734,N_13888);
nor U17403 (N_17403,N_11945,N_12170);
nand U17404 (N_17404,N_13555,N_12165);
or U17405 (N_17405,N_14921,N_12900);
or U17406 (N_17406,N_11345,N_14735);
nand U17407 (N_17407,N_12912,N_14606);
nor U17408 (N_17408,N_13695,N_12179);
nand U17409 (N_17409,N_10464,N_11235);
or U17410 (N_17410,N_10539,N_12475);
nand U17411 (N_17411,N_12954,N_13371);
and U17412 (N_17412,N_12328,N_10649);
nand U17413 (N_17413,N_13386,N_12718);
and U17414 (N_17414,N_13434,N_14395);
and U17415 (N_17415,N_11236,N_11210);
nand U17416 (N_17416,N_10458,N_12153);
nor U17417 (N_17417,N_10112,N_11375);
nand U17418 (N_17418,N_14904,N_10613);
xor U17419 (N_17419,N_12703,N_13176);
or U17420 (N_17420,N_14837,N_13952);
nand U17421 (N_17421,N_12265,N_13289);
or U17422 (N_17422,N_11099,N_13365);
and U17423 (N_17423,N_12039,N_10901);
nor U17424 (N_17424,N_11926,N_14009);
or U17425 (N_17425,N_10246,N_13068);
xnor U17426 (N_17426,N_14382,N_11519);
nor U17427 (N_17427,N_12041,N_12031);
or U17428 (N_17428,N_11933,N_10836);
nor U17429 (N_17429,N_11429,N_13624);
and U17430 (N_17430,N_13663,N_13290);
nand U17431 (N_17431,N_12483,N_11234);
and U17432 (N_17432,N_10070,N_11869);
or U17433 (N_17433,N_13953,N_12525);
and U17434 (N_17434,N_12067,N_13286);
nor U17435 (N_17435,N_11779,N_10553);
xor U17436 (N_17436,N_13923,N_10922);
or U17437 (N_17437,N_13830,N_14734);
nor U17438 (N_17438,N_13811,N_11814);
nand U17439 (N_17439,N_10732,N_11439);
nand U17440 (N_17440,N_14281,N_11874);
and U17441 (N_17441,N_13271,N_12741);
nand U17442 (N_17442,N_12853,N_13234);
nand U17443 (N_17443,N_10088,N_13970);
nor U17444 (N_17444,N_14075,N_12035);
xnor U17445 (N_17445,N_13488,N_10840);
and U17446 (N_17446,N_14764,N_13596);
nor U17447 (N_17447,N_14637,N_12194);
nand U17448 (N_17448,N_12700,N_12974);
nand U17449 (N_17449,N_11894,N_14014);
or U17450 (N_17450,N_13667,N_11997);
or U17451 (N_17451,N_11239,N_12789);
nor U17452 (N_17452,N_11807,N_12270);
and U17453 (N_17453,N_13339,N_12692);
and U17454 (N_17454,N_14086,N_11986);
and U17455 (N_17455,N_12762,N_12271);
xor U17456 (N_17456,N_10550,N_14573);
nand U17457 (N_17457,N_14332,N_13845);
and U17458 (N_17458,N_13917,N_13890);
xor U17459 (N_17459,N_11173,N_12511);
or U17460 (N_17460,N_13231,N_14432);
nor U17461 (N_17461,N_13734,N_10324);
nor U17462 (N_17462,N_10949,N_11260);
xnor U17463 (N_17463,N_13042,N_10391);
nand U17464 (N_17464,N_10776,N_11714);
and U17465 (N_17465,N_11655,N_11222);
or U17466 (N_17466,N_12169,N_12399);
or U17467 (N_17467,N_11442,N_11363);
nand U17468 (N_17468,N_11999,N_12837);
or U17469 (N_17469,N_13931,N_14042);
and U17470 (N_17470,N_12548,N_10850);
nor U17471 (N_17471,N_12546,N_13921);
or U17472 (N_17472,N_12042,N_13648);
or U17473 (N_17473,N_14019,N_13026);
nand U17474 (N_17474,N_14749,N_12878);
nand U17475 (N_17475,N_10499,N_10341);
and U17476 (N_17476,N_13795,N_10233);
xor U17477 (N_17477,N_14515,N_12582);
xnor U17478 (N_17478,N_13014,N_12459);
or U17479 (N_17479,N_12534,N_10181);
or U17480 (N_17480,N_12972,N_11500);
and U17481 (N_17481,N_11397,N_14094);
nor U17482 (N_17482,N_11801,N_11650);
nand U17483 (N_17483,N_11879,N_13841);
xnor U17484 (N_17484,N_12496,N_13363);
and U17485 (N_17485,N_11664,N_11956);
and U17486 (N_17486,N_11756,N_12286);
xnor U17487 (N_17487,N_11567,N_11646);
and U17488 (N_17488,N_10125,N_10293);
and U17489 (N_17489,N_14617,N_14599);
nand U17490 (N_17490,N_13547,N_12653);
or U17491 (N_17491,N_10983,N_10903);
or U17492 (N_17492,N_13827,N_14144);
or U17493 (N_17493,N_11494,N_13028);
and U17494 (N_17494,N_13137,N_13874);
nand U17495 (N_17495,N_12722,N_14507);
nor U17496 (N_17496,N_10188,N_12793);
and U17497 (N_17497,N_12895,N_11765);
nand U17498 (N_17498,N_14909,N_11116);
nor U17499 (N_17499,N_11441,N_10042);
nand U17500 (N_17500,N_14360,N_12772);
or U17501 (N_17501,N_14151,N_13730);
nor U17502 (N_17502,N_11602,N_12880);
nor U17503 (N_17503,N_11391,N_11243);
xnor U17504 (N_17504,N_14618,N_14816);
nand U17505 (N_17505,N_10674,N_13397);
and U17506 (N_17506,N_10926,N_12002);
nor U17507 (N_17507,N_10611,N_12415);
and U17508 (N_17508,N_11820,N_13270);
or U17509 (N_17509,N_14588,N_13142);
and U17510 (N_17510,N_10752,N_13648);
or U17511 (N_17511,N_13479,N_13882);
or U17512 (N_17512,N_10026,N_13472);
nand U17513 (N_17513,N_13800,N_12582);
nand U17514 (N_17514,N_14212,N_14605);
nand U17515 (N_17515,N_11406,N_12137);
or U17516 (N_17516,N_14604,N_11949);
nand U17517 (N_17517,N_12690,N_12109);
or U17518 (N_17518,N_14793,N_14769);
and U17519 (N_17519,N_11132,N_12466);
nor U17520 (N_17520,N_10295,N_11893);
and U17521 (N_17521,N_12972,N_10523);
nor U17522 (N_17522,N_11293,N_11009);
nor U17523 (N_17523,N_14590,N_10357);
or U17524 (N_17524,N_10801,N_14993);
or U17525 (N_17525,N_13222,N_10657);
nor U17526 (N_17526,N_10850,N_12822);
or U17527 (N_17527,N_14146,N_10289);
or U17528 (N_17528,N_10879,N_14434);
nor U17529 (N_17529,N_11470,N_14201);
nor U17530 (N_17530,N_12388,N_13083);
nor U17531 (N_17531,N_10973,N_13418);
nand U17532 (N_17532,N_14457,N_11634);
nand U17533 (N_17533,N_14934,N_14541);
nand U17534 (N_17534,N_12906,N_11560);
nand U17535 (N_17535,N_11106,N_13557);
nand U17536 (N_17536,N_13080,N_10525);
nand U17537 (N_17537,N_13651,N_13541);
and U17538 (N_17538,N_14910,N_11292);
or U17539 (N_17539,N_14389,N_11128);
or U17540 (N_17540,N_14657,N_10674);
xor U17541 (N_17541,N_14141,N_13505);
and U17542 (N_17542,N_13571,N_14531);
and U17543 (N_17543,N_14744,N_13686);
xnor U17544 (N_17544,N_14570,N_11220);
nand U17545 (N_17545,N_13419,N_12620);
or U17546 (N_17546,N_14940,N_10967);
nor U17547 (N_17547,N_12153,N_12470);
nor U17548 (N_17548,N_14906,N_13782);
or U17549 (N_17549,N_12031,N_14832);
nor U17550 (N_17550,N_13260,N_12776);
and U17551 (N_17551,N_13619,N_13337);
nor U17552 (N_17552,N_11772,N_10768);
nand U17553 (N_17553,N_12523,N_12197);
and U17554 (N_17554,N_12292,N_11968);
xor U17555 (N_17555,N_11285,N_12744);
nand U17556 (N_17556,N_13194,N_10878);
nand U17557 (N_17557,N_10122,N_13225);
nor U17558 (N_17558,N_13567,N_12865);
and U17559 (N_17559,N_11145,N_10209);
and U17560 (N_17560,N_14092,N_14113);
nor U17561 (N_17561,N_10431,N_12344);
nand U17562 (N_17562,N_13585,N_10591);
xor U17563 (N_17563,N_13115,N_13506);
and U17564 (N_17564,N_10719,N_12129);
nand U17565 (N_17565,N_12185,N_10258);
or U17566 (N_17566,N_10281,N_11897);
and U17567 (N_17567,N_10997,N_13586);
nor U17568 (N_17568,N_14259,N_12665);
nand U17569 (N_17569,N_11780,N_13941);
xor U17570 (N_17570,N_13986,N_13709);
or U17571 (N_17571,N_12356,N_11327);
or U17572 (N_17572,N_13585,N_12831);
or U17573 (N_17573,N_13354,N_12101);
nand U17574 (N_17574,N_14244,N_10453);
or U17575 (N_17575,N_10937,N_13291);
nor U17576 (N_17576,N_14644,N_14035);
nand U17577 (N_17577,N_11264,N_13823);
nand U17578 (N_17578,N_13478,N_14996);
nor U17579 (N_17579,N_11000,N_10035);
nand U17580 (N_17580,N_13350,N_11293);
nand U17581 (N_17581,N_14869,N_10637);
nor U17582 (N_17582,N_10484,N_10436);
or U17583 (N_17583,N_14212,N_12478);
or U17584 (N_17584,N_11337,N_14748);
and U17585 (N_17585,N_12706,N_11291);
xor U17586 (N_17586,N_10712,N_13752);
and U17587 (N_17587,N_11475,N_13035);
nor U17588 (N_17588,N_13945,N_11099);
or U17589 (N_17589,N_10264,N_13802);
or U17590 (N_17590,N_14209,N_14416);
xor U17591 (N_17591,N_12335,N_13999);
nand U17592 (N_17592,N_14667,N_12864);
and U17593 (N_17593,N_10578,N_11400);
nor U17594 (N_17594,N_10652,N_12993);
and U17595 (N_17595,N_13862,N_10283);
nand U17596 (N_17596,N_14383,N_10778);
and U17597 (N_17597,N_11595,N_12052);
or U17598 (N_17598,N_12711,N_14484);
nand U17599 (N_17599,N_11034,N_12461);
or U17600 (N_17600,N_12985,N_12213);
or U17601 (N_17601,N_10931,N_11179);
nor U17602 (N_17602,N_11785,N_12282);
nor U17603 (N_17603,N_13078,N_12131);
nand U17604 (N_17604,N_11541,N_12301);
or U17605 (N_17605,N_14318,N_12130);
or U17606 (N_17606,N_13941,N_14103);
and U17607 (N_17607,N_12866,N_10518);
nand U17608 (N_17608,N_12818,N_11723);
nor U17609 (N_17609,N_11583,N_13993);
xor U17610 (N_17610,N_13902,N_12436);
nor U17611 (N_17611,N_13338,N_14283);
nand U17612 (N_17612,N_12551,N_11549);
or U17613 (N_17613,N_13729,N_13266);
nor U17614 (N_17614,N_11413,N_10464);
and U17615 (N_17615,N_14479,N_13910);
or U17616 (N_17616,N_10889,N_14861);
nand U17617 (N_17617,N_12730,N_13425);
or U17618 (N_17618,N_12686,N_11420);
and U17619 (N_17619,N_13297,N_12752);
nor U17620 (N_17620,N_13818,N_11487);
or U17621 (N_17621,N_13217,N_14552);
and U17622 (N_17622,N_12625,N_13864);
nor U17623 (N_17623,N_10849,N_14693);
and U17624 (N_17624,N_11254,N_12720);
nor U17625 (N_17625,N_14085,N_12214);
or U17626 (N_17626,N_14174,N_13126);
nor U17627 (N_17627,N_10066,N_12467);
nor U17628 (N_17628,N_11142,N_14017);
or U17629 (N_17629,N_12511,N_10302);
or U17630 (N_17630,N_11377,N_10631);
nand U17631 (N_17631,N_14973,N_11986);
nand U17632 (N_17632,N_12696,N_11126);
nand U17633 (N_17633,N_13251,N_12994);
or U17634 (N_17634,N_13502,N_10780);
xnor U17635 (N_17635,N_12479,N_12791);
nor U17636 (N_17636,N_14217,N_11198);
or U17637 (N_17637,N_12510,N_13595);
or U17638 (N_17638,N_12512,N_13588);
nor U17639 (N_17639,N_10496,N_11899);
xnor U17640 (N_17640,N_11331,N_10188);
and U17641 (N_17641,N_12081,N_14688);
or U17642 (N_17642,N_13464,N_10531);
nand U17643 (N_17643,N_14596,N_14403);
or U17644 (N_17644,N_14398,N_14152);
or U17645 (N_17645,N_11173,N_12117);
nor U17646 (N_17646,N_14548,N_13775);
nor U17647 (N_17647,N_14597,N_13546);
and U17648 (N_17648,N_12999,N_13514);
or U17649 (N_17649,N_11707,N_12229);
and U17650 (N_17650,N_13397,N_11883);
nor U17651 (N_17651,N_13095,N_14315);
nand U17652 (N_17652,N_12657,N_13869);
nand U17653 (N_17653,N_11321,N_12528);
and U17654 (N_17654,N_10837,N_10962);
nor U17655 (N_17655,N_12282,N_12461);
or U17656 (N_17656,N_12456,N_14328);
nor U17657 (N_17657,N_11138,N_11701);
and U17658 (N_17658,N_11723,N_11930);
nor U17659 (N_17659,N_13201,N_10002);
and U17660 (N_17660,N_14444,N_14278);
and U17661 (N_17661,N_13159,N_10493);
or U17662 (N_17662,N_14884,N_10004);
and U17663 (N_17663,N_13989,N_13716);
xnor U17664 (N_17664,N_13962,N_14209);
nor U17665 (N_17665,N_10930,N_10462);
nor U17666 (N_17666,N_12577,N_12165);
nor U17667 (N_17667,N_10342,N_10416);
xnor U17668 (N_17668,N_13554,N_14563);
and U17669 (N_17669,N_12473,N_14302);
nand U17670 (N_17670,N_13280,N_14842);
and U17671 (N_17671,N_10474,N_10165);
nor U17672 (N_17672,N_11572,N_13121);
nor U17673 (N_17673,N_12382,N_14737);
nand U17674 (N_17674,N_10142,N_12835);
nor U17675 (N_17675,N_13678,N_14029);
nor U17676 (N_17676,N_13255,N_11125);
nor U17677 (N_17677,N_12520,N_13804);
nor U17678 (N_17678,N_10600,N_11942);
nand U17679 (N_17679,N_10047,N_12083);
or U17680 (N_17680,N_13534,N_11408);
and U17681 (N_17681,N_10957,N_10027);
and U17682 (N_17682,N_12664,N_13572);
nor U17683 (N_17683,N_13667,N_14344);
nand U17684 (N_17684,N_14933,N_14520);
and U17685 (N_17685,N_14360,N_13797);
nor U17686 (N_17686,N_14927,N_12729);
and U17687 (N_17687,N_12238,N_10506);
nand U17688 (N_17688,N_12214,N_14697);
nand U17689 (N_17689,N_11895,N_14714);
xor U17690 (N_17690,N_13391,N_14586);
nor U17691 (N_17691,N_12551,N_13016);
and U17692 (N_17692,N_11003,N_14607);
nand U17693 (N_17693,N_13395,N_13844);
xnor U17694 (N_17694,N_14086,N_11916);
nor U17695 (N_17695,N_13746,N_12655);
or U17696 (N_17696,N_11402,N_14751);
xor U17697 (N_17697,N_13676,N_10832);
and U17698 (N_17698,N_13677,N_10417);
and U17699 (N_17699,N_11690,N_14103);
nand U17700 (N_17700,N_11623,N_11108);
and U17701 (N_17701,N_10341,N_11442);
nand U17702 (N_17702,N_14462,N_14948);
nand U17703 (N_17703,N_14487,N_13852);
or U17704 (N_17704,N_13753,N_11846);
nand U17705 (N_17705,N_13574,N_14304);
nand U17706 (N_17706,N_14055,N_12588);
nor U17707 (N_17707,N_13177,N_11951);
nand U17708 (N_17708,N_14279,N_11172);
xor U17709 (N_17709,N_10511,N_13389);
nor U17710 (N_17710,N_11434,N_14026);
or U17711 (N_17711,N_10984,N_11008);
or U17712 (N_17712,N_14819,N_11346);
and U17713 (N_17713,N_12617,N_12080);
nor U17714 (N_17714,N_12228,N_12827);
nand U17715 (N_17715,N_13534,N_13511);
or U17716 (N_17716,N_10373,N_14419);
and U17717 (N_17717,N_11237,N_11474);
nor U17718 (N_17718,N_14765,N_13492);
nor U17719 (N_17719,N_14707,N_11483);
nand U17720 (N_17720,N_10611,N_13923);
and U17721 (N_17721,N_10238,N_11435);
xnor U17722 (N_17722,N_14925,N_13585);
nor U17723 (N_17723,N_11871,N_12517);
or U17724 (N_17724,N_10725,N_11111);
or U17725 (N_17725,N_12696,N_11893);
and U17726 (N_17726,N_13161,N_14231);
nand U17727 (N_17727,N_12242,N_12780);
and U17728 (N_17728,N_13354,N_13359);
and U17729 (N_17729,N_13612,N_11085);
or U17730 (N_17730,N_14946,N_11564);
or U17731 (N_17731,N_14615,N_13988);
xnor U17732 (N_17732,N_14399,N_14487);
and U17733 (N_17733,N_10928,N_13587);
xnor U17734 (N_17734,N_14981,N_12784);
nor U17735 (N_17735,N_10119,N_12406);
or U17736 (N_17736,N_12516,N_11897);
nor U17737 (N_17737,N_13621,N_10634);
or U17738 (N_17738,N_12700,N_11063);
or U17739 (N_17739,N_12325,N_13160);
nand U17740 (N_17740,N_12966,N_11172);
and U17741 (N_17741,N_12395,N_10305);
or U17742 (N_17742,N_14748,N_12621);
xor U17743 (N_17743,N_12330,N_12732);
nor U17744 (N_17744,N_12588,N_10640);
nor U17745 (N_17745,N_13733,N_11961);
and U17746 (N_17746,N_13276,N_11578);
or U17747 (N_17747,N_11969,N_12903);
or U17748 (N_17748,N_12589,N_12369);
xor U17749 (N_17749,N_11942,N_12919);
nand U17750 (N_17750,N_13823,N_12548);
xor U17751 (N_17751,N_11476,N_11511);
nor U17752 (N_17752,N_11962,N_11343);
or U17753 (N_17753,N_11018,N_10331);
and U17754 (N_17754,N_11797,N_13032);
or U17755 (N_17755,N_11675,N_11031);
nor U17756 (N_17756,N_12172,N_11888);
nand U17757 (N_17757,N_14477,N_13563);
or U17758 (N_17758,N_11992,N_14215);
nand U17759 (N_17759,N_14843,N_11600);
or U17760 (N_17760,N_11676,N_13557);
or U17761 (N_17761,N_12410,N_14210);
or U17762 (N_17762,N_10516,N_10042);
or U17763 (N_17763,N_13198,N_10858);
or U17764 (N_17764,N_10333,N_12891);
nand U17765 (N_17765,N_10799,N_11085);
nand U17766 (N_17766,N_11139,N_13255);
or U17767 (N_17767,N_11603,N_13193);
nor U17768 (N_17768,N_14631,N_14237);
nand U17769 (N_17769,N_12711,N_10318);
and U17770 (N_17770,N_10121,N_10533);
nor U17771 (N_17771,N_14608,N_14612);
or U17772 (N_17772,N_14681,N_12064);
and U17773 (N_17773,N_14109,N_10411);
or U17774 (N_17774,N_11597,N_13997);
or U17775 (N_17775,N_10113,N_13323);
and U17776 (N_17776,N_12789,N_12324);
nor U17777 (N_17777,N_10527,N_10494);
or U17778 (N_17778,N_10402,N_13177);
xnor U17779 (N_17779,N_12910,N_10261);
nor U17780 (N_17780,N_10606,N_13751);
and U17781 (N_17781,N_14894,N_13736);
nor U17782 (N_17782,N_14404,N_13391);
or U17783 (N_17783,N_13535,N_13667);
or U17784 (N_17784,N_13369,N_13221);
nand U17785 (N_17785,N_12492,N_11347);
nand U17786 (N_17786,N_11017,N_10269);
and U17787 (N_17787,N_14875,N_10079);
nand U17788 (N_17788,N_10025,N_14433);
xnor U17789 (N_17789,N_10244,N_12182);
xnor U17790 (N_17790,N_12959,N_14050);
or U17791 (N_17791,N_11928,N_13293);
nor U17792 (N_17792,N_13853,N_10977);
or U17793 (N_17793,N_12179,N_10726);
nand U17794 (N_17794,N_10669,N_12591);
xor U17795 (N_17795,N_11954,N_12966);
and U17796 (N_17796,N_10700,N_12511);
and U17797 (N_17797,N_12239,N_13071);
nand U17798 (N_17798,N_12768,N_13392);
nor U17799 (N_17799,N_12237,N_11211);
or U17800 (N_17800,N_10587,N_14906);
or U17801 (N_17801,N_10221,N_14208);
nand U17802 (N_17802,N_11761,N_11768);
nand U17803 (N_17803,N_12376,N_13467);
nand U17804 (N_17804,N_14771,N_10722);
nor U17805 (N_17805,N_12387,N_12180);
and U17806 (N_17806,N_12241,N_13484);
nor U17807 (N_17807,N_12590,N_13979);
nand U17808 (N_17808,N_13101,N_11915);
nand U17809 (N_17809,N_10502,N_14855);
xor U17810 (N_17810,N_14836,N_13638);
nand U17811 (N_17811,N_12992,N_10766);
or U17812 (N_17812,N_13132,N_12443);
or U17813 (N_17813,N_13368,N_11694);
and U17814 (N_17814,N_11774,N_11336);
nor U17815 (N_17815,N_10628,N_12000);
nor U17816 (N_17816,N_13778,N_12807);
and U17817 (N_17817,N_12039,N_12422);
or U17818 (N_17818,N_13178,N_14426);
nand U17819 (N_17819,N_13138,N_10085);
nand U17820 (N_17820,N_13153,N_14624);
and U17821 (N_17821,N_11003,N_10527);
nor U17822 (N_17822,N_12795,N_13252);
nor U17823 (N_17823,N_10985,N_10337);
and U17824 (N_17824,N_12704,N_12739);
nor U17825 (N_17825,N_13049,N_13702);
nand U17826 (N_17826,N_12489,N_11365);
or U17827 (N_17827,N_11820,N_10521);
nor U17828 (N_17828,N_10387,N_11879);
and U17829 (N_17829,N_11888,N_14015);
xor U17830 (N_17830,N_12720,N_12205);
or U17831 (N_17831,N_10370,N_10929);
nand U17832 (N_17832,N_11512,N_10514);
nor U17833 (N_17833,N_12654,N_11754);
xor U17834 (N_17834,N_14771,N_12971);
and U17835 (N_17835,N_13144,N_12525);
or U17836 (N_17836,N_10201,N_13950);
nor U17837 (N_17837,N_12258,N_13472);
nand U17838 (N_17838,N_10656,N_11900);
nor U17839 (N_17839,N_13749,N_10002);
and U17840 (N_17840,N_10137,N_10891);
nand U17841 (N_17841,N_12385,N_14489);
and U17842 (N_17842,N_10115,N_14530);
and U17843 (N_17843,N_11668,N_10353);
and U17844 (N_17844,N_12098,N_11334);
and U17845 (N_17845,N_13268,N_13874);
or U17846 (N_17846,N_11052,N_13135);
nor U17847 (N_17847,N_13694,N_13418);
xor U17848 (N_17848,N_10423,N_10315);
nor U17849 (N_17849,N_12768,N_14254);
and U17850 (N_17850,N_13267,N_12084);
or U17851 (N_17851,N_11535,N_14972);
and U17852 (N_17852,N_10294,N_13228);
or U17853 (N_17853,N_11651,N_13599);
or U17854 (N_17854,N_10640,N_11220);
or U17855 (N_17855,N_11757,N_10087);
nor U17856 (N_17856,N_13696,N_12834);
or U17857 (N_17857,N_13694,N_13770);
and U17858 (N_17858,N_11895,N_12040);
or U17859 (N_17859,N_10941,N_13537);
and U17860 (N_17860,N_13867,N_11229);
nor U17861 (N_17861,N_12712,N_10399);
and U17862 (N_17862,N_11385,N_10238);
and U17863 (N_17863,N_13004,N_12468);
and U17864 (N_17864,N_13615,N_13632);
nor U17865 (N_17865,N_12670,N_12600);
or U17866 (N_17866,N_12749,N_14540);
nor U17867 (N_17867,N_14396,N_12492);
nand U17868 (N_17868,N_11275,N_12677);
nor U17869 (N_17869,N_10673,N_13815);
and U17870 (N_17870,N_14296,N_10164);
nor U17871 (N_17871,N_12597,N_13843);
and U17872 (N_17872,N_14624,N_10011);
nor U17873 (N_17873,N_14228,N_11006);
nand U17874 (N_17874,N_14814,N_13428);
nor U17875 (N_17875,N_13273,N_10811);
nor U17876 (N_17876,N_14419,N_14851);
nor U17877 (N_17877,N_10455,N_10863);
and U17878 (N_17878,N_14331,N_10598);
nand U17879 (N_17879,N_14534,N_10632);
and U17880 (N_17880,N_13242,N_12175);
nor U17881 (N_17881,N_10434,N_12129);
nor U17882 (N_17882,N_10983,N_13030);
nor U17883 (N_17883,N_13232,N_11428);
and U17884 (N_17884,N_13058,N_11409);
or U17885 (N_17885,N_12682,N_14245);
and U17886 (N_17886,N_11266,N_13151);
xor U17887 (N_17887,N_12938,N_11371);
and U17888 (N_17888,N_10427,N_11718);
nand U17889 (N_17889,N_12824,N_12223);
nand U17890 (N_17890,N_10087,N_10923);
nand U17891 (N_17891,N_12208,N_12787);
nand U17892 (N_17892,N_12223,N_10298);
nor U17893 (N_17893,N_13540,N_10840);
and U17894 (N_17894,N_11467,N_12350);
and U17895 (N_17895,N_13120,N_11281);
nor U17896 (N_17896,N_14281,N_13690);
nor U17897 (N_17897,N_10096,N_13894);
and U17898 (N_17898,N_13526,N_14578);
and U17899 (N_17899,N_10375,N_14990);
and U17900 (N_17900,N_10461,N_12011);
nand U17901 (N_17901,N_11397,N_10365);
and U17902 (N_17902,N_11826,N_11978);
nand U17903 (N_17903,N_13047,N_14841);
nand U17904 (N_17904,N_11101,N_13007);
xnor U17905 (N_17905,N_10906,N_11509);
nor U17906 (N_17906,N_10671,N_13736);
and U17907 (N_17907,N_13926,N_13399);
or U17908 (N_17908,N_12282,N_14884);
or U17909 (N_17909,N_10814,N_12928);
nor U17910 (N_17910,N_13094,N_11940);
and U17911 (N_17911,N_12340,N_14658);
nand U17912 (N_17912,N_11477,N_11382);
nand U17913 (N_17913,N_10767,N_11697);
nand U17914 (N_17914,N_12988,N_14028);
nand U17915 (N_17915,N_12837,N_14502);
or U17916 (N_17916,N_10014,N_14661);
nor U17917 (N_17917,N_10511,N_13385);
and U17918 (N_17918,N_13033,N_10362);
or U17919 (N_17919,N_10655,N_14172);
nor U17920 (N_17920,N_14295,N_13288);
or U17921 (N_17921,N_10622,N_10894);
nand U17922 (N_17922,N_12639,N_10157);
nor U17923 (N_17923,N_10501,N_12955);
or U17924 (N_17924,N_13934,N_12601);
and U17925 (N_17925,N_11149,N_10492);
or U17926 (N_17926,N_11745,N_12497);
nand U17927 (N_17927,N_11724,N_11221);
nand U17928 (N_17928,N_10446,N_12309);
nand U17929 (N_17929,N_14326,N_14976);
and U17930 (N_17930,N_11226,N_14396);
nand U17931 (N_17931,N_10193,N_12397);
or U17932 (N_17932,N_11653,N_10305);
and U17933 (N_17933,N_10067,N_10806);
or U17934 (N_17934,N_14818,N_11129);
and U17935 (N_17935,N_13289,N_11943);
or U17936 (N_17936,N_14180,N_10019);
nand U17937 (N_17937,N_13408,N_10875);
nor U17938 (N_17938,N_10532,N_11483);
nor U17939 (N_17939,N_11686,N_10566);
and U17940 (N_17940,N_13864,N_14131);
nand U17941 (N_17941,N_13206,N_14980);
xor U17942 (N_17942,N_11525,N_13727);
nor U17943 (N_17943,N_12077,N_11480);
xnor U17944 (N_17944,N_11306,N_11580);
nand U17945 (N_17945,N_11077,N_12530);
and U17946 (N_17946,N_14161,N_11633);
and U17947 (N_17947,N_12413,N_11025);
nand U17948 (N_17948,N_11450,N_11264);
or U17949 (N_17949,N_13584,N_10519);
and U17950 (N_17950,N_10898,N_12410);
or U17951 (N_17951,N_14395,N_12711);
or U17952 (N_17952,N_12393,N_11479);
nand U17953 (N_17953,N_13674,N_11925);
nor U17954 (N_17954,N_12046,N_10320);
and U17955 (N_17955,N_10785,N_14991);
xor U17956 (N_17956,N_11063,N_12050);
or U17957 (N_17957,N_11104,N_14913);
or U17958 (N_17958,N_13034,N_12581);
xnor U17959 (N_17959,N_11411,N_12578);
xnor U17960 (N_17960,N_10650,N_11196);
nand U17961 (N_17961,N_12371,N_10334);
or U17962 (N_17962,N_10985,N_10465);
xnor U17963 (N_17963,N_14879,N_10866);
nor U17964 (N_17964,N_11408,N_10373);
and U17965 (N_17965,N_11966,N_13403);
nor U17966 (N_17966,N_11281,N_12584);
or U17967 (N_17967,N_11869,N_11155);
and U17968 (N_17968,N_14416,N_14750);
or U17969 (N_17969,N_13260,N_12692);
nand U17970 (N_17970,N_13824,N_14463);
nor U17971 (N_17971,N_11363,N_10650);
and U17972 (N_17972,N_12871,N_14509);
nor U17973 (N_17973,N_10049,N_13453);
nor U17974 (N_17974,N_10640,N_12771);
nor U17975 (N_17975,N_10438,N_10939);
and U17976 (N_17976,N_13004,N_14747);
nor U17977 (N_17977,N_13257,N_12188);
nor U17978 (N_17978,N_11817,N_13910);
nor U17979 (N_17979,N_11857,N_14077);
and U17980 (N_17980,N_10361,N_11340);
and U17981 (N_17981,N_10115,N_10748);
and U17982 (N_17982,N_13928,N_13710);
nand U17983 (N_17983,N_14944,N_14258);
or U17984 (N_17984,N_14837,N_14730);
or U17985 (N_17985,N_13980,N_10163);
xor U17986 (N_17986,N_14885,N_13972);
or U17987 (N_17987,N_10683,N_12671);
nand U17988 (N_17988,N_13007,N_14583);
nor U17989 (N_17989,N_14312,N_13467);
and U17990 (N_17990,N_11033,N_14406);
nor U17991 (N_17991,N_14002,N_10036);
or U17992 (N_17992,N_10665,N_13482);
and U17993 (N_17993,N_14618,N_13094);
or U17994 (N_17994,N_12750,N_14730);
nand U17995 (N_17995,N_14152,N_10769);
and U17996 (N_17996,N_14625,N_12423);
nor U17997 (N_17997,N_10376,N_14142);
xor U17998 (N_17998,N_13106,N_14978);
nor U17999 (N_17999,N_10858,N_11557);
nor U18000 (N_18000,N_11847,N_13572);
or U18001 (N_18001,N_11890,N_12186);
and U18002 (N_18002,N_11020,N_11739);
nand U18003 (N_18003,N_11628,N_13083);
nor U18004 (N_18004,N_11380,N_14352);
nand U18005 (N_18005,N_12191,N_13066);
and U18006 (N_18006,N_10814,N_11349);
or U18007 (N_18007,N_10603,N_13231);
nor U18008 (N_18008,N_12478,N_10824);
or U18009 (N_18009,N_10314,N_12686);
nand U18010 (N_18010,N_12168,N_11068);
or U18011 (N_18011,N_11299,N_10549);
xor U18012 (N_18012,N_10984,N_12206);
nor U18013 (N_18013,N_12395,N_10659);
nand U18014 (N_18014,N_14917,N_13004);
and U18015 (N_18015,N_14792,N_11146);
nand U18016 (N_18016,N_13877,N_14316);
xnor U18017 (N_18017,N_14530,N_11550);
and U18018 (N_18018,N_13968,N_10475);
nand U18019 (N_18019,N_14845,N_13600);
nor U18020 (N_18020,N_14510,N_12277);
nor U18021 (N_18021,N_12202,N_14609);
and U18022 (N_18022,N_12658,N_12043);
and U18023 (N_18023,N_13666,N_14179);
and U18024 (N_18024,N_10169,N_10797);
nand U18025 (N_18025,N_14571,N_10770);
nor U18026 (N_18026,N_10315,N_12356);
nand U18027 (N_18027,N_11396,N_14828);
nand U18028 (N_18028,N_11446,N_13989);
nand U18029 (N_18029,N_11565,N_12375);
or U18030 (N_18030,N_11922,N_10438);
and U18031 (N_18031,N_13147,N_12591);
nand U18032 (N_18032,N_14053,N_10636);
xnor U18033 (N_18033,N_10679,N_14130);
xor U18034 (N_18034,N_10133,N_13977);
or U18035 (N_18035,N_10418,N_11414);
and U18036 (N_18036,N_11981,N_14604);
or U18037 (N_18037,N_14634,N_13615);
or U18038 (N_18038,N_14132,N_13987);
and U18039 (N_18039,N_13929,N_14336);
and U18040 (N_18040,N_13806,N_10215);
xor U18041 (N_18041,N_10447,N_12236);
and U18042 (N_18042,N_12689,N_10473);
or U18043 (N_18043,N_14941,N_12283);
or U18044 (N_18044,N_13953,N_10217);
and U18045 (N_18045,N_10848,N_14715);
or U18046 (N_18046,N_11097,N_11307);
and U18047 (N_18047,N_14688,N_12245);
xor U18048 (N_18048,N_10668,N_14624);
nor U18049 (N_18049,N_10448,N_13930);
nand U18050 (N_18050,N_11139,N_11652);
nor U18051 (N_18051,N_13064,N_10370);
or U18052 (N_18052,N_10534,N_12510);
or U18053 (N_18053,N_13556,N_13852);
nand U18054 (N_18054,N_10790,N_12553);
xnor U18055 (N_18055,N_10418,N_12878);
or U18056 (N_18056,N_11886,N_14402);
nand U18057 (N_18057,N_12770,N_11807);
nand U18058 (N_18058,N_10883,N_14985);
and U18059 (N_18059,N_13719,N_10404);
or U18060 (N_18060,N_12005,N_12491);
and U18061 (N_18061,N_13242,N_12730);
nand U18062 (N_18062,N_11492,N_11949);
nand U18063 (N_18063,N_12258,N_10719);
nor U18064 (N_18064,N_11406,N_14014);
nand U18065 (N_18065,N_10768,N_12042);
xnor U18066 (N_18066,N_11058,N_14101);
nor U18067 (N_18067,N_14576,N_10897);
nand U18068 (N_18068,N_13859,N_11295);
xnor U18069 (N_18069,N_12049,N_13395);
nor U18070 (N_18070,N_11297,N_11421);
nor U18071 (N_18071,N_14722,N_10710);
or U18072 (N_18072,N_13456,N_13001);
nand U18073 (N_18073,N_13980,N_14088);
and U18074 (N_18074,N_12304,N_11347);
nand U18075 (N_18075,N_14195,N_14755);
and U18076 (N_18076,N_14932,N_13123);
or U18077 (N_18077,N_11424,N_11022);
and U18078 (N_18078,N_10807,N_13046);
nand U18079 (N_18079,N_11631,N_13409);
and U18080 (N_18080,N_11404,N_10344);
nand U18081 (N_18081,N_12058,N_13225);
or U18082 (N_18082,N_13726,N_11897);
and U18083 (N_18083,N_13517,N_12700);
or U18084 (N_18084,N_12388,N_13133);
and U18085 (N_18085,N_14916,N_10834);
nor U18086 (N_18086,N_14130,N_13249);
xor U18087 (N_18087,N_10571,N_11236);
and U18088 (N_18088,N_12869,N_13251);
nor U18089 (N_18089,N_12144,N_11977);
and U18090 (N_18090,N_12763,N_11600);
xnor U18091 (N_18091,N_11864,N_11977);
nor U18092 (N_18092,N_12995,N_14595);
nand U18093 (N_18093,N_11856,N_12711);
and U18094 (N_18094,N_14327,N_10939);
and U18095 (N_18095,N_13178,N_12295);
nor U18096 (N_18096,N_13672,N_11815);
nor U18097 (N_18097,N_13708,N_14380);
and U18098 (N_18098,N_11483,N_13619);
nand U18099 (N_18099,N_11160,N_11445);
nand U18100 (N_18100,N_12940,N_13986);
and U18101 (N_18101,N_10757,N_12529);
and U18102 (N_18102,N_13888,N_11180);
xnor U18103 (N_18103,N_10704,N_11097);
or U18104 (N_18104,N_14577,N_13329);
nand U18105 (N_18105,N_12129,N_13913);
and U18106 (N_18106,N_12007,N_10251);
nand U18107 (N_18107,N_10713,N_14440);
nor U18108 (N_18108,N_11367,N_11832);
nor U18109 (N_18109,N_12712,N_12571);
or U18110 (N_18110,N_14264,N_12523);
nor U18111 (N_18111,N_11695,N_11654);
xnor U18112 (N_18112,N_10413,N_13729);
nand U18113 (N_18113,N_12346,N_13438);
and U18114 (N_18114,N_10337,N_13038);
nand U18115 (N_18115,N_12171,N_13871);
nand U18116 (N_18116,N_10426,N_10475);
xnor U18117 (N_18117,N_11557,N_13127);
or U18118 (N_18118,N_10878,N_14722);
nand U18119 (N_18119,N_13585,N_12101);
and U18120 (N_18120,N_14637,N_12303);
or U18121 (N_18121,N_10329,N_14776);
and U18122 (N_18122,N_13994,N_14160);
nor U18123 (N_18123,N_12389,N_10420);
or U18124 (N_18124,N_12670,N_14665);
nor U18125 (N_18125,N_12206,N_10497);
nand U18126 (N_18126,N_11264,N_14374);
nand U18127 (N_18127,N_12864,N_13074);
or U18128 (N_18128,N_14808,N_12224);
or U18129 (N_18129,N_11333,N_12417);
nor U18130 (N_18130,N_10722,N_14679);
nor U18131 (N_18131,N_11088,N_12933);
nor U18132 (N_18132,N_11538,N_10520);
and U18133 (N_18133,N_10178,N_13136);
nand U18134 (N_18134,N_14239,N_13281);
and U18135 (N_18135,N_14355,N_11552);
or U18136 (N_18136,N_14564,N_13164);
nand U18137 (N_18137,N_13659,N_10885);
or U18138 (N_18138,N_10155,N_12059);
xnor U18139 (N_18139,N_14934,N_12959);
nor U18140 (N_18140,N_10762,N_14926);
and U18141 (N_18141,N_10080,N_11165);
xnor U18142 (N_18142,N_10922,N_11324);
or U18143 (N_18143,N_13779,N_13786);
nor U18144 (N_18144,N_13450,N_10590);
and U18145 (N_18145,N_12703,N_12965);
and U18146 (N_18146,N_13268,N_10535);
nand U18147 (N_18147,N_12585,N_14474);
or U18148 (N_18148,N_13280,N_13949);
nor U18149 (N_18149,N_13450,N_14085);
and U18150 (N_18150,N_12079,N_10548);
xnor U18151 (N_18151,N_13886,N_11884);
nand U18152 (N_18152,N_11399,N_10365);
nor U18153 (N_18153,N_10664,N_14300);
and U18154 (N_18154,N_10340,N_13649);
nand U18155 (N_18155,N_11079,N_13519);
nor U18156 (N_18156,N_12045,N_12536);
nor U18157 (N_18157,N_12992,N_10390);
and U18158 (N_18158,N_14051,N_12500);
nand U18159 (N_18159,N_13976,N_13778);
or U18160 (N_18160,N_12857,N_13875);
nor U18161 (N_18161,N_11678,N_11399);
nand U18162 (N_18162,N_13112,N_12560);
nor U18163 (N_18163,N_13758,N_11772);
or U18164 (N_18164,N_11577,N_13539);
nand U18165 (N_18165,N_14866,N_14720);
nand U18166 (N_18166,N_14620,N_13386);
and U18167 (N_18167,N_10438,N_14791);
and U18168 (N_18168,N_11147,N_14095);
nand U18169 (N_18169,N_10025,N_11545);
nand U18170 (N_18170,N_14438,N_11458);
xnor U18171 (N_18171,N_14395,N_10902);
nand U18172 (N_18172,N_14033,N_14886);
or U18173 (N_18173,N_14234,N_13126);
or U18174 (N_18174,N_14711,N_14621);
and U18175 (N_18175,N_14983,N_12817);
xnor U18176 (N_18176,N_14471,N_11265);
or U18177 (N_18177,N_13199,N_13197);
nor U18178 (N_18178,N_11219,N_13619);
or U18179 (N_18179,N_12967,N_11915);
or U18180 (N_18180,N_10655,N_10665);
nand U18181 (N_18181,N_10388,N_14658);
xor U18182 (N_18182,N_11546,N_13848);
nand U18183 (N_18183,N_10151,N_10238);
and U18184 (N_18184,N_13869,N_11623);
and U18185 (N_18185,N_12661,N_10558);
or U18186 (N_18186,N_11894,N_10537);
or U18187 (N_18187,N_14264,N_12941);
nand U18188 (N_18188,N_13102,N_10620);
or U18189 (N_18189,N_11549,N_14457);
nand U18190 (N_18190,N_11694,N_12672);
nor U18191 (N_18191,N_14361,N_14779);
nor U18192 (N_18192,N_12563,N_10693);
or U18193 (N_18193,N_13965,N_13439);
nand U18194 (N_18194,N_12170,N_10532);
or U18195 (N_18195,N_11860,N_13109);
nand U18196 (N_18196,N_13211,N_12785);
xnor U18197 (N_18197,N_12260,N_12196);
xor U18198 (N_18198,N_14490,N_11258);
or U18199 (N_18199,N_14339,N_11977);
nor U18200 (N_18200,N_14618,N_11476);
nand U18201 (N_18201,N_14083,N_14279);
and U18202 (N_18202,N_11428,N_13450);
nor U18203 (N_18203,N_11950,N_13244);
or U18204 (N_18204,N_10123,N_11683);
xnor U18205 (N_18205,N_14121,N_11267);
nor U18206 (N_18206,N_14550,N_11684);
or U18207 (N_18207,N_11345,N_13359);
or U18208 (N_18208,N_14637,N_13892);
and U18209 (N_18209,N_14265,N_11284);
or U18210 (N_18210,N_14544,N_14307);
or U18211 (N_18211,N_14549,N_14391);
or U18212 (N_18212,N_10827,N_14733);
xor U18213 (N_18213,N_12065,N_13510);
or U18214 (N_18214,N_14064,N_10110);
or U18215 (N_18215,N_10591,N_13179);
or U18216 (N_18216,N_13680,N_14649);
xor U18217 (N_18217,N_10154,N_11792);
nand U18218 (N_18218,N_13001,N_14251);
nor U18219 (N_18219,N_12183,N_11908);
xnor U18220 (N_18220,N_13245,N_10021);
nor U18221 (N_18221,N_10793,N_12986);
nand U18222 (N_18222,N_11405,N_12003);
or U18223 (N_18223,N_10082,N_12881);
nand U18224 (N_18224,N_12932,N_11715);
nand U18225 (N_18225,N_11684,N_11683);
nand U18226 (N_18226,N_13646,N_12734);
and U18227 (N_18227,N_11686,N_13729);
nand U18228 (N_18228,N_10037,N_13714);
xnor U18229 (N_18229,N_10307,N_12097);
nand U18230 (N_18230,N_10071,N_13106);
nand U18231 (N_18231,N_12010,N_11381);
or U18232 (N_18232,N_10481,N_13624);
nor U18233 (N_18233,N_14322,N_10482);
nand U18234 (N_18234,N_14255,N_10328);
nand U18235 (N_18235,N_11762,N_12451);
and U18236 (N_18236,N_11400,N_13095);
nor U18237 (N_18237,N_12441,N_13799);
and U18238 (N_18238,N_12423,N_11088);
or U18239 (N_18239,N_11258,N_10163);
and U18240 (N_18240,N_13576,N_10625);
or U18241 (N_18241,N_11131,N_13099);
xor U18242 (N_18242,N_12528,N_11876);
nor U18243 (N_18243,N_11392,N_10761);
and U18244 (N_18244,N_10450,N_13118);
nand U18245 (N_18245,N_10427,N_10064);
nor U18246 (N_18246,N_14633,N_12199);
and U18247 (N_18247,N_12022,N_13063);
or U18248 (N_18248,N_14646,N_13333);
xnor U18249 (N_18249,N_10714,N_14017);
nand U18250 (N_18250,N_14785,N_13085);
nor U18251 (N_18251,N_13440,N_14908);
and U18252 (N_18252,N_10228,N_11513);
or U18253 (N_18253,N_11719,N_10705);
nor U18254 (N_18254,N_11930,N_13642);
and U18255 (N_18255,N_13801,N_14819);
xnor U18256 (N_18256,N_14996,N_11823);
and U18257 (N_18257,N_11595,N_13385);
nand U18258 (N_18258,N_10977,N_13094);
and U18259 (N_18259,N_11964,N_12245);
nor U18260 (N_18260,N_12223,N_13639);
and U18261 (N_18261,N_13909,N_10459);
and U18262 (N_18262,N_13275,N_14541);
or U18263 (N_18263,N_14310,N_11733);
nor U18264 (N_18264,N_14593,N_11411);
nand U18265 (N_18265,N_13304,N_13768);
nor U18266 (N_18266,N_10225,N_14568);
nand U18267 (N_18267,N_13924,N_13714);
and U18268 (N_18268,N_14909,N_12831);
xor U18269 (N_18269,N_14328,N_11451);
or U18270 (N_18270,N_13587,N_13862);
nor U18271 (N_18271,N_10803,N_13826);
and U18272 (N_18272,N_12944,N_10784);
nand U18273 (N_18273,N_11976,N_12141);
nand U18274 (N_18274,N_10462,N_14005);
nand U18275 (N_18275,N_14683,N_10294);
and U18276 (N_18276,N_13435,N_14335);
and U18277 (N_18277,N_11959,N_11155);
nand U18278 (N_18278,N_11015,N_11098);
or U18279 (N_18279,N_14391,N_11523);
nor U18280 (N_18280,N_12912,N_14980);
and U18281 (N_18281,N_13115,N_11686);
nand U18282 (N_18282,N_10123,N_13750);
and U18283 (N_18283,N_14484,N_13653);
nor U18284 (N_18284,N_12944,N_13329);
and U18285 (N_18285,N_13301,N_10458);
or U18286 (N_18286,N_13707,N_11728);
nor U18287 (N_18287,N_13483,N_12757);
and U18288 (N_18288,N_14703,N_12059);
and U18289 (N_18289,N_14726,N_13657);
nor U18290 (N_18290,N_14165,N_12306);
nand U18291 (N_18291,N_10414,N_14882);
and U18292 (N_18292,N_12571,N_13371);
xor U18293 (N_18293,N_11144,N_10222);
nand U18294 (N_18294,N_10954,N_13433);
or U18295 (N_18295,N_12744,N_10633);
and U18296 (N_18296,N_14038,N_14339);
nand U18297 (N_18297,N_10207,N_11205);
nor U18298 (N_18298,N_11386,N_11140);
nand U18299 (N_18299,N_11916,N_11425);
nand U18300 (N_18300,N_13868,N_13414);
nand U18301 (N_18301,N_10219,N_12170);
or U18302 (N_18302,N_13144,N_10177);
and U18303 (N_18303,N_11611,N_13637);
nand U18304 (N_18304,N_12191,N_11005);
nand U18305 (N_18305,N_11713,N_10323);
nand U18306 (N_18306,N_12319,N_10341);
nand U18307 (N_18307,N_14173,N_11617);
nor U18308 (N_18308,N_10792,N_13998);
nand U18309 (N_18309,N_14748,N_13039);
or U18310 (N_18310,N_13021,N_12658);
or U18311 (N_18311,N_12758,N_14847);
nand U18312 (N_18312,N_14874,N_10968);
nand U18313 (N_18313,N_14259,N_11805);
and U18314 (N_18314,N_11075,N_10159);
nor U18315 (N_18315,N_10290,N_10083);
or U18316 (N_18316,N_12172,N_12160);
nor U18317 (N_18317,N_13232,N_10293);
and U18318 (N_18318,N_11046,N_10103);
or U18319 (N_18319,N_11000,N_14550);
xnor U18320 (N_18320,N_12188,N_12750);
nor U18321 (N_18321,N_13145,N_14122);
or U18322 (N_18322,N_12894,N_10558);
nand U18323 (N_18323,N_13380,N_12576);
nor U18324 (N_18324,N_10933,N_14682);
nand U18325 (N_18325,N_10086,N_12922);
nor U18326 (N_18326,N_10322,N_13829);
and U18327 (N_18327,N_11147,N_12075);
xor U18328 (N_18328,N_13764,N_10635);
and U18329 (N_18329,N_10041,N_10174);
nor U18330 (N_18330,N_12392,N_11855);
nor U18331 (N_18331,N_11048,N_11401);
and U18332 (N_18332,N_13882,N_10979);
xnor U18333 (N_18333,N_14034,N_13752);
or U18334 (N_18334,N_10162,N_10851);
nor U18335 (N_18335,N_10751,N_14356);
and U18336 (N_18336,N_10235,N_13988);
and U18337 (N_18337,N_10620,N_13702);
xor U18338 (N_18338,N_10304,N_12766);
and U18339 (N_18339,N_14365,N_14820);
nor U18340 (N_18340,N_13675,N_13241);
and U18341 (N_18341,N_11888,N_10904);
xnor U18342 (N_18342,N_12735,N_13476);
nand U18343 (N_18343,N_14296,N_12273);
nand U18344 (N_18344,N_12072,N_13811);
nor U18345 (N_18345,N_10537,N_12013);
nor U18346 (N_18346,N_10469,N_14251);
xnor U18347 (N_18347,N_13869,N_11300);
and U18348 (N_18348,N_11485,N_10121);
nor U18349 (N_18349,N_14209,N_14830);
or U18350 (N_18350,N_12521,N_12752);
nand U18351 (N_18351,N_13256,N_11237);
and U18352 (N_18352,N_13999,N_13301);
nor U18353 (N_18353,N_14898,N_14770);
or U18354 (N_18354,N_14995,N_13999);
nand U18355 (N_18355,N_12887,N_10953);
and U18356 (N_18356,N_13324,N_14304);
nor U18357 (N_18357,N_11711,N_10296);
or U18358 (N_18358,N_11291,N_14123);
nor U18359 (N_18359,N_14644,N_13260);
nand U18360 (N_18360,N_12034,N_10083);
and U18361 (N_18361,N_11152,N_13575);
nand U18362 (N_18362,N_11975,N_12776);
nor U18363 (N_18363,N_14839,N_11801);
nor U18364 (N_18364,N_14257,N_14408);
nand U18365 (N_18365,N_14221,N_14243);
nand U18366 (N_18366,N_12952,N_13667);
nor U18367 (N_18367,N_10991,N_11410);
or U18368 (N_18368,N_13593,N_12965);
nand U18369 (N_18369,N_10071,N_13047);
nor U18370 (N_18370,N_11526,N_14155);
nand U18371 (N_18371,N_10684,N_12208);
and U18372 (N_18372,N_14946,N_14766);
nand U18373 (N_18373,N_10156,N_12906);
nor U18374 (N_18374,N_10252,N_10305);
xor U18375 (N_18375,N_13817,N_10665);
nor U18376 (N_18376,N_14895,N_13133);
and U18377 (N_18377,N_11973,N_10908);
or U18378 (N_18378,N_13902,N_10911);
or U18379 (N_18379,N_14049,N_12351);
nand U18380 (N_18380,N_13773,N_13902);
or U18381 (N_18381,N_11747,N_10724);
nand U18382 (N_18382,N_13546,N_10263);
nor U18383 (N_18383,N_14127,N_14425);
nand U18384 (N_18384,N_13213,N_10453);
and U18385 (N_18385,N_11115,N_14967);
or U18386 (N_18386,N_13893,N_12600);
nand U18387 (N_18387,N_14095,N_13150);
and U18388 (N_18388,N_10541,N_14988);
xnor U18389 (N_18389,N_14122,N_10785);
and U18390 (N_18390,N_11562,N_12986);
nand U18391 (N_18391,N_10969,N_13948);
xor U18392 (N_18392,N_13228,N_14252);
xnor U18393 (N_18393,N_10106,N_11093);
xnor U18394 (N_18394,N_13273,N_13317);
nand U18395 (N_18395,N_12813,N_13431);
nand U18396 (N_18396,N_10133,N_11280);
nor U18397 (N_18397,N_10895,N_14291);
nand U18398 (N_18398,N_10419,N_10107);
nor U18399 (N_18399,N_14448,N_12749);
and U18400 (N_18400,N_14313,N_12992);
nor U18401 (N_18401,N_11990,N_10741);
nor U18402 (N_18402,N_13612,N_12828);
or U18403 (N_18403,N_13041,N_12463);
xor U18404 (N_18404,N_13625,N_12985);
xnor U18405 (N_18405,N_10752,N_10861);
and U18406 (N_18406,N_13024,N_13057);
nor U18407 (N_18407,N_12467,N_14796);
nor U18408 (N_18408,N_10909,N_14323);
and U18409 (N_18409,N_10119,N_10559);
or U18410 (N_18410,N_14151,N_10966);
nand U18411 (N_18411,N_13260,N_11632);
or U18412 (N_18412,N_11574,N_13216);
and U18413 (N_18413,N_11395,N_13424);
and U18414 (N_18414,N_12740,N_12153);
nand U18415 (N_18415,N_11638,N_10046);
nor U18416 (N_18416,N_14425,N_14788);
and U18417 (N_18417,N_13230,N_12324);
or U18418 (N_18418,N_13723,N_14374);
nor U18419 (N_18419,N_11768,N_10620);
nand U18420 (N_18420,N_13500,N_10301);
and U18421 (N_18421,N_13401,N_10993);
and U18422 (N_18422,N_11798,N_14728);
nor U18423 (N_18423,N_14599,N_12802);
and U18424 (N_18424,N_11819,N_13161);
and U18425 (N_18425,N_12880,N_13530);
xnor U18426 (N_18426,N_12082,N_11637);
or U18427 (N_18427,N_13303,N_13208);
nand U18428 (N_18428,N_12924,N_10335);
nand U18429 (N_18429,N_12696,N_13473);
nand U18430 (N_18430,N_10629,N_11980);
or U18431 (N_18431,N_11631,N_12937);
or U18432 (N_18432,N_13379,N_12771);
xnor U18433 (N_18433,N_11861,N_11491);
and U18434 (N_18434,N_12174,N_14259);
nor U18435 (N_18435,N_14704,N_14767);
xor U18436 (N_18436,N_12139,N_14210);
nor U18437 (N_18437,N_14010,N_10721);
or U18438 (N_18438,N_12610,N_14254);
nand U18439 (N_18439,N_13853,N_11139);
nor U18440 (N_18440,N_14464,N_10431);
nand U18441 (N_18441,N_10689,N_13657);
nand U18442 (N_18442,N_10280,N_13163);
or U18443 (N_18443,N_14687,N_12212);
or U18444 (N_18444,N_11664,N_14286);
or U18445 (N_18445,N_13991,N_13892);
and U18446 (N_18446,N_12475,N_13799);
nor U18447 (N_18447,N_13489,N_11226);
or U18448 (N_18448,N_14971,N_14019);
nand U18449 (N_18449,N_12099,N_13193);
or U18450 (N_18450,N_13358,N_12278);
nand U18451 (N_18451,N_11346,N_14389);
and U18452 (N_18452,N_10105,N_11509);
nand U18453 (N_18453,N_13900,N_14578);
or U18454 (N_18454,N_13253,N_13756);
or U18455 (N_18455,N_13074,N_12753);
or U18456 (N_18456,N_12628,N_14589);
nor U18457 (N_18457,N_13170,N_12876);
nand U18458 (N_18458,N_14671,N_10158);
or U18459 (N_18459,N_10779,N_14759);
xnor U18460 (N_18460,N_11860,N_13891);
nor U18461 (N_18461,N_10266,N_13427);
and U18462 (N_18462,N_13953,N_12319);
or U18463 (N_18463,N_13068,N_11276);
xnor U18464 (N_18464,N_12646,N_12270);
nand U18465 (N_18465,N_12497,N_12678);
nand U18466 (N_18466,N_13225,N_14721);
nor U18467 (N_18467,N_12755,N_10387);
or U18468 (N_18468,N_13296,N_14534);
and U18469 (N_18469,N_14425,N_13187);
nand U18470 (N_18470,N_12999,N_11404);
nand U18471 (N_18471,N_14678,N_13972);
or U18472 (N_18472,N_11346,N_10335);
nand U18473 (N_18473,N_14656,N_12546);
and U18474 (N_18474,N_12136,N_14662);
or U18475 (N_18475,N_13293,N_11752);
and U18476 (N_18476,N_11240,N_13376);
and U18477 (N_18477,N_14344,N_14093);
and U18478 (N_18478,N_10625,N_12223);
and U18479 (N_18479,N_13156,N_13027);
and U18480 (N_18480,N_13131,N_11432);
and U18481 (N_18481,N_12428,N_11537);
and U18482 (N_18482,N_14847,N_14334);
nor U18483 (N_18483,N_14871,N_13893);
nor U18484 (N_18484,N_11439,N_14799);
or U18485 (N_18485,N_10112,N_14680);
nand U18486 (N_18486,N_10479,N_11059);
and U18487 (N_18487,N_11774,N_10369);
or U18488 (N_18488,N_14597,N_10616);
or U18489 (N_18489,N_11404,N_14677);
or U18490 (N_18490,N_12251,N_10568);
or U18491 (N_18491,N_11501,N_13572);
and U18492 (N_18492,N_13196,N_11264);
or U18493 (N_18493,N_11357,N_11160);
or U18494 (N_18494,N_10425,N_10080);
nor U18495 (N_18495,N_10634,N_12168);
and U18496 (N_18496,N_14389,N_14782);
nor U18497 (N_18497,N_11666,N_11578);
or U18498 (N_18498,N_11281,N_12852);
nand U18499 (N_18499,N_11859,N_10218);
nor U18500 (N_18500,N_13461,N_11439);
xnor U18501 (N_18501,N_10461,N_12079);
xnor U18502 (N_18502,N_14346,N_14895);
nand U18503 (N_18503,N_11002,N_11673);
nor U18504 (N_18504,N_14872,N_12992);
and U18505 (N_18505,N_12416,N_14743);
and U18506 (N_18506,N_13184,N_12292);
xor U18507 (N_18507,N_11327,N_13532);
nand U18508 (N_18508,N_13654,N_13230);
nand U18509 (N_18509,N_11081,N_10797);
xor U18510 (N_18510,N_13058,N_12187);
nand U18511 (N_18511,N_10825,N_11484);
or U18512 (N_18512,N_10213,N_14197);
nor U18513 (N_18513,N_14039,N_13063);
nor U18514 (N_18514,N_10968,N_11016);
xor U18515 (N_18515,N_11417,N_10105);
xor U18516 (N_18516,N_14917,N_13918);
and U18517 (N_18517,N_10863,N_12664);
and U18518 (N_18518,N_10577,N_12160);
nor U18519 (N_18519,N_11049,N_13931);
or U18520 (N_18520,N_11820,N_13022);
nand U18521 (N_18521,N_13461,N_10642);
nor U18522 (N_18522,N_14298,N_13157);
nand U18523 (N_18523,N_13804,N_11488);
nor U18524 (N_18524,N_13555,N_14595);
and U18525 (N_18525,N_13272,N_10808);
or U18526 (N_18526,N_12821,N_12423);
nand U18527 (N_18527,N_11718,N_14574);
xnor U18528 (N_18528,N_14496,N_10451);
or U18529 (N_18529,N_13735,N_11822);
or U18530 (N_18530,N_13031,N_10939);
nand U18531 (N_18531,N_12139,N_10425);
and U18532 (N_18532,N_10907,N_14120);
and U18533 (N_18533,N_14799,N_12807);
nand U18534 (N_18534,N_11278,N_11853);
and U18535 (N_18535,N_12488,N_11907);
and U18536 (N_18536,N_14236,N_14264);
nand U18537 (N_18537,N_14700,N_13140);
or U18538 (N_18538,N_11159,N_11807);
nor U18539 (N_18539,N_11270,N_12277);
nand U18540 (N_18540,N_14306,N_13306);
nor U18541 (N_18541,N_10047,N_12311);
and U18542 (N_18542,N_11399,N_11665);
nand U18543 (N_18543,N_12299,N_14606);
or U18544 (N_18544,N_13018,N_11069);
and U18545 (N_18545,N_11678,N_13009);
and U18546 (N_18546,N_10904,N_14845);
nand U18547 (N_18547,N_11868,N_10263);
and U18548 (N_18548,N_14313,N_11308);
nand U18549 (N_18549,N_10513,N_13131);
or U18550 (N_18550,N_12733,N_13747);
nor U18551 (N_18551,N_10516,N_11536);
and U18552 (N_18552,N_10009,N_10978);
and U18553 (N_18553,N_10506,N_14849);
and U18554 (N_18554,N_13300,N_11595);
nor U18555 (N_18555,N_11815,N_12122);
or U18556 (N_18556,N_10077,N_14415);
or U18557 (N_18557,N_11424,N_11653);
nand U18558 (N_18558,N_10737,N_13847);
nor U18559 (N_18559,N_10080,N_10728);
or U18560 (N_18560,N_12493,N_14488);
or U18561 (N_18561,N_14571,N_11055);
and U18562 (N_18562,N_12302,N_11679);
and U18563 (N_18563,N_13987,N_10985);
nand U18564 (N_18564,N_14160,N_13001);
nand U18565 (N_18565,N_12014,N_11014);
xor U18566 (N_18566,N_14173,N_14923);
and U18567 (N_18567,N_10782,N_10715);
or U18568 (N_18568,N_10944,N_14006);
nor U18569 (N_18569,N_10498,N_10258);
nand U18570 (N_18570,N_10085,N_10666);
or U18571 (N_18571,N_14263,N_12774);
and U18572 (N_18572,N_10327,N_13524);
and U18573 (N_18573,N_12197,N_14928);
and U18574 (N_18574,N_10428,N_11151);
or U18575 (N_18575,N_14261,N_14419);
or U18576 (N_18576,N_11122,N_10133);
nand U18577 (N_18577,N_10705,N_11336);
nor U18578 (N_18578,N_14347,N_12499);
or U18579 (N_18579,N_10103,N_14459);
and U18580 (N_18580,N_13064,N_13768);
nand U18581 (N_18581,N_13035,N_14134);
nor U18582 (N_18582,N_11065,N_10989);
xnor U18583 (N_18583,N_13449,N_11412);
nor U18584 (N_18584,N_13202,N_14987);
and U18585 (N_18585,N_12111,N_11760);
or U18586 (N_18586,N_12960,N_13515);
and U18587 (N_18587,N_10454,N_10490);
nor U18588 (N_18588,N_11614,N_10746);
nand U18589 (N_18589,N_12444,N_13557);
nor U18590 (N_18590,N_13860,N_12347);
nor U18591 (N_18591,N_12371,N_10494);
nor U18592 (N_18592,N_11796,N_10044);
and U18593 (N_18593,N_12967,N_13586);
and U18594 (N_18594,N_14247,N_11999);
and U18595 (N_18595,N_12263,N_13546);
or U18596 (N_18596,N_13403,N_13239);
nor U18597 (N_18597,N_11073,N_11787);
or U18598 (N_18598,N_14052,N_14343);
or U18599 (N_18599,N_10115,N_14148);
nor U18600 (N_18600,N_13431,N_12096);
or U18601 (N_18601,N_11760,N_11054);
xor U18602 (N_18602,N_12909,N_12750);
and U18603 (N_18603,N_12153,N_14669);
and U18604 (N_18604,N_13104,N_10259);
xor U18605 (N_18605,N_14308,N_14465);
and U18606 (N_18606,N_13192,N_11091);
xor U18607 (N_18607,N_14317,N_12711);
nand U18608 (N_18608,N_10868,N_14634);
nor U18609 (N_18609,N_11546,N_13621);
nand U18610 (N_18610,N_11862,N_10182);
nor U18611 (N_18611,N_10547,N_13126);
or U18612 (N_18612,N_11787,N_11009);
nor U18613 (N_18613,N_13260,N_13913);
and U18614 (N_18614,N_13119,N_14538);
nor U18615 (N_18615,N_12841,N_10131);
nand U18616 (N_18616,N_11044,N_10559);
nand U18617 (N_18617,N_14660,N_13850);
or U18618 (N_18618,N_10885,N_13681);
or U18619 (N_18619,N_14683,N_12969);
xor U18620 (N_18620,N_13287,N_12310);
nand U18621 (N_18621,N_11970,N_11340);
nand U18622 (N_18622,N_10819,N_14408);
and U18623 (N_18623,N_10554,N_10406);
and U18624 (N_18624,N_10896,N_13185);
and U18625 (N_18625,N_10064,N_10418);
and U18626 (N_18626,N_13953,N_13963);
and U18627 (N_18627,N_13873,N_12193);
xnor U18628 (N_18628,N_13092,N_14226);
and U18629 (N_18629,N_10376,N_10580);
or U18630 (N_18630,N_12219,N_10387);
nor U18631 (N_18631,N_12342,N_12094);
nand U18632 (N_18632,N_13479,N_11551);
or U18633 (N_18633,N_14227,N_14735);
nor U18634 (N_18634,N_14773,N_14392);
and U18635 (N_18635,N_10354,N_12349);
or U18636 (N_18636,N_12347,N_10015);
and U18637 (N_18637,N_10528,N_10177);
nand U18638 (N_18638,N_11717,N_10948);
or U18639 (N_18639,N_13196,N_12354);
or U18640 (N_18640,N_14041,N_12044);
nor U18641 (N_18641,N_14796,N_13978);
nand U18642 (N_18642,N_10767,N_14589);
nor U18643 (N_18643,N_11933,N_12602);
or U18644 (N_18644,N_10912,N_12183);
and U18645 (N_18645,N_10730,N_12137);
nor U18646 (N_18646,N_13605,N_12689);
and U18647 (N_18647,N_11683,N_12497);
and U18648 (N_18648,N_13914,N_11076);
and U18649 (N_18649,N_14017,N_12860);
and U18650 (N_18650,N_13514,N_13314);
or U18651 (N_18651,N_13556,N_12218);
or U18652 (N_18652,N_10105,N_13754);
or U18653 (N_18653,N_10081,N_10487);
or U18654 (N_18654,N_11882,N_12134);
or U18655 (N_18655,N_11574,N_10992);
nand U18656 (N_18656,N_10708,N_10498);
or U18657 (N_18657,N_11213,N_13490);
xor U18658 (N_18658,N_12702,N_11370);
nand U18659 (N_18659,N_13909,N_12284);
nor U18660 (N_18660,N_12869,N_12011);
nor U18661 (N_18661,N_13849,N_11781);
or U18662 (N_18662,N_14729,N_14062);
nand U18663 (N_18663,N_10350,N_14510);
nor U18664 (N_18664,N_10593,N_13146);
and U18665 (N_18665,N_10815,N_10170);
nand U18666 (N_18666,N_10961,N_10964);
nand U18667 (N_18667,N_10061,N_14407);
nor U18668 (N_18668,N_13348,N_14388);
nand U18669 (N_18669,N_14784,N_14902);
and U18670 (N_18670,N_11178,N_11039);
nand U18671 (N_18671,N_14309,N_11345);
nand U18672 (N_18672,N_12450,N_13914);
nor U18673 (N_18673,N_12506,N_12957);
nand U18674 (N_18674,N_13008,N_14892);
nor U18675 (N_18675,N_14188,N_12118);
or U18676 (N_18676,N_14577,N_14784);
nor U18677 (N_18677,N_11952,N_10534);
or U18678 (N_18678,N_12551,N_14386);
nor U18679 (N_18679,N_14290,N_11000);
nor U18680 (N_18680,N_11877,N_11778);
nand U18681 (N_18681,N_14091,N_10474);
or U18682 (N_18682,N_10656,N_14763);
or U18683 (N_18683,N_11904,N_11229);
nand U18684 (N_18684,N_14834,N_14619);
nor U18685 (N_18685,N_12498,N_14600);
and U18686 (N_18686,N_11325,N_14960);
nor U18687 (N_18687,N_11182,N_14243);
xnor U18688 (N_18688,N_11681,N_13533);
or U18689 (N_18689,N_12889,N_10611);
nand U18690 (N_18690,N_11286,N_10145);
and U18691 (N_18691,N_14934,N_10624);
and U18692 (N_18692,N_12957,N_10541);
nand U18693 (N_18693,N_11810,N_11146);
and U18694 (N_18694,N_14847,N_13044);
nand U18695 (N_18695,N_10911,N_10214);
and U18696 (N_18696,N_12609,N_10956);
nand U18697 (N_18697,N_12258,N_12795);
nor U18698 (N_18698,N_11331,N_14500);
and U18699 (N_18699,N_10541,N_10724);
and U18700 (N_18700,N_12788,N_12859);
and U18701 (N_18701,N_13267,N_10483);
nand U18702 (N_18702,N_10913,N_11961);
xor U18703 (N_18703,N_14791,N_11233);
and U18704 (N_18704,N_10984,N_14522);
and U18705 (N_18705,N_12526,N_13623);
or U18706 (N_18706,N_10561,N_11903);
and U18707 (N_18707,N_12992,N_10169);
and U18708 (N_18708,N_14816,N_10403);
or U18709 (N_18709,N_11584,N_11535);
xnor U18710 (N_18710,N_12659,N_10073);
xor U18711 (N_18711,N_11989,N_11982);
nand U18712 (N_18712,N_11596,N_10441);
nor U18713 (N_18713,N_10993,N_11547);
and U18714 (N_18714,N_13998,N_14202);
or U18715 (N_18715,N_13118,N_14434);
or U18716 (N_18716,N_14827,N_14313);
or U18717 (N_18717,N_13013,N_11453);
and U18718 (N_18718,N_13003,N_10867);
nand U18719 (N_18719,N_12365,N_10945);
or U18720 (N_18720,N_10561,N_10854);
nor U18721 (N_18721,N_10386,N_11613);
and U18722 (N_18722,N_11635,N_14341);
or U18723 (N_18723,N_12555,N_10619);
nor U18724 (N_18724,N_11979,N_11894);
and U18725 (N_18725,N_14397,N_13366);
nand U18726 (N_18726,N_11313,N_12484);
nand U18727 (N_18727,N_10633,N_11571);
nor U18728 (N_18728,N_10140,N_12674);
nor U18729 (N_18729,N_10118,N_11165);
and U18730 (N_18730,N_14365,N_11079);
or U18731 (N_18731,N_12548,N_10613);
or U18732 (N_18732,N_10640,N_14787);
nor U18733 (N_18733,N_14357,N_12863);
and U18734 (N_18734,N_13296,N_14713);
xor U18735 (N_18735,N_13327,N_12268);
nand U18736 (N_18736,N_12724,N_12301);
nor U18737 (N_18737,N_10437,N_13228);
or U18738 (N_18738,N_14979,N_11041);
nor U18739 (N_18739,N_12899,N_11437);
nor U18740 (N_18740,N_10471,N_13793);
nor U18741 (N_18741,N_10045,N_12936);
nand U18742 (N_18742,N_11611,N_12076);
and U18743 (N_18743,N_10644,N_10623);
or U18744 (N_18744,N_10136,N_11815);
nor U18745 (N_18745,N_10311,N_12865);
or U18746 (N_18746,N_10986,N_13457);
nand U18747 (N_18747,N_14594,N_11915);
nor U18748 (N_18748,N_10086,N_10180);
nor U18749 (N_18749,N_12397,N_14525);
and U18750 (N_18750,N_12997,N_13009);
xor U18751 (N_18751,N_14100,N_10480);
or U18752 (N_18752,N_10239,N_12228);
and U18753 (N_18753,N_11587,N_12531);
nor U18754 (N_18754,N_10129,N_14206);
or U18755 (N_18755,N_10473,N_14792);
nand U18756 (N_18756,N_10383,N_13669);
nand U18757 (N_18757,N_13400,N_11947);
nor U18758 (N_18758,N_14755,N_14585);
and U18759 (N_18759,N_14294,N_13825);
nand U18760 (N_18760,N_12050,N_12445);
and U18761 (N_18761,N_13147,N_12179);
or U18762 (N_18762,N_10032,N_12599);
nor U18763 (N_18763,N_14955,N_10061);
or U18764 (N_18764,N_12930,N_10001);
nand U18765 (N_18765,N_11759,N_14709);
nand U18766 (N_18766,N_11796,N_11025);
nor U18767 (N_18767,N_12994,N_10180);
and U18768 (N_18768,N_11725,N_12590);
nor U18769 (N_18769,N_13071,N_14902);
nor U18770 (N_18770,N_14568,N_13680);
nand U18771 (N_18771,N_14532,N_14276);
nand U18772 (N_18772,N_12542,N_13322);
or U18773 (N_18773,N_14879,N_11219);
nand U18774 (N_18774,N_12381,N_14447);
nor U18775 (N_18775,N_13550,N_12615);
and U18776 (N_18776,N_10368,N_13218);
or U18777 (N_18777,N_10839,N_13235);
or U18778 (N_18778,N_11959,N_10420);
and U18779 (N_18779,N_10959,N_11883);
xnor U18780 (N_18780,N_13931,N_10813);
or U18781 (N_18781,N_10191,N_10312);
xor U18782 (N_18782,N_14606,N_10585);
nor U18783 (N_18783,N_13797,N_10282);
xnor U18784 (N_18784,N_14307,N_14296);
nand U18785 (N_18785,N_14925,N_10116);
nor U18786 (N_18786,N_14089,N_10580);
or U18787 (N_18787,N_12762,N_12692);
and U18788 (N_18788,N_11491,N_14052);
nor U18789 (N_18789,N_14374,N_13619);
nand U18790 (N_18790,N_14441,N_14149);
nand U18791 (N_18791,N_14645,N_14814);
nand U18792 (N_18792,N_14120,N_10541);
nor U18793 (N_18793,N_13997,N_13351);
nor U18794 (N_18794,N_13206,N_11942);
nor U18795 (N_18795,N_10516,N_12960);
and U18796 (N_18796,N_11591,N_10894);
or U18797 (N_18797,N_11759,N_13971);
nor U18798 (N_18798,N_11435,N_13698);
nor U18799 (N_18799,N_13995,N_12344);
or U18800 (N_18800,N_13162,N_11098);
or U18801 (N_18801,N_11011,N_14128);
and U18802 (N_18802,N_10284,N_11649);
nor U18803 (N_18803,N_13539,N_11197);
and U18804 (N_18804,N_14536,N_13229);
or U18805 (N_18805,N_10617,N_13560);
or U18806 (N_18806,N_14807,N_13049);
nor U18807 (N_18807,N_12929,N_10106);
nand U18808 (N_18808,N_11117,N_13541);
xor U18809 (N_18809,N_11752,N_14519);
and U18810 (N_18810,N_12826,N_10250);
and U18811 (N_18811,N_12400,N_13547);
or U18812 (N_18812,N_10516,N_14067);
and U18813 (N_18813,N_10800,N_11366);
nor U18814 (N_18814,N_12211,N_14843);
and U18815 (N_18815,N_10427,N_14063);
and U18816 (N_18816,N_10541,N_13610);
nand U18817 (N_18817,N_12670,N_14736);
and U18818 (N_18818,N_11784,N_13564);
or U18819 (N_18819,N_13636,N_14675);
nand U18820 (N_18820,N_14639,N_10655);
nor U18821 (N_18821,N_10540,N_11405);
or U18822 (N_18822,N_13473,N_13343);
nand U18823 (N_18823,N_14497,N_12218);
xor U18824 (N_18824,N_13536,N_14551);
and U18825 (N_18825,N_11850,N_10086);
nand U18826 (N_18826,N_12465,N_13042);
or U18827 (N_18827,N_11207,N_13113);
and U18828 (N_18828,N_13180,N_13838);
nand U18829 (N_18829,N_11473,N_14458);
and U18830 (N_18830,N_12220,N_13882);
or U18831 (N_18831,N_11504,N_10227);
or U18832 (N_18832,N_11118,N_11930);
nand U18833 (N_18833,N_13762,N_13393);
nor U18834 (N_18834,N_14799,N_10492);
xor U18835 (N_18835,N_11142,N_12087);
nor U18836 (N_18836,N_14841,N_12345);
nor U18837 (N_18837,N_14046,N_12735);
nor U18838 (N_18838,N_14320,N_12236);
nor U18839 (N_18839,N_11326,N_12411);
and U18840 (N_18840,N_12903,N_10367);
or U18841 (N_18841,N_10719,N_10703);
and U18842 (N_18842,N_14358,N_12971);
or U18843 (N_18843,N_10778,N_11049);
and U18844 (N_18844,N_12425,N_14017);
and U18845 (N_18845,N_11495,N_11416);
nand U18846 (N_18846,N_13584,N_12338);
nand U18847 (N_18847,N_11796,N_13686);
nor U18848 (N_18848,N_10809,N_10712);
nand U18849 (N_18849,N_10040,N_12378);
and U18850 (N_18850,N_14973,N_10656);
and U18851 (N_18851,N_14150,N_11492);
nand U18852 (N_18852,N_10950,N_14555);
and U18853 (N_18853,N_13924,N_11802);
nor U18854 (N_18854,N_10851,N_11796);
or U18855 (N_18855,N_12629,N_12527);
or U18856 (N_18856,N_12018,N_14799);
or U18857 (N_18857,N_11052,N_14705);
nand U18858 (N_18858,N_10453,N_11897);
nor U18859 (N_18859,N_10016,N_13676);
or U18860 (N_18860,N_13356,N_11291);
and U18861 (N_18861,N_11171,N_12392);
and U18862 (N_18862,N_14969,N_10150);
nor U18863 (N_18863,N_11366,N_14509);
xor U18864 (N_18864,N_10316,N_10704);
or U18865 (N_18865,N_11269,N_10184);
nand U18866 (N_18866,N_11071,N_13595);
or U18867 (N_18867,N_14697,N_13527);
xnor U18868 (N_18868,N_12171,N_11268);
and U18869 (N_18869,N_12019,N_13908);
nor U18870 (N_18870,N_10419,N_12452);
and U18871 (N_18871,N_11415,N_12539);
or U18872 (N_18872,N_10971,N_13317);
or U18873 (N_18873,N_10096,N_12168);
nor U18874 (N_18874,N_10233,N_12834);
and U18875 (N_18875,N_14447,N_10073);
nor U18876 (N_18876,N_14150,N_14393);
nor U18877 (N_18877,N_14538,N_13661);
xor U18878 (N_18878,N_12561,N_14408);
or U18879 (N_18879,N_12762,N_10020);
nand U18880 (N_18880,N_11240,N_11616);
nand U18881 (N_18881,N_10519,N_12329);
nand U18882 (N_18882,N_10199,N_12085);
and U18883 (N_18883,N_11647,N_11118);
and U18884 (N_18884,N_11501,N_13275);
nor U18885 (N_18885,N_13817,N_13438);
nand U18886 (N_18886,N_13160,N_13297);
nor U18887 (N_18887,N_11436,N_14954);
nor U18888 (N_18888,N_14978,N_12814);
xor U18889 (N_18889,N_14099,N_10479);
and U18890 (N_18890,N_10183,N_10932);
or U18891 (N_18891,N_14622,N_14687);
and U18892 (N_18892,N_12048,N_11026);
nand U18893 (N_18893,N_11650,N_14909);
xor U18894 (N_18894,N_11062,N_11206);
nor U18895 (N_18895,N_12871,N_14125);
or U18896 (N_18896,N_12673,N_11013);
and U18897 (N_18897,N_14102,N_12972);
nand U18898 (N_18898,N_14546,N_10617);
or U18899 (N_18899,N_11206,N_12440);
xnor U18900 (N_18900,N_10700,N_14908);
or U18901 (N_18901,N_11120,N_13980);
and U18902 (N_18902,N_13507,N_13423);
nor U18903 (N_18903,N_11858,N_11183);
and U18904 (N_18904,N_13139,N_11872);
nor U18905 (N_18905,N_13159,N_12051);
or U18906 (N_18906,N_10397,N_14533);
and U18907 (N_18907,N_14544,N_14178);
and U18908 (N_18908,N_14340,N_10405);
nand U18909 (N_18909,N_12938,N_13571);
nor U18910 (N_18910,N_13691,N_14780);
nand U18911 (N_18911,N_11345,N_10242);
nor U18912 (N_18912,N_14067,N_13237);
or U18913 (N_18913,N_13956,N_10548);
xor U18914 (N_18914,N_13414,N_10002);
and U18915 (N_18915,N_13423,N_11787);
and U18916 (N_18916,N_11884,N_11601);
nand U18917 (N_18917,N_10248,N_13159);
nor U18918 (N_18918,N_13378,N_10528);
nand U18919 (N_18919,N_12226,N_14287);
and U18920 (N_18920,N_10217,N_13629);
and U18921 (N_18921,N_13317,N_10993);
and U18922 (N_18922,N_12127,N_12106);
and U18923 (N_18923,N_13905,N_13039);
or U18924 (N_18924,N_11920,N_13283);
xor U18925 (N_18925,N_13326,N_14269);
nand U18926 (N_18926,N_12608,N_10509);
or U18927 (N_18927,N_12019,N_13579);
xor U18928 (N_18928,N_12284,N_12535);
nor U18929 (N_18929,N_13392,N_11069);
nand U18930 (N_18930,N_13740,N_12616);
and U18931 (N_18931,N_13411,N_11751);
xor U18932 (N_18932,N_13737,N_12385);
xor U18933 (N_18933,N_12612,N_13654);
xor U18934 (N_18934,N_12783,N_10729);
and U18935 (N_18935,N_10557,N_12302);
and U18936 (N_18936,N_11972,N_10378);
nor U18937 (N_18937,N_12707,N_12590);
or U18938 (N_18938,N_12303,N_11561);
and U18939 (N_18939,N_11482,N_11367);
nand U18940 (N_18940,N_10557,N_13964);
nor U18941 (N_18941,N_11534,N_10393);
xnor U18942 (N_18942,N_12628,N_12870);
nor U18943 (N_18943,N_12066,N_11695);
nand U18944 (N_18944,N_12227,N_10214);
or U18945 (N_18945,N_10154,N_10839);
or U18946 (N_18946,N_10140,N_14506);
and U18947 (N_18947,N_11285,N_10665);
and U18948 (N_18948,N_14477,N_10442);
or U18949 (N_18949,N_13134,N_13465);
or U18950 (N_18950,N_14029,N_10711);
nor U18951 (N_18951,N_11476,N_10467);
nor U18952 (N_18952,N_11680,N_11083);
xor U18953 (N_18953,N_11884,N_11576);
nand U18954 (N_18954,N_11075,N_11735);
and U18955 (N_18955,N_12196,N_13591);
nor U18956 (N_18956,N_14442,N_14109);
and U18957 (N_18957,N_13742,N_10520);
or U18958 (N_18958,N_13703,N_14232);
xnor U18959 (N_18959,N_12370,N_10814);
xor U18960 (N_18960,N_12048,N_11953);
nor U18961 (N_18961,N_11784,N_10217);
nand U18962 (N_18962,N_10046,N_10708);
and U18963 (N_18963,N_12214,N_14057);
xor U18964 (N_18964,N_12862,N_12076);
or U18965 (N_18965,N_11726,N_11160);
and U18966 (N_18966,N_12562,N_11332);
xor U18967 (N_18967,N_11944,N_13313);
and U18968 (N_18968,N_13818,N_12245);
nand U18969 (N_18969,N_12151,N_13895);
nand U18970 (N_18970,N_10034,N_13480);
nand U18971 (N_18971,N_13175,N_10310);
nand U18972 (N_18972,N_12749,N_10063);
nand U18973 (N_18973,N_12374,N_13084);
xor U18974 (N_18974,N_13477,N_12559);
or U18975 (N_18975,N_10249,N_13155);
and U18976 (N_18976,N_10843,N_13889);
nor U18977 (N_18977,N_12130,N_11263);
or U18978 (N_18978,N_11242,N_10186);
nor U18979 (N_18979,N_12555,N_14054);
and U18980 (N_18980,N_13500,N_10508);
nand U18981 (N_18981,N_10041,N_10692);
xnor U18982 (N_18982,N_10145,N_12069);
xor U18983 (N_18983,N_10118,N_12222);
xnor U18984 (N_18984,N_10250,N_10820);
xnor U18985 (N_18985,N_13324,N_14565);
and U18986 (N_18986,N_10702,N_11764);
or U18987 (N_18987,N_11987,N_11935);
xnor U18988 (N_18988,N_13266,N_14800);
nand U18989 (N_18989,N_11229,N_14283);
and U18990 (N_18990,N_11473,N_12546);
nor U18991 (N_18991,N_12159,N_13291);
nand U18992 (N_18992,N_11087,N_13156);
or U18993 (N_18993,N_11072,N_11513);
nand U18994 (N_18994,N_10230,N_13072);
nor U18995 (N_18995,N_10126,N_10833);
xnor U18996 (N_18996,N_10998,N_11880);
nand U18997 (N_18997,N_10371,N_13062);
nor U18998 (N_18998,N_12193,N_12546);
and U18999 (N_18999,N_13998,N_13036);
or U19000 (N_19000,N_12880,N_11018);
and U19001 (N_19001,N_10736,N_12965);
nor U19002 (N_19002,N_13968,N_11925);
or U19003 (N_19003,N_10018,N_14885);
nand U19004 (N_19004,N_11355,N_11792);
and U19005 (N_19005,N_12986,N_14956);
and U19006 (N_19006,N_12509,N_10305);
nor U19007 (N_19007,N_12690,N_14989);
and U19008 (N_19008,N_12613,N_12949);
nand U19009 (N_19009,N_11252,N_14599);
or U19010 (N_19010,N_12734,N_14128);
or U19011 (N_19011,N_13203,N_12285);
or U19012 (N_19012,N_13237,N_12834);
and U19013 (N_19013,N_10131,N_11627);
nor U19014 (N_19014,N_12091,N_10674);
nand U19015 (N_19015,N_10723,N_10698);
and U19016 (N_19016,N_13765,N_13355);
and U19017 (N_19017,N_10784,N_14848);
xor U19018 (N_19018,N_12218,N_12066);
and U19019 (N_19019,N_11031,N_14070);
and U19020 (N_19020,N_14734,N_10894);
nor U19021 (N_19021,N_12233,N_11914);
nand U19022 (N_19022,N_13419,N_12457);
or U19023 (N_19023,N_11905,N_13829);
and U19024 (N_19024,N_14202,N_13805);
nand U19025 (N_19025,N_10296,N_11026);
or U19026 (N_19026,N_10892,N_10199);
or U19027 (N_19027,N_12030,N_11483);
xor U19028 (N_19028,N_11741,N_11307);
or U19029 (N_19029,N_14377,N_11566);
or U19030 (N_19030,N_14535,N_13861);
or U19031 (N_19031,N_14501,N_12839);
nand U19032 (N_19032,N_13860,N_12246);
nor U19033 (N_19033,N_12483,N_13381);
nor U19034 (N_19034,N_13284,N_11439);
nand U19035 (N_19035,N_13501,N_10364);
or U19036 (N_19036,N_11492,N_11092);
nor U19037 (N_19037,N_10129,N_14183);
and U19038 (N_19038,N_13558,N_10369);
nor U19039 (N_19039,N_13220,N_11942);
and U19040 (N_19040,N_13164,N_10823);
or U19041 (N_19041,N_12933,N_11406);
nand U19042 (N_19042,N_11567,N_11790);
and U19043 (N_19043,N_13443,N_12636);
nand U19044 (N_19044,N_10189,N_12974);
or U19045 (N_19045,N_13985,N_13195);
or U19046 (N_19046,N_10216,N_14096);
nand U19047 (N_19047,N_12569,N_14461);
or U19048 (N_19048,N_12379,N_12321);
xor U19049 (N_19049,N_13706,N_14200);
nor U19050 (N_19050,N_13446,N_14614);
or U19051 (N_19051,N_11559,N_10307);
nor U19052 (N_19052,N_11561,N_10845);
nor U19053 (N_19053,N_10989,N_12289);
nand U19054 (N_19054,N_13148,N_13922);
xnor U19055 (N_19055,N_14582,N_13654);
or U19056 (N_19056,N_10615,N_12481);
nand U19057 (N_19057,N_13376,N_11220);
and U19058 (N_19058,N_13240,N_10933);
nor U19059 (N_19059,N_14887,N_12432);
or U19060 (N_19060,N_14376,N_11798);
nand U19061 (N_19061,N_13136,N_13964);
or U19062 (N_19062,N_13429,N_13746);
and U19063 (N_19063,N_10924,N_12575);
or U19064 (N_19064,N_13999,N_14180);
nor U19065 (N_19065,N_14914,N_12558);
and U19066 (N_19066,N_13912,N_11563);
and U19067 (N_19067,N_12307,N_12047);
and U19068 (N_19068,N_10648,N_14155);
nor U19069 (N_19069,N_11718,N_12494);
and U19070 (N_19070,N_11681,N_11214);
nor U19071 (N_19071,N_13624,N_11298);
and U19072 (N_19072,N_12884,N_13531);
xor U19073 (N_19073,N_12948,N_14438);
nor U19074 (N_19074,N_13065,N_13643);
nand U19075 (N_19075,N_13597,N_13462);
and U19076 (N_19076,N_11430,N_14950);
and U19077 (N_19077,N_10710,N_13631);
nand U19078 (N_19078,N_13673,N_11179);
nand U19079 (N_19079,N_11521,N_13814);
nor U19080 (N_19080,N_14898,N_10521);
xnor U19081 (N_19081,N_13506,N_11831);
nand U19082 (N_19082,N_12815,N_12915);
nor U19083 (N_19083,N_11103,N_13589);
xnor U19084 (N_19084,N_12093,N_12307);
nor U19085 (N_19085,N_12489,N_14675);
or U19086 (N_19086,N_14200,N_11121);
nand U19087 (N_19087,N_12938,N_14245);
nand U19088 (N_19088,N_11106,N_10703);
or U19089 (N_19089,N_13125,N_13208);
or U19090 (N_19090,N_14731,N_11777);
nand U19091 (N_19091,N_12115,N_14359);
and U19092 (N_19092,N_11350,N_14614);
nor U19093 (N_19093,N_13017,N_10710);
or U19094 (N_19094,N_14150,N_10562);
or U19095 (N_19095,N_13413,N_12733);
nand U19096 (N_19096,N_14815,N_14215);
nand U19097 (N_19097,N_14217,N_14958);
xnor U19098 (N_19098,N_13708,N_10408);
or U19099 (N_19099,N_13576,N_10481);
xor U19100 (N_19100,N_12610,N_10078);
nor U19101 (N_19101,N_12561,N_14473);
nand U19102 (N_19102,N_10578,N_11489);
and U19103 (N_19103,N_10008,N_11847);
nor U19104 (N_19104,N_12887,N_12546);
nand U19105 (N_19105,N_11109,N_14089);
or U19106 (N_19106,N_10028,N_13402);
nor U19107 (N_19107,N_14813,N_13399);
nand U19108 (N_19108,N_11321,N_13415);
nand U19109 (N_19109,N_13615,N_11962);
nand U19110 (N_19110,N_10046,N_10782);
or U19111 (N_19111,N_12268,N_12723);
and U19112 (N_19112,N_11381,N_14730);
and U19113 (N_19113,N_10982,N_12034);
nand U19114 (N_19114,N_12752,N_10117);
or U19115 (N_19115,N_13723,N_10386);
nor U19116 (N_19116,N_12263,N_13003);
and U19117 (N_19117,N_12556,N_10121);
nand U19118 (N_19118,N_12478,N_10334);
or U19119 (N_19119,N_14813,N_11136);
nor U19120 (N_19120,N_14030,N_12091);
or U19121 (N_19121,N_10385,N_14192);
and U19122 (N_19122,N_14748,N_13243);
nand U19123 (N_19123,N_12342,N_14117);
nor U19124 (N_19124,N_14785,N_14895);
nand U19125 (N_19125,N_10601,N_14825);
or U19126 (N_19126,N_13769,N_11983);
nand U19127 (N_19127,N_10434,N_13772);
nand U19128 (N_19128,N_12575,N_13668);
nor U19129 (N_19129,N_13283,N_14623);
or U19130 (N_19130,N_13061,N_10154);
and U19131 (N_19131,N_10724,N_12564);
xor U19132 (N_19132,N_10956,N_11131);
nand U19133 (N_19133,N_13791,N_13509);
nand U19134 (N_19134,N_12546,N_12438);
nor U19135 (N_19135,N_11881,N_11293);
nor U19136 (N_19136,N_12144,N_10925);
or U19137 (N_19137,N_14140,N_12213);
or U19138 (N_19138,N_13738,N_11258);
or U19139 (N_19139,N_10841,N_14452);
and U19140 (N_19140,N_11962,N_13933);
or U19141 (N_19141,N_14792,N_13002);
and U19142 (N_19142,N_12521,N_14437);
and U19143 (N_19143,N_10183,N_14253);
nor U19144 (N_19144,N_12530,N_10397);
nor U19145 (N_19145,N_12872,N_11886);
or U19146 (N_19146,N_11614,N_10772);
nor U19147 (N_19147,N_12296,N_10364);
nand U19148 (N_19148,N_12969,N_11084);
or U19149 (N_19149,N_11097,N_10334);
xor U19150 (N_19150,N_10483,N_10342);
xnor U19151 (N_19151,N_13196,N_12563);
nor U19152 (N_19152,N_10162,N_11143);
xnor U19153 (N_19153,N_14262,N_10354);
nor U19154 (N_19154,N_12422,N_11420);
xnor U19155 (N_19155,N_12679,N_13815);
nand U19156 (N_19156,N_14909,N_10106);
and U19157 (N_19157,N_13041,N_10908);
and U19158 (N_19158,N_13065,N_10375);
and U19159 (N_19159,N_11306,N_11715);
nor U19160 (N_19160,N_14623,N_12130);
and U19161 (N_19161,N_10176,N_14001);
and U19162 (N_19162,N_10962,N_10241);
and U19163 (N_19163,N_14199,N_12469);
or U19164 (N_19164,N_13089,N_12605);
or U19165 (N_19165,N_13723,N_12749);
nand U19166 (N_19166,N_11116,N_12765);
nor U19167 (N_19167,N_10951,N_12334);
xor U19168 (N_19168,N_11303,N_10289);
and U19169 (N_19169,N_10453,N_12916);
or U19170 (N_19170,N_10873,N_10708);
or U19171 (N_19171,N_11859,N_14117);
and U19172 (N_19172,N_11499,N_11580);
and U19173 (N_19173,N_13929,N_10228);
and U19174 (N_19174,N_13513,N_14561);
xnor U19175 (N_19175,N_11812,N_10772);
nand U19176 (N_19176,N_12830,N_12042);
and U19177 (N_19177,N_10643,N_14785);
nor U19178 (N_19178,N_12279,N_14884);
or U19179 (N_19179,N_12657,N_11149);
and U19180 (N_19180,N_11105,N_11863);
or U19181 (N_19181,N_11107,N_12316);
or U19182 (N_19182,N_14373,N_14174);
or U19183 (N_19183,N_10943,N_13707);
nor U19184 (N_19184,N_11755,N_14162);
and U19185 (N_19185,N_10322,N_14926);
or U19186 (N_19186,N_11205,N_12007);
xor U19187 (N_19187,N_14087,N_12697);
or U19188 (N_19188,N_14879,N_13721);
nand U19189 (N_19189,N_12584,N_10295);
nor U19190 (N_19190,N_12606,N_11054);
nor U19191 (N_19191,N_10808,N_10323);
nand U19192 (N_19192,N_13173,N_12501);
and U19193 (N_19193,N_11762,N_10421);
and U19194 (N_19194,N_10748,N_11436);
and U19195 (N_19195,N_13297,N_14161);
or U19196 (N_19196,N_14721,N_10646);
nand U19197 (N_19197,N_10488,N_13561);
or U19198 (N_19198,N_11322,N_11904);
nor U19199 (N_19199,N_13471,N_10416);
nor U19200 (N_19200,N_10709,N_13808);
and U19201 (N_19201,N_11856,N_11184);
nand U19202 (N_19202,N_11494,N_13672);
nand U19203 (N_19203,N_11605,N_11546);
xnor U19204 (N_19204,N_10376,N_13101);
nor U19205 (N_19205,N_12846,N_12158);
or U19206 (N_19206,N_13797,N_13137);
or U19207 (N_19207,N_13968,N_12296);
nor U19208 (N_19208,N_11978,N_14056);
and U19209 (N_19209,N_12905,N_14338);
nor U19210 (N_19210,N_11856,N_12843);
and U19211 (N_19211,N_10266,N_10467);
and U19212 (N_19212,N_13490,N_11251);
or U19213 (N_19213,N_14710,N_11908);
nand U19214 (N_19214,N_11322,N_14899);
nor U19215 (N_19215,N_10087,N_10336);
nand U19216 (N_19216,N_12138,N_11053);
nand U19217 (N_19217,N_11213,N_10429);
or U19218 (N_19218,N_14417,N_13793);
or U19219 (N_19219,N_12120,N_11930);
nor U19220 (N_19220,N_12731,N_13889);
nand U19221 (N_19221,N_12154,N_14493);
and U19222 (N_19222,N_11987,N_11671);
nor U19223 (N_19223,N_14975,N_12921);
nand U19224 (N_19224,N_12698,N_12172);
nand U19225 (N_19225,N_11893,N_11170);
and U19226 (N_19226,N_11269,N_11935);
xor U19227 (N_19227,N_14399,N_14860);
nand U19228 (N_19228,N_10553,N_12268);
and U19229 (N_19229,N_14510,N_11666);
and U19230 (N_19230,N_14381,N_13413);
nor U19231 (N_19231,N_10591,N_10454);
or U19232 (N_19232,N_11125,N_14955);
or U19233 (N_19233,N_12420,N_11516);
and U19234 (N_19234,N_12565,N_11540);
nor U19235 (N_19235,N_10817,N_14603);
nand U19236 (N_19236,N_14198,N_11271);
and U19237 (N_19237,N_13025,N_10726);
nand U19238 (N_19238,N_13161,N_12004);
nor U19239 (N_19239,N_11074,N_13850);
xor U19240 (N_19240,N_11687,N_11733);
or U19241 (N_19241,N_12453,N_13919);
nand U19242 (N_19242,N_12024,N_12021);
nand U19243 (N_19243,N_14628,N_10673);
and U19244 (N_19244,N_12911,N_14901);
xnor U19245 (N_19245,N_12569,N_11942);
and U19246 (N_19246,N_11761,N_13469);
nand U19247 (N_19247,N_14272,N_10746);
nand U19248 (N_19248,N_12805,N_12468);
xor U19249 (N_19249,N_12056,N_10238);
xor U19250 (N_19250,N_14128,N_13197);
nand U19251 (N_19251,N_13335,N_12523);
or U19252 (N_19252,N_11761,N_10007);
and U19253 (N_19253,N_12412,N_11833);
nand U19254 (N_19254,N_13047,N_12758);
nand U19255 (N_19255,N_11428,N_13985);
or U19256 (N_19256,N_11332,N_10239);
or U19257 (N_19257,N_13937,N_13730);
nor U19258 (N_19258,N_10335,N_11805);
nor U19259 (N_19259,N_14645,N_12786);
or U19260 (N_19260,N_10039,N_11459);
and U19261 (N_19261,N_13149,N_12530);
or U19262 (N_19262,N_10145,N_10664);
and U19263 (N_19263,N_13813,N_14620);
or U19264 (N_19264,N_13028,N_10854);
nor U19265 (N_19265,N_11981,N_12633);
nor U19266 (N_19266,N_13160,N_11225);
nand U19267 (N_19267,N_14688,N_11820);
nor U19268 (N_19268,N_12628,N_14372);
and U19269 (N_19269,N_10128,N_13215);
nand U19270 (N_19270,N_10951,N_14198);
nor U19271 (N_19271,N_12249,N_13835);
nand U19272 (N_19272,N_11794,N_12142);
nand U19273 (N_19273,N_12163,N_10819);
nand U19274 (N_19274,N_12973,N_11808);
nand U19275 (N_19275,N_14864,N_11626);
and U19276 (N_19276,N_10475,N_11062);
nand U19277 (N_19277,N_12994,N_10710);
nor U19278 (N_19278,N_10054,N_12992);
nand U19279 (N_19279,N_11618,N_11082);
or U19280 (N_19280,N_10004,N_10255);
xor U19281 (N_19281,N_11142,N_10036);
and U19282 (N_19282,N_13665,N_12212);
or U19283 (N_19283,N_10331,N_10614);
and U19284 (N_19284,N_10914,N_13456);
xor U19285 (N_19285,N_13270,N_11365);
nor U19286 (N_19286,N_12590,N_11573);
nand U19287 (N_19287,N_14058,N_12366);
and U19288 (N_19288,N_10559,N_11573);
and U19289 (N_19289,N_12551,N_12916);
and U19290 (N_19290,N_11977,N_11189);
and U19291 (N_19291,N_12298,N_11253);
or U19292 (N_19292,N_13556,N_12889);
nor U19293 (N_19293,N_11568,N_11103);
and U19294 (N_19294,N_12825,N_11069);
nand U19295 (N_19295,N_13198,N_12538);
nor U19296 (N_19296,N_13448,N_12073);
and U19297 (N_19297,N_12926,N_13684);
and U19298 (N_19298,N_12754,N_10983);
xnor U19299 (N_19299,N_13256,N_13095);
nand U19300 (N_19300,N_10278,N_14840);
nand U19301 (N_19301,N_10309,N_13490);
xor U19302 (N_19302,N_12890,N_11880);
and U19303 (N_19303,N_14826,N_13404);
nand U19304 (N_19304,N_12968,N_13558);
xnor U19305 (N_19305,N_14300,N_13736);
nand U19306 (N_19306,N_12876,N_10149);
nor U19307 (N_19307,N_14125,N_12187);
nor U19308 (N_19308,N_10427,N_11878);
xor U19309 (N_19309,N_12514,N_14430);
and U19310 (N_19310,N_12146,N_12604);
and U19311 (N_19311,N_10881,N_14436);
nor U19312 (N_19312,N_14103,N_14391);
xnor U19313 (N_19313,N_11011,N_14119);
nand U19314 (N_19314,N_13535,N_12376);
or U19315 (N_19315,N_10911,N_12978);
nor U19316 (N_19316,N_12786,N_12327);
nor U19317 (N_19317,N_10278,N_11546);
nand U19318 (N_19318,N_13341,N_14611);
or U19319 (N_19319,N_12711,N_11501);
nor U19320 (N_19320,N_11488,N_10142);
nand U19321 (N_19321,N_13657,N_11136);
nand U19322 (N_19322,N_12460,N_14300);
nor U19323 (N_19323,N_13250,N_13536);
and U19324 (N_19324,N_11895,N_14359);
nor U19325 (N_19325,N_10807,N_13481);
nor U19326 (N_19326,N_14092,N_12021);
nand U19327 (N_19327,N_12645,N_11846);
nand U19328 (N_19328,N_12667,N_10868);
and U19329 (N_19329,N_12374,N_12137);
or U19330 (N_19330,N_13530,N_11967);
or U19331 (N_19331,N_12496,N_14138);
nor U19332 (N_19332,N_11011,N_11102);
and U19333 (N_19333,N_10519,N_14071);
xor U19334 (N_19334,N_13505,N_13818);
nand U19335 (N_19335,N_11755,N_14734);
and U19336 (N_19336,N_14080,N_11776);
and U19337 (N_19337,N_13181,N_14991);
nor U19338 (N_19338,N_11750,N_10215);
nor U19339 (N_19339,N_12586,N_11016);
and U19340 (N_19340,N_14136,N_10423);
nand U19341 (N_19341,N_10566,N_10919);
and U19342 (N_19342,N_14401,N_13047);
and U19343 (N_19343,N_14495,N_11776);
nand U19344 (N_19344,N_13513,N_11307);
and U19345 (N_19345,N_12975,N_10636);
and U19346 (N_19346,N_10142,N_11838);
and U19347 (N_19347,N_11042,N_13693);
or U19348 (N_19348,N_10797,N_14601);
nor U19349 (N_19349,N_13570,N_13765);
nand U19350 (N_19350,N_13590,N_14420);
and U19351 (N_19351,N_11588,N_13302);
nand U19352 (N_19352,N_14970,N_14065);
nor U19353 (N_19353,N_10547,N_14724);
nor U19354 (N_19354,N_12692,N_13063);
and U19355 (N_19355,N_13132,N_11845);
and U19356 (N_19356,N_12597,N_11494);
or U19357 (N_19357,N_12657,N_12061);
and U19358 (N_19358,N_13892,N_12161);
or U19359 (N_19359,N_10411,N_10916);
and U19360 (N_19360,N_14142,N_14648);
or U19361 (N_19361,N_10665,N_11233);
nand U19362 (N_19362,N_13102,N_12234);
or U19363 (N_19363,N_11650,N_10599);
nor U19364 (N_19364,N_13661,N_10472);
nand U19365 (N_19365,N_13385,N_13322);
nor U19366 (N_19366,N_10608,N_13398);
nor U19367 (N_19367,N_14856,N_11729);
nor U19368 (N_19368,N_10758,N_12905);
nand U19369 (N_19369,N_13186,N_12880);
xnor U19370 (N_19370,N_10018,N_12712);
or U19371 (N_19371,N_12958,N_11967);
nand U19372 (N_19372,N_14607,N_10668);
nand U19373 (N_19373,N_11395,N_10759);
or U19374 (N_19374,N_10183,N_11327);
and U19375 (N_19375,N_10710,N_12535);
or U19376 (N_19376,N_14333,N_11479);
nand U19377 (N_19377,N_11971,N_13939);
nor U19378 (N_19378,N_13247,N_10965);
nand U19379 (N_19379,N_12318,N_12653);
or U19380 (N_19380,N_13945,N_11951);
nor U19381 (N_19381,N_10076,N_12239);
and U19382 (N_19382,N_11841,N_12564);
nor U19383 (N_19383,N_11328,N_10558);
and U19384 (N_19384,N_10785,N_10767);
nand U19385 (N_19385,N_11396,N_14055);
or U19386 (N_19386,N_13381,N_10370);
and U19387 (N_19387,N_11595,N_13819);
nand U19388 (N_19388,N_12434,N_14361);
or U19389 (N_19389,N_11822,N_13486);
and U19390 (N_19390,N_12244,N_11056);
nand U19391 (N_19391,N_12647,N_14331);
xnor U19392 (N_19392,N_10079,N_12496);
nand U19393 (N_19393,N_13841,N_10618);
nand U19394 (N_19394,N_12583,N_10830);
or U19395 (N_19395,N_11349,N_13818);
nand U19396 (N_19396,N_14556,N_11764);
and U19397 (N_19397,N_12610,N_13975);
xnor U19398 (N_19398,N_13017,N_10549);
and U19399 (N_19399,N_13792,N_12475);
and U19400 (N_19400,N_13727,N_10265);
or U19401 (N_19401,N_13010,N_12221);
nor U19402 (N_19402,N_14391,N_14242);
and U19403 (N_19403,N_10819,N_10543);
nor U19404 (N_19404,N_12044,N_13172);
and U19405 (N_19405,N_10943,N_10937);
or U19406 (N_19406,N_10872,N_11153);
nor U19407 (N_19407,N_13455,N_14357);
xnor U19408 (N_19408,N_11065,N_12400);
nor U19409 (N_19409,N_14602,N_14914);
nand U19410 (N_19410,N_10178,N_11221);
and U19411 (N_19411,N_12730,N_11819);
nand U19412 (N_19412,N_14982,N_14776);
and U19413 (N_19413,N_10151,N_12590);
and U19414 (N_19414,N_10419,N_14931);
nor U19415 (N_19415,N_14577,N_13697);
nor U19416 (N_19416,N_11212,N_13103);
xnor U19417 (N_19417,N_13930,N_13988);
and U19418 (N_19418,N_14039,N_12530);
nor U19419 (N_19419,N_11672,N_12511);
nand U19420 (N_19420,N_11952,N_13754);
nand U19421 (N_19421,N_11942,N_12078);
nor U19422 (N_19422,N_14904,N_12996);
or U19423 (N_19423,N_10940,N_12728);
nand U19424 (N_19424,N_11557,N_10463);
or U19425 (N_19425,N_12324,N_10483);
or U19426 (N_19426,N_10889,N_13335);
and U19427 (N_19427,N_11432,N_11847);
nor U19428 (N_19428,N_11039,N_11348);
nor U19429 (N_19429,N_12076,N_14173);
and U19430 (N_19430,N_13421,N_10145);
nand U19431 (N_19431,N_10989,N_14388);
nor U19432 (N_19432,N_14167,N_12343);
and U19433 (N_19433,N_13214,N_10795);
and U19434 (N_19434,N_14312,N_14195);
nor U19435 (N_19435,N_14695,N_10180);
nor U19436 (N_19436,N_10179,N_14206);
xor U19437 (N_19437,N_10819,N_11238);
nor U19438 (N_19438,N_11953,N_13142);
nor U19439 (N_19439,N_11395,N_11977);
nor U19440 (N_19440,N_11980,N_13490);
nor U19441 (N_19441,N_12406,N_12946);
or U19442 (N_19442,N_13746,N_11103);
nor U19443 (N_19443,N_10043,N_14925);
and U19444 (N_19444,N_11200,N_12949);
xnor U19445 (N_19445,N_12300,N_11021);
or U19446 (N_19446,N_13248,N_10296);
nand U19447 (N_19447,N_13429,N_10506);
nand U19448 (N_19448,N_11060,N_13981);
xor U19449 (N_19449,N_12777,N_14523);
nand U19450 (N_19450,N_14415,N_12151);
nor U19451 (N_19451,N_11961,N_13403);
and U19452 (N_19452,N_13377,N_11753);
nand U19453 (N_19453,N_13544,N_14395);
nor U19454 (N_19454,N_13490,N_11745);
and U19455 (N_19455,N_12980,N_14956);
and U19456 (N_19456,N_12503,N_12365);
or U19457 (N_19457,N_13418,N_13950);
or U19458 (N_19458,N_12774,N_11877);
and U19459 (N_19459,N_10744,N_12551);
nor U19460 (N_19460,N_13353,N_14388);
or U19461 (N_19461,N_12839,N_13818);
nand U19462 (N_19462,N_14116,N_13168);
xnor U19463 (N_19463,N_14561,N_10460);
nor U19464 (N_19464,N_14461,N_11696);
nor U19465 (N_19465,N_10223,N_14688);
and U19466 (N_19466,N_13770,N_12241);
or U19467 (N_19467,N_10098,N_10659);
nor U19468 (N_19468,N_11967,N_12825);
or U19469 (N_19469,N_12059,N_12918);
xnor U19470 (N_19470,N_10780,N_14278);
and U19471 (N_19471,N_14505,N_14148);
or U19472 (N_19472,N_11329,N_11228);
nor U19473 (N_19473,N_13831,N_10444);
nand U19474 (N_19474,N_10574,N_12619);
nand U19475 (N_19475,N_10805,N_14592);
or U19476 (N_19476,N_13753,N_14176);
xnor U19477 (N_19477,N_12630,N_10738);
xor U19478 (N_19478,N_14460,N_12524);
xnor U19479 (N_19479,N_13115,N_12242);
or U19480 (N_19480,N_14995,N_10627);
nor U19481 (N_19481,N_12269,N_13128);
nor U19482 (N_19482,N_11587,N_14845);
and U19483 (N_19483,N_12471,N_13834);
xnor U19484 (N_19484,N_13802,N_14872);
nand U19485 (N_19485,N_14630,N_13805);
nor U19486 (N_19486,N_12940,N_11019);
nand U19487 (N_19487,N_10013,N_11855);
and U19488 (N_19488,N_12029,N_12661);
or U19489 (N_19489,N_11371,N_13995);
nand U19490 (N_19490,N_10593,N_13117);
xor U19491 (N_19491,N_11764,N_12282);
nor U19492 (N_19492,N_10621,N_14122);
xor U19493 (N_19493,N_13101,N_10868);
nor U19494 (N_19494,N_11265,N_13867);
nand U19495 (N_19495,N_12783,N_14191);
or U19496 (N_19496,N_10962,N_11949);
or U19497 (N_19497,N_10838,N_12231);
or U19498 (N_19498,N_10972,N_13966);
nand U19499 (N_19499,N_14608,N_11792);
nor U19500 (N_19500,N_14064,N_13733);
and U19501 (N_19501,N_12969,N_14117);
nand U19502 (N_19502,N_13131,N_10119);
or U19503 (N_19503,N_14231,N_12907);
or U19504 (N_19504,N_14367,N_13287);
nand U19505 (N_19505,N_12981,N_11444);
or U19506 (N_19506,N_11715,N_11034);
nor U19507 (N_19507,N_14311,N_14064);
or U19508 (N_19508,N_11995,N_12420);
nor U19509 (N_19509,N_14869,N_14510);
or U19510 (N_19510,N_11772,N_13708);
and U19511 (N_19511,N_10234,N_11267);
nand U19512 (N_19512,N_14261,N_11362);
or U19513 (N_19513,N_14017,N_14862);
and U19514 (N_19514,N_11650,N_10236);
and U19515 (N_19515,N_11790,N_13116);
nor U19516 (N_19516,N_12318,N_10885);
and U19517 (N_19517,N_10051,N_11974);
xnor U19518 (N_19518,N_14104,N_12577);
xnor U19519 (N_19519,N_12071,N_14337);
and U19520 (N_19520,N_10467,N_12755);
or U19521 (N_19521,N_14555,N_12612);
nor U19522 (N_19522,N_14503,N_11129);
nor U19523 (N_19523,N_13100,N_12222);
and U19524 (N_19524,N_14958,N_10375);
or U19525 (N_19525,N_10179,N_12004);
or U19526 (N_19526,N_10244,N_11905);
or U19527 (N_19527,N_10271,N_13061);
nand U19528 (N_19528,N_10016,N_12196);
nor U19529 (N_19529,N_11207,N_14797);
nor U19530 (N_19530,N_10571,N_13882);
and U19531 (N_19531,N_13864,N_10217);
nand U19532 (N_19532,N_14985,N_14649);
nor U19533 (N_19533,N_12783,N_14538);
nor U19534 (N_19534,N_12358,N_12194);
or U19535 (N_19535,N_11383,N_10646);
and U19536 (N_19536,N_12096,N_10922);
and U19537 (N_19537,N_13108,N_10766);
xnor U19538 (N_19538,N_14478,N_12352);
or U19539 (N_19539,N_10323,N_13925);
nor U19540 (N_19540,N_11962,N_10460);
or U19541 (N_19541,N_11848,N_11681);
nor U19542 (N_19542,N_13555,N_14058);
and U19543 (N_19543,N_13462,N_12767);
and U19544 (N_19544,N_10608,N_11730);
nor U19545 (N_19545,N_14652,N_13606);
nand U19546 (N_19546,N_13829,N_13081);
or U19547 (N_19547,N_13517,N_10413);
and U19548 (N_19548,N_14307,N_10944);
nand U19549 (N_19549,N_11346,N_14926);
nor U19550 (N_19550,N_10353,N_13748);
and U19551 (N_19551,N_12698,N_12948);
and U19552 (N_19552,N_12797,N_13038);
xor U19553 (N_19553,N_10767,N_14703);
nand U19554 (N_19554,N_11449,N_12546);
xor U19555 (N_19555,N_12125,N_13088);
xnor U19556 (N_19556,N_11897,N_13411);
nand U19557 (N_19557,N_10932,N_13661);
and U19558 (N_19558,N_10601,N_11397);
xor U19559 (N_19559,N_11033,N_10415);
nor U19560 (N_19560,N_14937,N_14337);
nand U19561 (N_19561,N_13193,N_11764);
or U19562 (N_19562,N_14926,N_12413);
nor U19563 (N_19563,N_10268,N_10063);
nor U19564 (N_19564,N_14899,N_14817);
nand U19565 (N_19565,N_14447,N_12828);
nand U19566 (N_19566,N_11211,N_11245);
nand U19567 (N_19567,N_11817,N_10788);
nor U19568 (N_19568,N_12412,N_10993);
nand U19569 (N_19569,N_11602,N_14321);
and U19570 (N_19570,N_12004,N_14179);
or U19571 (N_19571,N_14277,N_13947);
and U19572 (N_19572,N_13412,N_14407);
and U19573 (N_19573,N_14176,N_12310);
nor U19574 (N_19574,N_12805,N_12762);
or U19575 (N_19575,N_10147,N_12063);
and U19576 (N_19576,N_12163,N_10470);
nor U19577 (N_19577,N_12326,N_11807);
nand U19578 (N_19578,N_14124,N_13509);
and U19579 (N_19579,N_10076,N_10534);
or U19580 (N_19580,N_14295,N_11610);
nand U19581 (N_19581,N_14687,N_13130);
and U19582 (N_19582,N_14550,N_11137);
nor U19583 (N_19583,N_12361,N_11215);
and U19584 (N_19584,N_14081,N_12455);
or U19585 (N_19585,N_11512,N_11862);
xor U19586 (N_19586,N_11909,N_10608);
and U19587 (N_19587,N_14847,N_10280);
nor U19588 (N_19588,N_11247,N_11673);
nand U19589 (N_19589,N_10770,N_12106);
nor U19590 (N_19590,N_11459,N_12362);
or U19591 (N_19591,N_14258,N_10469);
nand U19592 (N_19592,N_14384,N_12882);
or U19593 (N_19593,N_12600,N_14340);
or U19594 (N_19594,N_11297,N_13138);
nor U19595 (N_19595,N_11045,N_14616);
and U19596 (N_19596,N_14677,N_11976);
nand U19597 (N_19597,N_13296,N_11133);
xor U19598 (N_19598,N_14443,N_11440);
or U19599 (N_19599,N_11867,N_12057);
or U19600 (N_19600,N_14904,N_10071);
nand U19601 (N_19601,N_11174,N_14280);
or U19602 (N_19602,N_10995,N_12312);
nand U19603 (N_19603,N_12625,N_10322);
nor U19604 (N_19604,N_10842,N_11207);
nor U19605 (N_19605,N_11084,N_11805);
or U19606 (N_19606,N_11686,N_11086);
and U19607 (N_19607,N_11775,N_13756);
nand U19608 (N_19608,N_10736,N_11850);
and U19609 (N_19609,N_13882,N_11393);
and U19610 (N_19610,N_12710,N_14368);
or U19611 (N_19611,N_12393,N_12882);
or U19612 (N_19612,N_11443,N_13992);
or U19613 (N_19613,N_10543,N_14320);
or U19614 (N_19614,N_10418,N_14756);
nor U19615 (N_19615,N_12078,N_11640);
or U19616 (N_19616,N_12528,N_11119);
or U19617 (N_19617,N_14755,N_11358);
nand U19618 (N_19618,N_12463,N_13154);
nand U19619 (N_19619,N_12507,N_10372);
or U19620 (N_19620,N_10253,N_13996);
xor U19621 (N_19621,N_12398,N_12307);
and U19622 (N_19622,N_14053,N_14545);
nor U19623 (N_19623,N_12088,N_13525);
or U19624 (N_19624,N_13452,N_11808);
and U19625 (N_19625,N_10809,N_11376);
or U19626 (N_19626,N_12491,N_13336);
nor U19627 (N_19627,N_10982,N_12229);
nand U19628 (N_19628,N_11506,N_12686);
nor U19629 (N_19629,N_12633,N_11946);
nand U19630 (N_19630,N_14651,N_11093);
or U19631 (N_19631,N_13411,N_11609);
and U19632 (N_19632,N_12519,N_13032);
nor U19633 (N_19633,N_10084,N_12667);
or U19634 (N_19634,N_10578,N_10053);
nand U19635 (N_19635,N_13763,N_11070);
nor U19636 (N_19636,N_12711,N_10882);
nand U19637 (N_19637,N_11458,N_11730);
or U19638 (N_19638,N_13665,N_12760);
nor U19639 (N_19639,N_10450,N_10284);
or U19640 (N_19640,N_11354,N_10747);
nand U19641 (N_19641,N_10801,N_11689);
nor U19642 (N_19642,N_11207,N_12088);
nor U19643 (N_19643,N_11228,N_12977);
xnor U19644 (N_19644,N_11098,N_14834);
or U19645 (N_19645,N_11755,N_13273);
and U19646 (N_19646,N_10874,N_12521);
and U19647 (N_19647,N_13474,N_13451);
or U19648 (N_19648,N_13005,N_12981);
nand U19649 (N_19649,N_11489,N_14138);
and U19650 (N_19650,N_11279,N_14649);
nor U19651 (N_19651,N_12152,N_14431);
and U19652 (N_19652,N_11346,N_11189);
or U19653 (N_19653,N_12426,N_12086);
or U19654 (N_19654,N_14503,N_12268);
or U19655 (N_19655,N_10690,N_13246);
or U19656 (N_19656,N_14049,N_14610);
nand U19657 (N_19657,N_14483,N_12095);
or U19658 (N_19658,N_14618,N_10280);
and U19659 (N_19659,N_11740,N_14113);
nor U19660 (N_19660,N_13927,N_13712);
and U19661 (N_19661,N_10674,N_10583);
nand U19662 (N_19662,N_12474,N_12710);
nor U19663 (N_19663,N_12906,N_14158);
or U19664 (N_19664,N_14023,N_10618);
xnor U19665 (N_19665,N_14774,N_13930);
nor U19666 (N_19666,N_12817,N_10710);
or U19667 (N_19667,N_14326,N_14303);
and U19668 (N_19668,N_13514,N_12384);
nand U19669 (N_19669,N_11465,N_13688);
or U19670 (N_19670,N_10364,N_11882);
nor U19671 (N_19671,N_11115,N_13591);
and U19672 (N_19672,N_10045,N_14411);
nor U19673 (N_19673,N_14297,N_14506);
nor U19674 (N_19674,N_12240,N_14525);
or U19675 (N_19675,N_10698,N_10540);
and U19676 (N_19676,N_13255,N_14395);
and U19677 (N_19677,N_12056,N_14338);
xor U19678 (N_19678,N_11158,N_11031);
nor U19679 (N_19679,N_11881,N_10364);
and U19680 (N_19680,N_12110,N_12397);
and U19681 (N_19681,N_10460,N_14333);
and U19682 (N_19682,N_12807,N_10815);
nor U19683 (N_19683,N_11375,N_10496);
or U19684 (N_19684,N_10027,N_11278);
nand U19685 (N_19685,N_13040,N_10263);
xnor U19686 (N_19686,N_12089,N_11253);
or U19687 (N_19687,N_13781,N_13387);
or U19688 (N_19688,N_13572,N_11256);
xor U19689 (N_19689,N_12938,N_12984);
nand U19690 (N_19690,N_11657,N_14435);
or U19691 (N_19691,N_11981,N_11941);
nand U19692 (N_19692,N_11451,N_13182);
and U19693 (N_19693,N_12023,N_13081);
nand U19694 (N_19694,N_12125,N_10309);
and U19695 (N_19695,N_12273,N_12678);
or U19696 (N_19696,N_11550,N_11901);
and U19697 (N_19697,N_14775,N_10787);
and U19698 (N_19698,N_10064,N_10380);
and U19699 (N_19699,N_13862,N_14676);
nor U19700 (N_19700,N_11354,N_12675);
xnor U19701 (N_19701,N_12897,N_13009);
nand U19702 (N_19702,N_14185,N_11717);
xnor U19703 (N_19703,N_10595,N_12304);
xor U19704 (N_19704,N_14719,N_11719);
xor U19705 (N_19705,N_10921,N_10929);
nor U19706 (N_19706,N_10400,N_12047);
or U19707 (N_19707,N_14036,N_13973);
and U19708 (N_19708,N_13387,N_12792);
xnor U19709 (N_19709,N_14541,N_11020);
or U19710 (N_19710,N_14826,N_10921);
xnor U19711 (N_19711,N_14791,N_10221);
and U19712 (N_19712,N_13846,N_10272);
nor U19713 (N_19713,N_10285,N_14512);
or U19714 (N_19714,N_12076,N_13194);
nand U19715 (N_19715,N_11168,N_13388);
nor U19716 (N_19716,N_10593,N_13735);
and U19717 (N_19717,N_10013,N_11544);
xor U19718 (N_19718,N_11556,N_12347);
or U19719 (N_19719,N_11197,N_13344);
or U19720 (N_19720,N_10605,N_11070);
and U19721 (N_19721,N_14228,N_11629);
or U19722 (N_19722,N_10549,N_12937);
xnor U19723 (N_19723,N_11381,N_13526);
and U19724 (N_19724,N_12743,N_11891);
or U19725 (N_19725,N_10849,N_10239);
xnor U19726 (N_19726,N_11929,N_13933);
nand U19727 (N_19727,N_14324,N_10675);
nor U19728 (N_19728,N_13536,N_14152);
and U19729 (N_19729,N_10476,N_12814);
and U19730 (N_19730,N_13178,N_12304);
or U19731 (N_19731,N_12133,N_13693);
nor U19732 (N_19732,N_13435,N_11146);
and U19733 (N_19733,N_14431,N_13979);
and U19734 (N_19734,N_10894,N_10769);
or U19735 (N_19735,N_11150,N_13444);
nand U19736 (N_19736,N_14124,N_14128);
xor U19737 (N_19737,N_13210,N_13371);
xor U19738 (N_19738,N_12001,N_13902);
nor U19739 (N_19739,N_12066,N_13177);
or U19740 (N_19740,N_10102,N_13957);
nor U19741 (N_19741,N_14586,N_11727);
nand U19742 (N_19742,N_10128,N_12956);
nand U19743 (N_19743,N_10362,N_11400);
or U19744 (N_19744,N_12835,N_10412);
and U19745 (N_19745,N_13802,N_14021);
xor U19746 (N_19746,N_14453,N_11587);
and U19747 (N_19747,N_10204,N_14869);
and U19748 (N_19748,N_14270,N_13674);
nor U19749 (N_19749,N_10188,N_14236);
and U19750 (N_19750,N_12709,N_13367);
and U19751 (N_19751,N_10343,N_14498);
nand U19752 (N_19752,N_14019,N_13628);
or U19753 (N_19753,N_12232,N_13527);
nand U19754 (N_19754,N_10649,N_11513);
nor U19755 (N_19755,N_13606,N_13684);
xor U19756 (N_19756,N_11388,N_10740);
and U19757 (N_19757,N_11503,N_11234);
nor U19758 (N_19758,N_12544,N_11390);
or U19759 (N_19759,N_14553,N_11820);
and U19760 (N_19760,N_13553,N_14012);
nor U19761 (N_19761,N_11704,N_12552);
or U19762 (N_19762,N_12019,N_14774);
nor U19763 (N_19763,N_13478,N_10864);
and U19764 (N_19764,N_14984,N_12201);
and U19765 (N_19765,N_10789,N_13912);
xnor U19766 (N_19766,N_12998,N_10556);
nand U19767 (N_19767,N_12102,N_11814);
or U19768 (N_19768,N_12538,N_10311);
nand U19769 (N_19769,N_13049,N_11699);
and U19770 (N_19770,N_12555,N_12566);
nand U19771 (N_19771,N_13138,N_13708);
xnor U19772 (N_19772,N_13868,N_13067);
nand U19773 (N_19773,N_14823,N_12106);
or U19774 (N_19774,N_11093,N_10973);
nand U19775 (N_19775,N_11914,N_10620);
and U19776 (N_19776,N_10241,N_10052);
xor U19777 (N_19777,N_10631,N_10053);
and U19778 (N_19778,N_11944,N_12365);
nand U19779 (N_19779,N_14336,N_14823);
nand U19780 (N_19780,N_13441,N_10887);
and U19781 (N_19781,N_11246,N_12402);
and U19782 (N_19782,N_12569,N_10849);
xnor U19783 (N_19783,N_12202,N_13309);
and U19784 (N_19784,N_11674,N_12536);
nand U19785 (N_19785,N_12960,N_13270);
or U19786 (N_19786,N_13357,N_11702);
or U19787 (N_19787,N_14783,N_11942);
nand U19788 (N_19788,N_13959,N_10831);
nand U19789 (N_19789,N_12988,N_14260);
nand U19790 (N_19790,N_11665,N_10704);
xnor U19791 (N_19791,N_11100,N_11762);
nor U19792 (N_19792,N_11361,N_14298);
and U19793 (N_19793,N_12963,N_12666);
nor U19794 (N_19794,N_11694,N_12973);
nand U19795 (N_19795,N_10293,N_13749);
xor U19796 (N_19796,N_11019,N_10581);
and U19797 (N_19797,N_10861,N_10974);
nor U19798 (N_19798,N_10435,N_14090);
xor U19799 (N_19799,N_10777,N_13139);
or U19800 (N_19800,N_13330,N_12913);
nand U19801 (N_19801,N_14951,N_14512);
and U19802 (N_19802,N_12630,N_10045);
and U19803 (N_19803,N_10842,N_10814);
nand U19804 (N_19804,N_13059,N_11297);
xnor U19805 (N_19805,N_11327,N_14539);
and U19806 (N_19806,N_10612,N_13626);
nor U19807 (N_19807,N_11961,N_14332);
xnor U19808 (N_19808,N_11187,N_13018);
xor U19809 (N_19809,N_13610,N_13989);
nand U19810 (N_19810,N_10046,N_12335);
and U19811 (N_19811,N_12130,N_11917);
nor U19812 (N_19812,N_12274,N_13579);
and U19813 (N_19813,N_13681,N_12455);
and U19814 (N_19814,N_10609,N_10751);
nor U19815 (N_19815,N_14591,N_13303);
or U19816 (N_19816,N_11474,N_10549);
xnor U19817 (N_19817,N_12920,N_10045);
or U19818 (N_19818,N_12724,N_14796);
and U19819 (N_19819,N_11990,N_12773);
xor U19820 (N_19820,N_11738,N_14259);
and U19821 (N_19821,N_12571,N_10936);
nand U19822 (N_19822,N_14113,N_14558);
and U19823 (N_19823,N_13509,N_12458);
nor U19824 (N_19824,N_10913,N_13005);
nand U19825 (N_19825,N_12814,N_13642);
and U19826 (N_19826,N_11189,N_13056);
or U19827 (N_19827,N_11277,N_10283);
and U19828 (N_19828,N_10615,N_10620);
nor U19829 (N_19829,N_11729,N_12134);
nor U19830 (N_19830,N_11759,N_13521);
and U19831 (N_19831,N_14647,N_10729);
or U19832 (N_19832,N_10700,N_11860);
and U19833 (N_19833,N_10952,N_10103);
nand U19834 (N_19834,N_10648,N_10051);
nand U19835 (N_19835,N_11351,N_14911);
nor U19836 (N_19836,N_11813,N_10242);
or U19837 (N_19837,N_10783,N_14637);
nor U19838 (N_19838,N_13186,N_11862);
nand U19839 (N_19839,N_10606,N_11410);
nor U19840 (N_19840,N_14675,N_14635);
and U19841 (N_19841,N_12169,N_13240);
nor U19842 (N_19842,N_14046,N_10930);
nor U19843 (N_19843,N_10166,N_11122);
and U19844 (N_19844,N_14613,N_10911);
or U19845 (N_19845,N_13672,N_12539);
nand U19846 (N_19846,N_12702,N_10354);
nor U19847 (N_19847,N_12015,N_13781);
and U19848 (N_19848,N_12201,N_13939);
nor U19849 (N_19849,N_11739,N_11558);
xor U19850 (N_19850,N_12736,N_10090);
or U19851 (N_19851,N_10505,N_12767);
or U19852 (N_19852,N_14688,N_14550);
or U19853 (N_19853,N_12164,N_10268);
or U19854 (N_19854,N_11064,N_12337);
nor U19855 (N_19855,N_14893,N_14189);
or U19856 (N_19856,N_14259,N_13862);
xor U19857 (N_19857,N_12525,N_14417);
and U19858 (N_19858,N_11862,N_12835);
nand U19859 (N_19859,N_10793,N_12080);
nor U19860 (N_19860,N_12417,N_14734);
xnor U19861 (N_19861,N_13885,N_13005);
or U19862 (N_19862,N_14129,N_12405);
nor U19863 (N_19863,N_12223,N_14621);
xor U19864 (N_19864,N_12848,N_14830);
or U19865 (N_19865,N_14504,N_11252);
or U19866 (N_19866,N_14881,N_14260);
and U19867 (N_19867,N_10359,N_12670);
xnor U19868 (N_19868,N_11338,N_10630);
nor U19869 (N_19869,N_14502,N_14363);
nor U19870 (N_19870,N_14151,N_12088);
nor U19871 (N_19871,N_11817,N_12914);
nand U19872 (N_19872,N_13046,N_14630);
or U19873 (N_19873,N_12597,N_14220);
nor U19874 (N_19874,N_12487,N_10950);
nor U19875 (N_19875,N_10168,N_14454);
and U19876 (N_19876,N_12049,N_10917);
and U19877 (N_19877,N_12410,N_13092);
and U19878 (N_19878,N_12370,N_10995);
nor U19879 (N_19879,N_13803,N_13426);
and U19880 (N_19880,N_14273,N_12297);
nand U19881 (N_19881,N_11297,N_10012);
nand U19882 (N_19882,N_11230,N_10796);
nor U19883 (N_19883,N_14872,N_10351);
or U19884 (N_19884,N_12119,N_14052);
or U19885 (N_19885,N_14943,N_11299);
nor U19886 (N_19886,N_13486,N_10385);
nand U19887 (N_19887,N_12381,N_12996);
and U19888 (N_19888,N_14189,N_11879);
nor U19889 (N_19889,N_14610,N_14130);
or U19890 (N_19890,N_11785,N_14887);
nor U19891 (N_19891,N_13149,N_12040);
nand U19892 (N_19892,N_11244,N_13966);
and U19893 (N_19893,N_14579,N_10677);
nor U19894 (N_19894,N_13428,N_14455);
nor U19895 (N_19895,N_14020,N_12595);
nand U19896 (N_19896,N_10724,N_11948);
or U19897 (N_19897,N_14395,N_14841);
xnor U19898 (N_19898,N_10707,N_13600);
nor U19899 (N_19899,N_14367,N_13267);
or U19900 (N_19900,N_11953,N_12862);
nand U19901 (N_19901,N_13154,N_10235);
or U19902 (N_19902,N_11691,N_10662);
nand U19903 (N_19903,N_12927,N_10094);
nand U19904 (N_19904,N_13415,N_14626);
nor U19905 (N_19905,N_14574,N_12281);
and U19906 (N_19906,N_12732,N_11269);
and U19907 (N_19907,N_11510,N_12611);
or U19908 (N_19908,N_10525,N_12934);
nand U19909 (N_19909,N_14224,N_10053);
nor U19910 (N_19910,N_12633,N_14571);
or U19911 (N_19911,N_14536,N_10148);
xor U19912 (N_19912,N_12199,N_14326);
nor U19913 (N_19913,N_14912,N_12897);
xnor U19914 (N_19914,N_11995,N_14464);
nor U19915 (N_19915,N_10578,N_13668);
and U19916 (N_19916,N_13322,N_10851);
and U19917 (N_19917,N_11190,N_11970);
and U19918 (N_19918,N_13472,N_14392);
nor U19919 (N_19919,N_13168,N_13428);
nand U19920 (N_19920,N_10588,N_11844);
nand U19921 (N_19921,N_14637,N_14091);
or U19922 (N_19922,N_10990,N_11879);
and U19923 (N_19923,N_10064,N_11278);
nor U19924 (N_19924,N_11248,N_14042);
and U19925 (N_19925,N_11616,N_13289);
and U19926 (N_19926,N_11574,N_13850);
nand U19927 (N_19927,N_12812,N_13741);
nand U19928 (N_19928,N_10733,N_14103);
nand U19929 (N_19929,N_10833,N_13631);
or U19930 (N_19930,N_11049,N_12651);
nand U19931 (N_19931,N_10178,N_10236);
or U19932 (N_19932,N_13946,N_11949);
and U19933 (N_19933,N_10422,N_11339);
xor U19934 (N_19934,N_11806,N_12972);
and U19935 (N_19935,N_13105,N_10885);
nor U19936 (N_19936,N_14221,N_10367);
nor U19937 (N_19937,N_13318,N_11205);
or U19938 (N_19938,N_13778,N_12649);
and U19939 (N_19939,N_13599,N_12912);
and U19940 (N_19940,N_12774,N_10679);
nand U19941 (N_19941,N_11493,N_12696);
nor U19942 (N_19942,N_12725,N_10798);
and U19943 (N_19943,N_13099,N_12712);
or U19944 (N_19944,N_10440,N_14773);
nor U19945 (N_19945,N_14122,N_14171);
nor U19946 (N_19946,N_11615,N_14003);
xnor U19947 (N_19947,N_14462,N_12360);
and U19948 (N_19948,N_12514,N_10713);
nor U19949 (N_19949,N_14963,N_14523);
nand U19950 (N_19950,N_10261,N_11677);
and U19951 (N_19951,N_11690,N_13427);
xnor U19952 (N_19952,N_11177,N_12597);
xnor U19953 (N_19953,N_13494,N_10815);
and U19954 (N_19954,N_11971,N_11886);
nand U19955 (N_19955,N_10844,N_10012);
nor U19956 (N_19956,N_13668,N_14231);
nand U19957 (N_19957,N_11487,N_11746);
nand U19958 (N_19958,N_13465,N_11808);
and U19959 (N_19959,N_10920,N_12803);
and U19960 (N_19960,N_13031,N_11756);
or U19961 (N_19961,N_12206,N_13539);
xor U19962 (N_19962,N_10895,N_13384);
nor U19963 (N_19963,N_10238,N_14326);
and U19964 (N_19964,N_13928,N_13360);
nor U19965 (N_19965,N_10138,N_12707);
nor U19966 (N_19966,N_10344,N_14716);
xor U19967 (N_19967,N_12059,N_14275);
xor U19968 (N_19968,N_12489,N_13138);
and U19969 (N_19969,N_13877,N_11114);
xor U19970 (N_19970,N_12426,N_14465);
or U19971 (N_19971,N_13080,N_11900);
nor U19972 (N_19972,N_14182,N_10000);
nand U19973 (N_19973,N_10264,N_12705);
nand U19974 (N_19974,N_13106,N_13768);
xnor U19975 (N_19975,N_14283,N_11135);
nor U19976 (N_19976,N_12241,N_14512);
nor U19977 (N_19977,N_12699,N_14389);
nor U19978 (N_19978,N_13123,N_13164);
and U19979 (N_19979,N_12490,N_12866);
and U19980 (N_19980,N_12369,N_14109);
nor U19981 (N_19981,N_11317,N_12982);
nand U19982 (N_19982,N_13515,N_14245);
nor U19983 (N_19983,N_13855,N_10679);
nor U19984 (N_19984,N_11360,N_11983);
and U19985 (N_19985,N_10681,N_14733);
nand U19986 (N_19986,N_13406,N_11503);
nor U19987 (N_19987,N_11072,N_10914);
and U19988 (N_19988,N_12976,N_13635);
nand U19989 (N_19989,N_14425,N_13488);
and U19990 (N_19990,N_13420,N_12374);
or U19991 (N_19991,N_13102,N_11548);
and U19992 (N_19992,N_14299,N_10076);
nor U19993 (N_19993,N_10682,N_14854);
and U19994 (N_19994,N_14323,N_14196);
or U19995 (N_19995,N_12162,N_13283);
nand U19996 (N_19996,N_10503,N_13838);
nor U19997 (N_19997,N_10861,N_10445);
or U19998 (N_19998,N_10136,N_10875);
xor U19999 (N_19999,N_10155,N_12821);
nor U20000 (N_20000,N_19483,N_15533);
xnor U20001 (N_20001,N_15358,N_18623);
xnor U20002 (N_20002,N_18005,N_17126);
nand U20003 (N_20003,N_16132,N_15334);
and U20004 (N_20004,N_17852,N_16762);
xnor U20005 (N_20005,N_17951,N_17456);
xnor U20006 (N_20006,N_17525,N_16451);
xor U20007 (N_20007,N_19811,N_18122);
xor U20008 (N_20008,N_19621,N_17026);
or U20009 (N_20009,N_19590,N_17289);
nor U20010 (N_20010,N_18772,N_15231);
xor U20011 (N_20011,N_18564,N_19508);
nor U20012 (N_20012,N_16917,N_15725);
nand U20013 (N_20013,N_17959,N_16565);
and U20014 (N_20014,N_16033,N_18668);
or U20015 (N_20015,N_17813,N_19850);
or U20016 (N_20016,N_15246,N_17036);
and U20017 (N_20017,N_18933,N_15761);
nor U20018 (N_20018,N_16648,N_15735);
nor U20019 (N_20019,N_19977,N_19486);
and U20020 (N_20020,N_15925,N_16478);
and U20021 (N_20021,N_15798,N_18027);
nor U20022 (N_20022,N_18388,N_16413);
or U20023 (N_20023,N_16150,N_17915);
or U20024 (N_20024,N_18171,N_17090);
nand U20025 (N_20025,N_18379,N_18768);
nand U20026 (N_20026,N_15411,N_18999);
nor U20027 (N_20027,N_16819,N_16402);
or U20028 (N_20028,N_17069,N_19313);
nand U20029 (N_20029,N_17777,N_16484);
nand U20030 (N_20030,N_19064,N_17055);
nand U20031 (N_20031,N_19749,N_16259);
nand U20032 (N_20032,N_16324,N_18694);
or U20033 (N_20033,N_16652,N_18914);
nand U20034 (N_20034,N_17560,N_17874);
and U20035 (N_20035,N_15991,N_18524);
and U20036 (N_20036,N_18634,N_18296);
nand U20037 (N_20037,N_15897,N_17783);
nand U20038 (N_20038,N_19192,N_19118);
nor U20039 (N_20039,N_16381,N_18012);
or U20040 (N_20040,N_15819,N_15372);
nand U20041 (N_20041,N_19880,N_19305);
and U20042 (N_20042,N_17942,N_15091);
nor U20043 (N_20043,N_15715,N_16627);
and U20044 (N_20044,N_18087,N_19241);
nor U20045 (N_20045,N_16383,N_19316);
nor U20046 (N_20046,N_18294,N_18231);
nand U20047 (N_20047,N_18261,N_15392);
nand U20048 (N_20048,N_18497,N_16338);
nand U20049 (N_20049,N_17535,N_16277);
and U20050 (N_20050,N_15693,N_15047);
or U20051 (N_20051,N_16911,N_16349);
nor U20052 (N_20052,N_19351,N_15135);
and U20053 (N_20053,N_17624,N_15900);
nand U20054 (N_20054,N_15766,N_16171);
nor U20055 (N_20055,N_19526,N_16571);
nand U20056 (N_20056,N_15016,N_15563);
and U20057 (N_20057,N_19831,N_16689);
xor U20058 (N_20058,N_17475,N_15967);
xor U20059 (N_20059,N_15311,N_15399);
or U20060 (N_20060,N_15892,N_18046);
nor U20061 (N_20061,N_19204,N_15041);
nand U20062 (N_20062,N_17792,N_16084);
or U20063 (N_20063,N_17365,N_19746);
nand U20064 (N_20064,N_16116,N_16808);
nand U20065 (N_20065,N_19068,N_15888);
nand U20066 (N_20066,N_18055,N_18340);
and U20067 (N_20067,N_16497,N_17423);
nor U20068 (N_20068,N_19866,N_19368);
and U20069 (N_20069,N_19112,N_18154);
and U20070 (N_20070,N_16682,N_18977);
or U20071 (N_20071,N_19145,N_18582);
and U20072 (N_20072,N_16011,N_16832);
or U20073 (N_20073,N_19232,N_18830);
or U20074 (N_20074,N_16303,N_18786);
xor U20075 (N_20075,N_17745,N_19246);
nand U20076 (N_20076,N_19604,N_18007);
xnor U20077 (N_20077,N_17484,N_19176);
and U20078 (N_20078,N_17164,N_17327);
or U20079 (N_20079,N_18511,N_19071);
nand U20080 (N_20080,N_17808,N_19763);
nand U20081 (N_20081,N_16115,N_16583);
xor U20082 (N_20082,N_15444,N_19581);
and U20083 (N_20083,N_17501,N_18916);
or U20084 (N_20084,N_17502,N_19827);
xor U20085 (N_20085,N_19747,N_18872);
nor U20086 (N_20086,N_17408,N_19967);
and U20087 (N_20087,N_16097,N_16811);
and U20088 (N_20088,N_17006,N_16218);
and U20089 (N_20089,N_16248,N_17601);
nor U20090 (N_20090,N_17884,N_18286);
or U20091 (N_20091,N_19292,N_18319);
nor U20092 (N_20092,N_18120,N_16817);
nor U20093 (N_20093,N_16765,N_19655);
nor U20094 (N_20094,N_17835,N_16535);
nand U20095 (N_20095,N_17450,N_16877);
or U20096 (N_20096,N_18644,N_19341);
and U20097 (N_20097,N_16386,N_17531);
nand U20098 (N_20098,N_16058,N_19537);
or U20099 (N_20099,N_15579,N_16049);
nand U20100 (N_20100,N_15926,N_18841);
and U20101 (N_20101,N_19276,N_17492);
nor U20102 (N_20102,N_16982,N_16697);
or U20103 (N_20103,N_19667,N_19730);
or U20104 (N_20104,N_15241,N_19512);
and U20105 (N_20105,N_17779,N_19309);
and U20106 (N_20106,N_15238,N_15218);
nor U20107 (N_20107,N_19251,N_16939);
nand U20108 (N_20108,N_16184,N_18443);
xor U20109 (N_20109,N_19138,N_15596);
and U20110 (N_20110,N_16918,N_17538);
nor U20111 (N_20111,N_19732,N_17756);
xnor U20112 (N_20112,N_18606,N_17115);
nor U20113 (N_20113,N_19668,N_15100);
nand U20114 (N_20114,N_19430,N_15065);
and U20115 (N_20115,N_18718,N_16858);
nand U20116 (N_20116,N_18331,N_18085);
nand U20117 (N_20117,N_17628,N_17367);
nor U20118 (N_20118,N_16030,N_19008);
nand U20119 (N_20119,N_15629,N_17710);
and U20120 (N_20120,N_17195,N_16806);
nand U20121 (N_20121,N_17165,N_15318);
xnor U20122 (N_20122,N_17578,N_19653);
nand U20123 (N_20123,N_16938,N_18690);
nand U20124 (N_20124,N_19713,N_18291);
or U20125 (N_20125,N_17795,N_16999);
nor U20126 (N_20126,N_17843,N_19834);
nor U20127 (N_20127,N_15966,N_16691);
nand U20128 (N_20128,N_15811,N_19685);
xor U20129 (N_20129,N_19283,N_18566);
xnor U20130 (N_20130,N_17615,N_16659);
xor U20131 (N_20131,N_17645,N_15657);
or U20132 (N_20132,N_17857,N_18325);
or U20133 (N_20133,N_19933,N_16569);
nand U20134 (N_20134,N_16540,N_16421);
or U20135 (N_20135,N_19051,N_17943);
or U20136 (N_20136,N_18874,N_17461);
or U20137 (N_20137,N_16521,N_19433);
nand U20138 (N_20138,N_16371,N_19652);
xnor U20139 (N_20139,N_18762,N_19139);
and U20140 (N_20140,N_15731,N_15574);
xnor U20141 (N_20141,N_15712,N_16483);
xor U20142 (N_20142,N_15010,N_17198);
xor U20143 (N_20143,N_19388,N_17332);
and U20144 (N_20144,N_17944,N_19677);
and U20145 (N_20145,N_17184,N_16807);
or U20146 (N_20146,N_19669,N_15433);
or U20147 (N_20147,N_15542,N_17337);
nor U20148 (N_20148,N_16404,N_16065);
and U20149 (N_20149,N_16680,N_15872);
nor U20150 (N_20150,N_15415,N_17839);
xnor U20151 (N_20151,N_17070,N_15868);
and U20152 (N_20152,N_15664,N_15632);
nor U20153 (N_20153,N_16137,N_19625);
or U20154 (N_20154,N_18676,N_17127);
nand U20155 (N_20155,N_17189,N_19729);
and U20156 (N_20156,N_17802,N_16945);
or U20157 (N_20157,N_16743,N_19644);
or U20158 (N_20158,N_15572,N_16125);
nor U20159 (N_20159,N_15177,N_15964);
nor U20160 (N_20160,N_17956,N_18769);
nand U20161 (N_20161,N_18513,N_16334);
or U20162 (N_20162,N_15600,N_17292);
nand U20163 (N_20163,N_18732,N_19521);
nand U20164 (N_20164,N_16859,N_18745);
nand U20165 (N_20165,N_15654,N_16310);
and U20166 (N_20166,N_16455,N_19528);
nand U20167 (N_20167,N_16002,N_15219);
or U20168 (N_20168,N_19603,N_18833);
nand U20169 (N_20169,N_19498,N_15960);
nor U20170 (N_20170,N_16387,N_18402);
nor U20171 (N_20171,N_16431,N_16653);
and U20172 (N_20172,N_19432,N_17003);
or U20173 (N_20173,N_17606,N_16306);
nand U20174 (N_20174,N_19001,N_17633);
nand U20175 (N_20175,N_16021,N_19801);
nor U20176 (N_20176,N_15906,N_19796);
nor U20177 (N_20177,N_15578,N_15267);
and U20178 (N_20178,N_17474,N_16572);
nor U20179 (N_20179,N_19331,N_17350);
or U20180 (N_20180,N_15175,N_18061);
and U20181 (N_20181,N_15208,N_17417);
and U20182 (N_20182,N_18801,N_16606);
or U20183 (N_20183,N_15557,N_18896);
nand U20184 (N_20184,N_16007,N_16703);
and U20185 (N_20185,N_17506,N_15640);
and U20186 (N_20186,N_19724,N_18195);
and U20187 (N_20187,N_18950,N_15148);
xnor U20188 (N_20188,N_17149,N_19995);
nor U20189 (N_20189,N_17362,N_18685);
or U20190 (N_20190,N_16201,N_18078);
nor U20191 (N_20191,N_17746,N_18561);
nand U20192 (N_20192,N_17677,N_19375);
and U20193 (N_20193,N_16827,N_19396);
nor U20194 (N_20194,N_15366,N_17211);
and U20195 (N_20195,N_19689,N_15593);
and U20196 (N_20196,N_15069,N_15333);
or U20197 (N_20197,N_16824,N_18799);
nand U20198 (N_20198,N_19456,N_17557);
nor U20199 (N_20199,N_19089,N_16599);
nor U20200 (N_20200,N_16062,N_17158);
nor U20201 (N_20201,N_15723,N_17715);
and U20202 (N_20202,N_16401,N_18670);
or U20203 (N_20203,N_17285,N_15133);
or U20204 (N_20204,N_16373,N_15841);
xnor U20205 (N_20205,N_15276,N_19848);
or U20206 (N_20206,N_17768,N_17094);
nor U20207 (N_20207,N_16803,N_16332);
and U20208 (N_20208,N_18604,N_19244);
nand U20209 (N_20209,N_17559,N_19836);
and U20210 (N_20210,N_19018,N_15245);
and U20211 (N_20211,N_16623,N_17390);
nor U20212 (N_20212,N_17237,N_17229);
nand U20213 (N_20213,N_19981,N_19570);
nand U20214 (N_20214,N_18678,N_17170);
xor U20215 (N_20215,N_17296,N_15081);
nand U20216 (N_20216,N_18708,N_15565);
and U20217 (N_20217,N_19136,N_16793);
nand U20218 (N_20218,N_18996,N_15022);
and U20219 (N_20219,N_15695,N_15834);
nand U20220 (N_20220,N_18568,N_18642);
nor U20221 (N_20221,N_19318,N_19906);
nand U20222 (N_20222,N_16908,N_19262);
and U20223 (N_20223,N_17886,N_16503);
or U20224 (N_20224,N_16544,N_15298);
nand U20225 (N_20225,N_18264,N_17828);
or U20226 (N_20226,N_15988,N_19355);
nor U20227 (N_20227,N_18305,N_18461);
or U20228 (N_20228,N_16414,N_17622);
xnor U20229 (N_20229,N_16094,N_17632);
nand U20230 (N_20230,N_19543,N_18973);
and U20231 (N_20231,N_15226,N_18393);
nand U20232 (N_20232,N_16640,N_19260);
or U20233 (N_20233,N_19564,N_18562);
nand U20234 (N_20234,N_16751,N_19594);
nor U20235 (N_20235,N_17105,N_17772);
and U20236 (N_20236,N_18449,N_16822);
and U20237 (N_20237,N_18834,N_19364);
nor U20238 (N_20238,N_19562,N_19243);
or U20239 (N_20239,N_15409,N_18533);
xor U20240 (N_20240,N_16081,N_16103);
nor U20241 (N_20241,N_18948,N_16212);
nor U20242 (N_20242,N_18653,N_18376);
xor U20243 (N_20243,N_16673,N_18677);
or U20244 (N_20244,N_15437,N_15113);
nand U20245 (N_20245,N_15387,N_15580);
nor U20246 (N_20246,N_15271,N_19602);
nand U20247 (N_20247,N_18238,N_18060);
or U20248 (N_20248,N_19908,N_17549);
nand U20249 (N_20249,N_16355,N_19037);
nand U20250 (N_20250,N_18754,N_15537);
nand U20251 (N_20251,N_18185,N_15531);
nand U20252 (N_20252,N_17979,N_15252);
and U20253 (N_20253,N_15195,N_17311);
nor U20254 (N_20254,N_17752,N_15495);
nor U20255 (N_20255,N_17716,N_18995);
nand U20256 (N_20256,N_16067,N_16183);
nor U20257 (N_20257,N_15173,N_16821);
nand U20258 (N_20258,N_17890,N_18468);
nand U20259 (N_20259,N_15240,N_19670);
nand U20260 (N_20260,N_16816,N_15518);
and U20261 (N_20261,N_19042,N_17460);
and U20262 (N_20262,N_16319,N_15273);
and U20263 (N_20263,N_18155,N_19301);
and U20264 (N_20264,N_18050,N_15452);
nor U20265 (N_20265,N_15131,N_16744);
nor U20266 (N_20266,N_19783,N_17751);
nor U20267 (N_20267,N_19159,N_16992);
nor U20268 (N_20268,N_18086,N_18332);
nand U20269 (N_20269,N_18974,N_17861);
and U20270 (N_20270,N_17883,N_17352);
and U20271 (N_20271,N_19354,N_18913);
or U20272 (N_20272,N_17736,N_16469);
and U20273 (N_20273,N_16168,N_19210);
nor U20274 (N_20274,N_17592,N_17353);
or U20275 (N_20275,N_19366,N_17398);
xnor U20276 (N_20276,N_17396,N_19288);
or U20277 (N_20277,N_18981,N_18550);
or U20278 (N_20278,N_18146,N_15303);
and U20279 (N_20279,N_18997,N_17190);
nor U20280 (N_20280,N_17975,N_15752);
nor U20281 (N_20281,N_15386,N_18720);
nor U20282 (N_20282,N_17550,N_17041);
and U20283 (N_20283,N_16080,N_19764);
nor U20284 (N_20284,N_16295,N_18970);
nand U20285 (N_20285,N_17790,N_15205);
xnor U20286 (N_20286,N_16029,N_19511);
nand U20287 (N_20287,N_19807,N_17383);
xor U20288 (N_20288,N_18093,N_19868);
and U20289 (N_20289,N_17998,N_18647);
or U20290 (N_20290,N_19891,N_16485);
nand U20291 (N_20291,N_15522,N_15957);
or U20292 (N_20292,N_18897,N_16318);
and U20293 (N_20293,N_17274,N_17899);
or U20294 (N_20294,N_18496,N_17496);
nor U20295 (N_20295,N_18277,N_16126);
xnor U20296 (N_20296,N_16186,N_16281);
and U20297 (N_20297,N_18139,N_16441);
nand U20298 (N_20298,N_16985,N_19907);
and U20299 (N_20299,N_18457,N_18035);
or U20300 (N_20300,N_17574,N_18875);
nor U20301 (N_20301,N_18289,N_17160);
xnor U20302 (N_20302,N_17737,N_19381);
nor U20303 (N_20303,N_16085,N_15706);
nand U20304 (N_20304,N_16669,N_18303);
nor U20305 (N_20305,N_16388,N_15086);
or U20306 (N_20306,N_18447,N_17679);
or U20307 (N_20307,N_17970,N_15281);
and U20308 (N_20308,N_19916,N_19654);
and U20309 (N_20309,N_17321,N_17960);
and U20310 (N_20310,N_18115,N_19416);
or U20311 (N_20311,N_17222,N_16952);
nand U20312 (N_20312,N_19736,N_15662);
nand U20313 (N_20313,N_16051,N_17056);
nor U20314 (N_20314,N_19255,N_15032);
or U20315 (N_20315,N_18083,N_19338);
nor U20316 (N_20316,N_15744,N_17940);
nor U20317 (N_20317,N_15756,N_16475);
nand U20318 (N_20318,N_19424,N_17984);
nand U20319 (N_20319,N_19769,N_18490);
or U20320 (N_20320,N_17136,N_15652);
and U20321 (N_20321,N_17604,N_16548);
nor U20322 (N_20322,N_17258,N_19889);
and U20323 (N_20323,N_19675,N_16501);
xor U20324 (N_20324,N_18193,N_16439);
or U20325 (N_20325,N_19153,N_15064);
or U20326 (N_20326,N_16601,N_17084);
nor U20327 (N_20327,N_17010,N_15944);
xnor U20328 (N_20328,N_16275,N_16003);
nand U20329 (N_20329,N_15448,N_19558);
nor U20330 (N_20330,N_16273,N_19871);
nor U20331 (N_20331,N_19083,N_18858);
nand U20332 (N_20332,N_18586,N_17878);
and U20333 (N_20333,N_19943,N_17262);
nor U20334 (N_20334,N_19403,N_16289);
xor U20335 (N_20335,N_15581,N_15855);
nand U20336 (N_20336,N_18505,N_18437);
and U20337 (N_20337,N_18523,N_18222);
nor U20338 (N_20338,N_19325,N_15806);
or U20339 (N_20339,N_17185,N_16156);
xor U20340 (N_20340,N_17335,N_16780);
nand U20341 (N_20341,N_18181,N_18752);
or U20342 (N_20342,N_16586,N_17071);
nor U20343 (N_20343,N_17401,N_19428);
nand U20344 (N_20344,N_18165,N_16643);
and U20345 (N_20345,N_19830,N_17188);
nor U20346 (N_20346,N_18326,N_18508);
or U20347 (N_20347,N_16860,N_19990);
xor U20348 (N_20348,N_15485,N_17697);
nor U20349 (N_20349,N_17570,N_17836);
and U20350 (N_20350,N_18502,N_17405);
and U20351 (N_20351,N_16869,N_19296);
nand U20352 (N_20352,N_18282,N_18389);
and U20353 (N_20353,N_15543,N_17114);
or U20354 (N_20354,N_15021,N_15324);
nor U20355 (N_20355,N_16700,N_16943);
nor U20356 (N_20356,N_15176,N_15994);
nor U20357 (N_20357,N_18483,N_18386);
xnor U20358 (N_20358,N_17938,N_19046);
nand U20359 (N_20359,N_19593,N_16795);
nand U20360 (N_20360,N_15292,N_16340);
or U20361 (N_20361,N_19953,N_19883);
nand U20362 (N_20362,N_16106,N_15122);
nor U20363 (N_20363,N_15685,N_15555);
or U20364 (N_20364,N_19169,N_15521);
xor U20365 (N_20365,N_16757,N_18709);
and U20366 (N_20366,N_16797,N_18549);
or U20367 (N_20367,N_18293,N_17742);
nand U20368 (N_20368,N_15611,N_18401);
nor U20369 (N_20369,N_15152,N_19931);
and U20370 (N_20370,N_16786,N_17850);
or U20371 (N_20371,N_18074,N_16684);
and U20372 (N_20372,N_17007,N_19004);
nor U20373 (N_20373,N_18956,N_19006);
or U20374 (N_20374,N_17186,N_18879);
xor U20375 (N_20375,N_19612,N_16424);
xnor U20376 (N_20376,N_15373,N_19909);
xor U20377 (N_20377,N_16818,N_19853);
nor U20378 (N_20378,N_15732,N_17430);
or U20379 (N_20379,N_19865,N_15038);
and U20380 (N_20380,N_18863,N_17636);
or U20381 (N_20381,N_17767,N_19532);
and U20382 (N_20382,N_19888,N_19849);
and U20383 (N_20383,N_19487,N_19024);
and U20384 (N_20384,N_18899,N_17786);
nor U20385 (N_20385,N_15034,N_17272);
nor U20386 (N_20386,N_19266,N_18721);
and U20387 (N_20387,N_19267,N_19328);
xnor U20388 (N_20388,N_17647,N_16846);
nand U20389 (N_20389,N_18605,N_15181);
or U20390 (N_20390,N_15345,N_18664);
nor U20391 (N_20391,N_15105,N_15026);
or U20392 (N_20392,N_19440,N_18592);
nand U20393 (N_20393,N_19845,N_19220);
or U20394 (N_20394,N_18894,N_19125);
nand U20395 (N_20395,N_16864,N_17286);
nand U20396 (N_20396,N_19884,N_18761);
nor U20397 (N_20397,N_15633,N_15954);
and U20398 (N_20398,N_16668,N_17470);
and U20399 (N_20399,N_19559,N_16365);
and U20400 (N_20400,N_17031,N_17200);
nand U20401 (N_20401,N_17051,N_17851);
and U20402 (N_20402,N_19439,N_16268);
nor U20403 (N_20403,N_17968,N_15714);
and U20404 (N_20404,N_18104,N_19207);
nor U20405 (N_20405,N_19582,N_15953);
nor U20406 (N_20406,N_19182,N_18785);
and U20407 (N_20407,N_15673,N_16050);
xnor U20408 (N_20408,N_19921,N_18444);
xnor U20409 (N_20409,N_18972,N_17387);
and U20410 (N_20410,N_15943,N_19007);
nand U20411 (N_20411,N_16769,N_18110);
xor U20412 (N_20412,N_19516,N_18022);
and U20413 (N_20413,N_18740,N_15214);
or U20414 (N_20414,N_19838,N_19402);
or U20415 (N_20415,N_18780,N_16981);
and U20416 (N_20416,N_19344,N_19641);
xor U20417 (N_20417,N_17301,N_15802);
nor U20418 (N_20418,N_16874,N_15489);
xor U20419 (N_20419,N_16852,N_18425);
and U20420 (N_20420,N_16873,N_18691);
nand U20421 (N_20421,N_18254,N_18633);
and U20422 (N_20422,N_16921,N_16069);
nor U20423 (N_20423,N_15655,N_18111);
or U20424 (N_20424,N_15566,N_16899);
xor U20425 (N_20425,N_19467,N_19275);
nand U20426 (N_20426,N_16986,N_16603);
or U20427 (N_20427,N_15102,N_19055);
nand U20428 (N_20428,N_18407,N_18667);
nor U20429 (N_20429,N_16492,N_16124);
nand U20430 (N_20430,N_16542,N_17937);
or U20431 (N_20431,N_17512,N_17244);
and U20432 (N_20432,N_16031,N_17718);
nor U20433 (N_20433,N_17175,N_18900);
or U20434 (N_20434,N_19787,N_19158);
nor U20435 (N_20435,N_17923,N_17782);
and U20436 (N_20436,N_18924,N_16882);
or U20437 (N_20437,N_17816,N_18126);
or U20438 (N_20438,N_18025,N_17214);
nand U20439 (N_20439,N_18395,N_17844);
or U20440 (N_20440,N_15337,N_15962);
and U20441 (N_20441,N_19134,N_18787);
nor U20442 (N_20442,N_17120,N_15264);
and U20443 (N_20443,N_17670,N_18499);
and U20444 (N_20444,N_15427,N_16393);
nand U20445 (N_20445,N_19754,N_15742);
nand U20446 (N_20446,N_19445,N_18696);
nand U20447 (N_20447,N_18756,N_15999);
or U20448 (N_20448,N_18335,N_18703);
and U20449 (N_20449,N_16975,N_17825);
xor U20450 (N_20450,N_17278,N_16678);
and U20451 (N_20451,N_16733,N_15046);
nor U20452 (N_20452,N_19666,N_16105);
nand U20453 (N_20453,N_17226,N_18419);
and U20454 (N_20454,N_17065,N_17279);
xor U20455 (N_20455,N_19099,N_15143);
or U20456 (N_20456,N_17325,N_16670);
nor U20457 (N_20457,N_19144,N_18689);
nand U20458 (N_20458,N_16907,N_16457);
or U20459 (N_20459,N_18250,N_18882);
and U20460 (N_20460,N_17391,N_18228);
nand U20461 (N_20461,N_17011,N_17762);
nand U20462 (N_20462,N_16160,N_19130);
nor U20463 (N_20463,N_17174,N_16887);
nand U20464 (N_20464,N_17681,N_19930);
xnor U20465 (N_20465,N_15827,N_15586);
nand U20466 (N_20466,N_16375,N_16174);
nand U20467 (N_20467,N_15776,N_18351);
xnor U20468 (N_20468,N_19237,N_15865);
nand U20469 (N_20469,N_19829,N_16432);
or U20470 (N_20470,N_15391,N_18224);
or U20471 (N_20471,N_18192,N_15426);
nand U20472 (N_20472,N_16395,N_18959);
and U20473 (N_20473,N_17038,N_15220);
nor U20474 (N_20474,N_17607,N_17465);
nand U20475 (N_20475,N_16913,N_18920);
and U20476 (N_20476,N_17564,N_16785);
or U20477 (N_20477,N_16876,N_17173);
nand U20478 (N_20478,N_15359,N_17263);
xnor U20479 (N_20479,N_15025,N_19098);
and U20480 (N_20480,N_15615,N_15383);
nor U20481 (N_20481,N_17449,N_18722);
nor U20482 (N_20482,N_16596,N_16088);
nor U20483 (N_20483,N_17515,N_17004);
and U20484 (N_20484,N_18966,N_16301);
nand U20485 (N_20485,N_18422,N_17819);
and U20486 (N_20486,N_18458,N_15526);
and U20487 (N_20487,N_17522,N_19026);
or U20488 (N_20488,N_19681,N_19234);
nor U20489 (N_20489,N_18861,N_18693);
or U20490 (N_20490,N_16686,N_18280);
xor U20491 (N_20491,N_18044,N_18229);
xor U20492 (N_20492,N_17658,N_17760);
or U20493 (N_20493,N_17872,N_19753);
nor U20494 (N_20494,N_16178,N_17823);
nor U20495 (N_20495,N_17714,N_15151);
or U20496 (N_20496,N_15733,N_17894);
and U20497 (N_20497,N_18257,N_17088);
and U20498 (N_20498,N_15326,N_15936);
xnor U20499 (N_20499,N_17478,N_18311);
and U20500 (N_20500,N_17623,N_16072);
xor U20501 (N_20501,N_15784,N_17324);
and U20502 (N_20502,N_19546,N_18725);
nand U20503 (N_20503,N_16920,N_17077);
or U20504 (N_20504,N_19073,N_15482);
nand U20505 (N_20505,N_15316,N_18715);
or U20506 (N_20506,N_18424,N_19306);
nand U20507 (N_20507,N_19745,N_17845);
xor U20508 (N_20508,N_16796,N_17566);
nor U20509 (N_20509,N_18128,N_17554);
nand U20510 (N_20510,N_18649,N_17734);
and U20511 (N_20511,N_15307,N_17193);
and U20512 (N_20512,N_15552,N_18453);
or U20513 (N_20513,N_17409,N_15302);
xnor U20514 (N_20514,N_16041,N_15509);
and U20515 (N_20515,N_15828,N_18251);
or U20516 (N_20516,N_19137,N_19706);
nand U20517 (N_20517,N_15523,N_17349);
and U20518 (N_20518,N_15335,N_18344);
or U20519 (N_20519,N_18454,N_17447);
and U20520 (N_20520,N_18770,N_18072);
xor U20521 (N_20521,N_19837,N_19705);
and U20522 (N_20522,N_15486,N_19287);
nand U20523 (N_20523,N_15475,N_17122);
nand U20524 (N_20524,N_19910,N_18153);
nand U20525 (N_20525,N_18501,N_18608);
nor U20526 (N_20526,N_16136,N_18829);
nor U20527 (N_20527,N_18797,N_19143);
nand U20528 (N_20528,N_18176,N_19541);
nor U20529 (N_20529,N_15560,N_16690);
and U20530 (N_20530,N_18609,N_16006);
and U20531 (N_20531,N_19751,N_18047);
nor U20532 (N_20532,N_19514,N_19828);
nand U20533 (N_20533,N_18356,N_15450);
nand U20534 (N_20534,N_15182,N_18382);
or U20535 (N_20535,N_19423,N_16988);
or U20536 (N_20536,N_17686,N_17925);
and U20537 (N_20537,N_17139,N_18982);
nor U20538 (N_20538,N_17799,N_16834);
or U20539 (N_20539,N_16181,N_18004);
nand U20540 (N_20540,N_17131,N_16237);
nor U20541 (N_20541,N_15727,N_18706);
or U20542 (N_20542,N_18704,N_17129);
nand U20543 (N_20543,N_19536,N_19460);
and U20544 (N_20544,N_16253,N_15539);
or U20545 (N_20545,N_18320,N_18075);
or U20546 (N_20546,N_17360,N_15384);
and U20547 (N_20547,N_17513,N_19506);
nand U20548 (N_20548,N_19999,N_16947);
or U20549 (N_20549,N_17420,N_17896);
xnor U20550 (N_20550,N_19864,N_15494);
and U20551 (N_20551,N_17903,N_17249);
xnor U20552 (N_20552,N_18987,N_15099);
nand U20553 (N_20553,N_17521,N_18838);
and U20554 (N_20554,N_17112,N_15288);
nand U20555 (N_20555,N_19488,N_19619);
nor U20556 (N_20556,N_18641,N_18934);
or U20557 (N_20557,N_18593,N_15382);
xnor U20558 (N_20558,N_16294,N_15885);
nor U20559 (N_20559,N_18921,N_15179);
nand U20560 (N_20560,N_18548,N_17921);
or U20561 (N_20561,N_18852,N_15389);
or U20562 (N_20562,N_19554,N_18324);
nand U20563 (N_20563,N_16931,N_19474);
xnor U20564 (N_20564,N_16598,N_17858);
or U20565 (N_20565,N_15136,N_15441);
or U20566 (N_20566,N_19459,N_18576);
nand U20567 (N_20567,N_17057,N_16725);
nor U20568 (N_20568,N_16256,N_19606);
or U20569 (N_20569,N_17250,N_19785);
or U20570 (N_20570,N_15544,N_17066);
or U20571 (N_20571,N_15434,N_16791);
or U20572 (N_20572,N_19567,N_18017);
or U20573 (N_20573,N_17744,N_17708);
or U20574 (N_20574,N_17345,N_19223);
or U20575 (N_20575,N_16957,N_17377);
nand U20576 (N_20576,N_15846,N_15689);
and U20577 (N_20577,N_17797,N_19175);
and U20578 (N_20578,N_15582,N_18162);
or U20579 (N_20579,N_17466,N_17880);
nor U20580 (N_20580,N_18269,N_16070);
nor U20581 (N_20581,N_18810,N_15757);
nand U20582 (N_20582,N_15870,N_15183);
nand U20583 (N_20583,N_19683,N_19963);
nor U20584 (N_20584,N_19304,N_19072);
nor U20585 (N_20585,N_17024,N_18711);
nand U20586 (N_20586,N_18825,N_17240);
nor U20587 (N_20587,N_15919,N_18065);
nor U20588 (N_20588,N_18610,N_18002);
and U20589 (N_20589,N_15913,N_16098);
nand U20590 (N_20590,N_18476,N_19154);
and U20591 (N_20591,N_17600,N_16498);
nand U20592 (N_20592,N_17093,N_18329);
or U20593 (N_20593,N_19697,N_16090);
nand U20594 (N_20594,N_18849,N_19116);
or U20595 (N_20595,N_15212,N_19561);
xor U20596 (N_20596,N_18355,N_16650);
and U20597 (N_20597,N_16154,N_17358);
nor U20598 (N_20598,N_18767,N_15146);
nor U20599 (N_20599,N_19240,N_16651);
or U20600 (N_20600,N_18178,N_18300);
or U20601 (N_20601,N_19998,N_15156);
nand U20602 (N_20602,N_19942,N_17817);
and U20603 (N_20603,N_17558,N_18308);
and U20604 (N_20604,N_18125,N_16843);
and U20605 (N_20605,N_16454,N_16418);
or U20606 (N_20606,N_18509,N_17609);
nand U20607 (N_20607,N_19509,N_16428);
nor U20608 (N_20608,N_15660,N_18544);
and U20609 (N_20609,N_15818,N_18137);
and U20610 (N_20610,N_17505,N_17110);
or U20611 (N_20611,N_16159,N_19194);
xor U20612 (N_20612,N_17910,N_15262);
or U20613 (N_20613,N_15844,N_16604);
and U20614 (N_20614,N_16883,N_19455);
and U20615 (N_20615,N_15638,N_15251);
nand U20616 (N_20616,N_16100,N_19412);
and U20617 (N_20617,N_19927,N_16035);
and U20618 (N_20618,N_16267,N_16587);
or U20619 (N_20619,N_17688,N_17882);
xor U20620 (N_20620,N_19452,N_17168);
xnor U20621 (N_20621,N_18431,N_16292);
and U20622 (N_20622,N_17841,N_16694);
or U20623 (N_20623,N_16463,N_17997);
nor U20624 (N_20624,N_15416,N_16073);
or U20625 (N_20625,N_18698,N_19700);
or U20626 (N_20626,N_16025,N_16642);
or U20627 (N_20627,N_16037,N_16513);
xor U20628 (N_20628,N_15829,N_18485);
or U20629 (N_20629,N_15569,N_18478);
and U20630 (N_20630,N_18854,N_16896);
xnor U20631 (N_20631,N_16551,N_19851);
xnor U20632 (N_20632,N_15369,N_19507);
nor U20633 (N_20633,N_16634,N_17354);
and U20634 (N_20634,N_16406,N_15420);
nor U20635 (N_20635,N_17154,N_17276);
or U20636 (N_20636,N_15339,N_17412);
nor U20637 (N_20637,N_16014,N_19350);
xnor U20638 (N_20638,N_18353,N_18926);
nand U20639 (N_20639,N_16577,N_17419);
nand U20640 (N_20640,N_17640,N_19367);
and U20641 (N_20641,N_16442,N_19189);
and U20642 (N_20642,N_18258,N_16430);
nor U20643 (N_20643,N_16143,N_15741);
nor U20644 (N_20644,N_19174,N_17853);
nor U20645 (N_20645,N_15104,N_18152);
or U20646 (N_20646,N_16429,N_17794);
nor U20647 (N_20647,N_17012,N_15728);
and U20648 (N_20648,N_15990,N_15656);
and U20649 (N_20649,N_16120,N_18656);
or U20650 (N_20650,N_16345,N_16749);
or U20651 (N_20651,N_18119,N_19302);
and U20652 (N_20652,N_19515,N_19221);
nand U20653 (N_20653,N_19816,N_16089);
xnor U20654 (N_20654,N_19274,N_18188);
and U20655 (N_20655,N_18723,N_18570);
or U20656 (N_20656,N_18716,N_19788);
nand U20657 (N_20657,N_18650,N_17869);
and U20658 (N_20658,N_19336,N_19826);
nor U20659 (N_20659,N_16713,N_18954);
nor U20660 (N_20660,N_15472,N_15950);
nor U20661 (N_20661,N_18039,N_17017);
or U20662 (N_20662,N_17133,N_15896);
or U20663 (N_20663,N_19896,N_17348);
nor U20664 (N_20664,N_18739,N_18038);
nor U20665 (N_20665,N_15467,N_17556);
or U20666 (N_20666,N_17508,N_19822);
and U20667 (N_20667,N_15556,N_16104);
or U20668 (N_20668,N_15037,N_17180);
xnor U20669 (N_20669,N_15598,N_18179);
nand U20670 (N_20670,N_17520,N_16760);
nand U20671 (N_20671,N_15202,N_17150);
xnor U20672 (N_20672,N_15406,N_17494);
or U20673 (N_20673,N_16052,N_16842);
xor U20674 (N_20674,N_17643,N_16265);
nor U20675 (N_20675,N_18871,N_18901);
and U20676 (N_20676,N_17781,N_17818);
nand U20677 (N_20677,N_17308,N_18287);
or U20678 (N_20678,N_17411,N_16930);
nand U20679 (N_20679,N_17873,N_17192);
or U20680 (N_20680,N_16767,N_17924);
nor U20681 (N_20681,N_15681,N_19155);
xnor U20682 (N_20682,N_18775,N_16830);
and U20683 (N_20683,N_18412,N_16674);
and U20684 (N_20684,N_19172,N_19285);
or U20685 (N_20685,N_15862,N_15825);
nor U20686 (N_20686,N_17072,N_16644);
and U20687 (N_20687,N_18015,N_18821);
nor U20688 (N_20688,N_15998,N_16529);
or U20689 (N_20689,N_17394,N_18631);
and U20690 (N_20690,N_18132,N_19721);
or U20691 (N_20691,N_18687,N_17182);
nor U20692 (N_20692,N_16854,N_18199);
nor U20693 (N_20693,N_15395,N_15431);
nor U20694 (N_20694,N_17062,N_17699);
xor U20695 (N_20695,N_17711,N_15207);
nor U20696 (N_20696,N_17934,N_18191);
and U20697 (N_20697,N_17462,N_17680);
nand U20698 (N_20698,N_15055,N_18077);
or U20699 (N_20699,N_15045,N_19264);
nand U20700 (N_20700,N_15294,N_15350);
or U20701 (N_20701,N_19679,N_16494);
nand U20702 (N_20702,N_17108,N_17141);
and U20703 (N_20703,N_18348,N_18585);
nor U20704 (N_20704,N_17008,N_16527);
and U20705 (N_20705,N_16624,N_18611);
and U20706 (N_20706,N_15261,N_18338);
nand U20707 (N_20707,N_16379,N_19349);
or U20708 (N_20708,N_15746,N_16940);
nor U20709 (N_20709,N_17236,N_19298);
nor U20710 (N_20710,N_18366,N_18688);
or U20711 (N_20711,N_15328,N_16157);
and U20712 (N_20712,N_17510,N_16766);
or U20713 (N_20713,N_15782,N_18594);
nor U20714 (N_20714,N_17376,N_15670);
nand U20715 (N_20715,N_17271,N_16139);
nand U20716 (N_20716,N_18657,N_18963);
nand U20717 (N_20717,N_16480,N_17207);
xnor U20718 (N_20718,N_17741,N_18521);
nor U20719 (N_20719,N_16914,N_17895);
and U20720 (N_20720,N_16433,N_15368);
nand U20721 (N_20721,N_15203,N_15401);
or U20722 (N_20722,N_15348,N_17831);
nand U20723 (N_20723,N_18532,N_17963);
nand U20724 (N_20724,N_15044,N_19530);
or U20725 (N_20725,N_18406,N_18314);
nand U20726 (N_20726,N_19672,N_18885);
and U20727 (N_20727,N_16191,N_19087);
nor U20728 (N_20728,N_17611,N_19245);
and U20729 (N_20729,N_17864,N_19229);
nor U20730 (N_20730,N_16851,N_19053);
nand U20731 (N_20731,N_16337,N_17871);
nor U20732 (N_20732,N_16974,N_16728);
xor U20733 (N_20733,N_15891,N_18213);
xnor U20734 (N_20734,N_15097,N_16969);
xnor U20735 (N_20735,N_19772,N_17381);
nor U20736 (N_20736,N_18547,N_15772);
and U20737 (N_20737,N_17364,N_19741);
and U20738 (N_20738,N_16723,N_19086);
nand U20739 (N_20739,N_17665,N_17148);
nor U20740 (N_20740,N_15650,N_15805);
nand U20741 (N_20741,N_15137,N_15935);
nor U20742 (N_20742,N_17602,N_15464);
nor U20743 (N_20743,N_15649,N_15473);
and U20744 (N_20744,N_16382,N_18985);
or U20745 (N_20745,N_18232,N_15667);
or U20746 (N_20746,N_19627,N_16708);
or U20747 (N_20747,N_19595,N_19370);
nand U20748 (N_20748,N_19188,N_19231);
nor U20749 (N_20749,N_15738,N_19263);
and U20750 (N_20750,N_17913,N_18734);
nand U20751 (N_20751,N_16384,N_18612);
and U20752 (N_20752,N_18742,N_17594);
and U20753 (N_20753,N_16176,N_15200);
nor U20754 (N_20754,N_17442,N_16667);
nand U20755 (N_20755,N_17785,N_15669);
nor U20756 (N_20756,N_15213,N_15374);
or U20757 (N_20757,N_15947,N_17109);
nand U20758 (N_20758,N_16192,N_19002);
and U20759 (N_20759,N_17993,N_16942);
nand U20760 (N_20760,N_18219,N_17261);
xor U20761 (N_20761,N_15106,N_16108);
nor U20762 (N_20762,N_19185,N_19841);
xor U20763 (N_20763,N_17724,N_18815);
xnor U20764 (N_20764,N_19710,N_17743);
nand U20765 (N_20765,N_15506,N_16066);
nor U20766 (N_20766,N_17631,N_19357);
xnor U20767 (N_20767,N_15436,N_15166);
nor U20768 (N_20768,N_17827,N_18860);
xnor U20769 (N_20769,N_18559,N_17656);
nor U20770 (N_20770,N_15643,N_18665);
nor U20771 (N_20771,N_18971,N_17761);
nor U20772 (N_20772,N_15070,N_16397);
nor U20773 (N_20773,N_15894,N_15561);
or U20774 (N_20774,N_15004,N_19734);
and U20775 (N_20775,N_17455,N_16368);
or U20776 (N_20776,N_17932,N_17701);
or U20777 (N_20777,N_16520,N_16217);
and U20778 (N_20778,N_18470,N_16812);
nand U20779 (N_20779,N_18962,N_16950);
nor U20780 (N_20780,N_16517,N_19310);
or U20781 (N_20781,N_16436,N_19997);
nor U20782 (N_20782,N_17952,N_17317);
nand U20783 (N_20783,N_16016,N_18563);
or U20784 (N_20784,N_19794,N_18522);
and U20785 (N_20785,N_18405,N_17342);
nor U20786 (N_20786,N_18823,N_16288);
or U20787 (N_20787,N_15254,N_18855);
and U20788 (N_20788,N_19166,N_18053);
or U20789 (N_20789,N_18518,N_19108);
nand U20790 (N_20790,N_18263,N_17162);
and U20791 (N_20791,N_16250,N_16411);
or U20792 (N_20792,N_15610,N_18262);
nand U20793 (N_20793,N_16980,N_16568);
nor U20794 (N_20794,N_15597,N_15979);
nand U20795 (N_20795,N_19352,N_19805);
nor U20796 (N_20796,N_16496,N_17338);
nor U20797 (N_20797,N_17804,N_19353);
xor U20798 (N_20798,N_17463,N_16440);
or U20799 (N_20799,N_17941,N_15289);
nor U20800 (N_20800,N_15992,N_15909);
nand U20801 (N_20801,N_15729,N_19472);
nor U20802 (N_20802,N_16302,N_17936);
xnor U20803 (N_20803,N_15229,N_19315);
or U20804 (N_20804,N_17225,N_18990);
xor U20805 (N_20805,N_17598,N_15807);
or U20806 (N_20806,N_17595,N_16801);
or U20807 (N_20807,N_16438,N_16792);
nor U20808 (N_20808,N_19230,N_17204);
or U20809 (N_20809,N_18931,N_19571);
or U20810 (N_20810,N_15164,N_18961);
xnor U20811 (N_20811,N_18952,N_15110);
nor U20812 (N_20812,N_16755,N_18474);
or U20813 (N_20813,N_15490,N_15683);
nand U20814 (N_20814,N_15063,N_16707);
and U20815 (N_20815,N_19035,N_15821);
nand U20816 (N_20816,N_16199,N_19505);
and U20817 (N_20817,N_16077,N_19572);
nor U20818 (N_20818,N_16177,N_16515);
xor U20819 (N_20819,N_18828,N_15634);
or U20820 (N_20820,N_15300,N_17480);
or U20821 (N_20821,N_16699,N_18968);
and U20822 (N_20822,N_18655,N_19107);
or U20823 (N_20823,N_17511,N_18891);
nand U20824 (N_20824,N_16745,N_17682);
nand U20825 (N_20825,N_18878,N_16752);
and U20826 (N_20826,N_16425,N_16448);
or U20827 (N_20827,N_19598,N_16234);
and U20828 (N_20828,N_16042,N_17692);
or U20829 (N_20829,N_16677,N_16203);
xnor U20830 (N_20830,N_16367,N_19184);
nand U20831 (N_20831,N_17722,N_19762);
or U20832 (N_20832,N_19473,N_16317);
and U20833 (N_20833,N_15702,N_16180);
nand U20834 (N_20834,N_17696,N_15549);
xor U20835 (N_20835,N_16632,N_16357);
nor U20836 (N_20836,N_15647,N_18747);
and U20837 (N_20837,N_17231,N_17107);
and U20838 (N_20838,N_18743,N_18226);
nor U20839 (N_20839,N_16631,N_16190);
and U20840 (N_20840,N_19163,N_18208);
or U20841 (N_20841,N_15743,N_15959);
and U20842 (N_20842,N_15253,N_18068);
nor U20843 (N_20843,N_18928,N_17732);
and U20844 (N_20844,N_15266,N_16101);
nand U20845 (N_20845,N_15414,N_17497);
nor U20846 (N_20846,N_17571,N_15432);
nand U20847 (N_20847,N_15057,N_17982);
nand U20848 (N_20848,N_16380,N_17404);
or U20849 (N_20849,N_18297,N_16506);
and U20850 (N_20850,N_18599,N_18295);
nor U20851 (N_20851,N_19513,N_16427);
and U20852 (N_20852,N_15532,N_19329);
or U20853 (N_20853,N_17672,N_16993);
xor U20854 (N_20854,N_18373,N_15816);
and U20855 (N_20855,N_15653,N_19041);
nand U20856 (N_20856,N_18826,N_18345);
and U20857 (N_20857,N_19991,N_19012);
or U20858 (N_20858,N_19434,N_17034);
nand U20859 (N_20859,N_15792,N_19191);
nand U20860 (N_20860,N_19579,N_15376);
or U20861 (N_20861,N_18148,N_18492);
nand U20862 (N_20862,N_18883,N_17740);
or U20863 (N_20863,N_15487,N_17955);
or U20864 (N_20864,N_18992,N_18957);
and U20865 (N_20865,N_16112,N_18000);
or U20866 (N_20866,N_18575,N_16839);
xnor U20867 (N_20867,N_15832,N_17403);
and U20868 (N_20868,N_15354,N_19911);
and U20869 (N_20869,N_18283,N_15849);
nor U20870 (N_20870,N_19248,N_19454);
or U20871 (N_20871,N_17617,N_19628);
or U20872 (N_20872,N_16955,N_17908);
or U20873 (N_20873,N_18753,N_18041);
or U20874 (N_20874,N_16279,N_19956);
nand U20875 (N_20875,N_19339,N_16394);
nand U20876 (N_20876,N_18542,N_16679);
nand U20877 (N_20877,N_16998,N_18019);
and U20878 (N_20878,N_15028,N_17290);
or U20879 (N_20879,N_15768,N_18674);
nand U20880 (N_20880,N_16774,N_19321);
or U20881 (N_20881,N_19045,N_15939);
nand U20882 (N_20882,N_19170,N_16584);
and U20883 (N_20883,N_16731,N_18462);
nor U20884 (N_20884,N_16398,N_15684);
nand U20885 (N_20885,N_19899,N_19015);
nor U20886 (N_20886,N_18958,N_18321);
and U20887 (N_20887,N_19996,N_19925);
or U20888 (N_20888,N_17833,N_17319);
nand U20889 (N_20889,N_15758,N_15621);
nor U20890 (N_20890,N_17916,N_19960);
nand U20891 (N_20891,N_17329,N_15478);
or U20892 (N_20892,N_15901,N_16471);
or U20893 (N_20893,N_15385,N_17177);
nor U20894 (N_20894,N_16473,N_15793);
nand U20895 (N_20895,N_19551,N_15236);
nand U20896 (N_20896,N_17651,N_15546);
or U20897 (N_20897,N_15899,N_18285);
nor U20898 (N_20898,N_15142,N_16835);
or U20899 (N_20899,N_19520,N_19250);
nand U20900 (N_20900,N_18459,N_15644);
and U20901 (N_20901,N_19019,N_15424);
nand U20902 (N_20902,N_18984,N_18031);
xnor U20903 (N_20903,N_18080,N_18095);
and U20904 (N_20904,N_16360,N_16537);
nor U20905 (N_20905,N_15759,N_16554);
or U20906 (N_20906,N_16526,N_17253);
nand U20907 (N_20907,N_17729,N_16719);
nand U20908 (N_20908,N_19613,N_16778);
nand U20909 (N_20909,N_16884,N_19660);
and U20910 (N_20910,N_18198,N_19611);
and U20911 (N_20911,N_16300,N_15974);
and U20912 (N_20912,N_19813,N_17426);
xor U20913 (N_20913,N_16350,N_18941);
or U20914 (N_20914,N_17978,N_18370);
and U20915 (N_20915,N_19695,N_17117);
nor U20916 (N_20916,N_17642,N_19299);
and U20917 (N_20917,N_17320,N_16960);
or U20918 (N_20918,N_17788,N_18136);
nand U20919 (N_20919,N_19723,N_19120);
nor U20920 (N_20920,N_19972,N_15648);
nor U20921 (N_20921,N_16343,N_15515);
nor U20922 (N_20922,N_17422,N_18755);
nor U20923 (N_20923,N_18975,N_17683);
nand U20924 (N_20924,N_17773,N_17553);
and U20925 (N_20925,N_15513,N_18565);
nand U20926 (N_20926,N_18018,N_19379);
or U20927 (N_20927,N_18052,N_18731);
nand U20928 (N_20928,N_16505,N_18571);
or U20929 (N_20929,N_15011,N_17668);
nand U20930 (N_20930,N_15837,N_18411);
xnor U20931 (N_20931,N_16514,N_19020);
xnor U20932 (N_20932,N_16567,N_19330);
nand U20933 (N_20933,N_19121,N_18045);
or U20934 (N_20934,N_15603,N_17614);
nand U20935 (N_20935,N_16452,N_16434);
nand U20936 (N_20936,N_17846,N_18777);
and U20937 (N_20937,N_19183,N_19386);
and U20938 (N_20938,N_18408,N_19726);
nor U20939 (N_20939,N_19795,N_18309);
or U20940 (N_20940,N_19010,N_18096);
and U20941 (N_20941,N_19254,N_16114);
or U20942 (N_20942,N_18781,N_16820);
nand U20943 (N_20943,N_16847,N_18372);
nor U20944 (N_20944,N_19481,N_18235);
xor U20945 (N_20945,N_16739,N_16964);
and U20946 (N_20946,N_17351,N_18400);
nor U20947 (N_20947,N_18116,N_17013);
and U20948 (N_20948,N_19043,N_18118);
xnor U20949 (N_20949,N_16499,N_16293);
or U20950 (N_20950,N_19499,N_19817);
nand U20951 (N_20951,N_19959,N_17787);
and U20952 (N_20952,N_15263,N_15422);
or U20953 (N_20953,N_18652,N_16467);
nor U20954 (N_20954,N_19623,N_17907);
and U20955 (N_20955,N_16758,N_15801);
or U20956 (N_20956,N_16676,N_17927);
nand U20957 (N_20957,N_16996,N_18583);
or U20958 (N_20958,N_15842,N_19738);
or U20959 (N_20959,N_17220,N_19270);
nor U20960 (N_20960,N_16865,N_19596);
nand U20961 (N_20961,N_18988,N_15704);
or U20962 (N_20962,N_16356,N_19502);
nor U20963 (N_20963,N_16607,N_19227);
and U20964 (N_20964,N_18794,N_16464);
and U20965 (N_20965,N_17488,N_15257);
nand U20966 (N_20966,N_15380,N_17309);
and U20967 (N_20967,N_15465,N_19633);
xor U20968 (N_20968,N_19063,N_18377);
nand U20969 (N_20969,N_15061,N_19195);
and U20970 (N_20970,N_19577,N_16582);
nand U20971 (N_20971,N_19156,N_19097);
and U20972 (N_20972,N_19265,N_15018);
xnor U20973 (N_20973,N_15559,N_15039);
nor U20974 (N_20974,N_18350,N_17482);
or U20975 (N_20975,N_17621,N_19077);
or U20976 (N_20976,N_19414,N_19662);
nand U20977 (N_20977,N_15986,N_15084);
nor U20978 (N_20978,N_18368,N_19970);
or U20979 (N_20979,N_19067,N_18079);
xnor U20980 (N_20980,N_18249,N_15428);
xnor U20981 (N_20981,N_17676,N_18955);
and U20982 (N_20982,N_15843,N_19476);
nand U20983 (N_20983,N_19206,N_15126);
nand U20984 (N_20984,N_17856,N_19969);
or U20985 (N_20985,N_15550,N_18624);
nand U20986 (N_20986,N_16346,N_19766);
or U20987 (N_20987,N_16948,N_18218);
xor U20988 (N_20988,N_19531,N_17493);
nand U20989 (N_20989,N_17375,N_19090);
and U20990 (N_20990,N_19676,N_19219);
and U20991 (N_20991,N_15810,N_18034);
nand U20992 (N_20992,N_15255,N_16923);
nor U20993 (N_20993,N_17102,N_18660);
or U20994 (N_20994,N_15360,N_15573);
nor U20995 (N_20995,N_17958,N_18629);
or U20996 (N_20996,N_15687,N_16850);
and U20997 (N_20997,N_18040,N_16770);
xnor U20998 (N_20998,N_16534,N_18069);
nor U20999 (N_20999,N_18847,N_18866);
nand U21000 (N_21000,N_19802,N_15783);
and U21001 (N_21001,N_16995,N_19197);
or U21002 (N_21002,N_16193,N_15796);
nand U21003 (N_21003,N_19610,N_19093);
nand U21004 (N_21004,N_19180,N_15547);
nor U21005 (N_21005,N_19922,N_16595);
and U21006 (N_21006,N_18201,N_16602);
or U21007 (N_21007,N_18683,N_17314);
nor U21008 (N_21008,N_18084,N_15158);
nor U21009 (N_21009,N_18489,N_19983);
and U21010 (N_21010,N_19984,N_18960);
and U21011 (N_21011,N_19588,N_18526);
and U21012 (N_21012,N_19583,N_19975);
nand U21013 (N_21013,N_19435,N_18013);
nand U21014 (N_21014,N_16965,N_15864);
nand U21015 (N_21015,N_16721,N_18186);
and U21016 (N_21016,N_18744,N_15571);
xnor U21017 (N_21017,N_19291,N_16142);
and U21018 (N_21018,N_15447,N_18848);
and U21019 (N_21019,N_19463,N_18932);
or U21020 (N_21020,N_19737,N_18134);
or U21021 (N_21021,N_15390,N_15777);
or U21022 (N_21022,N_17784,N_16158);
nor U21023 (N_21023,N_15501,N_18100);
and U21024 (N_21024,N_15278,N_19132);
nand U21025 (N_21025,N_19994,N_19091);
xnor U21026 (N_21026,N_17029,N_17060);
nand U21027 (N_21027,N_16543,N_15408);
nand U21028 (N_21028,N_17969,N_16251);
nand U21029 (N_21029,N_19141,N_19645);
xor U21030 (N_21030,N_19557,N_19784);
nand U21031 (N_21031,N_18635,N_18719);
nor U21032 (N_21032,N_16880,N_16347);
or U21033 (N_21033,N_17002,N_18600);
and U21034 (N_21034,N_18273,N_19890);
and U21035 (N_21035,N_16688,N_18671);
nor U21036 (N_21036,N_17495,N_17946);
xor U21037 (N_21037,N_17648,N_18197);
nand U21038 (N_21038,N_18042,N_17464);
nor U21039 (N_21039,N_18519,N_15162);
nand U21040 (N_21040,N_19599,N_17764);
or U21041 (N_21041,N_15795,N_15698);
xor U21042 (N_21042,N_19982,N_17930);
and U21043 (N_21043,N_15088,N_18144);
xor U21044 (N_21044,N_16221,N_18271);
xnor U21045 (N_21045,N_19814,N_15995);
nand U21046 (N_21046,N_17675,N_18233);
xnor U21047 (N_21047,N_19810,N_17499);
and U21048 (N_21048,N_16692,N_15239);
nor U21049 (N_21049,N_15312,N_15498);
or U21050 (N_21050,N_19773,N_15601);
nand U21051 (N_21051,N_18230,N_16219);
nor U21052 (N_21052,N_18940,N_16207);
nor U21053 (N_21053,N_18140,N_19952);
nand U21054 (N_21054,N_15635,N_15138);
xnor U21055 (N_21055,N_16696,N_18157);
and U21056 (N_21056,N_19578,N_19709);
nor U21057 (N_21057,N_18591,N_17906);
or U21058 (N_21058,N_17678,N_16407);
xnor U21059 (N_21059,N_17074,N_19748);
or U21060 (N_21060,N_19059,N_16063);
nor U21061 (N_21061,N_18836,N_16672);
nor U21062 (N_21062,N_16038,N_15403);
and U21063 (N_21063,N_18637,N_15558);
xor U21064 (N_21064,N_17436,N_17563);
or U21065 (N_21065,N_16550,N_15838);
nor U21066 (N_21066,N_17639,N_18816);
nand U21067 (N_21067,N_18220,N_18679);
and U21068 (N_21068,N_19324,N_19986);
nand U21069 (N_21069,N_19992,N_19651);
or U21070 (N_21070,N_19044,N_15442);
or U21071 (N_21071,N_16576,N_18661);
nand U21072 (N_21072,N_18935,N_15496);
or U21073 (N_21073,N_17081,N_17961);
xor U21074 (N_21074,N_18145,N_18021);
nand U21075 (N_21075,N_18923,N_19879);
xor U21076 (N_21076,N_19239,N_16637);
nor U21077 (N_21077,N_18536,N_16563);
or U21078 (N_21078,N_15187,N_15343);
nand U21079 (N_21079,N_17242,N_18880);
and U21080 (N_21080,N_17241,N_15456);
nor U21081 (N_21081,N_15071,N_15808);
nand U21082 (N_21082,N_17080,N_15349);
xnor U21083 (N_21083,N_16000,N_16118);
or U21084 (N_21084,N_15908,N_15060);
or U21085 (N_21085,N_16935,N_18248);
nand U21086 (N_21086,N_15594,N_17664);
and U21087 (N_21087,N_19756,N_17868);
and U21088 (N_21088,N_16264,N_16656);
or U21089 (N_21089,N_15651,N_15696);
and U21090 (N_21090,N_15794,N_15584);
nand U21091 (N_21091,N_15357,N_16553);
nor U21092 (N_21092,N_17197,N_15305);
nor U21093 (N_21093,N_15588,N_18030);
nor U21094 (N_21094,N_17954,N_15375);
and U21095 (N_21095,N_17694,N_18746);
or U21096 (N_21096,N_18352,N_15367);
nand U21097 (N_21097,N_19744,N_16701);
nand U21098 (N_21098,N_16655,N_15914);
or U21099 (N_21099,N_19465,N_17048);
or U21100 (N_21100,N_18404,N_18654);
nand U21101 (N_21101,N_18101,N_16312);
nand U21102 (N_21102,N_17005,N_16169);
nor U21103 (N_21103,N_17976,N_18011);
nand U21104 (N_21104,N_16764,N_19469);
and U21105 (N_21105,N_16330,N_16875);
or U21106 (N_21106,N_18491,N_15050);
nand U21107 (N_21107,N_16446,N_19742);
or U21108 (N_21108,N_15009,N_19096);
xor U21109 (N_21109,N_15108,N_16560);
nand U21110 (N_21110,N_16519,N_16323);
nor U21111 (N_21111,N_17985,N_15708);
nand U21112 (N_21112,N_19378,N_15730);
or U21113 (N_21113,N_19939,N_17905);
or U21114 (N_21114,N_16490,N_17366);
nor U21115 (N_21115,N_16060,N_17124);
nand U21116 (N_21116,N_15812,N_17859);
nor U21117 (N_21117,N_16161,N_19376);
nor U21118 (N_21118,N_17451,N_17500);
and U21119 (N_21119,N_18313,N_15404);
nor U21120 (N_21120,N_19190,N_18026);
or U21121 (N_21121,N_19347,N_15809);
or U21122 (N_21122,N_17083,N_18349);
nand U21123 (N_21123,N_18090,N_15154);
or U21124 (N_21124,N_17671,N_16726);
or U21125 (N_21125,N_19856,N_18196);
and U21126 (N_21126,N_15658,N_17234);
xor U21127 (N_21127,N_17974,N_16815);
or U21128 (N_21128,N_15144,N_17706);
nand U21129 (N_21129,N_16370,N_15951);
or U21130 (N_21130,N_17085,N_15170);
or U21131 (N_21131,N_19383,N_17281);
or U21132 (N_21132,N_15799,N_17318);
nand U21133 (N_21133,N_17720,N_19360);
nand U21134 (N_21134,N_15755,N_17087);
nand U21135 (N_21135,N_18737,N_15265);
and U21136 (N_21136,N_15538,N_17565);
and U21137 (N_21137,N_15989,N_18415);
xor U21138 (N_21138,N_17726,N_17266);
xor U21139 (N_21139,N_17287,N_16057);
nand U21140 (N_21140,N_18534,N_15127);
nand U21141 (N_21141,N_17949,N_15364);
nand U21142 (N_21142,N_19029,N_18113);
nor U21143 (N_21143,N_18862,N_19179);
nor U21144 (N_21144,N_16925,N_19034);
and U21145 (N_21145,N_17378,N_16507);
or U21146 (N_21146,N_17257,N_17775);
nor U21147 (N_21147,N_16666,N_15027);
nor U21148 (N_21148,N_17568,N_19269);
nand U21149 (N_21149,N_17569,N_18288);
or U21150 (N_21150,N_18427,N_17669);
or U21151 (N_21151,N_18036,N_15243);
nand U21152 (N_21152,N_17770,N_18615);
nand U21153 (N_21153,N_17705,N_16220);
nand U21154 (N_21154,N_18054,N_18048);
or U21155 (N_21155,N_15886,N_19224);
nand U21156 (N_21156,N_16048,N_16783);
nor U21157 (N_21157,N_17517,N_17840);
or U21158 (N_21158,N_19759,N_18105);
nor U21159 (N_21159,N_19525,N_16771);
and U21160 (N_21160,N_16776,N_18616);
or U21161 (N_21161,N_16333,N_18626);
nand U21162 (N_21162,N_17990,N_18023);
and U21163 (N_21163,N_17616,N_17948);
nand U21164 (N_21164,N_16892,N_19393);
nor U21165 (N_21165,N_16741,N_19203);
or U21166 (N_21166,N_17299,N_16284);
and U21167 (N_21167,N_17086,N_19940);
and U21168 (N_21168,N_16722,N_18697);
nor U21169 (N_21169,N_16502,N_18813);
or U21170 (N_21170,N_17848,N_19253);
and U21171 (N_21171,N_17888,N_18525);
or U21172 (N_21172,N_17698,N_16130);
nor U21173 (N_21173,N_17238,N_18791);
and U21174 (N_21174,N_17765,N_19779);
xor U21175 (N_21175,N_19835,N_16541);
nor U21176 (N_21176,N_18601,N_18466);
nand U21177 (N_21177,N_19047,N_17400);
nand U21178 (N_21178,N_15530,N_15668);
and U21179 (N_21179,N_18658,N_15778);
xnor U21180 (N_21180,N_15163,N_19437);
nor U21181 (N_21181,N_18252,N_19201);
nor U21182 (N_21182,N_17738,N_18029);
nor U21183 (N_21183,N_18169,N_19934);
nor U21184 (N_21184,N_15215,N_17392);
or U21185 (N_21185,N_15665,N_19519);
and U21186 (N_21186,N_16516,N_17725);
nor U21187 (N_21187,N_15997,N_18367);
or U21188 (N_21188,N_15139,N_18937);
nor U21189 (N_21189,N_15471,N_16249);
or U21190 (N_21190,N_16466,N_19646);
nand U21191 (N_21191,N_19418,N_18099);
nor U21192 (N_21192,N_16552,N_16376);
nand U21193 (N_21193,N_17900,N_19202);
and U21194 (N_21194,N_16664,N_19069);
nor U21195 (N_21195,N_15451,N_17749);
and U21196 (N_21196,N_17476,N_16366);
or U21197 (N_21197,N_18337,N_17530);
and U21198 (N_21198,N_16358,N_15968);
nor U21199 (N_21199,N_17100,N_17687);
nor U21200 (N_21200,N_16556,N_15627);
nor U21201 (N_21201,N_15153,N_15342);
and U21202 (N_21202,N_17176,N_15293);
xnor U21203 (N_21203,N_15462,N_15234);
or U21204 (N_21204,N_18766,N_17491);
or U21205 (N_21205,N_19809,N_15898);
nand U21206 (N_21206,N_18590,N_19718);
or U21207 (N_21207,N_19533,N_18451);
nor U21208 (N_21208,N_15739,N_18989);
nor U21209 (N_21209,N_16518,N_19147);
nand U21210 (N_21210,N_19957,N_19656);
nor U21211 (N_21211,N_18818,N_18357);
nand U21212 (N_21212,N_18699,N_19941);
nor U21213 (N_21213,N_19171,N_19894);
or U21214 (N_21214,N_18481,N_15287);
or U21215 (N_21215,N_17999,N_17421);
nand U21216 (N_21216,N_15320,N_18947);
nand U21217 (N_21217,N_17322,N_17750);
and U21218 (N_21218,N_16837,N_17707);
nand U21219 (N_21219,N_17646,N_15858);
nand U21220 (N_21220,N_19771,N_15053);
nand U21221 (N_21221,N_15089,N_19877);
nand U21222 (N_21222,N_17487,N_17655);
or U21223 (N_21223,N_17847,N_16508);
nor U21224 (N_21224,N_17357,N_19038);
nand U21225 (N_21225,N_17904,N_15659);
nor U21226 (N_21226,N_15429,N_15871);
nor U21227 (N_21227,N_18520,N_15985);
or U21228 (N_21228,N_15941,N_17438);
nand U21229 (N_21229,N_18779,N_16862);
nor U21230 (N_21230,N_15323,N_19033);
nor U21231 (N_21231,N_15248,N_16597);
nor U21232 (N_21232,N_17933,N_19634);
nand U21233 (N_21233,N_16777,N_18784);
nor U21234 (N_21234,N_15259,N_16912);
nor U21235 (N_21235,N_18865,N_19870);
or U21236 (N_21236,N_17971,N_15824);
nand U21237 (N_21237,N_15945,N_17516);
nor U21238 (N_21238,N_16951,N_19271);
or U21239 (N_21239,N_16244,N_16468);
and U21240 (N_21240,N_18418,N_15800);
or U21241 (N_21241,N_19152,N_19222);
nand U21242 (N_21242,N_15929,N_15724);
xnor U21243 (N_21243,N_18194,N_17425);
and U21244 (N_21244,N_16967,N_15244);
and U21245 (N_21245,N_15915,N_16493);
and U21246 (N_21246,N_18908,N_18423);
nor U21247 (N_21247,N_17977,N_15512);
nand U21248 (N_21248,N_18255,N_15677);
nand U21249 (N_21249,N_15817,N_15815);
or U21250 (N_21250,N_18014,N_17371);
and U21251 (N_21251,N_17800,N_19682);
nor U21252 (N_21252,N_19752,N_16309);
nor U21253 (N_21253,N_18733,N_17551);
nand U21254 (N_21254,N_19218,N_17562);
or U21255 (N_21255,N_18421,N_19944);
and U21256 (N_21256,N_18301,N_16809);
and U21257 (N_21257,N_18976,N_18529);
and U21258 (N_21258,N_19458,N_18588);
and U21259 (N_21259,N_16710,N_16086);
nand U21260 (N_21260,N_17213,N_18245);
nor U21261 (N_21261,N_16665,N_18843);
xor U21262 (N_21262,N_19494,N_17099);
and U21263 (N_21263,N_15511,N_16290);
and U21264 (N_21264,N_17230,N_19031);
nand U21265 (N_21265,N_18705,N_16276);
nand U21266 (N_21266,N_19401,N_17739);
or U21267 (N_21267,N_19446,N_19936);
and U21268 (N_21268,N_19573,N_15789);
xnor U21269 (N_21269,N_17849,N_19768);
nor U21270 (N_21270,N_16638,N_18817);
or U21271 (N_21271,N_16905,N_15430);
xnor U21272 (N_21272,N_15520,N_15984);
nand U21273 (N_21273,N_15310,N_15517);
nor U21274 (N_21274,N_16231,N_18385);
or U21275 (N_21275,N_19678,N_15180);
or U21276 (N_21276,N_19539,N_15094);
and U21277 (N_21277,N_19078,N_17597);
nor U21278 (N_21278,N_19056,N_17277);
and U21279 (N_21279,N_18215,N_16714);
and U21280 (N_21280,N_17581,N_18059);
nor U21281 (N_21281,N_15851,N_15412);
or U21282 (N_21282,N_19361,N_16831);
nor U21283 (N_21283,N_15924,N_18089);
and U21284 (N_21284,N_16222,N_19070);
xor U21285 (N_21285,N_19566,N_17577);
or U21286 (N_21286,N_17202,N_16871);
nand U21287 (N_21287,N_17385,N_17251);
and U21288 (N_21288,N_16736,N_16354);
and U21289 (N_21289,N_18409,N_18949);
or U21290 (N_21290,N_16894,N_16236);
nor U21291 (N_21291,N_17811,N_15942);
nor U21292 (N_21292,N_17395,N_19177);
nand U21293 (N_21293,N_18429,N_17344);
nand U21294 (N_21294,N_17567,N_16420);
nor U21295 (N_21295,N_18158,N_15775);
nor U21296 (N_21296,N_15189,N_17473);
and U21297 (N_21297,N_18207,N_17898);
nand U21298 (N_21298,N_17113,N_16863);
or U21299 (N_21299,N_16546,N_16990);
or U21300 (N_21300,N_19547,N_18094);
or U21301 (N_21301,N_19576,N_19903);
or U21302 (N_21302,N_16958,N_19568);
nand U21303 (N_21303,N_19833,N_18870);
xor U21304 (N_21304,N_15624,N_17766);
and U21305 (N_21305,N_16617,N_19032);
nor U21306 (N_21306,N_19639,N_19128);
and U21307 (N_21307,N_18246,N_15466);
nor U21308 (N_21308,N_18918,N_18384);
or U21309 (N_21309,N_16511,N_17429);
and U21310 (N_21310,N_17537,N_15748);
or U21311 (N_21311,N_16660,N_15223);
nor U21312 (N_21312,N_17917,N_15614);
nor U21313 (N_21313,N_18795,N_17247);
or U21314 (N_21314,N_15058,N_17183);
or U21315 (N_21315,N_18890,N_19765);
nand U21316 (N_21316,N_18919,N_15854);
or U21317 (N_21317,N_17860,N_16910);
or U21318 (N_21318,N_19337,N_16922);
xnor U21319 (N_21319,N_19343,N_17644);
nand U21320 (N_21320,N_17591,N_19692);
nand U21321 (N_21321,N_19824,N_17330);
nand U21322 (N_21322,N_18528,N_17929);
nand U21323 (N_21323,N_19421,N_16260);
or U21324 (N_21324,N_17897,N_18487);
or U21325 (N_21325,N_18790,N_19966);
or U21326 (N_21326,N_15035,N_16102);
or U21327 (N_21327,N_17346,N_19490);
nor U21328 (N_21328,N_19804,N_16693);
or U21329 (N_21329,N_19164,N_17270);
nor U21330 (N_21330,N_17044,N_18302);
xor U21331 (N_21331,N_15927,N_17045);
or U21332 (N_21332,N_18256,N_15646);
and U21333 (N_21333,N_19392,N_19102);
nor U21334 (N_21334,N_15980,N_15121);
nor U21335 (N_21335,N_16509,N_19778);
nor U21336 (N_21336,N_16110,N_18009);
or U21337 (N_21337,N_17388,N_15973);
or U21338 (N_21338,N_19592,N_15297);
or U21339 (N_21339,N_15920,N_19165);
or U21340 (N_21340,N_18112,N_19205);
or U21341 (N_21341,N_18174,N_16971);
nand U21342 (N_21342,N_17201,N_17265);
nand U21343 (N_21343,N_15194,N_19278);
nand U21344 (N_21344,N_19586,N_18789);
nor U21345 (N_21345,N_15230,N_19947);
or U21346 (N_21346,N_16729,N_15605);
nor U21347 (N_21347,N_15675,N_19114);
nand U21348 (N_21348,N_15604,N_16844);
and U21349 (N_21349,N_16878,N_19688);
and U21350 (N_21350,N_16335,N_16681);
and U21351 (N_21351,N_15132,N_16476);
xor U21352 (N_21352,N_18803,N_15269);
or U21353 (N_21353,N_15351,N_19825);
nor U21354 (N_21354,N_15840,N_16024);
or U21355 (N_21355,N_15587,N_16131);
xor U21356 (N_21356,N_16590,N_17691);
nand U21357 (N_21357,N_19397,N_15260);
nor U21358 (N_21358,N_17393,N_15956);
and U21359 (N_21359,N_17922,N_19529);
nand U21360 (N_21360,N_19127,N_16146);
nor U21361 (N_21361,N_19495,N_19003);
and U21362 (N_21362,N_16616,N_16200);
nor U21363 (N_21363,N_15201,N_15445);
nor U21364 (N_21364,N_17135,N_15306);
nor U21365 (N_21365,N_16487,N_19466);
xor U21366 (N_21366,N_16197,N_19587);
or U21367 (N_21367,N_15500,N_18217);
nor U21368 (N_21368,N_18221,N_15082);
or U21369 (N_21369,N_19881,N_19140);
nand U21370 (N_21370,N_19358,N_15680);
nand U21371 (N_21371,N_19048,N_16445);
nand U21372 (N_21372,N_16165,N_15321);
nand U21373 (N_21373,N_16763,N_18484);
or U21374 (N_21374,N_17661,N_17454);
nand U21375 (N_21375,N_15413,N_19415);
and U21376 (N_21376,N_15642,N_16465);
nand U21377 (N_21377,N_19775,N_16241);
nand U21378 (N_21378,N_16372,N_18358);
or U21379 (N_21379,N_15388,N_16979);
and U21380 (N_21380,N_18776,N_15833);
nand U21381 (N_21381,N_17914,N_18008);
nand U21382 (N_21382,N_15469,N_19308);
or U21383 (N_21383,N_17019,N_15876);
or U21384 (N_21384,N_19198,N_19740);
xor U21385 (N_21385,N_18160,N_15933);
nand U21386 (N_21386,N_19601,N_15690);
nand U21387 (N_21387,N_19919,N_16412);
nor U21388 (N_21388,N_16902,N_17909);
nand U21389 (N_21389,N_16954,N_17334);
or U21390 (N_21390,N_15457,N_16470);
or U21391 (N_21391,N_18807,N_17243);
and U21392 (N_21392,N_16976,N_16861);
nand U21393 (N_21393,N_17439,N_15754);
nor U21394 (N_21394,N_18081,N_18596);
nor U21395 (N_21395,N_18619,N_17151);
nor U21396 (N_21396,N_19215,N_18636);
nor U21397 (N_21397,N_19964,N_19549);
nor U21398 (N_21398,N_18839,N_17331);
nor U21399 (N_21399,N_19923,N_17733);
nor U21400 (N_21400,N_19968,N_15785);
xnor U21401 (N_21401,N_15459,N_17254);
nor U21402 (N_21402,N_19082,N_18237);
nand U21403 (N_21403,N_17443,N_19372);
nand U21404 (N_21404,N_18467,N_15963);
or U21405 (N_21405,N_16589,N_17379);
or U21406 (N_21406,N_16390,N_19342);
and U21407 (N_21407,N_15859,N_16151);
and U21408 (N_21408,N_18392,N_19750);
and U21409 (N_21409,N_15080,N_16227);
nor U21410 (N_21410,N_15996,N_16408);
xnor U21411 (N_21411,N_19482,N_17076);
nand U21412 (N_21412,N_16630,N_16243);
nor U21413 (N_21413,N_17382,N_16615);
and U21414 (N_21414,N_15527,N_16304);
nand U21415 (N_21415,N_18259,N_18728);
nand U21416 (N_21416,N_15699,N_18903);
nor U21417 (N_21417,N_19151,N_15875);
nand U21418 (N_21418,N_16339,N_19958);
and U21419 (N_21419,N_15848,N_18341);
or U21420 (N_21420,N_18538,N_19563);
nor U21421 (N_21421,N_18617,N_17584);
or U21422 (N_21422,N_15309,N_19200);
nor U21423 (N_21423,N_17981,N_15174);
nand U21424 (N_21424,N_17269,N_18558);
nor U21425 (N_21425,N_16889,N_18930);
or U21426 (N_21426,N_18873,N_15052);
and U21427 (N_21427,N_17596,N_15606);
nand U21428 (N_21428,N_19217,N_15423);
and U21429 (N_21429,N_16056,N_16657);
nand U21430 (N_21430,N_19258,N_19993);
xnor U21431 (N_21431,N_19133,N_16299);
nand U21432 (N_21432,N_18106,N_17629);
nand U21433 (N_21433,N_19671,N_18147);
or U21434 (N_21434,N_16001,N_16152);
xor U21435 (N_21435,N_19384,N_16074);
nor U21436 (N_21436,N_17798,N_15008);
xor U21437 (N_21437,N_17424,N_18673);
nand U21438 (N_21438,N_15721,N_19113);
and U21439 (N_21439,N_18710,N_16229);
xor U21440 (N_21440,N_17988,N_15165);
nor U21441 (N_21441,N_17774,N_15617);
and U21442 (N_21442,N_16919,N_15014);
nor U21443 (N_21443,N_16005,N_19808);
nor U21444 (N_21444,N_18651,N_19609);
or U21445 (N_21445,N_17194,N_16695);
or U21446 (N_21446,N_17807,N_18516);
or U21447 (N_21447,N_16247,N_18692);
or U21448 (N_21448,N_17996,N_17875);
nand U21449 (N_21449,N_17313,N_19249);
nor U21450 (N_21450,N_17965,N_15167);
nor U21451 (N_21451,N_19095,N_16730);
or U21452 (N_21452,N_15051,N_16210);
or U21453 (N_21453,N_18730,N_16833);
or U21454 (N_21454,N_16444,N_19701);
and U21455 (N_21455,N_18103,N_17605);
and U21456 (N_21456,N_19312,N_18618);
and U21457 (N_21457,N_18572,N_19643);
xor U21458 (N_21458,N_18788,N_15224);
xor U21459 (N_21459,N_16916,N_19569);
and U21460 (N_21460,N_18760,N_16495);
or U21461 (N_21461,N_16904,N_16622);
nor U21462 (N_21462,N_19334,N_15272);
nand U21463 (N_21463,N_16374,N_17406);
or U21464 (N_21464,N_18151,N_15519);
and U21465 (N_21465,N_18556,N_15001);
or U21466 (N_21466,N_15510,N_19119);
nor U21467 (N_21467,N_15553,N_15676);
nand U21468 (N_21468,N_16933,N_17599);
and U21469 (N_21469,N_17283,N_18336);
nand U21470 (N_21470,N_19782,N_18378);
and U21471 (N_21471,N_19115,N_15107);
or U21472 (N_21472,N_19902,N_17821);
or U21473 (N_21473,N_15336,N_15697);
xor U21474 (N_21474,N_18527,N_18175);
nor U21475 (N_21475,N_16987,N_19389);
nor U21476 (N_21476,N_15410,N_17082);
nand U21477 (N_21477,N_16953,N_16122);
or U21478 (N_21478,N_18598,N_15313);
xnor U21479 (N_21479,N_19039,N_19560);
or U21480 (N_21480,N_19451,N_17042);
nor U21481 (N_21481,N_17826,N_16570);
xnor U21482 (N_21482,N_15781,N_19900);
or U21483 (N_21483,N_19973,N_19052);
nand U21484 (N_21484,N_18108,N_16423);
or U21485 (N_21485,N_19694,N_17972);
nor U21486 (N_21486,N_18020,N_17171);
nand U21487 (N_21487,N_19649,N_19399);
and U21488 (N_21488,N_18835,N_16718);
nor U21489 (N_21489,N_18857,N_16311);
nor U21490 (N_21490,N_15169,N_19160);
and U21491 (N_21491,N_19979,N_15023);
and U21492 (N_21492,N_18669,N_16017);
or U21493 (N_21493,N_15946,N_16605);
and U21494 (N_21494,N_18227,N_19504);
and U21495 (N_21495,N_15402,N_19385);
or U21496 (N_21496,N_15912,N_16798);
or U21497 (N_21497,N_16252,N_16322);
nor U21498 (N_21498,N_19314,N_16153);
or U21499 (N_21499,N_18266,N_16857);
nand U21500 (N_21500,N_15911,N_17428);
or U21501 (N_21501,N_16486,N_19162);
nor U21502 (N_21502,N_19534,N_16204);
and U21503 (N_21503,N_15903,N_17620);
nor U21504 (N_21504,N_18951,N_16867);
nand U21505 (N_21505,N_18553,N_17147);
or U21506 (N_21506,N_19471,N_15686);
and U21507 (N_21507,N_17575,N_17049);
or U21508 (N_21508,N_19442,N_18212);
or U21509 (N_21509,N_18270,N_15978);
nor U21510 (N_21510,N_18567,N_15767);
nor U21511 (N_21511,N_18805,N_17295);
nand U21512 (N_21512,N_19273,N_16790);
xor U21513 (N_21513,N_17096,N_18206);
nor U21514 (N_21514,N_16784,N_16566);
or U21515 (N_21515,N_16799,N_18822);
nor U21516 (N_21516,N_19674,N_19449);
and U21517 (N_21517,N_17526,N_16639);
and U21518 (N_21518,N_17064,N_19470);
xnor U21519 (N_21519,N_18622,N_19286);
nor U21520 (N_21520,N_18680,N_17918);
or U21521 (N_21521,N_15718,N_16141);
nand U21522 (N_21522,N_15470,N_19663);
and U21523 (N_21523,N_17304,N_18893);
nor U21524 (N_21524,N_15592,N_19300);
nor U21525 (N_21525,N_19491,N_19377);
nor U21526 (N_21526,N_15691,N_18944);
or U21527 (N_21527,N_15120,N_17498);
and U21528 (N_21528,N_18643,N_15119);
and U21529 (N_21529,N_17248,N_16187);
and U21530 (N_21530,N_15206,N_16078);
xor U21531 (N_21531,N_16320,N_18058);
nand U21532 (N_21532,N_18274,N_16019);
or U21533 (N_21533,N_16064,N_19009);
nor U21534 (N_21534,N_18028,N_19441);
xor U21535 (N_21535,N_18183,N_17399);
nand U21536 (N_21536,N_18757,N_17103);
xor U21537 (N_21537,N_16327,N_18056);
or U21538 (N_21538,N_16155,N_15720);
nand U21539 (N_21539,N_19496,N_15857);
nor U21540 (N_21540,N_17704,N_18479);
nor U21541 (N_21541,N_18763,N_17291);
or U21542 (N_21542,N_19699,N_19425);
and U21543 (N_21543,N_16573,N_15548);
nor U21544 (N_21544,N_15290,N_17310);
and U21545 (N_21545,N_17469,N_16459);
and U21546 (N_21546,N_16989,N_16488);
xor U21547 (N_21547,N_17040,N_19303);
or U21548 (N_21548,N_19149,N_19186);
and U21549 (N_21549,N_16362,N_17928);
nand U21550 (N_21550,N_19080,N_18354);
nor U21551 (N_21551,N_19632,N_19060);
or U21552 (N_21552,N_15631,N_15740);
nand U21553 (N_21553,N_15779,N_15860);
nand U21554 (N_21554,N_16997,N_18312);
nor U21555 (N_21555,N_16266,N_17994);
or U21556 (N_21556,N_16140,N_17075);
and U21557 (N_21557,N_18831,N_18812);
nand U21558 (N_21558,N_15692,N_17091);
or U21559 (N_21559,N_16261,N_17132);
xnor U21560 (N_21560,N_18032,N_16329);
nand U21561 (N_21561,N_16972,N_19049);
and U21562 (N_21562,N_16004,N_16613);
and U21563 (N_21563,N_17441,N_17453);
or U21564 (N_21564,N_15172,N_17793);
and U21565 (N_21565,N_15711,N_19289);
and U21566 (N_21566,N_15256,N_18774);
nor U21567 (N_21567,N_16419,N_19391);
or U21568 (N_21568,N_19484,N_19394);
nand U21569 (N_21569,N_15836,N_16594);
or U21570 (N_21570,N_19126,N_16198);
and U21571 (N_21571,N_16010,N_15625);
xor U21572 (N_21572,N_17166,N_15130);
nor U21573 (N_21573,N_18450,N_19630);
nor U21574 (N_21574,N_16255,N_15488);
nand U21575 (N_21575,N_18749,N_19938);
nand U21576 (N_21576,N_18504,N_19054);
and U21577 (N_21577,N_18574,N_17221);
nor U21578 (N_21578,N_18517,N_19092);
and U21579 (N_21579,N_18049,N_16702);
or U21580 (N_21580,N_15850,N_19111);
or U21581 (N_21581,N_19929,N_15446);
nor U21582 (N_21582,N_18602,N_18603);
or U21583 (N_21583,N_18712,N_18953);
or U21584 (N_21584,N_15330,N_16076);
and U21585 (N_21585,N_16202,N_18597);
nor U21586 (N_21586,N_17693,N_18832);
nand U21587 (N_21587,N_15332,N_18493);
nor U21588 (N_21588,N_18247,N_18541);
and U21589 (N_21589,N_18625,N_19199);
nor U21590 (N_21590,N_15717,N_16578);
xnor U21591 (N_21591,N_15524,N_16015);
and U21592 (N_21592,N_16133,N_18998);
or U21593 (N_21593,N_16223,N_19213);
or U21594 (N_21594,N_18980,N_19556);
nand U21595 (N_21595,N_18531,N_19233);
nand U21596 (N_21596,N_15232,N_18589);
nand U21597 (N_21597,N_19363,N_15666);
xor U21598 (N_21598,N_15845,N_19373);
and U21599 (N_21599,N_15753,N_16903);
nand U21600 (N_21600,N_15461,N_16838);
or U21601 (N_21601,N_17161,N_16230);
and U21602 (N_21602,N_18759,N_15040);
nor U21603 (N_21603,N_18420,N_18906);
nand U21604 (N_21604,N_18488,N_16341);
or U21605 (N_21605,N_15619,N_16611);
and U21606 (N_21606,N_17199,N_16872);
or U21607 (N_21607,N_15736,N_18738);
nand U21608 (N_21608,N_19659,N_15377);
nand U21609 (N_21609,N_16977,N_16166);
nor U21610 (N_21610,N_15190,N_16359);
nor U21611 (N_21611,N_17728,N_15277);
nand U21612 (N_21612,N_19332,N_19419);
and U21613 (N_21613,N_15048,N_18902);
nand U21614 (N_21614,N_18543,N_17759);
or U21615 (N_21615,N_17073,N_17747);
xor U21616 (N_21616,N_18506,N_19150);
or U21617 (N_21617,N_15567,N_18102);
and U21618 (N_21618,N_18498,N_17297);
nand U21619 (N_21619,N_18627,N_17445);
or U21620 (N_21620,N_17134,N_17268);
or U21621 (N_21621,N_17187,N_16458);
nor U21622 (N_21622,N_18578,N_15419);
nand U21623 (N_21623,N_16600,N_15031);
and U21624 (N_21624,N_17529,N_18682);
and U21625 (N_21625,N_19535,N_16881);
xnor U21626 (N_21626,N_15331,N_15371);
and U21627 (N_21627,N_16352,N_17389);
or U21628 (N_21628,N_18276,N_15618);
nand U21629 (N_21629,N_16213,N_17758);
or U21630 (N_21630,N_16716,N_17730);
or U21631 (N_21631,N_17630,N_15716);
and U21632 (N_21632,N_19717,N_18109);
nand U21633 (N_21633,N_15134,N_15516);
nor U21634 (N_21634,N_19781,N_18545);
nand U21635 (N_21635,N_15049,N_17865);
nand U21636 (N_21636,N_19216,N_16053);
and U21637 (N_21637,N_17721,N_17298);
nor U21638 (N_21638,N_15813,N_18837);
and U21639 (N_21639,N_16403,N_15575);
xnor U21640 (N_21640,N_16206,N_19948);
xnor U21641 (N_21641,N_18495,N_19962);
xor U21642 (N_21642,N_18702,N_15541);
nand U21643 (N_21643,N_18557,N_16800);
nand U21644 (N_21644,N_18445,N_16524);
or U21645 (N_21645,N_18771,N_17333);
or U21646 (N_21646,N_16291,N_15076);
nor U21647 (N_21647,N_15054,N_17957);
nand U21648 (N_21648,N_16449,N_16047);
xor U21649 (N_21649,N_17866,N_17727);
or U21650 (N_21650,N_15551,N_17806);
nor U21651 (N_21651,N_19382,N_18346);
nand U21652 (N_21652,N_17667,N_19716);
nand U21653 (N_21653,N_19374,N_18782);
nor U21654 (N_21654,N_15932,N_17440);
xnor U21655 (N_21655,N_18383,N_15188);
or U21656 (N_21656,N_18279,N_15012);
nor U21657 (N_21657,N_17822,N_18792);
and U21658 (N_21658,N_19875,N_15141);
nor U21659 (N_21659,N_19555,N_19025);
and U21660 (N_21660,N_16836,N_17889);
or U21661 (N_21661,N_17650,N_18278);
and U21662 (N_21662,N_16732,N_18811);
xnor U21663 (N_21663,N_18868,N_19605);
and U21664 (N_21664,N_19122,N_19362);
nor U21665 (N_21665,N_16385,N_16761);
xnor U21666 (N_21666,N_15591,N_19493);
and U21667 (N_21667,N_17561,N_19319);
nand U21668 (N_21668,N_16829,N_15525);
nor U21669 (N_21669,N_18006,N_17181);
nand U21670 (N_21670,N_16263,N_19743);
nor U21671 (N_21671,N_17810,N_17893);
or U21672 (N_21672,N_16040,N_17152);
nand U21673 (N_21673,N_16461,N_15536);
nor U21674 (N_21674,N_18475,N_17467);
nor U21675 (N_21675,N_19450,N_16924);
and U21676 (N_21676,N_17252,N_18202);
or U21677 (N_21677,N_16099,N_15463);
and U21678 (N_21678,N_16782,N_16545);
nor U21679 (N_21679,N_15160,N_18946);
nor U21680 (N_21680,N_19212,N_18824);
and U21681 (N_21681,N_16794,N_17347);
nor U21682 (N_21682,N_19497,N_16841);
nand U21683 (N_21683,N_15863,N_18182);
or U21684 (N_21684,N_18546,N_17339);
or U21685 (N_21685,N_16107,N_19235);
nor U21686 (N_21686,N_19058,N_15007);
nand U21687 (N_21687,N_19867,N_19544);
nor U21688 (N_21688,N_19475,N_17514);
or U21689 (N_21689,N_16163,N_16282);
and U21690 (N_21690,N_17619,N_17169);
xnor U21691 (N_21691,N_15083,N_19257);
xnor U21692 (N_21692,N_16209,N_16039);
nand U21693 (N_21693,N_15937,N_17178);
xor U21694 (N_21694,N_16027,N_16773);
or U21695 (N_21695,N_16054,N_18070);
nand U21696 (N_21696,N_19110,N_16405);
nor U21697 (N_21697,N_18864,N_19698);
nor U21698 (N_21698,N_15713,N_18173);
and U21699 (N_21699,N_17919,N_15607);
and U21700 (N_21700,N_15159,N_19893);
nand U21701 (N_21701,N_19735,N_17966);
nor U21702 (N_21702,N_19413,N_18463);
and U21703 (N_21703,N_18460,N_15688);
nor U21704 (N_21704,N_16706,N_18477);
and U21705 (N_21705,N_16626,N_17452);
xor U21706 (N_21706,N_15780,N_15887);
nor U21707 (N_21707,N_15921,N_19242);
nor U21708 (N_21708,N_19803,N_15233);
nor U21709 (N_21709,N_17033,N_16574);
or U21710 (N_21710,N_18225,N_15938);
nor U21711 (N_21711,N_17016,N_19980);
and U21712 (N_21712,N_18798,N_16547);
or U21713 (N_21713,N_17300,N_17144);
or U21714 (N_21714,N_15616,N_19869);
and U21715 (N_21715,N_19798,N_17125);
or U21716 (N_21716,N_19214,N_16898);
and U21717 (N_21717,N_17275,N_17503);
xor U21718 (N_21718,N_19857,N_19852);
and U21719 (N_21719,N_16804,N_17228);
xor U21720 (N_21720,N_15005,N_17618);
and U21721 (N_21721,N_18439,N_15029);
nand U21722 (N_21722,N_17992,N_17532);
or U21723 (N_21723,N_18887,N_17987);
nor U21724 (N_21724,N_17209,N_15883);
nand U21725 (N_21725,N_16759,N_19638);
nand U21726 (N_21726,N_15024,N_16936);
and U21727 (N_21727,N_15682,N_15637);
or U21728 (N_21728,N_16724,N_16592);
nand U21729 (N_21729,N_15066,N_19226);
nand U21730 (N_21730,N_18428,N_19758);
nor U21731 (N_21731,N_18978,N_18881);
nand U21732 (N_21732,N_17021,N_16734);
or U21733 (N_21733,N_19398,N_16963);
and U21734 (N_21734,N_17116,N_16472);
nor U21735 (N_21735,N_15087,N_15476);
nand U21736 (N_21736,N_17964,N_19892);
or U21737 (N_21737,N_17137,N_19780);
xor U21738 (N_21738,N_17980,N_17437);
nor U21739 (N_21739,N_17572,N_19348);
nand U21740 (N_21740,N_19842,N_18091);
nor U21741 (N_21741,N_15249,N_16336);
or U21742 (N_21742,N_18473,N_15630);
nand U21743 (N_21743,N_16287,N_16717);
or U21744 (N_21744,N_15073,N_18184);
nand U21745 (N_21745,N_17146,N_18396);
and U21746 (N_21746,N_19129,N_15150);
or U21747 (N_21747,N_17356,N_18735);
and U21748 (N_21748,N_19793,N_15774);
nor U21749 (N_21749,N_15602,N_16196);
nand U21750 (N_21750,N_16868,N_16549);
and U21751 (N_21751,N_15453,N_15972);
nand U21752 (N_21752,N_15398,N_15204);
and U21753 (N_21753,N_15645,N_17590);
xor U21754 (N_21754,N_15987,N_17306);
nand U21755 (N_21755,N_17657,N_17444);
nand U21756 (N_21756,N_17862,N_16235);
nor U21757 (N_21757,N_18503,N_16555);
and U21758 (N_21758,N_17867,N_19585);
xor U21759 (N_21759,N_15791,N_18369);
nor U21760 (N_21760,N_19510,N_17205);
or U21761 (N_21761,N_18410,N_19124);
or U21762 (N_21762,N_16138,N_18554);
or U21763 (N_21763,N_18910,N_19920);
xnor U21764 (N_21764,N_16460,N_16961);
and U21765 (N_21765,N_16937,N_16523);
nand U21766 (N_21766,N_17809,N_17483);
and U21767 (N_21767,N_17068,N_18717);
xor U21768 (N_21768,N_19422,N_18500);
or U21769 (N_21769,N_15663,N_18555);
nand U21770 (N_21770,N_17206,N_19719);
and U21771 (N_21771,N_19050,N_17284);
and U21772 (N_21772,N_19839,N_16789);
nor U21773 (N_21773,N_18172,N_18334);
nand U21774 (N_21774,N_18177,N_16321);
xor U21775 (N_21775,N_17020,N_16891);
and U21776 (N_21776,N_18628,N_16043);
xnor U21777 (N_21777,N_19800,N_17063);
or U21778 (N_21778,N_16272,N_17157);
or U21779 (N_21779,N_18796,N_19618);
nand U21780 (N_21780,N_15483,N_17684);
nand U21781 (N_21781,N_15750,N_16612);
and U21782 (N_21782,N_15186,N_15356);
nand U21783 (N_21783,N_16079,N_15830);
nor U21784 (N_21784,N_17582,N_15344);
xnor U21785 (N_21785,N_18938,N_19961);
or U21786 (N_21786,N_15878,N_15199);
nand U21787 (N_21787,N_19974,N_18907);
nand U21788 (N_21788,N_18292,N_18579);
nor U21789 (N_21789,N_19323,N_18024);
nor U21790 (N_21790,N_19410,N_18239);
nor U21791 (N_21791,N_15861,N_17662);
nor U21792 (N_21792,N_19636,N_19913);
or U21793 (N_21793,N_18727,N_19228);
nor U21794 (N_21794,N_19074,N_17023);
or U21795 (N_21795,N_17092,N_17219);
and U21796 (N_21796,N_18037,N_16283);
nand U21797 (N_21797,N_15554,N_17427);
nand U21798 (N_21798,N_19311,N_19426);
or U21799 (N_21799,N_18888,N_19075);
nor U21800 (N_21800,N_15852,N_16750);
nor U21801 (N_21801,N_17123,N_18515);
nand U21802 (N_21802,N_15902,N_19168);
nand U21803 (N_21803,N_17920,N_16510);
and U21804 (N_21804,N_18724,N_19843);
or U21805 (N_21805,N_17336,N_15497);
nor U21806 (N_21806,N_19400,N_19365);
and U21807 (N_21807,N_18381,N_15338);
or U21808 (N_21808,N_18472,N_18398);
nor U21809 (N_21809,N_17748,N_15609);
and U21810 (N_21810,N_19550,N_15315);
nand U21811 (N_21811,N_19000,N_16662);
or U21812 (N_21812,N_17573,N_18359);
nor U21813 (N_21813,N_17543,N_18066);
or U21814 (N_21814,N_18330,N_17341);
nor U21815 (N_21815,N_16968,N_15970);
nand U21816 (N_21816,N_16941,N_19014);
xor U21817 (N_21817,N_18114,N_17032);
and U21818 (N_21818,N_16944,N_18819);
and U21819 (N_21819,N_15124,N_19901);
or U21820 (N_21820,N_17834,N_15595);
nand U21821 (N_21821,N_17039,N_18290);
or U21822 (N_21822,N_19935,N_17887);
nor U21823 (N_21823,N_19094,N_16845);
xor U21824 (N_21824,N_18001,N_15072);
or U21825 (N_21825,N_19799,N_15435);
nor U21826 (N_21826,N_15123,N_18242);
nand U21827 (N_21827,N_16147,N_15074);
and U21828 (N_21828,N_17541,N_18163);
nor U21829 (N_21829,N_15129,N_18343);
nor U21830 (N_21830,N_19142,N_17926);
nor U21831 (N_21831,N_19731,N_19062);
nand U21832 (N_21832,N_17953,N_18304);
xnor U21833 (N_21833,N_19390,N_16045);
nor U21834 (N_21834,N_19624,N_19340);
or U21835 (N_21835,N_19951,N_17224);
nand U21836 (N_21836,N_18241,N_19478);
or U21837 (N_21837,N_15477,N_19978);
nor U21838 (N_21838,N_15235,N_17771);
or U21839 (N_21839,N_15020,N_18107);
or U21840 (N_21840,N_15184,N_19686);
or U21841 (N_21841,N_16353,N_17613);
and U21842 (N_21842,N_16614,N_15209);
or U21843 (N_21843,N_16740,N_18804);
nor U21844 (N_21844,N_17583,N_16633);
or U21845 (N_21845,N_17218,N_17881);
nand U21846 (N_21846,N_19702,N_18853);
xnor U21847 (N_21847,N_18645,N_15361);
nor U21848 (N_21848,N_18240,N_19614);
nand U21849 (N_21849,N_16747,N_15502);
or U21850 (N_21850,N_17235,N_19333);
xnor U21851 (N_21851,N_18793,N_19776);
and U21852 (N_21852,N_19924,N_19985);
xnor U21853 (N_21853,N_15839,N_16959);
nor U21854 (N_21854,N_16675,N_17413);
nand U21855 (N_21855,N_17481,N_18363);
xnor U21856 (N_21856,N_18494,N_18211);
nand U21857 (N_21857,N_16316,N_17368);
or U21858 (N_21858,N_19932,N_16127);
nand U21859 (N_21859,N_15329,N_15873);
and U21860 (N_21860,N_18131,N_19720);
xnor U21861 (N_21861,N_17863,N_19387);
or U21862 (N_21862,N_17892,N_15678);
or U21863 (N_21863,N_16082,N_15661);
or U21864 (N_21864,N_15881,N_19687);
and U21865 (N_21865,N_18632,N_19616);
and U21866 (N_21866,N_15820,N_17663);
and U21867 (N_21867,N_17776,N_16453);
and U21868 (N_21868,N_19631,N_16698);
nand U21869 (N_21869,N_18869,N_19085);
nand U21870 (N_21870,N_19280,N_17789);
and U21871 (N_21871,N_17723,N_17479);
nand U21872 (N_21872,N_18765,N_17695);
xnor U21873 (N_21873,N_19167,N_19457);
nand U21874 (N_21874,N_18809,N_15145);
or U21875 (N_21875,N_17703,N_16629);
nor U21876 (N_21876,N_17014,N_15583);
xnor U21877 (N_21877,N_17104,N_19468);
nor U21878 (N_21878,N_15006,N_18062);
nand U21879 (N_21879,N_18315,N_17216);
nor U21880 (N_21880,N_19209,N_18876);
and U21881 (N_21881,N_18510,N_19131);
nand U21882 (N_21882,N_15111,N_19448);
or U21883 (N_21883,N_19178,N_17555);
and U21884 (N_21884,N_18686,N_18223);
nor U21885 (N_21885,N_16238,N_18867);
nand U21886 (N_21886,N_18275,N_15198);
nand U21887 (N_21887,N_18097,N_19016);
or U21888 (N_21888,N_19261,N_19225);
or U21889 (N_21889,N_17939,N_16331);
and U21890 (N_21890,N_16128,N_15363);
nand U21891 (N_21891,N_19281,N_15769);
nor U21892 (N_21892,N_17046,N_15327);
nand U21893 (N_21893,N_18808,N_18552);
and U21894 (N_21894,N_16308,N_17111);
and U21895 (N_21895,N_15981,N_18306);
nand U21896 (N_21896,N_16620,N_18438);
xnor U21897 (N_21897,N_16326,N_15831);
and U21898 (N_21898,N_17589,N_18945);
nor U21899 (N_21899,N_19905,N_19335);
nand U21900 (N_21900,N_18413,N_18253);
and U21901 (N_21901,N_17264,N_18639);
nor U21902 (N_21902,N_19196,N_19792);
or U21903 (N_21903,N_18707,N_17435);
or U21904 (N_21904,N_19658,N_16055);
nor U21905 (N_21905,N_17754,N_15455);
nor U21906 (N_21906,N_19664,N_15237);
nor U21907 (N_21907,N_18814,N_17267);
and U21908 (N_21908,N_17210,N_17468);
and U21909 (N_21909,N_16269,N_18433);
nor U21910 (N_21910,N_15242,N_18364);
or U21911 (N_21911,N_17576,N_19247);
and U21912 (N_21912,N_15479,N_18979);
nor U21913 (N_21913,N_18127,N_15965);
nand U21914 (N_21914,N_16705,N_15325);
or U21915 (N_21915,N_17288,N_19607);
nor U21916 (N_21916,N_16121,N_18323);
nor U21917 (N_21917,N_19635,N_17637);
nor U21918 (N_21918,N_17130,N_19438);
and U21919 (N_21919,N_17386,N_18043);
or U21920 (N_21920,N_18560,N_18581);
nor U21921 (N_21921,N_16435,N_19722);
or U21922 (N_21922,N_15210,N_18143);
nand U21923 (N_21923,N_19103,N_17755);
nor U21924 (N_21924,N_18455,N_16753);
xnor U21925 (N_21925,N_16409,N_17217);
nor U21926 (N_21926,N_18700,N_19500);
or U21927 (N_21927,N_19345,N_19406);
and U21928 (N_21928,N_17196,N_19797);
and U21929 (N_21929,N_17641,N_17540);
nor U21930 (N_21930,N_18339,N_15726);
xor U21931 (N_21931,N_16205,N_16539);
nor U21932 (N_21932,N_18904,N_15585);
or U21933 (N_21933,N_15407,N_19084);
nor U21934 (N_21934,N_17246,N_19862);
nor U21935 (N_21935,N_15178,N_16522);
nand U21936 (N_21936,N_16591,N_16813);
nand U21937 (N_21937,N_17233,N_15418);
or U21938 (N_21938,N_19322,N_18216);
and U21939 (N_21939,N_16558,N_17361);
xnor U21940 (N_21940,N_17101,N_15599);
or U21941 (N_21941,N_17814,N_17001);
nand U21942 (N_21942,N_16618,N_16417);
nor U21943 (N_21943,N_17059,N_17685);
and U21944 (N_21944,N_17876,N_17593);
nor U21945 (N_21945,N_17735,N_19820);
and U21946 (N_21946,N_16671,N_17138);
and U21947 (N_21947,N_17815,N_15869);
or U21948 (N_21948,N_19989,N_15112);
nor U21949 (N_21949,N_16028,N_17534);
nand U21950 (N_21950,N_17653,N_17588);
and U21951 (N_21951,N_18394,N_19522);
or U21952 (N_21952,N_16245,N_19545);
nor U21953 (N_21953,N_19912,N_16315);
xnor U21954 (N_21954,N_17947,N_18430);
or U21955 (N_21955,N_18142,N_16489);
nand U21956 (N_21956,N_15620,N_19640);
nand U21957 (N_21957,N_15340,N_19444);
and U21958 (N_21958,N_17416,N_18886);
xnor U21959 (N_21959,N_15362,N_18800);
nor U21960 (N_21960,N_18442,N_17402);
or U21961 (N_21961,N_19462,N_17626);
nor U21962 (N_21962,N_15529,N_15109);
nor U21963 (N_21963,N_16687,N_19703);
or U21964 (N_21964,N_15562,N_18167);
xnor U21965 (N_21965,N_17106,N_15077);
nor U21966 (N_21966,N_16270,N_19767);
nand U21967 (N_21967,N_19538,N_19882);
or U21968 (N_21968,N_18361,N_17542);
nor U21969 (N_21969,N_17418,N_17397);
nand U21970 (N_21970,N_16400,N_18621);
or U21971 (N_21971,N_18365,N_17212);
or U21972 (N_21972,N_16119,N_16991);
nor U21973 (N_21973,N_16096,N_15217);
nor U21974 (N_21974,N_19277,N_19135);
nor U21975 (N_21975,N_17545,N_16823);
nand U21976 (N_21976,N_16646,N_15443);
nor U21977 (N_21977,N_15961,N_17625);
and U21978 (N_21978,N_15274,N_15000);
nor U21979 (N_21979,N_19146,N_18214);
nand U21980 (N_21980,N_16879,N_16167);
nand U21981 (N_21981,N_19117,N_17259);
and U21982 (N_21982,N_17945,N_15955);
and U21983 (N_21983,N_15977,N_16491);
nor U21984 (N_21984,N_16342,N_17302);
or U21985 (N_21985,N_15540,N_17548);
and U21986 (N_21986,N_18236,N_19823);
and U21987 (N_21987,N_18033,N_15322);
or U21988 (N_21988,N_15378,N_16530);
nor U21989 (N_21989,N_17518,N_16978);
nand U21990 (N_21990,N_15514,N_18729);
and U21991 (N_21991,N_16361,N_17717);
nand U21992 (N_21992,N_18535,N_18580);
or U21993 (N_21993,N_17608,N_15679);
xor U21994 (N_21994,N_18170,N_18922);
nor U21995 (N_21995,N_15341,N_15285);
nor U21996 (N_21996,N_18845,N_18156);
or U21997 (N_21997,N_18802,N_16162);
nor U21998 (N_21998,N_18595,N_19408);
and U21999 (N_21999,N_18448,N_19477);
and U22000 (N_22000,N_19904,N_15917);
or U22001 (N_22001,N_16022,N_19100);
or U22002 (N_22002,N_16636,N_18965);
or U22003 (N_22003,N_19420,N_15737);
or U22004 (N_22004,N_18967,N_19915);
nor U22005 (N_22005,N_18551,N_16609);
and U22006 (N_22006,N_16278,N_19109);
nand U22007 (N_22007,N_19480,N_17328);
nand U22008 (N_22008,N_19580,N_17163);
nor U22009 (N_22009,N_16134,N_18806);
nand U22010 (N_22010,N_16727,N_18417);
xnor U22011 (N_22011,N_16647,N_15928);
nor U22012 (N_22012,N_18204,N_17227);
and U22013 (N_22013,N_17172,N_17763);
nor U22014 (N_22014,N_16683,N_19714);
nor U22015 (N_22015,N_15904,N_15639);
nor U22016 (N_22016,N_18895,N_15771);
xnor U22017 (N_22017,N_15352,N_15589);
nand U22018 (N_22018,N_19885,N_15440);
nor U22019 (N_22019,N_18764,N_16768);
or U22020 (N_22020,N_18133,N_16709);
nand U22021 (N_22021,N_17829,N_18773);
xor U22022 (N_22022,N_19757,N_17673);
and U22023 (N_22023,N_15258,N_16787);
or U22024 (N_22024,N_18064,N_18640);
nand U22025 (N_22025,N_19620,N_16754);
nand U22026 (N_22026,N_17989,N_19088);
nor U22027 (N_22027,N_16185,N_17027);
nor U22028 (N_22028,N_18912,N_19542);
or U22029 (N_22029,N_15098,N_15308);
xnor U22030 (N_22030,N_16305,N_19661);
nand U22031 (N_22031,N_18281,N_17232);
nand U22032 (N_22032,N_18915,N_16621);
or U22033 (N_22033,N_16443,N_16195);
nor U22034 (N_22034,N_19489,N_18284);
and U22035 (N_22035,N_19950,N_15499);
nor U22036 (N_22036,N_16711,N_19028);
or U22037 (N_22037,N_19395,N_15103);
or U22038 (N_22038,N_18856,N_15079);
and U22039 (N_22039,N_18135,N_16641);
and U22040 (N_22040,N_19629,N_16962);
nor U22041 (N_22041,N_17812,N_16504);
nor U22042 (N_22042,N_15067,N_16148);
nor U22043 (N_22043,N_17654,N_15275);
or U22044 (N_22044,N_17666,N_17282);
or U22045 (N_22045,N_17050,N_18911);
or U22046 (N_22046,N_17603,N_15705);
nor U22047 (N_22047,N_17991,N_17307);
nor U22048 (N_22048,N_15140,N_16564);
or U22049 (N_22049,N_19238,N_17459);
xor U22050 (N_22050,N_15013,N_15355);
and U22051 (N_22051,N_16092,N_17950);
nor U22052 (N_22052,N_17142,N_16188);
or U22053 (N_22053,N_15493,N_17255);
or U22054 (N_22054,N_15319,N_17431);
nor U22055 (N_22055,N_18530,N_19021);
or U22056 (N_22056,N_16928,N_15228);
nor U22057 (N_22057,N_16328,N_16886);
and U22058 (N_22058,N_15745,N_15480);
and U22059 (N_22059,N_17030,N_15765);
nand U22060 (N_22060,N_15722,N_16450);
nor U22061 (N_22061,N_17485,N_19637);
or U22062 (N_22062,N_15907,N_15484);
and U22063 (N_22063,N_16208,N_19027);
xor U22064 (N_22064,N_18844,N_17153);
and U22065 (N_22065,N_19023,N_18614);
or U22066 (N_22066,N_17191,N_15279);
or U22067 (N_22067,N_16848,N_17121);
xnor U22068 (N_22068,N_16257,N_17343);
nor U22069 (N_22069,N_15284,N_16856);
nand U22070 (N_22070,N_19293,N_16742);
and U22071 (N_22071,N_19657,N_16481);
nor U22072 (N_22072,N_18003,N_18092);
and U22073 (N_22073,N_15952,N_16900);
and U22074 (N_22074,N_15033,N_17523);
nor U22075 (N_22075,N_17118,N_17652);
and U22076 (N_22076,N_17054,N_19819);
nor U22077 (N_22077,N_18465,N_15250);
or U22078 (N_22078,N_18234,N_18210);
nor U22079 (N_22079,N_17524,N_17547);
or U22080 (N_22080,N_15763,N_15734);
or U22081 (N_22081,N_17471,N_19897);
and U22082 (N_22082,N_18630,N_15787);
nor U22083 (N_22083,N_15613,N_19600);
nand U22084 (N_22084,N_19272,N_17370);
xnor U22085 (N_22085,N_16927,N_16378);
and U22086 (N_22086,N_18310,N_19256);
or U22087 (N_22087,N_17986,N_16802);
nor U22088 (N_22088,N_16756,N_19518);
nor U22089 (N_22089,N_19976,N_19928);
and U22090 (N_22090,N_15612,N_19608);
nor U22091 (N_22091,N_17533,N_15564);
nand U22092 (N_22092,N_19626,N_17159);
and U22093 (N_22093,N_15458,N_15889);
nand U22094 (N_22094,N_18939,N_19854);
xor U22095 (N_22095,N_16046,N_15481);
nor U22096 (N_22096,N_16720,N_15570);
nor U22097 (N_22097,N_18414,N_18842);
nand U22098 (N_22098,N_17891,N_18071);
or U22099 (N_22099,N_17585,N_16068);
xor U22100 (N_22100,N_15641,N_19447);
and U22101 (N_22101,N_17312,N_17580);
nand U22102 (N_22102,N_18991,N_19527);
and U22103 (N_22103,N_19914,N_17842);
and U22104 (N_22104,N_19369,N_16805);
or U22105 (N_22105,N_16149,N_15577);
nor U22106 (N_22106,N_17155,N_16164);
or U22107 (N_22107,N_16109,N_16915);
and U22108 (N_22108,N_18672,N_15971);
and U22109 (N_22109,N_15826,N_17504);
nor U22110 (N_22110,N_19696,N_18164);
nor U22111 (N_22111,N_19622,N_16239);
or U22112 (N_22112,N_17028,N_17294);
nand U22113 (N_22113,N_19790,N_18057);
and U22114 (N_22114,N_17838,N_15460);
and U22115 (N_22115,N_15227,N_19844);
and U22116 (N_22116,N_17552,N_16619);
nor U22117 (N_22117,N_15867,N_18969);
nor U22118 (N_22118,N_16525,N_18840);
or U22119 (N_22119,N_18123,N_15085);
nand U22120 (N_22120,N_18150,N_18141);
nor U22121 (N_22121,N_16170,N_19173);
nand U22122 (N_22122,N_19279,N_16593);
or U22123 (N_22123,N_16855,N_17709);
xnor U22124 (N_22124,N_17612,N_16840);
and U22125 (N_22125,N_16274,N_15042);
nand U22126 (N_22126,N_16296,N_17458);
and U22127 (N_22127,N_15528,N_18695);
nand U22128 (N_22128,N_19259,N_17967);
nor U22129 (N_22129,N_19761,N_15128);
or U22130 (N_22130,N_16242,N_19949);
or U22131 (N_22131,N_16826,N_16189);
or U22132 (N_22132,N_18203,N_15918);
or U22133 (N_22133,N_17660,N_16145);
or U22134 (N_22134,N_17047,N_19650);
or U22135 (N_22135,N_15149,N_17260);
or U22136 (N_22136,N_18573,N_15880);
or U22137 (N_22137,N_15015,N_15890);
and U22138 (N_22138,N_16416,N_18507);
nand U22139 (N_22139,N_16983,N_16738);
and U22140 (N_22140,N_15983,N_18130);
nor U22141 (N_22141,N_16608,N_17885);
xnor U22142 (N_22142,N_18464,N_19863);
nor U22143 (N_22143,N_18265,N_15017);
nor U22144 (N_22144,N_19895,N_16258);
nor U22145 (N_22145,N_18322,N_17536);
nand U22146 (N_22146,N_19876,N_18200);
or U22147 (N_22147,N_18983,N_16091);
or U22148 (N_22148,N_18149,N_19106);
or U22149 (N_22149,N_15030,N_15770);
nand U22150 (N_22150,N_15710,N_18243);
nand U22151 (N_22151,N_19252,N_16746);
or U22152 (N_22152,N_19485,N_17315);
xnor U22153 (N_22153,N_18748,N_16966);
and U22154 (N_22154,N_18577,N_18943);
nand U22155 (N_22155,N_18205,N_18850);
and U22156 (N_22156,N_16036,N_18426);
nand U22157 (N_22157,N_18434,N_19777);
xor U22158 (N_22158,N_18391,N_16462);
or U22159 (N_22159,N_17098,N_17674);
nand U22160 (N_22160,N_19690,N_18390);
and U22161 (N_22161,N_15975,N_15438);
or U22162 (N_22162,N_19327,N_17380);
nor U22163 (N_22163,N_17507,N_15002);
nor U22164 (N_22164,N_16214,N_17778);
nand U22165 (N_22165,N_16890,N_16581);
or U22166 (N_22166,N_15056,N_18587);
xor U22167 (N_22167,N_17305,N_15397);
or U22168 (N_22168,N_15304,N_19597);
xnor U22169 (N_22169,N_19704,N_18701);
and U22170 (N_22170,N_19066,N_15115);
nand U22171 (N_22171,N_18342,N_19712);
nand U22172 (N_22172,N_17434,N_19443);
nor U22173 (N_22173,N_15823,N_16233);
and U22174 (N_22174,N_15700,N_17415);
or U22175 (N_22175,N_16929,N_18662);
or U22176 (N_22176,N_15116,N_16325);
nor U22177 (N_22177,N_18063,N_19193);
and U22178 (N_22178,N_17638,N_17855);
and U22179 (N_22179,N_19236,N_16984);
nand U22180 (N_22180,N_18088,N_18360);
and U22181 (N_22181,N_18684,N_16009);
and U22182 (N_22182,N_18917,N_18082);
nor U22183 (N_22183,N_16649,N_16363);
nor U22184 (N_22184,N_19022,N_15853);
nor U22185 (N_22185,N_16175,N_15270);
nor U22186 (N_22186,N_15396,N_18190);
and U22187 (N_22187,N_16456,N_16437);
or U22188 (N_22188,N_17757,N_18446);
nor U22189 (N_22189,N_16426,N_18416);
and U22190 (N_22190,N_16447,N_18569);
or U22191 (N_22191,N_19565,N_16888);
or U22192 (N_22192,N_19320,N_18327);
nand U22193 (N_22193,N_15895,N_19057);
nor U22194 (N_22194,N_16849,N_17702);
and U22195 (N_22195,N_15931,N_15421);
and U22196 (N_22196,N_19647,N_19181);
or U22197 (N_22197,N_15394,N_19297);
xnor U22198 (N_22198,N_18750,N_16901);
nand U22199 (N_22199,N_17239,N_17700);
or U22200 (N_22200,N_15608,N_19548);
and U22201 (N_22201,N_15866,N_15576);
nand U22202 (N_22202,N_15059,N_19918);
or U22203 (N_22203,N_15622,N_18362);
and U22204 (N_22204,N_18537,N_17140);
xnor U22205 (N_22205,N_15283,N_17128);
or U22206 (N_22206,N_16654,N_18317);
nand U22207 (N_22207,N_18877,N_17712);
or U22208 (N_22208,N_17490,N_16895);
nand U22209 (N_22209,N_15623,N_16271);
or U22210 (N_22210,N_18397,N_17690);
or U22211 (N_22211,N_16044,N_18540);
or U22212 (N_22212,N_18399,N_17830);
or U22213 (N_22213,N_19411,N_19846);
and U22214 (N_22214,N_18244,N_15222);
or U22215 (N_22215,N_16575,N_18117);
nand U22216 (N_22216,N_15003,N_19492);
or U22217 (N_22217,N_16232,N_15590);
xor U22218 (N_22218,N_19821,N_16737);
or U22219 (N_22219,N_18440,N_19017);
or U22220 (N_22220,N_17156,N_15365);
nor U22221 (N_22221,N_17854,N_15916);
nor U22222 (N_22222,N_19479,N_19786);
or U22223 (N_22223,N_17832,N_19815);
or U22224 (N_22224,N_16663,N_16926);
or U22225 (N_22225,N_15747,N_16825);
and U22226 (N_22226,N_16415,N_18403);
or U22227 (N_22227,N_18486,N_17472);
or U22228 (N_22228,N_17273,N_17634);
and U22229 (N_22229,N_19937,N_19407);
nand U22230 (N_22230,N_18736,N_17519);
and U22231 (N_22231,N_19417,N_19874);
nor U22232 (N_22232,N_17805,N_16579);
or U22233 (N_22233,N_19945,N_17544);
and U22234 (N_22234,N_19208,N_18884);
or U22235 (N_22235,N_15910,N_17769);
or U22236 (N_22236,N_15934,N_16182);
nor U22237 (N_22237,N_18067,N_18584);
or U22238 (N_22238,N_18469,N_19517);
and U22239 (N_22239,N_15882,N_16533);
nand U22240 (N_22240,N_15062,N_17061);
and U22241 (N_22241,N_19715,N_15507);
and U22242 (N_22242,N_15709,N_17303);
or U22243 (N_22243,N_17015,N_16012);
nand U22244 (N_22244,N_15535,N_16285);
or U22245 (N_22245,N_18298,N_15468);
nand U22246 (N_22246,N_18892,N_16956);
nor U22247 (N_22247,N_18783,N_19148);
nor U22248 (N_22248,N_19524,N_18435);
and U22249 (N_22249,N_15835,N_17753);
and U22250 (N_22250,N_17780,N_19708);
nand U22251 (N_22251,N_18124,N_18209);
nand U22252 (N_22252,N_16994,N_17962);
or U22253 (N_22253,N_16297,N_16479);
and U22254 (N_22254,N_17037,N_16389);
nor U22255 (N_22255,N_18659,N_19431);
nand U22256 (N_22256,N_17340,N_15117);
or U22257 (N_22257,N_16225,N_17877);
nor U22258 (N_22258,N_19926,N_19789);
or U22259 (N_22259,N_19123,N_19282);
or U22260 (N_22260,N_15247,N_17095);
or U22261 (N_22261,N_17796,N_16351);
and U22262 (N_22262,N_16866,N_17820);
nand U22263 (N_22263,N_15703,N_19725);
nand U22264 (N_22264,N_18851,N_15393);
and U22265 (N_22265,N_19728,N_16748);
or U22266 (N_22266,N_16934,N_19284);
and U22267 (N_22267,N_19317,N_16906);
nor U22268 (N_22268,N_17414,N_19552);
and U22269 (N_22269,N_16071,N_15969);
or U22270 (N_22270,N_17369,N_16585);
nor U22271 (N_22271,N_16172,N_16228);
xor U22272 (N_22272,N_19081,N_15068);
or U22273 (N_22273,N_17058,N_18646);
or U22274 (N_22274,N_17363,N_17067);
nand U22275 (N_22275,N_19847,N_16810);
nand U22276 (N_22276,N_16020,N_15425);
nand U22277 (N_22277,N_16909,N_16500);
or U22278 (N_22278,N_19553,N_18180);
or U22279 (N_22279,N_17316,N_16111);
nand U22280 (N_22280,N_18512,N_16254);
nor U22281 (N_22281,N_16828,N_17586);
and U22282 (N_22282,N_15503,N_16224);
or U22283 (N_22283,N_17610,N_19954);
nand U22284 (N_22284,N_16779,N_16625);
nor U22285 (N_22285,N_16897,N_16973);
or U22286 (N_22286,N_16173,N_15822);
and U22287 (N_22287,N_18387,N_15628);
and U22288 (N_22288,N_16588,N_15095);
and U22289 (N_22289,N_15216,N_15449);
nor U22290 (N_22290,N_17911,N_17457);
nand U22291 (N_22291,N_15568,N_18260);
nor U22292 (N_22292,N_17167,N_17509);
nor U22293 (N_22293,N_17870,N_15814);
and U22294 (N_22294,N_15191,N_17649);
or U22295 (N_22295,N_18333,N_17973);
nand U22296 (N_22296,N_15492,N_19860);
nor U22297 (N_22297,N_16735,N_18666);
nor U22298 (N_22298,N_16949,N_19727);
xor U22299 (N_22299,N_17035,N_15893);
nand U22300 (N_22300,N_18713,N_19346);
nor U22301 (N_22301,N_18909,N_17022);
or U22302 (N_22302,N_15804,N_15168);
nor U22303 (N_22303,N_15268,N_15185);
and U22304 (N_22304,N_18010,N_17713);
or U22305 (N_22305,N_18076,N_15671);
and U22306 (N_22306,N_18613,N_18620);
nand U22307 (N_22307,N_15295,N_17052);
xnor U22308 (N_22308,N_17374,N_19987);
xnor U22309 (N_22309,N_15760,N_16396);
nand U22310 (N_22310,N_16313,N_17931);
xnor U22311 (N_22311,N_15694,N_19693);
nor U22312 (N_22312,N_18778,N_18456);
or U22313 (N_22313,N_15674,N_19673);
xor U22314 (N_22314,N_18925,N_15439);
nand U22315 (N_22315,N_19739,N_15379);
nand U22316 (N_22316,N_19988,N_19733);
or U22317 (N_22317,N_16482,N_19061);
nor U22318 (N_22318,N_16536,N_17018);
xor U22319 (N_22319,N_19840,N_19648);
nor U22320 (N_22320,N_15280,N_19404);
and U22321 (N_22321,N_16512,N_19707);
or U22322 (N_22322,N_16240,N_18648);
nand U22323 (N_22323,N_16008,N_16561);
and U22324 (N_22324,N_17203,N_18663);
or U22325 (N_22325,N_19307,N_15211);
xor U22326 (N_22326,N_19105,N_18161);
and U22327 (N_22327,N_18607,N_19523);
and U22328 (N_22328,N_15719,N_17527);
or U22329 (N_22329,N_16059,N_15125);
nor U22330 (N_22330,N_16123,N_18051);
xnor U22331 (N_22331,N_17902,N_19955);
or U22332 (N_22332,N_16477,N_19887);
or U22333 (N_22333,N_16410,N_15192);
nor U22334 (N_22334,N_19013,N_17791);
or U22335 (N_22335,N_18098,N_18994);
nor U22336 (N_22336,N_16628,N_19665);
or U22337 (N_22337,N_17689,N_16364);
nor U22338 (N_22338,N_17143,N_16557);
nand U22339 (N_22339,N_19104,N_15672);
nor U22340 (N_22340,N_18307,N_15751);
xnor U22341 (N_22341,N_15036,N_16246);
and U22342 (N_22342,N_16392,N_15474);
and U22343 (N_22343,N_18889,N_17486);
nor U22344 (N_22344,N_15291,N_19429);
nor U22345 (N_22345,N_15147,N_18936);
xor U22346 (N_22346,N_19326,N_15982);
or U22347 (N_22347,N_15790,N_17359);
and U22348 (N_22348,N_17280,N_16715);
and U22349 (N_22349,N_19268,N_17215);
and U22350 (N_22350,N_18374,N_16307);
nand U22351 (N_22351,N_19161,N_16194);
nand U22352 (N_22352,N_15786,N_18827);
and U22353 (N_22353,N_19409,N_15090);
nor U22354 (N_22354,N_18726,N_19461);
nor U22355 (N_22355,N_18267,N_18187);
nor U22356 (N_22356,N_17837,N_17384);
and U22357 (N_22357,N_16348,N_15225);
and U22358 (N_22358,N_16075,N_19711);
nor U22359 (N_22359,N_18714,N_18751);
or U22360 (N_22360,N_19873,N_16391);
or U22361 (N_22361,N_16061,N_19211);
and U22362 (N_22362,N_18380,N_15940);
or U22363 (N_22363,N_15353,N_16870);
xnor U22364 (N_22364,N_18993,N_17659);
nand U22365 (N_22365,N_19356,N_15879);
nor U22366 (N_22366,N_18638,N_17983);
nor U22367 (N_22367,N_19965,N_16179);
or U22368 (N_22368,N_15884,N_19079);
or U22369 (N_22369,N_16562,N_18675);
nand U22370 (N_22370,N_18347,N_15317);
and U22371 (N_22371,N_15508,N_17448);
or U22372 (N_22372,N_16946,N_17824);
or U22373 (N_22373,N_15504,N_16095);
or U22374 (N_22374,N_15019,N_17223);
and U22375 (N_22375,N_17539,N_17879);
nor U22376 (N_22376,N_18073,N_17000);
nor U22377 (N_22377,N_19371,N_16704);
nand U22378 (N_22378,N_18820,N_19065);
and U22379 (N_22379,N_15197,N_15286);
nand U22380 (N_22380,N_19642,N_19917);
nor U22381 (N_22381,N_17635,N_19691);
or U22382 (N_22382,N_17256,N_17801);
nand U22383 (N_22383,N_19405,N_15534);
nor U22384 (N_22384,N_15381,N_18441);
or U22385 (N_22385,N_17208,N_16216);
or U22386 (N_22386,N_16788,N_16645);
nor U22387 (N_22387,N_15749,N_19011);
xor U22388 (N_22388,N_17043,N_15161);
xor U22389 (N_22389,N_16885,N_17489);
nor U22390 (N_22390,N_16215,N_15922);
and U22391 (N_22391,N_16474,N_19946);
and U22392 (N_22392,N_17119,N_18452);
and U22393 (N_22393,N_18986,N_15282);
nor U22394 (N_22394,N_17587,N_16814);
nor U22395 (N_22395,N_18758,N_17407);
xnor U22396 (N_22396,N_18129,N_19615);
or U22397 (N_22397,N_15874,N_16685);
nand U22398 (N_22398,N_16117,N_18272);
or U22399 (N_22399,N_17579,N_19076);
and U22400 (N_22400,N_18905,N_18859);
or U22401 (N_22401,N_18166,N_16658);
nand U22402 (N_22402,N_15847,N_16893);
xnor U22403 (N_22403,N_16932,N_15301);
nand U22404 (N_22404,N_16580,N_16144);
or U22405 (N_22405,N_19818,N_16422);
nand U22406 (N_22406,N_17803,N_15454);
nor U22407 (N_22407,N_16286,N_18539);
xor U22408 (N_22408,N_19540,N_19501);
nand U22409 (N_22409,N_19760,N_16211);
and U22410 (N_22410,N_17432,N_15764);
nor U22411 (N_22411,N_16369,N_15636);
or U22412 (N_22412,N_15505,N_15193);
nand U22413 (N_22413,N_15118,N_19774);
and U22414 (N_22414,N_16559,N_17089);
nand U22415 (N_22415,N_17433,N_19503);
xnor U22416 (N_22416,N_16093,N_18432);
or U22417 (N_22417,N_17731,N_19157);
nand U22418 (N_22418,N_16280,N_17078);
nand U22419 (N_22419,N_15803,N_15958);
or U22420 (N_22420,N_17446,N_16661);
and U22421 (N_22421,N_19859,N_18168);
nor U22422 (N_22422,N_15093,N_18681);
and U22423 (N_22423,N_15417,N_16772);
nand U22424 (N_22424,N_15762,N_19294);
nor U22425 (N_22425,N_15196,N_17528);
or U22426 (N_22426,N_19464,N_19574);
or U22427 (N_22427,N_16226,N_16018);
nor U22428 (N_22428,N_19858,N_17323);
nor U22429 (N_22429,N_18964,N_16377);
xnor U22430 (N_22430,N_19040,N_19187);
and U22431 (N_22431,N_19584,N_16129);
nand U22432 (N_22432,N_15092,N_18929);
nor U22433 (N_22433,N_15347,N_15856);
nor U22434 (N_22434,N_18121,N_15101);
nor U22435 (N_22435,N_17179,N_17245);
nand U22436 (N_22436,N_18375,N_19295);
and U22437 (N_22437,N_16083,N_17901);
or U22438 (N_22438,N_17355,N_15346);
xnor U22439 (N_22439,N_18189,N_19591);
xor U22440 (N_22440,N_18480,N_18318);
nor U22441 (N_22441,N_15157,N_15797);
xor U22442 (N_22442,N_18846,N_19806);
nor U22443 (N_22443,N_15155,N_19005);
and U22444 (N_22444,N_15877,N_15923);
nor U22445 (N_22445,N_18016,N_16781);
nor U22446 (N_22446,N_17477,N_19898);
nand U22447 (N_22447,N_16635,N_19101);
xor U22448 (N_22448,N_15043,N_19770);
nor U22449 (N_22449,N_19427,N_17627);
and U22450 (N_22450,N_15299,N_15114);
and U22451 (N_22451,N_18514,N_18942);
or U22452 (N_22452,N_15370,N_15949);
or U22453 (N_22453,N_16538,N_19036);
or U22454 (N_22454,N_16610,N_19380);
and U22455 (N_22455,N_17009,N_15221);
and U22456 (N_22456,N_18138,N_16532);
or U22457 (N_22457,N_18371,N_19755);
or U22458 (N_22458,N_17097,N_16528);
nor U22459 (N_22459,N_17719,N_18316);
nor U22460 (N_22460,N_15626,N_15296);
or U22461 (N_22461,N_16712,N_16344);
and U22462 (N_22462,N_19886,N_18741);
nor U22463 (N_22463,N_16032,N_19855);
xor U22464 (N_22464,N_15075,N_16970);
nand U22465 (N_22465,N_15400,N_16853);
nor U22466 (N_22466,N_17373,N_17053);
nor U22467 (N_22467,N_15773,N_16087);
xnor U22468 (N_22468,N_19680,N_19861);
or U22469 (N_22469,N_18898,N_15976);
nand U22470 (N_22470,N_18927,N_15993);
or U22471 (N_22471,N_16135,N_18299);
or U22472 (N_22472,N_16013,N_16026);
or U22473 (N_22473,N_19812,N_15171);
and U22474 (N_22474,N_15078,N_19872);
and U22475 (N_22475,N_17935,N_15405);
xnor U22476 (N_22476,N_16298,N_17995);
xnor U22477 (N_22477,N_18328,N_17293);
xnor U22478 (N_22478,N_19359,N_18159);
and U22479 (N_22479,N_15707,N_15491);
xnor U22480 (N_22480,N_17912,N_15701);
or U22481 (N_22481,N_17145,N_16023);
nor U22482 (N_22482,N_16775,N_16399);
xor U22483 (N_22483,N_19589,N_19971);
nor U22484 (N_22484,N_16314,N_19832);
nor U22485 (N_22485,N_17326,N_19030);
or U22486 (N_22486,N_18268,N_16531);
xor U22487 (N_22487,N_15905,N_18436);
or U22488 (N_22488,N_17410,N_15930);
nor U22489 (N_22489,N_18471,N_19684);
and U22490 (N_22490,N_16262,N_17025);
nand U22491 (N_22491,N_15948,N_15096);
and U22492 (N_22492,N_19453,N_16113);
xor U22493 (N_22493,N_17546,N_15788);
or U22494 (N_22494,N_15314,N_19791);
nor U22495 (N_22495,N_17372,N_18482);
nor U22496 (N_22496,N_15545,N_19575);
nand U22497 (N_22497,N_16034,N_19436);
or U22498 (N_22498,N_19617,N_19878);
and U22499 (N_22499,N_19290,N_17079);
nand U22500 (N_22500,N_19862,N_15173);
or U22501 (N_22501,N_16114,N_16365);
and U22502 (N_22502,N_15377,N_16150);
nor U22503 (N_22503,N_19586,N_15687);
nand U22504 (N_22504,N_15021,N_19979);
and U22505 (N_22505,N_15662,N_17794);
nand U22506 (N_22506,N_19947,N_16557);
or U22507 (N_22507,N_19867,N_15482);
and U22508 (N_22508,N_19654,N_19308);
and U22509 (N_22509,N_17356,N_16687);
nand U22510 (N_22510,N_15960,N_15852);
or U22511 (N_22511,N_15907,N_18084);
nand U22512 (N_22512,N_19959,N_19183);
xor U22513 (N_22513,N_15033,N_19101);
or U22514 (N_22514,N_15374,N_16748);
and U22515 (N_22515,N_19142,N_17713);
nor U22516 (N_22516,N_19961,N_15254);
or U22517 (N_22517,N_16975,N_19439);
nor U22518 (N_22518,N_18882,N_18571);
nor U22519 (N_22519,N_19452,N_15161);
nand U22520 (N_22520,N_15621,N_15570);
nor U22521 (N_22521,N_17081,N_19062);
xor U22522 (N_22522,N_15337,N_18514);
or U22523 (N_22523,N_18554,N_19953);
nor U22524 (N_22524,N_18368,N_17354);
or U22525 (N_22525,N_15497,N_16086);
nand U22526 (N_22526,N_18426,N_16381);
nand U22527 (N_22527,N_17730,N_15480);
and U22528 (N_22528,N_18846,N_15431);
or U22529 (N_22529,N_16512,N_16326);
nor U22530 (N_22530,N_16885,N_16906);
nor U22531 (N_22531,N_16325,N_18962);
and U22532 (N_22532,N_16864,N_18384);
nand U22533 (N_22533,N_18894,N_19319);
nand U22534 (N_22534,N_17583,N_17390);
and U22535 (N_22535,N_17490,N_16929);
nor U22536 (N_22536,N_17138,N_17554);
or U22537 (N_22537,N_18918,N_16074);
nand U22538 (N_22538,N_17430,N_17452);
or U22539 (N_22539,N_15417,N_19407);
or U22540 (N_22540,N_15385,N_18869);
or U22541 (N_22541,N_19188,N_16809);
nor U22542 (N_22542,N_15158,N_19846);
xor U22543 (N_22543,N_16036,N_18102);
and U22544 (N_22544,N_15090,N_17346);
nand U22545 (N_22545,N_19747,N_18569);
or U22546 (N_22546,N_16530,N_16366);
nor U22547 (N_22547,N_16499,N_19558);
or U22548 (N_22548,N_15424,N_19657);
and U22549 (N_22549,N_15891,N_16740);
nand U22550 (N_22550,N_15504,N_18909);
or U22551 (N_22551,N_18588,N_18969);
nand U22552 (N_22552,N_18110,N_17464);
or U22553 (N_22553,N_19830,N_18698);
and U22554 (N_22554,N_18379,N_15937);
nand U22555 (N_22555,N_17021,N_19998);
and U22556 (N_22556,N_17326,N_17676);
xor U22557 (N_22557,N_19647,N_16893);
nor U22558 (N_22558,N_17233,N_16725);
and U22559 (N_22559,N_18435,N_19181);
and U22560 (N_22560,N_18173,N_18601);
and U22561 (N_22561,N_18075,N_19326);
nand U22562 (N_22562,N_18441,N_16536);
nand U22563 (N_22563,N_19939,N_19935);
or U22564 (N_22564,N_17315,N_17895);
nor U22565 (N_22565,N_18625,N_16381);
nor U22566 (N_22566,N_17727,N_17584);
nand U22567 (N_22567,N_17741,N_18660);
or U22568 (N_22568,N_15112,N_15338);
and U22569 (N_22569,N_16674,N_16376);
or U22570 (N_22570,N_16242,N_19788);
nor U22571 (N_22571,N_19710,N_19524);
and U22572 (N_22572,N_17063,N_17481);
nor U22573 (N_22573,N_18499,N_19862);
or U22574 (N_22574,N_15880,N_16500);
and U22575 (N_22575,N_19779,N_16106);
and U22576 (N_22576,N_15979,N_19012);
nand U22577 (N_22577,N_15705,N_15234);
nor U22578 (N_22578,N_19183,N_15561);
and U22579 (N_22579,N_18088,N_15508);
and U22580 (N_22580,N_18957,N_19329);
nor U22581 (N_22581,N_17324,N_15996);
nand U22582 (N_22582,N_18582,N_16304);
or U22583 (N_22583,N_17808,N_18855);
and U22584 (N_22584,N_19131,N_17702);
nor U22585 (N_22585,N_19015,N_16336);
xor U22586 (N_22586,N_17101,N_16585);
xnor U22587 (N_22587,N_15192,N_15380);
nand U22588 (N_22588,N_17809,N_19706);
nand U22589 (N_22589,N_16663,N_16817);
and U22590 (N_22590,N_16369,N_18435);
or U22591 (N_22591,N_17529,N_17137);
nand U22592 (N_22592,N_17223,N_15758);
nand U22593 (N_22593,N_15673,N_18685);
nand U22594 (N_22594,N_17779,N_15749);
nor U22595 (N_22595,N_15215,N_17507);
nand U22596 (N_22596,N_19162,N_16987);
and U22597 (N_22597,N_18024,N_19527);
xor U22598 (N_22598,N_17889,N_15734);
or U22599 (N_22599,N_19217,N_15004);
or U22600 (N_22600,N_16233,N_17922);
nand U22601 (N_22601,N_19734,N_18786);
or U22602 (N_22602,N_15209,N_15555);
nand U22603 (N_22603,N_16210,N_17459);
nand U22604 (N_22604,N_16515,N_17443);
nand U22605 (N_22605,N_17090,N_15117);
and U22606 (N_22606,N_17752,N_15112);
or U22607 (N_22607,N_18935,N_15265);
nand U22608 (N_22608,N_19846,N_17071);
or U22609 (N_22609,N_17847,N_17771);
nand U22610 (N_22610,N_17333,N_15735);
nand U22611 (N_22611,N_15574,N_16749);
nor U22612 (N_22612,N_16742,N_17686);
and U22613 (N_22613,N_19651,N_19565);
and U22614 (N_22614,N_15505,N_18869);
and U22615 (N_22615,N_17013,N_19074);
and U22616 (N_22616,N_16148,N_15834);
nor U22617 (N_22617,N_19250,N_15879);
or U22618 (N_22618,N_16348,N_17705);
and U22619 (N_22619,N_15419,N_18463);
or U22620 (N_22620,N_17340,N_15029);
nor U22621 (N_22621,N_16765,N_15000);
nor U22622 (N_22622,N_15129,N_19997);
or U22623 (N_22623,N_17548,N_18400);
or U22624 (N_22624,N_19324,N_17981);
and U22625 (N_22625,N_17337,N_15493);
nor U22626 (N_22626,N_19113,N_17399);
xnor U22627 (N_22627,N_19067,N_17002);
nand U22628 (N_22628,N_15620,N_15630);
nor U22629 (N_22629,N_15871,N_15661);
nor U22630 (N_22630,N_16749,N_18253);
xnor U22631 (N_22631,N_15599,N_18699);
nand U22632 (N_22632,N_19118,N_18516);
nor U22633 (N_22633,N_15909,N_17455);
nor U22634 (N_22634,N_17743,N_15588);
or U22635 (N_22635,N_17587,N_18928);
or U22636 (N_22636,N_15446,N_17750);
nor U22637 (N_22637,N_15159,N_19898);
nand U22638 (N_22638,N_18329,N_16957);
xnor U22639 (N_22639,N_18928,N_16593);
nand U22640 (N_22640,N_18516,N_16516);
xnor U22641 (N_22641,N_17588,N_17070);
nand U22642 (N_22642,N_18939,N_19350);
or U22643 (N_22643,N_16283,N_16281);
and U22644 (N_22644,N_18861,N_15357);
nand U22645 (N_22645,N_16808,N_18344);
or U22646 (N_22646,N_18488,N_19703);
nor U22647 (N_22647,N_17091,N_15984);
and U22648 (N_22648,N_17705,N_16984);
nor U22649 (N_22649,N_17369,N_15305);
or U22650 (N_22650,N_17502,N_16779);
nand U22651 (N_22651,N_16249,N_16497);
nand U22652 (N_22652,N_18649,N_19248);
or U22653 (N_22653,N_15406,N_18306);
nor U22654 (N_22654,N_19262,N_16982);
nand U22655 (N_22655,N_18409,N_17743);
and U22656 (N_22656,N_15835,N_18213);
nor U22657 (N_22657,N_19039,N_19934);
or U22658 (N_22658,N_18129,N_19424);
and U22659 (N_22659,N_19237,N_16797);
or U22660 (N_22660,N_17747,N_18345);
nand U22661 (N_22661,N_18206,N_17126);
nand U22662 (N_22662,N_16479,N_16990);
or U22663 (N_22663,N_15265,N_17685);
and U22664 (N_22664,N_19568,N_15813);
nor U22665 (N_22665,N_16861,N_19747);
and U22666 (N_22666,N_15689,N_19247);
or U22667 (N_22667,N_17044,N_15534);
or U22668 (N_22668,N_19585,N_19084);
and U22669 (N_22669,N_15403,N_15355);
or U22670 (N_22670,N_17619,N_15791);
and U22671 (N_22671,N_18114,N_18223);
nand U22672 (N_22672,N_17432,N_18153);
nor U22673 (N_22673,N_18452,N_15768);
or U22674 (N_22674,N_18757,N_19560);
xnor U22675 (N_22675,N_19311,N_17142);
nand U22676 (N_22676,N_15957,N_15463);
and U22677 (N_22677,N_16367,N_18171);
nor U22678 (N_22678,N_15225,N_15572);
nand U22679 (N_22679,N_18991,N_18344);
and U22680 (N_22680,N_16648,N_16626);
nor U22681 (N_22681,N_19184,N_17016);
nand U22682 (N_22682,N_19094,N_19532);
xor U22683 (N_22683,N_16453,N_16867);
xnor U22684 (N_22684,N_19076,N_17270);
xor U22685 (N_22685,N_15269,N_17167);
xor U22686 (N_22686,N_19305,N_19690);
nand U22687 (N_22687,N_16315,N_18226);
nand U22688 (N_22688,N_18213,N_16413);
or U22689 (N_22689,N_16814,N_19946);
or U22690 (N_22690,N_17983,N_18231);
and U22691 (N_22691,N_17180,N_19535);
nor U22692 (N_22692,N_19194,N_19802);
and U22693 (N_22693,N_16373,N_17521);
and U22694 (N_22694,N_19556,N_19453);
nor U22695 (N_22695,N_15722,N_15713);
or U22696 (N_22696,N_15848,N_16071);
and U22697 (N_22697,N_16736,N_18227);
nor U22698 (N_22698,N_15140,N_16265);
nand U22699 (N_22699,N_19471,N_15534);
nor U22700 (N_22700,N_16928,N_18594);
nand U22701 (N_22701,N_17037,N_16478);
and U22702 (N_22702,N_16394,N_18071);
or U22703 (N_22703,N_17371,N_18063);
nand U22704 (N_22704,N_18080,N_18154);
or U22705 (N_22705,N_15158,N_18750);
nand U22706 (N_22706,N_16225,N_16740);
or U22707 (N_22707,N_16855,N_19417);
xor U22708 (N_22708,N_18941,N_19183);
or U22709 (N_22709,N_18663,N_17302);
or U22710 (N_22710,N_18858,N_18566);
xor U22711 (N_22711,N_16761,N_15213);
nand U22712 (N_22712,N_15248,N_16285);
or U22713 (N_22713,N_15948,N_16048);
nor U22714 (N_22714,N_19243,N_18810);
and U22715 (N_22715,N_18557,N_15344);
nand U22716 (N_22716,N_19241,N_17382);
or U22717 (N_22717,N_18401,N_19099);
nand U22718 (N_22718,N_17440,N_18110);
xor U22719 (N_22719,N_15779,N_18755);
xnor U22720 (N_22720,N_16195,N_18813);
or U22721 (N_22721,N_19021,N_19132);
nand U22722 (N_22722,N_18278,N_19480);
nand U22723 (N_22723,N_15947,N_15508);
nand U22724 (N_22724,N_17190,N_17876);
or U22725 (N_22725,N_17114,N_15823);
nand U22726 (N_22726,N_17409,N_18205);
or U22727 (N_22727,N_18491,N_15659);
nor U22728 (N_22728,N_18673,N_19826);
and U22729 (N_22729,N_15007,N_15728);
nand U22730 (N_22730,N_19594,N_17200);
and U22731 (N_22731,N_15985,N_16833);
or U22732 (N_22732,N_18675,N_18259);
nor U22733 (N_22733,N_15436,N_17413);
nand U22734 (N_22734,N_16402,N_16783);
and U22735 (N_22735,N_17907,N_15838);
xnor U22736 (N_22736,N_16007,N_18065);
nand U22737 (N_22737,N_18698,N_18357);
nor U22738 (N_22738,N_18571,N_19142);
nor U22739 (N_22739,N_18540,N_17580);
nand U22740 (N_22740,N_19231,N_16265);
nor U22741 (N_22741,N_15580,N_15066);
nor U22742 (N_22742,N_18517,N_15501);
nor U22743 (N_22743,N_19726,N_17697);
xor U22744 (N_22744,N_19114,N_17799);
nand U22745 (N_22745,N_17776,N_16930);
and U22746 (N_22746,N_17320,N_17005);
nand U22747 (N_22747,N_15818,N_19466);
and U22748 (N_22748,N_16458,N_15886);
or U22749 (N_22749,N_17858,N_19652);
or U22750 (N_22750,N_15934,N_15594);
nand U22751 (N_22751,N_17681,N_18069);
or U22752 (N_22752,N_16541,N_18947);
or U22753 (N_22753,N_15172,N_18958);
or U22754 (N_22754,N_19238,N_18240);
nand U22755 (N_22755,N_17338,N_16027);
nor U22756 (N_22756,N_18237,N_19854);
or U22757 (N_22757,N_18384,N_16601);
nor U22758 (N_22758,N_18894,N_19671);
nor U22759 (N_22759,N_15737,N_16121);
and U22760 (N_22760,N_17269,N_16182);
or U22761 (N_22761,N_15994,N_17178);
nor U22762 (N_22762,N_18257,N_19597);
nor U22763 (N_22763,N_19605,N_15282);
nor U22764 (N_22764,N_19350,N_19973);
nor U22765 (N_22765,N_17565,N_17002);
and U22766 (N_22766,N_15176,N_18482);
or U22767 (N_22767,N_15246,N_16010);
nand U22768 (N_22768,N_15309,N_17388);
and U22769 (N_22769,N_18498,N_19754);
and U22770 (N_22770,N_18606,N_18104);
nor U22771 (N_22771,N_17966,N_16525);
and U22772 (N_22772,N_17354,N_17323);
nand U22773 (N_22773,N_15862,N_15175);
and U22774 (N_22774,N_16229,N_18797);
nor U22775 (N_22775,N_15411,N_17363);
nor U22776 (N_22776,N_15618,N_16005);
nor U22777 (N_22777,N_19002,N_15565);
xnor U22778 (N_22778,N_18861,N_16634);
nor U22779 (N_22779,N_15281,N_15354);
and U22780 (N_22780,N_17813,N_19856);
or U22781 (N_22781,N_16557,N_18209);
and U22782 (N_22782,N_19171,N_19395);
nand U22783 (N_22783,N_19972,N_15794);
and U22784 (N_22784,N_19835,N_16447);
nor U22785 (N_22785,N_17650,N_16534);
and U22786 (N_22786,N_19903,N_16626);
and U22787 (N_22787,N_19962,N_18366);
nor U22788 (N_22788,N_17513,N_16110);
or U22789 (N_22789,N_17253,N_19463);
nor U22790 (N_22790,N_17440,N_17481);
or U22791 (N_22791,N_15388,N_15336);
or U22792 (N_22792,N_15578,N_18781);
and U22793 (N_22793,N_18164,N_19683);
and U22794 (N_22794,N_18527,N_16062);
nand U22795 (N_22795,N_17830,N_17003);
and U22796 (N_22796,N_17223,N_19947);
nor U22797 (N_22797,N_19076,N_19243);
and U22798 (N_22798,N_19022,N_15192);
nand U22799 (N_22799,N_19177,N_16226);
or U22800 (N_22800,N_16520,N_18932);
and U22801 (N_22801,N_15120,N_19883);
nand U22802 (N_22802,N_16758,N_17739);
or U22803 (N_22803,N_15687,N_19654);
nor U22804 (N_22804,N_19575,N_19265);
nor U22805 (N_22805,N_16451,N_17767);
and U22806 (N_22806,N_18872,N_17429);
xnor U22807 (N_22807,N_16152,N_17531);
nor U22808 (N_22808,N_18196,N_17109);
nand U22809 (N_22809,N_19866,N_18468);
nor U22810 (N_22810,N_15093,N_19857);
nand U22811 (N_22811,N_15490,N_18176);
and U22812 (N_22812,N_16867,N_15833);
and U22813 (N_22813,N_19382,N_19320);
or U22814 (N_22814,N_17319,N_19116);
nand U22815 (N_22815,N_15569,N_16964);
nand U22816 (N_22816,N_19183,N_19097);
and U22817 (N_22817,N_17680,N_17929);
or U22818 (N_22818,N_16037,N_15089);
xor U22819 (N_22819,N_16001,N_17021);
nand U22820 (N_22820,N_17856,N_18911);
and U22821 (N_22821,N_18264,N_16846);
nand U22822 (N_22822,N_16013,N_19977);
nand U22823 (N_22823,N_18509,N_17644);
xnor U22824 (N_22824,N_19025,N_18195);
or U22825 (N_22825,N_15771,N_18290);
nor U22826 (N_22826,N_16533,N_16105);
or U22827 (N_22827,N_15885,N_18445);
and U22828 (N_22828,N_17828,N_16754);
nor U22829 (N_22829,N_15546,N_17026);
and U22830 (N_22830,N_18327,N_17846);
or U22831 (N_22831,N_16602,N_15274);
xnor U22832 (N_22832,N_16539,N_16671);
nor U22833 (N_22833,N_19692,N_17898);
xor U22834 (N_22834,N_16485,N_17477);
nand U22835 (N_22835,N_17290,N_15165);
xnor U22836 (N_22836,N_15179,N_16793);
nand U22837 (N_22837,N_15777,N_16526);
or U22838 (N_22838,N_17416,N_18201);
xor U22839 (N_22839,N_19683,N_17663);
and U22840 (N_22840,N_16293,N_16228);
nor U22841 (N_22841,N_18210,N_15431);
nand U22842 (N_22842,N_15701,N_18802);
nor U22843 (N_22843,N_16348,N_19845);
nand U22844 (N_22844,N_19902,N_19147);
nor U22845 (N_22845,N_18918,N_19169);
and U22846 (N_22846,N_15572,N_16183);
and U22847 (N_22847,N_18604,N_18185);
and U22848 (N_22848,N_15298,N_19681);
xnor U22849 (N_22849,N_17997,N_16835);
or U22850 (N_22850,N_18599,N_18480);
and U22851 (N_22851,N_16257,N_16672);
or U22852 (N_22852,N_17611,N_18097);
xor U22853 (N_22853,N_17850,N_15217);
and U22854 (N_22854,N_19307,N_15537);
nand U22855 (N_22855,N_19255,N_15087);
nor U22856 (N_22856,N_17498,N_15707);
and U22857 (N_22857,N_15343,N_18009);
xor U22858 (N_22858,N_17042,N_15092);
and U22859 (N_22859,N_16992,N_16063);
and U22860 (N_22860,N_15385,N_15450);
or U22861 (N_22861,N_16006,N_18307);
nor U22862 (N_22862,N_19661,N_17566);
nor U22863 (N_22863,N_16333,N_18753);
and U22864 (N_22864,N_19620,N_19473);
and U22865 (N_22865,N_15774,N_17918);
nor U22866 (N_22866,N_18805,N_16162);
or U22867 (N_22867,N_17701,N_18204);
nor U22868 (N_22868,N_18462,N_19230);
and U22869 (N_22869,N_19119,N_18643);
nand U22870 (N_22870,N_19374,N_19997);
or U22871 (N_22871,N_19522,N_16748);
nand U22872 (N_22872,N_16988,N_16902);
or U22873 (N_22873,N_16218,N_19429);
nor U22874 (N_22874,N_17911,N_18796);
and U22875 (N_22875,N_17646,N_16930);
nor U22876 (N_22876,N_18849,N_16933);
nand U22877 (N_22877,N_15926,N_16396);
nand U22878 (N_22878,N_19435,N_19425);
xnor U22879 (N_22879,N_15189,N_15830);
and U22880 (N_22880,N_17380,N_17781);
and U22881 (N_22881,N_17643,N_17375);
or U22882 (N_22882,N_18756,N_18847);
nand U22883 (N_22883,N_18816,N_17232);
or U22884 (N_22884,N_19630,N_15757);
nor U22885 (N_22885,N_17119,N_15547);
nand U22886 (N_22886,N_16120,N_16569);
and U22887 (N_22887,N_19917,N_19130);
or U22888 (N_22888,N_17540,N_15139);
and U22889 (N_22889,N_17717,N_18467);
and U22890 (N_22890,N_19733,N_18630);
nand U22891 (N_22891,N_19430,N_18503);
or U22892 (N_22892,N_19955,N_15814);
or U22893 (N_22893,N_16185,N_15949);
and U22894 (N_22894,N_16956,N_15442);
nor U22895 (N_22895,N_16094,N_19413);
nor U22896 (N_22896,N_19109,N_16467);
or U22897 (N_22897,N_19109,N_16180);
and U22898 (N_22898,N_16146,N_18435);
xnor U22899 (N_22899,N_16969,N_15401);
or U22900 (N_22900,N_15854,N_17026);
nor U22901 (N_22901,N_17655,N_15623);
nor U22902 (N_22902,N_19672,N_17620);
or U22903 (N_22903,N_15011,N_17098);
xnor U22904 (N_22904,N_16101,N_16649);
or U22905 (N_22905,N_19647,N_15558);
nor U22906 (N_22906,N_15364,N_19310);
or U22907 (N_22907,N_19147,N_15130);
or U22908 (N_22908,N_18503,N_18947);
and U22909 (N_22909,N_15592,N_18802);
or U22910 (N_22910,N_18720,N_18669);
and U22911 (N_22911,N_18437,N_19210);
nor U22912 (N_22912,N_18424,N_17535);
nand U22913 (N_22913,N_16954,N_17517);
xnor U22914 (N_22914,N_17106,N_19336);
and U22915 (N_22915,N_15141,N_16455);
or U22916 (N_22916,N_19971,N_18762);
and U22917 (N_22917,N_16113,N_19966);
nor U22918 (N_22918,N_18012,N_18157);
nand U22919 (N_22919,N_17913,N_19356);
or U22920 (N_22920,N_17978,N_19716);
nor U22921 (N_22921,N_17645,N_16756);
or U22922 (N_22922,N_16355,N_19464);
and U22923 (N_22923,N_15964,N_19429);
and U22924 (N_22924,N_17674,N_16991);
and U22925 (N_22925,N_16671,N_16554);
and U22926 (N_22926,N_18635,N_19493);
nand U22927 (N_22927,N_19773,N_18856);
nor U22928 (N_22928,N_18391,N_18874);
nand U22929 (N_22929,N_19160,N_16248);
nor U22930 (N_22930,N_17522,N_19758);
nand U22931 (N_22931,N_15640,N_15022);
and U22932 (N_22932,N_17783,N_17716);
nor U22933 (N_22933,N_16436,N_19343);
or U22934 (N_22934,N_18722,N_16529);
xnor U22935 (N_22935,N_19355,N_18488);
xnor U22936 (N_22936,N_16270,N_18831);
or U22937 (N_22937,N_15315,N_19073);
or U22938 (N_22938,N_19038,N_19356);
nand U22939 (N_22939,N_17061,N_16865);
nand U22940 (N_22940,N_17960,N_15377);
nand U22941 (N_22941,N_19592,N_15809);
nor U22942 (N_22942,N_18177,N_17446);
and U22943 (N_22943,N_15584,N_15933);
and U22944 (N_22944,N_19403,N_16965);
or U22945 (N_22945,N_18420,N_16435);
and U22946 (N_22946,N_17134,N_19089);
nand U22947 (N_22947,N_18237,N_16288);
nand U22948 (N_22948,N_17181,N_16943);
nor U22949 (N_22949,N_17430,N_19136);
nor U22950 (N_22950,N_17095,N_17399);
and U22951 (N_22951,N_19660,N_16037);
and U22952 (N_22952,N_18223,N_19373);
nor U22953 (N_22953,N_18101,N_16523);
and U22954 (N_22954,N_16074,N_15834);
and U22955 (N_22955,N_15055,N_16226);
and U22956 (N_22956,N_15549,N_17334);
or U22957 (N_22957,N_17471,N_17585);
and U22958 (N_22958,N_19109,N_15393);
nand U22959 (N_22959,N_19681,N_16957);
nand U22960 (N_22960,N_16259,N_19945);
nand U22961 (N_22961,N_15483,N_16731);
and U22962 (N_22962,N_15835,N_15731);
or U22963 (N_22963,N_15500,N_17397);
or U22964 (N_22964,N_15580,N_17145);
nand U22965 (N_22965,N_16579,N_19304);
nor U22966 (N_22966,N_18536,N_16174);
or U22967 (N_22967,N_16302,N_17198);
or U22968 (N_22968,N_19623,N_19456);
or U22969 (N_22969,N_18978,N_19865);
or U22970 (N_22970,N_17537,N_18423);
nor U22971 (N_22971,N_16934,N_17186);
nand U22972 (N_22972,N_15496,N_18876);
nand U22973 (N_22973,N_16006,N_15314);
or U22974 (N_22974,N_16758,N_16323);
nand U22975 (N_22975,N_16321,N_18403);
nor U22976 (N_22976,N_17995,N_15133);
or U22977 (N_22977,N_16221,N_18923);
nor U22978 (N_22978,N_15046,N_15281);
nand U22979 (N_22979,N_16511,N_17091);
and U22980 (N_22980,N_15445,N_18995);
nor U22981 (N_22981,N_15327,N_16496);
nand U22982 (N_22982,N_16218,N_18745);
xnor U22983 (N_22983,N_19104,N_15162);
nand U22984 (N_22984,N_16740,N_17944);
or U22985 (N_22985,N_16825,N_15277);
nand U22986 (N_22986,N_15564,N_16312);
and U22987 (N_22987,N_15434,N_17462);
and U22988 (N_22988,N_17264,N_17585);
and U22989 (N_22989,N_16071,N_17973);
and U22990 (N_22990,N_18663,N_15297);
nor U22991 (N_22991,N_19618,N_15156);
xor U22992 (N_22992,N_18211,N_19947);
nand U22993 (N_22993,N_19177,N_16372);
nand U22994 (N_22994,N_15536,N_15338);
xor U22995 (N_22995,N_18778,N_19292);
nor U22996 (N_22996,N_19165,N_16134);
nand U22997 (N_22997,N_17909,N_16478);
nand U22998 (N_22998,N_19300,N_15839);
and U22999 (N_22999,N_16195,N_15696);
or U23000 (N_23000,N_16124,N_18785);
nor U23001 (N_23001,N_18927,N_16038);
and U23002 (N_23002,N_18699,N_16799);
nand U23003 (N_23003,N_18568,N_19870);
nor U23004 (N_23004,N_19225,N_16702);
and U23005 (N_23005,N_19332,N_16608);
nand U23006 (N_23006,N_19317,N_16556);
or U23007 (N_23007,N_18412,N_18420);
nand U23008 (N_23008,N_16509,N_18766);
nor U23009 (N_23009,N_17529,N_15713);
xnor U23010 (N_23010,N_18012,N_18045);
and U23011 (N_23011,N_15955,N_19432);
xnor U23012 (N_23012,N_19453,N_18031);
nand U23013 (N_23013,N_16988,N_18752);
nor U23014 (N_23014,N_17551,N_18416);
and U23015 (N_23015,N_17301,N_15330);
nor U23016 (N_23016,N_16694,N_19096);
or U23017 (N_23017,N_19803,N_19559);
and U23018 (N_23018,N_18916,N_19059);
nand U23019 (N_23019,N_19949,N_19051);
or U23020 (N_23020,N_17142,N_19972);
nand U23021 (N_23021,N_17631,N_18201);
nand U23022 (N_23022,N_15980,N_18586);
nor U23023 (N_23023,N_19067,N_18046);
nor U23024 (N_23024,N_15549,N_17592);
nand U23025 (N_23025,N_17905,N_19107);
nand U23026 (N_23026,N_16935,N_15570);
or U23027 (N_23027,N_18375,N_18875);
or U23028 (N_23028,N_18627,N_18715);
nor U23029 (N_23029,N_15562,N_16602);
nand U23030 (N_23030,N_18520,N_17183);
or U23031 (N_23031,N_17968,N_15959);
xnor U23032 (N_23032,N_15017,N_15999);
and U23033 (N_23033,N_18311,N_15033);
or U23034 (N_23034,N_17207,N_15683);
and U23035 (N_23035,N_16571,N_19851);
nor U23036 (N_23036,N_16484,N_15165);
or U23037 (N_23037,N_16896,N_15707);
and U23038 (N_23038,N_17322,N_15534);
nand U23039 (N_23039,N_17080,N_19770);
nor U23040 (N_23040,N_19236,N_15470);
nor U23041 (N_23041,N_16171,N_18474);
nand U23042 (N_23042,N_17557,N_19445);
or U23043 (N_23043,N_17576,N_18451);
xnor U23044 (N_23044,N_19915,N_16263);
or U23045 (N_23045,N_19277,N_15632);
nand U23046 (N_23046,N_17731,N_19733);
or U23047 (N_23047,N_15194,N_15009);
and U23048 (N_23048,N_19678,N_18300);
nand U23049 (N_23049,N_16729,N_17215);
or U23050 (N_23050,N_18365,N_16157);
and U23051 (N_23051,N_15911,N_17073);
nor U23052 (N_23052,N_16728,N_17463);
or U23053 (N_23053,N_19287,N_18782);
or U23054 (N_23054,N_15738,N_17409);
or U23055 (N_23055,N_19230,N_18846);
or U23056 (N_23056,N_17734,N_18263);
and U23057 (N_23057,N_15977,N_19916);
xor U23058 (N_23058,N_18959,N_16619);
and U23059 (N_23059,N_17650,N_16871);
or U23060 (N_23060,N_18534,N_15152);
or U23061 (N_23061,N_19655,N_15385);
and U23062 (N_23062,N_19195,N_17069);
or U23063 (N_23063,N_16530,N_17176);
or U23064 (N_23064,N_19850,N_19630);
nand U23065 (N_23065,N_19069,N_17780);
nand U23066 (N_23066,N_18632,N_16483);
and U23067 (N_23067,N_15417,N_16803);
or U23068 (N_23068,N_19267,N_18723);
and U23069 (N_23069,N_15899,N_18044);
or U23070 (N_23070,N_17950,N_17830);
nor U23071 (N_23071,N_19936,N_18123);
or U23072 (N_23072,N_18578,N_19721);
or U23073 (N_23073,N_18361,N_18233);
nor U23074 (N_23074,N_18650,N_18538);
or U23075 (N_23075,N_15581,N_16300);
and U23076 (N_23076,N_16374,N_17321);
nand U23077 (N_23077,N_19853,N_16069);
nand U23078 (N_23078,N_18697,N_18308);
nor U23079 (N_23079,N_15127,N_19393);
nand U23080 (N_23080,N_17693,N_17576);
and U23081 (N_23081,N_19585,N_16603);
nand U23082 (N_23082,N_18111,N_15410);
nand U23083 (N_23083,N_18445,N_16451);
nor U23084 (N_23084,N_19200,N_16676);
nor U23085 (N_23085,N_18679,N_19055);
nand U23086 (N_23086,N_19986,N_16707);
nor U23087 (N_23087,N_18523,N_17344);
nor U23088 (N_23088,N_17546,N_19851);
or U23089 (N_23089,N_19047,N_17803);
nor U23090 (N_23090,N_18528,N_17853);
nor U23091 (N_23091,N_17289,N_19615);
and U23092 (N_23092,N_18966,N_19025);
and U23093 (N_23093,N_15836,N_19740);
and U23094 (N_23094,N_16285,N_15267);
or U23095 (N_23095,N_15033,N_18211);
and U23096 (N_23096,N_16674,N_18477);
or U23097 (N_23097,N_17330,N_15772);
nor U23098 (N_23098,N_15858,N_18875);
nand U23099 (N_23099,N_16016,N_15055);
or U23100 (N_23100,N_19291,N_16244);
nor U23101 (N_23101,N_15920,N_15561);
or U23102 (N_23102,N_16625,N_19209);
xnor U23103 (N_23103,N_19017,N_18266);
nor U23104 (N_23104,N_15526,N_17658);
nor U23105 (N_23105,N_18631,N_16304);
and U23106 (N_23106,N_19930,N_18598);
nor U23107 (N_23107,N_18251,N_16261);
nand U23108 (N_23108,N_19957,N_19251);
nor U23109 (N_23109,N_18842,N_17219);
nand U23110 (N_23110,N_15776,N_17826);
nand U23111 (N_23111,N_16659,N_15099);
nand U23112 (N_23112,N_19534,N_17839);
nor U23113 (N_23113,N_15770,N_15540);
nand U23114 (N_23114,N_15065,N_17936);
nor U23115 (N_23115,N_19019,N_17748);
xnor U23116 (N_23116,N_15281,N_17236);
nor U23117 (N_23117,N_15091,N_18730);
and U23118 (N_23118,N_16444,N_17382);
nand U23119 (N_23119,N_17020,N_19587);
and U23120 (N_23120,N_15523,N_16877);
and U23121 (N_23121,N_19689,N_17469);
and U23122 (N_23122,N_16705,N_19702);
nor U23123 (N_23123,N_16342,N_17505);
nor U23124 (N_23124,N_17527,N_16831);
or U23125 (N_23125,N_19689,N_15935);
or U23126 (N_23126,N_15926,N_15804);
and U23127 (N_23127,N_18552,N_18923);
or U23128 (N_23128,N_18409,N_16003);
nand U23129 (N_23129,N_18649,N_17196);
nand U23130 (N_23130,N_19445,N_17011);
nor U23131 (N_23131,N_16304,N_15228);
nor U23132 (N_23132,N_17881,N_18102);
nand U23133 (N_23133,N_19185,N_18635);
and U23134 (N_23134,N_16332,N_17045);
or U23135 (N_23135,N_15404,N_18197);
or U23136 (N_23136,N_15927,N_15129);
and U23137 (N_23137,N_19312,N_18420);
or U23138 (N_23138,N_16875,N_19643);
nand U23139 (N_23139,N_16204,N_19617);
nand U23140 (N_23140,N_15571,N_19097);
and U23141 (N_23141,N_17287,N_15529);
or U23142 (N_23142,N_19079,N_17831);
or U23143 (N_23143,N_19385,N_19688);
or U23144 (N_23144,N_17696,N_19155);
and U23145 (N_23145,N_18462,N_15457);
and U23146 (N_23146,N_15119,N_18225);
or U23147 (N_23147,N_17321,N_17883);
nor U23148 (N_23148,N_16241,N_19373);
nand U23149 (N_23149,N_15615,N_19948);
nand U23150 (N_23150,N_16711,N_15933);
nor U23151 (N_23151,N_15653,N_17359);
or U23152 (N_23152,N_17666,N_18222);
and U23153 (N_23153,N_18490,N_19805);
and U23154 (N_23154,N_16410,N_17920);
nand U23155 (N_23155,N_17884,N_17386);
nand U23156 (N_23156,N_19521,N_17776);
nor U23157 (N_23157,N_18903,N_16305);
or U23158 (N_23158,N_19864,N_16299);
and U23159 (N_23159,N_19065,N_16452);
and U23160 (N_23160,N_19458,N_15265);
nand U23161 (N_23161,N_18502,N_17059);
and U23162 (N_23162,N_15921,N_17205);
nor U23163 (N_23163,N_15101,N_15153);
nor U23164 (N_23164,N_19693,N_15828);
nand U23165 (N_23165,N_15138,N_16686);
nor U23166 (N_23166,N_19355,N_18969);
and U23167 (N_23167,N_15526,N_17413);
or U23168 (N_23168,N_15158,N_18496);
or U23169 (N_23169,N_19598,N_15987);
and U23170 (N_23170,N_15111,N_16752);
or U23171 (N_23171,N_19213,N_15245);
nand U23172 (N_23172,N_17186,N_18961);
and U23173 (N_23173,N_15036,N_16616);
and U23174 (N_23174,N_17800,N_19073);
xor U23175 (N_23175,N_15806,N_17576);
nor U23176 (N_23176,N_15270,N_18110);
or U23177 (N_23177,N_15288,N_18518);
xor U23178 (N_23178,N_19795,N_18903);
nor U23179 (N_23179,N_19147,N_16620);
and U23180 (N_23180,N_17704,N_18537);
or U23181 (N_23181,N_15898,N_16495);
or U23182 (N_23182,N_19609,N_16506);
nor U23183 (N_23183,N_19206,N_19583);
nand U23184 (N_23184,N_15763,N_15482);
xor U23185 (N_23185,N_18169,N_18748);
nand U23186 (N_23186,N_17489,N_18540);
nand U23187 (N_23187,N_15869,N_19580);
nor U23188 (N_23188,N_15229,N_17239);
nand U23189 (N_23189,N_19607,N_15608);
or U23190 (N_23190,N_18032,N_18508);
and U23191 (N_23191,N_17010,N_17331);
nor U23192 (N_23192,N_15684,N_19344);
xnor U23193 (N_23193,N_19434,N_16121);
and U23194 (N_23194,N_16828,N_19016);
nor U23195 (N_23195,N_17278,N_16920);
nor U23196 (N_23196,N_15471,N_15104);
nand U23197 (N_23197,N_15527,N_16920);
or U23198 (N_23198,N_17828,N_16429);
nand U23199 (N_23199,N_15249,N_17671);
nor U23200 (N_23200,N_17896,N_17856);
nand U23201 (N_23201,N_19488,N_19557);
nand U23202 (N_23202,N_15586,N_15378);
or U23203 (N_23203,N_17777,N_19149);
and U23204 (N_23204,N_17734,N_15250);
nand U23205 (N_23205,N_16138,N_16312);
xnor U23206 (N_23206,N_16565,N_17922);
xor U23207 (N_23207,N_17680,N_17375);
and U23208 (N_23208,N_15968,N_18785);
and U23209 (N_23209,N_16127,N_15980);
nor U23210 (N_23210,N_18000,N_18617);
nand U23211 (N_23211,N_16265,N_19149);
nand U23212 (N_23212,N_16205,N_17708);
xnor U23213 (N_23213,N_17976,N_16701);
nand U23214 (N_23214,N_16479,N_19146);
or U23215 (N_23215,N_18272,N_16614);
nor U23216 (N_23216,N_15325,N_16126);
nor U23217 (N_23217,N_17443,N_16067);
and U23218 (N_23218,N_15513,N_17706);
or U23219 (N_23219,N_16290,N_19806);
and U23220 (N_23220,N_18315,N_18321);
or U23221 (N_23221,N_16654,N_19439);
nand U23222 (N_23222,N_17682,N_15940);
nand U23223 (N_23223,N_18707,N_18322);
and U23224 (N_23224,N_18060,N_19987);
nand U23225 (N_23225,N_19692,N_17680);
nor U23226 (N_23226,N_17135,N_16479);
nor U23227 (N_23227,N_15267,N_19449);
nand U23228 (N_23228,N_15439,N_18780);
xor U23229 (N_23229,N_19536,N_18057);
or U23230 (N_23230,N_19970,N_18241);
and U23231 (N_23231,N_16961,N_15689);
xor U23232 (N_23232,N_19345,N_17272);
or U23233 (N_23233,N_19996,N_19843);
or U23234 (N_23234,N_18615,N_17755);
nor U23235 (N_23235,N_19994,N_19059);
nand U23236 (N_23236,N_15634,N_18047);
xor U23237 (N_23237,N_15809,N_19413);
or U23238 (N_23238,N_16999,N_17758);
and U23239 (N_23239,N_16891,N_16083);
nor U23240 (N_23240,N_17244,N_16286);
nand U23241 (N_23241,N_15706,N_18700);
or U23242 (N_23242,N_19763,N_16840);
and U23243 (N_23243,N_17984,N_15198);
and U23244 (N_23244,N_16623,N_19385);
nand U23245 (N_23245,N_18138,N_16339);
nor U23246 (N_23246,N_19879,N_18053);
nand U23247 (N_23247,N_17896,N_16817);
nand U23248 (N_23248,N_18964,N_18931);
xor U23249 (N_23249,N_19029,N_19178);
nand U23250 (N_23250,N_16486,N_15624);
or U23251 (N_23251,N_17405,N_16084);
xor U23252 (N_23252,N_19713,N_17029);
and U23253 (N_23253,N_17108,N_16421);
nor U23254 (N_23254,N_19893,N_15136);
or U23255 (N_23255,N_16685,N_18579);
nand U23256 (N_23256,N_19642,N_18657);
nand U23257 (N_23257,N_17780,N_18670);
or U23258 (N_23258,N_18750,N_15237);
xor U23259 (N_23259,N_18329,N_19286);
nand U23260 (N_23260,N_15140,N_16285);
or U23261 (N_23261,N_17893,N_19647);
nand U23262 (N_23262,N_15390,N_19524);
or U23263 (N_23263,N_15731,N_16845);
or U23264 (N_23264,N_18963,N_15646);
nand U23265 (N_23265,N_18292,N_16478);
nand U23266 (N_23266,N_15778,N_15256);
and U23267 (N_23267,N_16701,N_17394);
nor U23268 (N_23268,N_17565,N_16892);
and U23269 (N_23269,N_15862,N_15130);
or U23270 (N_23270,N_19420,N_15187);
and U23271 (N_23271,N_16493,N_18655);
and U23272 (N_23272,N_19809,N_15427);
nor U23273 (N_23273,N_18181,N_19659);
and U23274 (N_23274,N_15872,N_16911);
and U23275 (N_23275,N_16101,N_19624);
or U23276 (N_23276,N_16426,N_19681);
nand U23277 (N_23277,N_15073,N_17888);
nor U23278 (N_23278,N_16312,N_19825);
nor U23279 (N_23279,N_17832,N_15361);
or U23280 (N_23280,N_17893,N_15151);
or U23281 (N_23281,N_18091,N_17754);
nand U23282 (N_23282,N_16940,N_17923);
nor U23283 (N_23283,N_17908,N_19942);
nor U23284 (N_23284,N_18570,N_17547);
nand U23285 (N_23285,N_18203,N_17059);
and U23286 (N_23286,N_18292,N_18964);
or U23287 (N_23287,N_16836,N_17362);
xnor U23288 (N_23288,N_19687,N_17806);
xor U23289 (N_23289,N_19685,N_15645);
xnor U23290 (N_23290,N_16521,N_18364);
nand U23291 (N_23291,N_18034,N_18915);
or U23292 (N_23292,N_19816,N_17840);
nor U23293 (N_23293,N_18007,N_17013);
xnor U23294 (N_23294,N_16637,N_18970);
and U23295 (N_23295,N_16364,N_15184);
nand U23296 (N_23296,N_19811,N_17953);
or U23297 (N_23297,N_16870,N_19837);
or U23298 (N_23298,N_18598,N_17420);
nand U23299 (N_23299,N_15504,N_18149);
nand U23300 (N_23300,N_16457,N_19440);
nor U23301 (N_23301,N_18798,N_17775);
nor U23302 (N_23302,N_17814,N_15447);
or U23303 (N_23303,N_19620,N_16164);
xor U23304 (N_23304,N_17209,N_19583);
and U23305 (N_23305,N_15989,N_16443);
or U23306 (N_23306,N_16247,N_17331);
nor U23307 (N_23307,N_18754,N_18373);
nor U23308 (N_23308,N_15500,N_18811);
nand U23309 (N_23309,N_15761,N_17971);
and U23310 (N_23310,N_16176,N_17635);
or U23311 (N_23311,N_16607,N_18944);
or U23312 (N_23312,N_17324,N_19917);
and U23313 (N_23313,N_17358,N_17252);
and U23314 (N_23314,N_17502,N_15382);
nand U23315 (N_23315,N_15090,N_16903);
and U23316 (N_23316,N_19208,N_15950);
xor U23317 (N_23317,N_17951,N_17612);
or U23318 (N_23318,N_15664,N_15229);
nor U23319 (N_23319,N_19409,N_16392);
or U23320 (N_23320,N_18014,N_19630);
or U23321 (N_23321,N_19697,N_18797);
xor U23322 (N_23322,N_15288,N_18457);
nand U23323 (N_23323,N_17246,N_15826);
or U23324 (N_23324,N_15195,N_19473);
xnor U23325 (N_23325,N_16378,N_19652);
nand U23326 (N_23326,N_16225,N_16055);
nand U23327 (N_23327,N_16278,N_18102);
nor U23328 (N_23328,N_19404,N_18189);
and U23329 (N_23329,N_18327,N_17473);
xnor U23330 (N_23330,N_18055,N_19597);
and U23331 (N_23331,N_18053,N_17898);
or U23332 (N_23332,N_19198,N_19448);
nand U23333 (N_23333,N_18164,N_15469);
and U23334 (N_23334,N_17915,N_15958);
nor U23335 (N_23335,N_16652,N_17350);
nand U23336 (N_23336,N_17677,N_18412);
or U23337 (N_23337,N_15380,N_15877);
or U23338 (N_23338,N_15590,N_18879);
nor U23339 (N_23339,N_19817,N_18861);
nand U23340 (N_23340,N_16181,N_18775);
or U23341 (N_23341,N_16168,N_16907);
or U23342 (N_23342,N_15825,N_18670);
nand U23343 (N_23343,N_19111,N_19809);
nand U23344 (N_23344,N_17368,N_15232);
or U23345 (N_23345,N_17972,N_19574);
and U23346 (N_23346,N_17086,N_19998);
xor U23347 (N_23347,N_16042,N_17286);
or U23348 (N_23348,N_17408,N_19467);
xor U23349 (N_23349,N_17582,N_15837);
and U23350 (N_23350,N_15446,N_19433);
or U23351 (N_23351,N_19777,N_15679);
nor U23352 (N_23352,N_17896,N_19764);
nor U23353 (N_23353,N_16220,N_19763);
or U23354 (N_23354,N_18468,N_15808);
nor U23355 (N_23355,N_18754,N_19703);
and U23356 (N_23356,N_15704,N_19407);
nand U23357 (N_23357,N_15877,N_18236);
nor U23358 (N_23358,N_19305,N_18158);
and U23359 (N_23359,N_18613,N_19071);
or U23360 (N_23360,N_19138,N_16148);
nand U23361 (N_23361,N_16987,N_16584);
or U23362 (N_23362,N_15471,N_17496);
and U23363 (N_23363,N_16384,N_15107);
nor U23364 (N_23364,N_16546,N_15328);
nand U23365 (N_23365,N_18125,N_19940);
or U23366 (N_23366,N_16553,N_19532);
nand U23367 (N_23367,N_16591,N_17340);
nor U23368 (N_23368,N_15218,N_19302);
nand U23369 (N_23369,N_16933,N_17365);
nor U23370 (N_23370,N_15805,N_15848);
xor U23371 (N_23371,N_19631,N_17543);
or U23372 (N_23372,N_19560,N_19479);
xnor U23373 (N_23373,N_18157,N_18990);
nand U23374 (N_23374,N_17638,N_16250);
or U23375 (N_23375,N_19457,N_15816);
nand U23376 (N_23376,N_16254,N_19090);
and U23377 (N_23377,N_18852,N_15368);
nand U23378 (N_23378,N_16657,N_16117);
nand U23379 (N_23379,N_16672,N_16436);
xor U23380 (N_23380,N_15071,N_16564);
nand U23381 (N_23381,N_19389,N_15748);
or U23382 (N_23382,N_19620,N_18297);
xor U23383 (N_23383,N_15145,N_15747);
or U23384 (N_23384,N_17031,N_16531);
nand U23385 (N_23385,N_17517,N_19771);
and U23386 (N_23386,N_16572,N_17200);
or U23387 (N_23387,N_18470,N_18788);
and U23388 (N_23388,N_16547,N_19101);
nor U23389 (N_23389,N_19621,N_19455);
nand U23390 (N_23390,N_17627,N_15662);
nor U23391 (N_23391,N_17456,N_18575);
and U23392 (N_23392,N_15324,N_18209);
or U23393 (N_23393,N_18482,N_15517);
xor U23394 (N_23394,N_17350,N_17062);
or U23395 (N_23395,N_15171,N_19995);
or U23396 (N_23396,N_19715,N_19868);
nand U23397 (N_23397,N_19129,N_16101);
nand U23398 (N_23398,N_15546,N_15389);
or U23399 (N_23399,N_17356,N_17332);
nor U23400 (N_23400,N_18416,N_15051);
nand U23401 (N_23401,N_16350,N_17916);
nand U23402 (N_23402,N_16402,N_16471);
nor U23403 (N_23403,N_17742,N_18748);
nand U23404 (N_23404,N_16337,N_18511);
and U23405 (N_23405,N_17560,N_19731);
nand U23406 (N_23406,N_16646,N_17178);
nand U23407 (N_23407,N_18440,N_18829);
or U23408 (N_23408,N_16158,N_16656);
xnor U23409 (N_23409,N_17315,N_15438);
and U23410 (N_23410,N_18913,N_15704);
or U23411 (N_23411,N_15311,N_19925);
and U23412 (N_23412,N_19188,N_17756);
and U23413 (N_23413,N_19959,N_19111);
and U23414 (N_23414,N_18434,N_17516);
nor U23415 (N_23415,N_18941,N_17108);
nor U23416 (N_23416,N_15294,N_16805);
nor U23417 (N_23417,N_17497,N_17300);
and U23418 (N_23418,N_19615,N_16903);
nand U23419 (N_23419,N_18681,N_18369);
nor U23420 (N_23420,N_17069,N_17614);
nand U23421 (N_23421,N_17485,N_19255);
and U23422 (N_23422,N_15175,N_17525);
xnor U23423 (N_23423,N_15528,N_15392);
and U23424 (N_23424,N_18526,N_16030);
xnor U23425 (N_23425,N_18867,N_17410);
and U23426 (N_23426,N_19995,N_18285);
and U23427 (N_23427,N_19706,N_19722);
nand U23428 (N_23428,N_19940,N_15201);
and U23429 (N_23429,N_17150,N_17919);
nor U23430 (N_23430,N_18072,N_16357);
xnor U23431 (N_23431,N_15702,N_19311);
xnor U23432 (N_23432,N_19081,N_15395);
xor U23433 (N_23433,N_15281,N_19279);
xnor U23434 (N_23434,N_18731,N_19544);
nor U23435 (N_23435,N_15631,N_16891);
nor U23436 (N_23436,N_16932,N_15556);
nand U23437 (N_23437,N_17799,N_15574);
and U23438 (N_23438,N_15730,N_16862);
nand U23439 (N_23439,N_15447,N_17841);
nor U23440 (N_23440,N_16409,N_18641);
and U23441 (N_23441,N_18911,N_18848);
or U23442 (N_23442,N_19609,N_19036);
and U23443 (N_23443,N_19443,N_17679);
nor U23444 (N_23444,N_17586,N_19390);
nand U23445 (N_23445,N_15096,N_15479);
or U23446 (N_23446,N_15518,N_18508);
and U23447 (N_23447,N_16122,N_15375);
nand U23448 (N_23448,N_16119,N_18743);
or U23449 (N_23449,N_19140,N_16113);
xnor U23450 (N_23450,N_16142,N_17673);
and U23451 (N_23451,N_18202,N_18789);
nor U23452 (N_23452,N_15704,N_19017);
or U23453 (N_23453,N_16068,N_15937);
nand U23454 (N_23454,N_18434,N_16146);
nand U23455 (N_23455,N_19339,N_17264);
or U23456 (N_23456,N_19804,N_17785);
and U23457 (N_23457,N_18261,N_15971);
xor U23458 (N_23458,N_16207,N_19457);
or U23459 (N_23459,N_19105,N_18960);
xnor U23460 (N_23460,N_19567,N_16672);
or U23461 (N_23461,N_16327,N_15470);
nand U23462 (N_23462,N_19749,N_17409);
and U23463 (N_23463,N_19442,N_16770);
nor U23464 (N_23464,N_15883,N_17326);
and U23465 (N_23465,N_17516,N_18105);
nand U23466 (N_23466,N_15839,N_19323);
nor U23467 (N_23467,N_17800,N_19865);
xnor U23468 (N_23468,N_17041,N_17555);
nand U23469 (N_23469,N_17528,N_17544);
or U23470 (N_23470,N_15127,N_18314);
nand U23471 (N_23471,N_18403,N_17536);
nor U23472 (N_23472,N_18281,N_18176);
nand U23473 (N_23473,N_18877,N_16614);
and U23474 (N_23474,N_18916,N_16291);
nand U23475 (N_23475,N_17797,N_19355);
nand U23476 (N_23476,N_19699,N_17505);
or U23477 (N_23477,N_15859,N_16540);
nor U23478 (N_23478,N_15542,N_18797);
nand U23479 (N_23479,N_19350,N_18258);
nand U23480 (N_23480,N_16467,N_18107);
nor U23481 (N_23481,N_17074,N_16476);
or U23482 (N_23482,N_16556,N_15510);
or U23483 (N_23483,N_17982,N_18779);
or U23484 (N_23484,N_16626,N_18915);
or U23485 (N_23485,N_17551,N_19373);
nand U23486 (N_23486,N_15431,N_17586);
xor U23487 (N_23487,N_15781,N_19207);
nand U23488 (N_23488,N_18322,N_15923);
or U23489 (N_23489,N_15780,N_19017);
and U23490 (N_23490,N_17469,N_16076);
and U23491 (N_23491,N_16024,N_17357);
and U23492 (N_23492,N_18180,N_15244);
nor U23493 (N_23493,N_18374,N_16652);
and U23494 (N_23494,N_15677,N_16857);
nand U23495 (N_23495,N_15175,N_19792);
or U23496 (N_23496,N_15460,N_15311);
and U23497 (N_23497,N_17663,N_18666);
nand U23498 (N_23498,N_19439,N_18693);
nand U23499 (N_23499,N_17651,N_16928);
xnor U23500 (N_23500,N_16744,N_15605);
nor U23501 (N_23501,N_17466,N_15299);
or U23502 (N_23502,N_16913,N_17774);
and U23503 (N_23503,N_18338,N_18054);
nand U23504 (N_23504,N_19731,N_16555);
or U23505 (N_23505,N_15615,N_16661);
and U23506 (N_23506,N_15712,N_16819);
and U23507 (N_23507,N_15360,N_16287);
nand U23508 (N_23508,N_16168,N_17771);
or U23509 (N_23509,N_17446,N_16872);
nand U23510 (N_23510,N_16640,N_15377);
nand U23511 (N_23511,N_15043,N_16854);
xnor U23512 (N_23512,N_16368,N_19141);
nand U23513 (N_23513,N_15978,N_18852);
or U23514 (N_23514,N_15363,N_19610);
nor U23515 (N_23515,N_18306,N_16496);
or U23516 (N_23516,N_19140,N_15186);
nor U23517 (N_23517,N_17655,N_17736);
nor U23518 (N_23518,N_18758,N_16932);
or U23519 (N_23519,N_15548,N_17384);
and U23520 (N_23520,N_17230,N_17747);
and U23521 (N_23521,N_18235,N_17374);
nand U23522 (N_23522,N_19893,N_17157);
nor U23523 (N_23523,N_15342,N_15980);
xnor U23524 (N_23524,N_16201,N_16799);
or U23525 (N_23525,N_15819,N_16984);
xor U23526 (N_23526,N_15384,N_18559);
nand U23527 (N_23527,N_17150,N_16648);
nor U23528 (N_23528,N_17024,N_15120);
and U23529 (N_23529,N_17597,N_18432);
or U23530 (N_23530,N_15482,N_16408);
xor U23531 (N_23531,N_17158,N_19696);
nand U23532 (N_23532,N_19836,N_17112);
nor U23533 (N_23533,N_18424,N_16672);
xor U23534 (N_23534,N_15407,N_17204);
and U23535 (N_23535,N_15647,N_17482);
or U23536 (N_23536,N_15084,N_19962);
nand U23537 (N_23537,N_18027,N_16731);
nor U23538 (N_23538,N_19226,N_18892);
nor U23539 (N_23539,N_17086,N_16819);
or U23540 (N_23540,N_18387,N_15306);
and U23541 (N_23541,N_18458,N_17065);
nand U23542 (N_23542,N_19643,N_16315);
nand U23543 (N_23543,N_15640,N_19290);
nand U23544 (N_23544,N_19858,N_15039);
nor U23545 (N_23545,N_18469,N_17544);
and U23546 (N_23546,N_19885,N_18818);
nor U23547 (N_23547,N_17724,N_15216);
nor U23548 (N_23548,N_16636,N_17458);
nor U23549 (N_23549,N_19492,N_19558);
or U23550 (N_23550,N_15879,N_16250);
nand U23551 (N_23551,N_15985,N_15799);
or U23552 (N_23552,N_15076,N_19912);
and U23553 (N_23553,N_17583,N_19205);
xor U23554 (N_23554,N_16215,N_16824);
or U23555 (N_23555,N_16944,N_17502);
or U23556 (N_23556,N_16175,N_17501);
nand U23557 (N_23557,N_16391,N_18184);
or U23558 (N_23558,N_17347,N_17666);
nor U23559 (N_23559,N_15141,N_16797);
or U23560 (N_23560,N_16360,N_17503);
and U23561 (N_23561,N_15586,N_18401);
and U23562 (N_23562,N_15448,N_17500);
nand U23563 (N_23563,N_17942,N_18476);
and U23564 (N_23564,N_15040,N_16517);
and U23565 (N_23565,N_17025,N_15178);
and U23566 (N_23566,N_17061,N_15153);
nor U23567 (N_23567,N_17783,N_15099);
nor U23568 (N_23568,N_18760,N_18754);
or U23569 (N_23569,N_18309,N_15721);
nor U23570 (N_23570,N_17516,N_19743);
xnor U23571 (N_23571,N_16880,N_19845);
or U23572 (N_23572,N_17645,N_15165);
nand U23573 (N_23573,N_18299,N_15204);
nor U23574 (N_23574,N_19288,N_18112);
and U23575 (N_23575,N_17569,N_15907);
or U23576 (N_23576,N_17230,N_19429);
nand U23577 (N_23577,N_18078,N_18200);
or U23578 (N_23578,N_15434,N_19526);
xor U23579 (N_23579,N_19368,N_17777);
nand U23580 (N_23580,N_18628,N_15755);
nor U23581 (N_23581,N_19807,N_18658);
nor U23582 (N_23582,N_18563,N_18957);
nand U23583 (N_23583,N_17216,N_18578);
or U23584 (N_23584,N_15590,N_17955);
nand U23585 (N_23585,N_17349,N_15986);
nand U23586 (N_23586,N_17347,N_17284);
nor U23587 (N_23587,N_18072,N_17128);
nor U23588 (N_23588,N_19917,N_16553);
nand U23589 (N_23589,N_17929,N_18226);
nand U23590 (N_23590,N_18444,N_16377);
or U23591 (N_23591,N_18962,N_16153);
nor U23592 (N_23592,N_18220,N_15970);
nand U23593 (N_23593,N_16595,N_16498);
nor U23594 (N_23594,N_17709,N_16180);
nor U23595 (N_23595,N_16719,N_15349);
and U23596 (N_23596,N_17488,N_16652);
nand U23597 (N_23597,N_16472,N_18560);
nor U23598 (N_23598,N_17561,N_17343);
nor U23599 (N_23599,N_16425,N_19153);
xor U23600 (N_23600,N_19671,N_17327);
nor U23601 (N_23601,N_18109,N_17260);
nand U23602 (N_23602,N_16415,N_16945);
or U23603 (N_23603,N_18515,N_16971);
or U23604 (N_23604,N_18959,N_16955);
nand U23605 (N_23605,N_18990,N_15485);
nor U23606 (N_23606,N_15278,N_17478);
nand U23607 (N_23607,N_19361,N_19058);
nor U23608 (N_23608,N_19538,N_17954);
nor U23609 (N_23609,N_16466,N_15920);
or U23610 (N_23610,N_15500,N_15699);
or U23611 (N_23611,N_15613,N_15492);
nor U23612 (N_23612,N_16735,N_18178);
xnor U23613 (N_23613,N_17262,N_15303);
or U23614 (N_23614,N_15627,N_16262);
nor U23615 (N_23615,N_16726,N_16583);
and U23616 (N_23616,N_18717,N_15875);
nor U23617 (N_23617,N_16347,N_19658);
nor U23618 (N_23618,N_17172,N_17956);
or U23619 (N_23619,N_15107,N_15321);
or U23620 (N_23620,N_16061,N_18649);
and U23621 (N_23621,N_15945,N_19873);
and U23622 (N_23622,N_19666,N_16857);
or U23623 (N_23623,N_16025,N_16801);
or U23624 (N_23624,N_18797,N_19196);
or U23625 (N_23625,N_15714,N_18573);
nor U23626 (N_23626,N_15945,N_16894);
nand U23627 (N_23627,N_18557,N_17041);
nor U23628 (N_23628,N_18619,N_18512);
nand U23629 (N_23629,N_16785,N_15975);
xnor U23630 (N_23630,N_18395,N_17336);
nand U23631 (N_23631,N_19423,N_16321);
and U23632 (N_23632,N_16050,N_17623);
xor U23633 (N_23633,N_16154,N_15849);
or U23634 (N_23634,N_17423,N_18599);
or U23635 (N_23635,N_18209,N_19513);
and U23636 (N_23636,N_19762,N_16926);
or U23637 (N_23637,N_15428,N_16294);
or U23638 (N_23638,N_17307,N_16202);
or U23639 (N_23639,N_16021,N_19087);
nand U23640 (N_23640,N_17142,N_17972);
nand U23641 (N_23641,N_17912,N_16518);
and U23642 (N_23642,N_18505,N_19086);
or U23643 (N_23643,N_17510,N_18727);
xor U23644 (N_23644,N_15870,N_17871);
nor U23645 (N_23645,N_17508,N_19941);
and U23646 (N_23646,N_19003,N_18072);
and U23647 (N_23647,N_19056,N_15678);
or U23648 (N_23648,N_18453,N_17721);
xnor U23649 (N_23649,N_16344,N_18078);
or U23650 (N_23650,N_17042,N_18262);
and U23651 (N_23651,N_19386,N_18104);
xnor U23652 (N_23652,N_15144,N_16000);
and U23653 (N_23653,N_16363,N_17170);
and U23654 (N_23654,N_17911,N_19576);
nor U23655 (N_23655,N_17630,N_16111);
nor U23656 (N_23656,N_15089,N_19148);
xnor U23657 (N_23657,N_16394,N_16534);
nand U23658 (N_23658,N_15178,N_17820);
and U23659 (N_23659,N_17461,N_16193);
or U23660 (N_23660,N_15603,N_18235);
nand U23661 (N_23661,N_19033,N_15395);
nor U23662 (N_23662,N_15817,N_17028);
and U23663 (N_23663,N_18092,N_15944);
nor U23664 (N_23664,N_17376,N_16421);
nand U23665 (N_23665,N_16191,N_19423);
or U23666 (N_23666,N_19643,N_15184);
nand U23667 (N_23667,N_19651,N_18514);
and U23668 (N_23668,N_16139,N_17538);
or U23669 (N_23669,N_19217,N_17481);
nand U23670 (N_23670,N_16769,N_18224);
nor U23671 (N_23671,N_17726,N_15391);
and U23672 (N_23672,N_17581,N_17999);
or U23673 (N_23673,N_16922,N_17119);
nor U23674 (N_23674,N_19292,N_15155);
or U23675 (N_23675,N_19661,N_16020);
or U23676 (N_23676,N_17827,N_17447);
nor U23677 (N_23677,N_17564,N_18881);
nand U23678 (N_23678,N_17131,N_16767);
and U23679 (N_23679,N_15738,N_19563);
or U23680 (N_23680,N_15998,N_16235);
nor U23681 (N_23681,N_17101,N_16349);
nor U23682 (N_23682,N_17551,N_15290);
and U23683 (N_23683,N_15102,N_17660);
and U23684 (N_23684,N_19276,N_15852);
or U23685 (N_23685,N_19509,N_19014);
xnor U23686 (N_23686,N_16100,N_18898);
nor U23687 (N_23687,N_19964,N_18212);
nor U23688 (N_23688,N_16247,N_17274);
nor U23689 (N_23689,N_16854,N_18020);
or U23690 (N_23690,N_16020,N_15770);
nand U23691 (N_23691,N_17335,N_15490);
or U23692 (N_23692,N_19048,N_15497);
nor U23693 (N_23693,N_18554,N_19122);
nor U23694 (N_23694,N_16093,N_18984);
or U23695 (N_23695,N_18834,N_18816);
and U23696 (N_23696,N_15227,N_19902);
nor U23697 (N_23697,N_19837,N_19056);
or U23698 (N_23698,N_15806,N_18295);
or U23699 (N_23699,N_15042,N_15948);
nor U23700 (N_23700,N_19191,N_19349);
nor U23701 (N_23701,N_17345,N_17524);
and U23702 (N_23702,N_16646,N_17733);
or U23703 (N_23703,N_18825,N_16573);
nor U23704 (N_23704,N_16548,N_15058);
nor U23705 (N_23705,N_15796,N_16560);
or U23706 (N_23706,N_19276,N_15085);
nand U23707 (N_23707,N_18766,N_16719);
and U23708 (N_23708,N_19161,N_16509);
or U23709 (N_23709,N_19997,N_17688);
or U23710 (N_23710,N_16248,N_16127);
or U23711 (N_23711,N_17893,N_16701);
xor U23712 (N_23712,N_15818,N_16545);
and U23713 (N_23713,N_18351,N_17357);
xnor U23714 (N_23714,N_19201,N_16427);
nand U23715 (N_23715,N_15077,N_17207);
xor U23716 (N_23716,N_15764,N_17799);
nand U23717 (N_23717,N_17368,N_18607);
or U23718 (N_23718,N_17101,N_16960);
and U23719 (N_23719,N_17957,N_17200);
nor U23720 (N_23720,N_19176,N_18607);
xnor U23721 (N_23721,N_16354,N_18254);
nand U23722 (N_23722,N_17284,N_16357);
or U23723 (N_23723,N_16484,N_18468);
nand U23724 (N_23724,N_17165,N_19128);
nand U23725 (N_23725,N_15167,N_19370);
and U23726 (N_23726,N_16425,N_15889);
or U23727 (N_23727,N_18547,N_16944);
nor U23728 (N_23728,N_17559,N_18346);
nor U23729 (N_23729,N_18795,N_19467);
nor U23730 (N_23730,N_18692,N_16274);
and U23731 (N_23731,N_18147,N_15177);
nand U23732 (N_23732,N_15116,N_15587);
nand U23733 (N_23733,N_19164,N_17749);
nor U23734 (N_23734,N_15192,N_18107);
nand U23735 (N_23735,N_15680,N_17379);
or U23736 (N_23736,N_17289,N_19655);
nor U23737 (N_23737,N_18008,N_18106);
and U23738 (N_23738,N_18202,N_18790);
or U23739 (N_23739,N_16311,N_15338);
or U23740 (N_23740,N_17289,N_18338);
and U23741 (N_23741,N_15636,N_15131);
nand U23742 (N_23742,N_17902,N_17800);
and U23743 (N_23743,N_15060,N_18181);
and U23744 (N_23744,N_18544,N_17442);
nor U23745 (N_23745,N_16392,N_15293);
xnor U23746 (N_23746,N_15125,N_16027);
nor U23747 (N_23747,N_19480,N_15134);
nor U23748 (N_23748,N_17802,N_19198);
and U23749 (N_23749,N_19602,N_18058);
nor U23750 (N_23750,N_16817,N_15840);
or U23751 (N_23751,N_18440,N_16895);
nand U23752 (N_23752,N_19401,N_19816);
xnor U23753 (N_23753,N_15024,N_17887);
or U23754 (N_23754,N_19627,N_18344);
nand U23755 (N_23755,N_18804,N_16873);
nor U23756 (N_23756,N_17004,N_17278);
and U23757 (N_23757,N_18504,N_16678);
nand U23758 (N_23758,N_16014,N_15003);
or U23759 (N_23759,N_17266,N_16022);
or U23760 (N_23760,N_17574,N_18454);
nand U23761 (N_23761,N_16189,N_16134);
nand U23762 (N_23762,N_16407,N_19286);
or U23763 (N_23763,N_16520,N_17356);
nor U23764 (N_23764,N_19461,N_16237);
nor U23765 (N_23765,N_17301,N_19531);
nor U23766 (N_23766,N_17856,N_15606);
nand U23767 (N_23767,N_17445,N_16055);
and U23768 (N_23768,N_16115,N_17781);
nand U23769 (N_23769,N_16013,N_19671);
nor U23770 (N_23770,N_16019,N_18762);
nor U23771 (N_23771,N_17387,N_18768);
or U23772 (N_23772,N_18731,N_17442);
nand U23773 (N_23773,N_15996,N_15433);
nand U23774 (N_23774,N_19531,N_18880);
and U23775 (N_23775,N_19908,N_15875);
nor U23776 (N_23776,N_16953,N_15839);
nand U23777 (N_23777,N_17097,N_18474);
nand U23778 (N_23778,N_19801,N_18572);
or U23779 (N_23779,N_17374,N_15232);
nor U23780 (N_23780,N_19660,N_15803);
nand U23781 (N_23781,N_18185,N_16425);
and U23782 (N_23782,N_18807,N_19115);
nand U23783 (N_23783,N_17950,N_16827);
xnor U23784 (N_23784,N_19559,N_19301);
and U23785 (N_23785,N_18001,N_17755);
or U23786 (N_23786,N_18034,N_16986);
xnor U23787 (N_23787,N_17755,N_17281);
nand U23788 (N_23788,N_18905,N_15693);
or U23789 (N_23789,N_17695,N_17818);
and U23790 (N_23790,N_19986,N_18960);
or U23791 (N_23791,N_19272,N_18768);
nor U23792 (N_23792,N_16237,N_16475);
nand U23793 (N_23793,N_17134,N_17407);
or U23794 (N_23794,N_18073,N_18979);
and U23795 (N_23795,N_16695,N_19845);
xnor U23796 (N_23796,N_15724,N_15636);
and U23797 (N_23797,N_18693,N_18085);
nor U23798 (N_23798,N_16088,N_19590);
nand U23799 (N_23799,N_15324,N_19814);
nand U23800 (N_23800,N_17110,N_17717);
nor U23801 (N_23801,N_17747,N_15755);
nor U23802 (N_23802,N_19551,N_17556);
nor U23803 (N_23803,N_15258,N_16462);
and U23804 (N_23804,N_19668,N_18245);
and U23805 (N_23805,N_18916,N_19619);
and U23806 (N_23806,N_17205,N_16238);
and U23807 (N_23807,N_17483,N_16669);
nor U23808 (N_23808,N_16498,N_16349);
and U23809 (N_23809,N_16385,N_15809);
and U23810 (N_23810,N_15320,N_16392);
nand U23811 (N_23811,N_18535,N_16855);
and U23812 (N_23812,N_17499,N_16756);
nand U23813 (N_23813,N_18461,N_15174);
and U23814 (N_23814,N_16207,N_19666);
nor U23815 (N_23815,N_15134,N_19224);
xor U23816 (N_23816,N_15145,N_16692);
nand U23817 (N_23817,N_19384,N_16835);
nand U23818 (N_23818,N_16631,N_15361);
nand U23819 (N_23819,N_18761,N_15119);
nor U23820 (N_23820,N_18875,N_19436);
or U23821 (N_23821,N_16288,N_19149);
and U23822 (N_23822,N_18391,N_17046);
nor U23823 (N_23823,N_17023,N_17718);
and U23824 (N_23824,N_16407,N_16506);
and U23825 (N_23825,N_18977,N_18081);
and U23826 (N_23826,N_19732,N_18588);
xor U23827 (N_23827,N_15313,N_18285);
nand U23828 (N_23828,N_16259,N_17168);
nor U23829 (N_23829,N_16660,N_19737);
nor U23830 (N_23830,N_17979,N_15037);
or U23831 (N_23831,N_15621,N_16163);
or U23832 (N_23832,N_17023,N_15715);
and U23833 (N_23833,N_15894,N_19095);
or U23834 (N_23834,N_15489,N_18340);
nand U23835 (N_23835,N_16172,N_18669);
or U23836 (N_23836,N_18114,N_17619);
or U23837 (N_23837,N_16035,N_17742);
or U23838 (N_23838,N_18101,N_19668);
nor U23839 (N_23839,N_19484,N_15915);
or U23840 (N_23840,N_18435,N_19751);
nor U23841 (N_23841,N_19811,N_17510);
and U23842 (N_23842,N_15384,N_19517);
or U23843 (N_23843,N_17571,N_18075);
nor U23844 (N_23844,N_15246,N_17910);
xnor U23845 (N_23845,N_16660,N_18571);
or U23846 (N_23846,N_19606,N_19301);
nor U23847 (N_23847,N_19146,N_16845);
and U23848 (N_23848,N_16441,N_17114);
nand U23849 (N_23849,N_17217,N_17051);
or U23850 (N_23850,N_17227,N_19795);
and U23851 (N_23851,N_18091,N_19792);
nor U23852 (N_23852,N_19994,N_19849);
nand U23853 (N_23853,N_15208,N_19095);
nand U23854 (N_23854,N_15190,N_17169);
and U23855 (N_23855,N_17356,N_15039);
nor U23856 (N_23856,N_17034,N_15428);
and U23857 (N_23857,N_16015,N_17662);
xnor U23858 (N_23858,N_18103,N_15878);
or U23859 (N_23859,N_15815,N_18876);
or U23860 (N_23860,N_17470,N_15143);
or U23861 (N_23861,N_16592,N_16328);
or U23862 (N_23862,N_16290,N_17203);
nor U23863 (N_23863,N_18869,N_16279);
xor U23864 (N_23864,N_18494,N_18107);
and U23865 (N_23865,N_19146,N_15125);
or U23866 (N_23866,N_16248,N_15508);
nor U23867 (N_23867,N_15006,N_15687);
nand U23868 (N_23868,N_16594,N_18233);
xor U23869 (N_23869,N_17734,N_18156);
and U23870 (N_23870,N_16960,N_17069);
nor U23871 (N_23871,N_19646,N_17028);
nand U23872 (N_23872,N_15539,N_15504);
nand U23873 (N_23873,N_15273,N_17088);
or U23874 (N_23874,N_15540,N_18487);
nor U23875 (N_23875,N_15023,N_16164);
xor U23876 (N_23876,N_15803,N_19796);
and U23877 (N_23877,N_18985,N_18301);
and U23878 (N_23878,N_18314,N_18783);
and U23879 (N_23879,N_15375,N_15233);
and U23880 (N_23880,N_19199,N_16431);
or U23881 (N_23881,N_19093,N_19884);
xnor U23882 (N_23882,N_16047,N_18962);
or U23883 (N_23883,N_17841,N_16263);
nor U23884 (N_23884,N_15080,N_18752);
nand U23885 (N_23885,N_17234,N_19544);
nand U23886 (N_23886,N_17284,N_15320);
or U23887 (N_23887,N_17338,N_19402);
nand U23888 (N_23888,N_17078,N_18772);
nor U23889 (N_23889,N_19617,N_19749);
nor U23890 (N_23890,N_15104,N_19747);
nor U23891 (N_23891,N_15980,N_16481);
nor U23892 (N_23892,N_19525,N_15990);
nor U23893 (N_23893,N_17686,N_15037);
or U23894 (N_23894,N_16993,N_16786);
or U23895 (N_23895,N_19566,N_18769);
and U23896 (N_23896,N_15155,N_15257);
nor U23897 (N_23897,N_17470,N_19491);
and U23898 (N_23898,N_15019,N_17145);
nor U23899 (N_23899,N_18590,N_17848);
nor U23900 (N_23900,N_18858,N_19139);
and U23901 (N_23901,N_18034,N_16554);
and U23902 (N_23902,N_18104,N_19173);
nand U23903 (N_23903,N_18741,N_16115);
nor U23904 (N_23904,N_18368,N_19940);
xnor U23905 (N_23905,N_15068,N_16771);
nand U23906 (N_23906,N_17745,N_18738);
and U23907 (N_23907,N_15949,N_19346);
or U23908 (N_23908,N_15005,N_18951);
or U23909 (N_23909,N_16576,N_17181);
nand U23910 (N_23910,N_18116,N_17391);
and U23911 (N_23911,N_19331,N_16744);
nor U23912 (N_23912,N_15311,N_18406);
xnor U23913 (N_23913,N_17186,N_17342);
xnor U23914 (N_23914,N_18093,N_17921);
or U23915 (N_23915,N_19339,N_18621);
nor U23916 (N_23916,N_17491,N_18536);
or U23917 (N_23917,N_17246,N_16526);
or U23918 (N_23918,N_15591,N_16482);
nor U23919 (N_23919,N_19202,N_19302);
nand U23920 (N_23920,N_19399,N_16054);
xor U23921 (N_23921,N_15607,N_16306);
and U23922 (N_23922,N_19732,N_19443);
or U23923 (N_23923,N_18707,N_15725);
nand U23924 (N_23924,N_15266,N_19943);
nor U23925 (N_23925,N_18771,N_16998);
xnor U23926 (N_23926,N_19488,N_16263);
nor U23927 (N_23927,N_19117,N_19196);
and U23928 (N_23928,N_19033,N_18692);
nor U23929 (N_23929,N_15019,N_18315);
nand U23930 (N_23930,N_19451,N_17271);
and U23931 (N_23931,N_16067,N_16509);
nor U23932 (N_23932,N_15277,N_15110);
or U23933 (N_23933,N_19416,N_15344);
xnor U23934 (N_23934,N_16495,N_19544);
nor U23935 (N_23935,N_15031,N_16426);
nor U23936 (N_23936,N_18136,N_16284);
and U23937 (N_23937,N_17989,N_15998);
xnor U23938 (N_23938,N_18700,N_19525);
and U23939 (N_23939,N_16246,N_19450);
or U23940 (N_23940,N_19483,N_19728);
and U23941 (N_23941,N_18094,N_18004);
nand U23942 (N_23942,N_16528,N_16595);
nand U23943 (N_23943,N_17787,N_15108);
and U23944 (N_23944,N_17144,N_19337);
nor U23945 (N_23945,N_18914,N_17126);
xnor U23946 (N_23946,N_17255,N_17662);
or U23947 (N_23947,N_16201,N_15160);
and U23948 (N_23948,N_17884,N_15965);
nand U23949 (N_23949,N_17706,N_15079);
and U23950 (N_23950,N_17016,N_15257);
xnor U23951 (N_23951,N_16935,N_18894);
nor U23952 (N_23952,N_18549,N_15574);
nor U23953 (N_23953,N_15967,N_16993);
or U23954 (N_23954,N_18427,N_15424);
or U23955 (N_23955,N_19117,N_16679);
nand U23956 (N_23956,N_17845,N_18845);
nor U23957 (N_23957,N_17225,N_16986);
xnor U23958 (N_23958,N_18556,N_17586);
nand U23959 (N_23959,N_19179,N_15101);
nand U23960 (N_23960,N_15129,N_17812);
or U23961 (N_23961,N_19045,N_18526);
nor U23962 (N_23962,N_19918,N_18968);
or U23963 (N_23963,N_18672,N_15635);
and U23964 (N_23964,N_17708,N_18461);
nand U23965 (N_23965,N_19449,N_18929);
and U23966 (N_23966,N_16897,N_18159);
nor U23967 (N_23967,N_15938,N_15991);
or U23968 (N_23968,N_19935,N_16531);
and U23969 (N_23969,N_17229,N_18831);
xor U23970 (N_23970,N_17691,N_17198);
or U23971 (N_23971,N_17118,N_19111);
nor U23972 (N_23972,N_18878,N_15019);
and U23973 (N_23973,N_19984,N_17713);
nand U23974 (N_23974,N_16784,N_15932);
nand U23975 (N_23975,N_17744,N_18734);
nor U23976 (N_23976,N_16200,N_17940);
nand U23977 (N_23977,N_16170,N_16245);
and U23978 (N_23978,N_15996,N_18463);
nand U23979 (N_23979,N_15179,N_19512);
and U23980 (N_23980,N_16053,N_19723);
or U23981 (N_23981,N_15765,N_19427);
or U23982 (N_23982,N_17801,N_17359);
xnor U23983 (N_23983,N_15089,N_18012);
xnor U23984 (N_23984,N_16968,N_15095);
or U23985 (N_23985,N_18863,N_15904);
nand U23986 (N_23986,N_18780,N_18128);
nand U23987 (N_23987,N_17089,N_15043);
or U23988 (N_23988,N_15744,N_15995);
or U23989 (N_23989,N_15937,N_15544);
and U23990 (N_23990,N_18333,N_18494);
nand U23991 (N_23991,N_17062,N_15933);
and U23992 (N_23992,N_16507,N_16440);
nor U23993 (N_23993,N_18171,N_19989);
nand U23994 (N_23994,N_17232,N_15400);
xnor U23995 (N_23995,N_17297,N_17207);
nand U23996 (N_23996,N_17365,N_18438);
and U23997 (N_23997,N_18433,N_19323);
nand U23998 (N_23998,N_16933,N_16231);
xnor U23999 (N_23999,N_18871,N_16466);
or U24000 (N_24000,N_16850,N_16558);
and U24001 (N_24001,N_16175,N_18402);
nand U24002 (N_24002,N_17562,N_16265);
and U24003 (N_24003,N_19930,N_17405);
or U24004 (N_24004,N_16251,N_17801);
or U24005 (N_24005,N_19044,N_18302);
or U24006 (N_24006,N_15089,N_19500);
nor U24007 (N_24007,N_18975,N_15422);
nand U24008 (N_24008,N_17885,N_19778);
and U24009 (N_24009,N_19049,N_18132);
or U24010 (N_24010,N_15388,N_19950);
xnor U24011 (N_24011,N_17684,N_17626);
xor U24012 (N_24012,N_19271,N_16394);
or U24013 (N_24013,N_18956,N_18723);
and U24014 (N_24014,N_16490,N_18438);
or U24015 (N_24015,N_18755,N_15538);
or U24016 (N_24016,N_16126,N_18552);
and U24017 (N_24017,N_16373,N_15389);
nor U24018 (N_24018,N_17792,N_18926);
and U24019 (N_24019,N_19727,N_19171);
nand U24020 (N_24020,N_19878,N_16348);
nor U24021 (N_24021,N_15116,N_15469);
or U24022 (N_24022,N_18807,N_16923);
and U24023 (N_24023,N_17415,N_15925);
nor U24024 (N_24024,N_16878,N_18530);
nor U24025 (N_24025,N_16903,N_17699);
and U24026 (N_24026,N_16507,N_18156);
or U24027 (N_24027,N_15646,N_19627);
and U24028 (N_24028,N_18328,N_19455);
nor U24029 (N_24029,N_17327,N_18662);
nor U24030 (N_24030,N_16330,N_17774);
and U24031 (N_24031,N_17145,N_18586);
nand U24032 (N_24032,N_16488,N_17750);
nand U24033 (N_24033,N_18161,N_15595);
nand U24034 (N_24034,N_16954,N_15967);
nand U24035 (N_24035,N_19411,N_16855);
nor U24036 (N_24036,N_19666,N_16096);
nor U24037 (N_24037,N_17482,N_17154);
nor U24038 (N_24038,N_15622,N_16452);
or U24039 (N_24039,N_15399,N_17821);
or U24040 (N_24040,N_18595,N_15172);
nor U24041 (N_24041,N_18087,N_15178);
nand U24042 (N_24042,N_15973,N_17380);
or U24043 (N_24043,N_19554,N_19424);
and U24044 (N_24044,N_18786,N_17393);
and U24045 (N_24045,N_16989,N_19019);
or U24046 (N_24046,N_16714,N_18813);
nand U24047 (N_24047,N_15766,N_17793);
nor U24048 (N_24048,N_16550,N_17445);
nand U24049 (N_24049,N_16285,N_15757);
and U24050 (N_24050,N_19744,N_15633);
or U24051 (N_24051,N_18812,N_17545);
and U24052 (N_24052,N_18281,N_18352);
nor U24053 (N_24053,N_16137,N_17677);
and U24054 (N_24054,N_18258,N_19432);
and U24055 (N_24055,N_16074,N_16800);
or U24056 (N_24056,N_17209,N_16994);
nor U24057 (N_24057,N_17329,N_18748);
nand U24058 (N_24058,N_17073,N_19843);
nand U24059 (N_24059,N_19933,N_16068);
or U24060 (N_24060,N_17929,N_15655);
and U24061 (N_24061,N_16833,N_15858);
nor U24062 (N_24062,N_17845,N_15702);
nor U24063 (N_24063,N_16006,N_17793);
xor U24064 (N_24064,N_18518,N_17095);
and U24065 (N_24065,N_18080,N_16006);
and U24066 (N_24066,N_15100,N_16163);
nand U24067 (N_24067,N_15132,N_15229);
or U24068 (N_24068,N_15750,N_17935);
xor U24069 (N_24069,N_18834,N_15791);
or U24070 (N_24070,N_15349,N_16304);
and U24071 (N_24071,N_19207,N_19060);
and U24072 (N_24072,N_17023,N_16553);
or U24073 (N_24073,N_19569,N_15014);
nand U24074 (N_24074,N_18855,N_16994);
nand U24075 (N_24075,N_15593,N_18536);
xnor U24076 (N_24076,N_19389,N_19289);
and U24077 (N_24077,N_19874,N_16163);
or U24078 (N_24078,N_17204,N_16984);
nor U24079 (N_24079,N_16037,N_17281);
and U24080 (N_24080,N_15450,N_15019);
nor U24081 (N_24081,N_16307,N_17688);
or U24082 (N_24082,N_16153,N_17463);
or U24083 (N_24083,N_18764,N_15783);
or U24084 (N_24084,N_15190,N_16483);
nand U24085 (N_24085,N_16400,N_18223);
nor U24086 (N_24086,N_18010,N_18881);
and U24087 (N_24087,N_17423,N_19039);
xnor U24088 (N_24088,N_19696,N_16299);
nand U24089 (N_24089,N_17236,N_19061);
nand U24090 (N_24090,N_16041,N_16872);
nand U24091 (N_24091,N_17462,N_17456);
or U24092 (N_24092,N_15224,N_18270);
nor U24093 (N_24093,N_19062,N_15690);
xnor U24094 (N_24094,N_17637,N_16780);
and U24095 (N_24095,N_19032,N_18031);
nand U24096 (N_24096,N_18149,N_17663);
xor U24097 (N_24097,N_18981,N_16825);
and U24098 (N_24098,N_15200,N_15340);
or U24099 (N_24099,N_19932,N_18919);
and U24100 (N_24100,N_15001,N_18071);
or U24101 (N_24101,N_16558,N_19336);
and U24102 (N_24102,N_16828,N_16766);
nand U24103 (N_24103,N_15729,N_15208);
and U24104 (N_24104,N_19824,N_15133);
nand U24105 (N_24105,N_16798,N_17692);
xnor U24106 (N_24106,N_19621,N_16663);
and U24107 (N_24107,N_19551,N_16451);
nor U24108 (N_24108,N_18173,N_17655);
xnor U24109 (N_24109,N_16854,N_19270);
nand U24110 (N_24110,N_15646,N_16753);
nor U24111 (N_24111,N_18818,N_17517);
nand U24112 (N_24112,N_17795,N_15901);
nor U24113 (N_24113,N_18004,N_19529);
and U24114 (N_24114,N_16257,N_16655);
or U24115 (N_24115,N_18122,N_19793);
nand U24116 (N_24116,N_16470,N_17627);
nand U24117 (N_24117,N_16006,N_15752);
and U24118 (N_24118,N_15362,N_18738);
nor U24119 (N_24119,N_15029,N_17960);
or U24120 (N_24120,N_18720,N_16543);
xnor U24121 (N_24121,N_17536,N_19321);
or U24122 (N_24122,N_17069,N_15529);
xnor U24123 (N_24123,N_15017,N_19004);
nor U24124 (N_24124,N_19422,N_18294);
or U24125 (N_24125,N_18344,N_17180);
or U24126 (N_24126,N_16986,N_18793);
nor U24127 (N_24127,N_15508,N_19392);
nand U24128 (N_24128,N_17444,N_17237);
nand U24129 (N_24129,N_19390,N_18950);
nand U24130 (N_24130,N_16867,N_16391);
nand U24131 (N_24131,N_19684,N_17040);
nor U24132 (N_24132,N_18657,N_18288);
or U24133 (N_24133,N_17505,N_17871);
or U24134 (N_24134,N_18925,N_17094);
or U24135 (N_24135,N_17446,N_19928);
nand U24136 (N_24136,N_16226,N_15576);
or U24137 (N_24137,N_15242,N_19132);
and U24138 (N_24138,N_17975,N_18241);
nor U24139 (N_24139,N_17292,N_16000);
nand U24140 (N_24140,N_18485,N_15593);
xor U24141 (N_24141,N_15549,N_15081);
nand U24142 (N_24142,N_19396,N_18174);
and U24143 (N_24143,N_18821,N_17995);
or U24144 (N_24144,N_18635,N_17336);
and U24145 (N_24145,N_15767,N_19429);
nand U24146 (N_24146,N_15554,N_19588);
and U24147 (N_24147,N_17168,N_15352);
nand U24148 (N_24148,N_15628,N_19820);
or U24149 (N_24149,N_15542,N_15862);
or U24150 (N_24150,N_15574,N_19435);
nor U24151 (N_24151,N_19559,N_17967);
nor U24152 (N_24152,N_19553,N_15084);
and U24153 (N_24153,N_19406,N_16040);
nor U24154 (N_24154,N_15552,N_16196);
nand U24155 (N_24155,N_17133,N_18371);
xor U24156 (N_24156,N_15138,N_17680);
and U24157 (N_24157,N_18435,N_16695);
nor U24158 (N_24158,N_17176,N_16817);
nand U24159 (N_24159,N_18951,N_15841);
nand U24160 (N_24160,N_19906,N_16279);
nor U24161 (N_24161,N_18708,N_17851);
or U24162 (N_24162,N_19041,N_19919);
or U24163 (N_24163,N_17134,N_17156);
nand U24164 (N_24164,N_15493,N_16667);
nor U24165 (N_24165,N_17941,N_19046);
nor U24166 (N_24166,N_18469,N_17643);
nor U24167 (N_24167,N_19259,N_16205);
or U24168 (N_24168,N_15858,N_19398);
xnor U24169 (N_24169,N_19454,N_18744);
nand U24170 (N_24170,N_15567,N_18815);
or U24171 (N_24171,N_16015,N_18792);
or U24172 (N_24172,N_18309,N_17987);
and U24173 (N_24173,N_16828,N_17406);
nor U24174 (N_24174,N_19215,N_15810);
and U24175 (N_24175,N_18070,N_15329);
or U24176 (N_24176,N_15421,N_16062);
or U24177 (N_24177,N_17953,N_17107);
xnor U24178 (N_24178,N_16126,N_18245);
or U24179 (N_24179,N_15166,N_16532);
and U24180 (N_24180,N_19737,N_17654);
nor U24181 (N_24181,N_16345,N_17713);
xor U24182 (N_24182,N_15505,N_17234);
and U24183 (N_24183,N_18742,N_19704);
nor U24184 (N_24184,N_17514,N_17430);
and U24185 (N_24185,N_17812,N_17476);
nand U24186 (N_24186,N_16343,N_15100);
and U24187 (N_24187,N_18333,N_16460);
and U24188 (N_24188,N_16913,N_17900);
or U24189 (N_24189,N_17029,N_19275);
or U24190 (N_24190,N_18119,N_15456);
nor U24191 (N_24191,N_18933,N_17749);
and U24192 (N_24192,N_15192,N_17288);
nor U24193 (N_24193,N_15344,N_17528);
and U24194 (N_24194,N_18338,N_19327);
and U24195 (N_24195,N_19621,N_18539);
nand U24196 (N_24196,N_17220,N_17052);
and U24197 (N_24197,N_19827,N_17686);
nand U24198 (N_24198,N_17493,N_18167);
and U24199 (N_24199,N_16248,N_17360);
nand U24200 (N_24200,N_15004,N_18770);
xor U24201 (N_24201,N_19734,N_16434);
and U24202 (N_24202,N_17109,N_19672);
nand U24203 (N_24203,N_15782,N_15800);
nand U24204 (N_24204,N_16628,N_18120);
and U24205 (N_24205,N_17905,N_18628);
nor U24206 (N_24206,N_15367,N_16618);
nor U24207 (N_24207,N_17757,N_16292);
and U24208 (N_24208,N_16379,N_15284);
and U24209 (N_24209,N_18985,N_15531);
nor U24210 (N_24210,N_18937,N_16017);
or U24211 (N_24211,N_16003,N_16191);
or U24212 (N_24212,N_15785,N_15848);
nand U24213 (N_24213,N_16333,N_17238);
nand U24214 (N_24214,N_16786,N_15548);
nor U24215 (N_24215,N_16540,N_17554);
xnor U24216 (N_24216,N_16886,N_19725);
and U24217 (N_24217,N_18232,N_17295);
or U24218 (N_24218,N_16697,N_16541);
nand U24219 (N_24219,N_16006,N_17957);
or U24220 (N_24220,N_19972,N_16804);
xnor U24221 (N_24221,N_18032,N_19524);
and U24222 (N_24222,N_18631,N_17268);
nand U24223 (N_24223,N_17740,N_18801);
and U24224 (N_24224,N_18354,N_19767);
xor U24225 (N_24225,N_18309,N_19470);
nor U24226 (N_24226,N_15508,N_18184);
nor U24227 (N_24227,N_18280,N_19173);
and U24228 (N_24228,N_16369,N_17011);
nor U24229 (N_24229,N_15537,N_15360);
nor U24230 (N_24230,N_16442,N_18876);
nand U24231 (N_24231,N_16689,N_18200);
and U24232 (N_24232,N_19044,N_15224);
xnor U24233 (N_24233,N_19310,N_17724);
and U24234 (N_24234,N_18506,N_15644);
nor U24235 (N_24235,N_17644,N_18334);
and U24236 (N_24236,N_15352,N_17069);
nor U24237 (N_24237,N_19247,N_18062);
nand U24238 (N_24238,N_15827,N_16870);
nor U24239 (N_24239,N_16031,N_17449);
and U24240 (N_24240,N_18707,N_15493);
nor U24241 (N_24241,N_18800,N_18107);
and U24242 (N_24242,N_19635,N_19115);
or U24243 (N_24243,N_18338,N_17097);
or U24244 (N_24244,N_16141,N_17010);
or U24245 (N_24245,N_16220,N_15195);
nor U24246 (N_24246,N_19135,N_18823);
nand U24247 (N_24247,N_15998,N_19027);
xnor U24248 (N_24248,N_15233,N_19060);
nand U24249 (N_24249,N_15877,N_17300);
xor U24250 (N_24250,N_18186,N_16946);
nor U24251 (N_24251,N_17739,N_17757);
nand U24252 (N_24252,N_18760,N_15773);
nand U24253 (N_24253,N_18180,N_16531);
nor U24254 (N_24254,N_16610,N_17083);
xor U24255 (N_24255,N_19175,N_18138);
and U24256 (N_24256,N_17520,N_19133);
nor U24257 (N_24257,N_16787,N_18787);
and U24258 (N_24258,N_16962,N_18334);
or U24259 (N_24259,N_16016,N_17993);
nor U24260 (N_24260,N_15531,N_15864);
nor U24261 (N_24261,N_15865,N_17076);
nor U24262 (N_24262,N_15669,N_16432);
or U24263 (N_24263,N_17201,N_16995);
nor U24264 (N_24264,N_17831,N_16371);
or U24265 (N_24265,N_19006,N_17905);
xnor U24266 (N_24266,N_15331,N_17225);
nor U24267 (N_24267,N_19948,N_16801);
or U24268 (N_24268,N_19669,N_16132);
or U24269 (N_24269,N_19632,N_18339);
and U24270 (N_24270,N_15707,N_19844);
nand U24271 (N_24271,N_19524,N_16345);
or U24272 (N_24272,N_18046,N_15994);
and U24273 (N_24273,N_16044,N_19115);
nor U24274 (N_24274,N_16874,N_16160);
or U24275 (N_24275,N_18163,N_18897);
nor U24276 (N_24276,N_15366,N_16082);
or U24277 (N_24277,N_16777,N_18312);
or U24278 (N_24278,N_15642,N_17176);
nor U24279 (N_24279,N_17610,N_17156);
nand U24280 (N_24280,N_15653,N_16719);
xnor U24281 (N_24281,N_19950,N_18086);
or U24282 (N_24282,N_15989,N_16932);
or U24283 (N_24283,N_17251,N_16743);
xnor U24284 (N_24284,N_16373,N_16020);
and U24285 (N_24285,N_15437,N_19888);
nand U24286 (N_24286,N_19671,N_19041);
and U24287 (N_24287,N_18611,N_19632);
and U24288 (N_24288,N_15478,N_18626);
nor U24289 (N_24289,N_17079,N_18719);
or U24290 (N_24290,N_15241,N_16707);
and U24291 (N_24291,N_17729,N_16744);
nor U24292 (N_24292,N_15202,N_16948);
nor U24293 (N_24293,N_17168,N_19924);
nor U24294 (N_24294,N_16390,N_18073);
xor U24295 (N_24295,N_17725,N_18705);
or U24296 (N_24296,N_17121,N_16549);
nand U24297 (N_24297,N_17961,N_18230);
or U24298 (N_24298,N_18498,N_17311);
nor U24299 (N_24299,N_17769,N_17958);
nand U24300 (N_24300,N_19784,N_18463);
xor U24301 (N_24301,N_17819,N_19056);
nor U24302 (N_24302,N_19942,N_19127);
nand U24303 (N_24303,N_18247,N_19397);
or U24304 (N_24304,N_17811,N_15388);
nand U24305 (N_24305,N_19943,N_16197);
xor U24306 (N_24306,N_16053,N_17209);
nor U24307 (N_24307,N_15919,N_18652);
or U24308 (N_24308,N_16583,N_18021);
or U24309 (N_24309,N_16450,N_19703);
nor U24310 (N_24310,N_16371,N_15676);
nor U24311 (N_24311,N_18377,N_19447);
nand U24312 (N_24312,N_15725,N_18019);
nor U24313 (N_24313,N_16288,N_16952);
nor U24314 (N_24314,N_19177,N_19184);
and U24315 (N_24315,N_19679,N_16264);
nor U24316 (N_24316,N_19003,N_17655);
and U24317 (N_24317,N_19590,N_19050);
nor U24318 (N_24318,N_17561,N_19413);
and U24319 (N_24319,N_17073,N_17130);
or U24320 (N_24320,N_18395,N_16845);
and U24321 (N_24321,N_15737,N_18150);
and U24322 (N_24322,N_17649,N_19885);
nand U24323 (N_24323,N_15582,N_18580);
xor U24324 (N_24324,N_16758,N_15066);
and U24325 (N_24325,N_15201,N_17789);
nor U24326 (N_24326,N_17552,N_15499);
nor U24327 (N_24327,N_19972,N_18231);
and U24328 (N_24328,N_16467,N_15046);
and U24329 (N_24329,N_17868,N_17540);
nand U24330 (N_24330,N_15028,N_16495);
nor U24331 (N_24331,N_18191,N_18480);
xor U24332 (N_24332,N_17352,N_18885);
nor U24333 (N_24333,N_17035,N_17414);
and U24334 (N_24334,N_15523,N_15127);
nand U24335 (N_24335,N_16254,N_18859);
nand U24336 (N_24336,N_16460,N_17866);
or U24337 (N_24337,N_15733,N_16965);
and U24338 (N_24338,N_19138,N_19562);
nor U24339 (N_24339,N_15734,N_18853);
and U24340 (N_24340,N_15765,N_15642);
nor U24341 (N_24341,N_15021,N_16271);
nor U24342 (N_24342,N_16275,N_18154);
nand U24343 (N_24343,N_16163,N_19428);
or U24344 (N_24344,N_16830,N_16646);
nor U24345 (N_24345,N_16103,N_17828);
and U24346 (N_24346,N_18951,N_19623);
nand U24347 (N_24347,N_17490,N_19990);
nand U24348 (N_24348,N_19073,N_18284);
xnor U24349 (N_24349,N_19331,N_15783);
and U24350 (N_24350,N_17972,N_15219);
xnor U24351 (N_24351,N_19675,N_18272);
nand U24352 (N_24352,N_19363,N_18366);
nor U24353 (N_24353,N_18699,N_17486);
or U24354 (N_24354,N_18991,N_16513);
or U24355 (N_24355,N_19085,N_18998);
nand U24356 (N_24356,N_19175,N_19809);
or U24357 (N_24357,N_16675,N_19261);
nand U24358 (N_24358,N_19996,N_18052);
nor U24359 (N_24359,N_19151,N_19371);
nor U24360 (N_24360,N_15163,N_19847);
and U24361 (N_24361,N_16749,N_19045);
nor U24362 (N_24362,N_16936,N_15980);
nor U24363 (N_24363,N_17040,N_19185);
nor U24364 (N_24364,N_17422,N_17984);
and U24365 (N_24365,N_17466,N_19365);
or U24366 (N_24366,N_17593,N_15004);
nand U24367 (N_24367,N_16711,N_16476);
and U24368 (N_24368,N_19761,N_19337);
nor U24369 (N_24369,N_15429,N_18581);
nor U24370 (N_24370,N_16158,N_19742);
and U24371 (N_24371,N_17618,N_18298);
nor U24372 (N_24372,N_18500,N_18972);
nor U24373 (N_24373,N_15487,N_15313);
or U24374 (N_24374,N_18419,N_17520);
or U24375 (N_24375,N_19922,N_18394);
or U24376 (N_24376,N_17589,N_19553);
and U24377 (N_24377,N_16347,N_18756);
and U24378 (N_24378,N_17086,N_19213);
or U24379 (N_24379,N_19029,N_18631);
and U24380 (N_24380,N_16206,N_18225);
nand U24381 (N_24381,N_19857,N_19865);
nor U24382 (N_24382,N_15024,N_19106);
xor U24383 (N_24383,N_18452,N_18717);
or U24384 (N_24384,N_19975,N_18829);
xnor U24385 (N_24385,N_17603,N_16386);
and U24386 (N_24386,N_16856,N_15641);
nor U24387 (N_24387,N_18412,N_15850);
or U24388 (N_24388,N_17860,N_18479);
or U24389 (N_24389,N_16760,N_18001);
and U24390 (N_24390,N_16935,N_17017);
and U24391 (N_24391,N_18359,N_17879);
nand U24392 (N_24392,N_16671,N_15947);
and U24393 (N_24393,N_19602,N_18250);
and U24394 (N_24394,N_16144,N_15638);
and U24395 (N_24395,N_18908,N_19665);
nand U24396 (N_24396,N_19369,N_18019);
and U24397 (N_24397,N_16894,N_17781);
nand U24398 (N_24398,N_19146,N_17311);
or U24399 (N_24399,N_16137,N_17627);
and U24400 (N_24400,N_17963,N_18360);
nand U24401 (N_24401,N_18688,N_16073);
nor U24402 (N_24402,N_19467,N_15629);
or U24403 (N_24403,N_16689,N_15773);
and U24404 (N_24404,N_19781,N_16845);
and U24405 (N_24405,N_18970,N_15820);
and U24406 (N_24406,N_16147,N_19548);
nor U24407 (N_24407,N_16982,N_16769);
or U24408 (N_24408,N_15524,N_18512);
or U24409 (N_24409,N_15774,N_16683);
nand U24410 (N_24410,N_18560,N_19544);
nand U24411 (N_24411,N_16289,N_17068);
nor U24412 (N_24412,N_17696,N_19837);
or U24413 (N_24413,N_16186,N_16571);
or U24414 (N_24414,N_18488,N_19345);
nand U24415 (N_24415,N_15379,N_18028);
and U24416 (N_24416,N_18790,N_19376);
nor U24417 (N_24417,N_16773,N_19771);
nor U24418 (N_24418,N_17303,N_16521);
nor U24419 (N_24419,N_16800,N_19805);
or U24420 (N_24420,N_17916,N_17140);
and U24421 (N_24421,N_19073,N_16070);
and U24422 (N_24422,N_16190,N_17850);
nor U24423 (N_24423,N_16994,N_17425);
xor U24424 (N_24424,N_17279,N_18752);
and U24425 (N_24425,N_16362,N_16599);
nand U24426 (N_24426,N_17065,N_16456);
nand U24427 (N_24427,N_16139,N_16974);
or U24428 (N_24428,N_19816,N_18278);
nand U24429 (N_24429,N_18892,N_15243);
or U24430 (N_24430,N_16115,N_16581);
nand U24431 (N_24431,N_17562,N_18277);
nand U24432 (N_24432,N_16605,N_19219);
nand U24433 (N_24433,N_15922,N_17252);
nand U24434 (N_24434,N_19587,N_18430);
nand U24435 (N_24435,N_15324,N_17828);
and U24436 (N_24436,N_15056,N_17141);
and U24437 (N_24437,N_19156,N_16995);
or U24438 (N_24438,N_17038,N_16151);
or U24439 (N_24439,N_19014,N_16236);
nand U24440 (N_24440,N_17795,N_18187);
nor U24441 (N_24441,N_19147,N_15035);
nor U24442 (N_24442,N_19283,N_18658);
or U24443 (N_24443,N_15829,N_16861);
xnor U24444 (N_24444,N_18998,N_19160);
or U24445 (N_24445,N_17706,N_17332);
and U24446 (N_24446,N_19757,N_19150);
nand U24447 (N_24447,N_16922,N_16782);
nor U24448 (N_24448,N_18894,N_16546);
or U24449 (N_24449,N_18214,N_16954);
nand U24450 (N_24450,N_19803,N_15644);
or U24451 (N_24451,N_18464,N_17349);
nand U24452 (N_24452,N_16250,N_17720);
and U24453 (N_24453,N_18188,N_16032);
and U24454 (N_24454,N_18827,N_15950);
and U24455 (N_24455,N_18205,N_16740);
and U24456 (N_24456,N_17694,N_17650);
nand U24457 (N_24457,N_19661,N_19681);
xnor U24458 (N_24458,N_16699,N_19192);
xnor U24459 (N_24459,N_17186,N_16604);
nor U24460 (N_24460,N_19779,N_18376);
or U24461 (N_24461,N_19879,N_17716);
nand U24462 (N_24462,N_19001,N_18572);
xor U24463 (N_24463,N_16728,N_15611);
and U24464 (N_24464,N_18796,N_16126);
nand U24465 (N_24465,N_18067,N_19254);
nor U24466 (N_24466,N_15774,N_17542);
nor U24467 (N_24467,N_16951,N_16441);
or U24468 (N_24468,N_19148,N_16289);
and U24469 (N_24469,N_16149,N_17321);
and U24470 (N_24470,N_17360,N_17224);
or U24471 (N_24471,N_17943,N_18876);
and U24472 (N_24472,N_17894,N_16091);
xor U24473 (N_24473,N_17245,N_15446);
nor U24474 (N_24474,N_15026,N_18067);
nand U24475 (N_24475,N_17615,N_15418);
nor U24476 (N_24476,N_17429,N_18659);
and U24477 (N_24477,N_17575,N_18021);
or U24478 (N_24478,N_16450,N_16048);
nor U24479 (N_24479,N_18407,N_18653);
nor U24480 (N_24480,N_15963,N_18986);
nor U24481 (N_24481,N_16206,N_18899);
xnor U24482 (N_24482,N_18153,N_16975);
and U24483 (N_24483,N_16545,N_18557);
and U24484 (N_24484,N_16971,N_19630);
or U24485 (N_24485,N_19444,N_18689);
or U24486 (N_24486,N_16268,N_17176);
or U24487 (N_24487,N_16169,N_19819);
nand U24488 (N_24488,N_15984,N_19202);
xnor U24489 (N_24489,N_19119,N_16789);
nor U24490 (N_24490,N_18229,N_16797);
or U24491 (N_24491,N_18776,N_15792);
nand U24492 (N_24492,N_17980,N_18115);
and U24493 (N_24493,N_16113,N_18466);
nand U24494 (N_24494,N_15178,N_16961);
nand U24495 (N_24495,N_19443,N_16424);
or U24496 (N_24496,N_18530,N_15424);
xnor U24497 (N_24497,N_16524,N_16258);
nand U24498 (N_24498,N_16414,N_18338);
nor U24499 (N_24499,N_19846,N_18866);
xor U24500 (N_24500,N_18310,N_17729);
or U24501 (N_24501,N_19942,N_15733);
nand U24502 (N_24502,N_15471,N_17015);
or U24503 (N_24503,N_15658,N_19927);
nor U24504 (N_24504,N_18540,N_18502);
nand U24505 (N_24505,N_17089,N_19799);
and U24506 (N_24506,N_15423,N_16627);
and U24507 (N_24507,N_18260,N_17183);
and U24508 (N_24508,N_18344,N_16550);
nor U24509 (N_24509,N_16369,N_16440);
or U24510 (N_24510,N_15477,N_16672);
and U24511 (N_24511,N_17582,N_18959);
and U24512 (N_24512,N_16835,N_18686);
and U24513 (N_24513,N_16726,N_18553);
and U24514 (N_24514,N_15068,N_18758);
nand U24515 (N_24515,N_18010,N_15488);
nand U24516 (N_24516,N_18204,N_15657);
xor U24517 (N_24517,N_16696,N_17744);
nor U24518 (N_24518,N_16829,N_19059);
nand U24519 (N_24519,N_16030,N_17335);
nor U24520 (N_24520,N_16296,N_16434);
nor U24521 (N_24521,N_19608,N_18282);
nor U24522 (N_24522,N_18521,N_19270);
nand U24523 (N_24523,N_18859,N_16241);
nand U24524 (N_24524,N_18686,N_18421);
and U24525 (N_24525,N_15978,N_18658);
or U24526 (N_24526,N_16352,N_16817);
nand U24527 (N_24527,N_15210,N_15370);
nor U24528 (N_24528,N_18174,N_17511);
nor U24529 (N_24529,N_16717,N_19051);
nor U24530 (N_24530,N_17929,N_15483);
xor U24531 (N_24531,N_17063,N_18229);
nand U24532 (N_24532,N_16288,N_15265);
nor U24533 (N_24533,N_16297,N_19410);
nand U24534 (N_24534,N_17162,N_15193);
xnor U24535 (N_24535,N_16983,N_15023);
nand U24536 (N_24536,N_18637,N_16739);
nor U24537 (N_24537,N_16120,N_17466);
nor U24538 (N_24538,N_17423,N_17106);
nand U24539 (N_24539,N_19206,N_17758);
or U24540 (N_24540,N_19511,N_18478);
nand U24541 (N_24541,N_19358,N_19060);
nand U24542 (N_24542,N_19045,N_18363);
xor U24543 (N_24543,N_19973,N_17197);
or U24544 (N_24544,N_17354,N_18966);
or U24545 (N_24545,N_19399,N_16254);
nand U24546 (N_24546,N_16358,N_17286);
nor U24547 (N_24547,N_19319,N_19833);
xor U24548 (N_24548,N_19539,N_19765);
and U24549 (N_24549,N_15611,N_19803);
and U24550 (N_24550,N_16281,N_19811);
nand U24551 (N_24551,N_15499,N_19341);
nor U24552 (N_24552,N_16169,N_19247);
xor U24553 (N_24553,N_17690,N_16902);
nor U24554 (N_24554,N_19970,N_17395);
or U24555 (N_24555,N_15367,N_17814);
and U24556 (N_24556,N_18467,N_15504);
nand U24557 (N_24557,N_16825,N_18630);
nor U24558 (N_24558,N_15218,N_18234);
nor U24559 (N_24559,N_19430,N_19540);
or U24560 (N_24560,N_16226,N_17473);
or U24561 (N_24561,N_16035,N_18120);
or U24562 (N_24562,N_16615,N_18657);
and U24563 (N_24563,N_19854,N_16423);
and U24564 (N_24564,N_17013,N_17789);
nand U24565 (N_24565,N_18310,N_18649);
nor U24566 (N_24566,N_18816,N_16684);
nor U24567 (N_24567,N_17501,N_17178);
nand U24568 (N_24568,N_18828,N_16201);
or U24569 (N_24569,N_17143,N_15847);
nor U24570 (N_24570,N_19382,N_18820);
nor U24571 (N_24571,N_18043,N_18944);
xnor U24572 (N_24572,N_19336,N_18304);
nor U24573 (N_24573,N_17315,N_18788);
nor U24574 (N_24574,N_19902,N_17857);
nand U24575 (N_24575,N_16154,N_16808);
nand U24576 (N_24576,N_17083,N_19028);
nand U24577 (N_24577,N_18258,N_18639);
and U24578 (N_24578,N_15155,N_16620);
nor U24579 (N_24579,N_19725,N_17718);
nor U24580 (N_24580,N_16182,N_15943);
or U24581 (N_24581,N_18315,N_19748);
or U24582 (N_24582,N_19953,N_18543);
nor U24583 (N_24583,N_18647,N_19330);
xor U24584 (N_24584,N_15444,N_19694);
xnor U24585 (N_24585,N_18597,N_18971);
and U24586 (N_24586,N_16613,N_17651);
xor U24587 (N_24587,N_16731,N_18178);
nand U24588 (N_24588,N_16506,N_16975);
and U24589 (N_24589,N_19326,N_17819);
nand U24590 (N_24590,N_18172,N_15649);
nand U24591 (N_24591,N_18317,N_16029);
or U24592 (N_24592,N_19849,N_15452);
nand U24593 (N_24593,N_19997,N_16144);
nor U24594 (N_24594,N_18341,N_17579);
or U24595 (N_24595,N_18702,N_17589);
nand U24596 (N_24596,N_19486,N_18704);
or U24597 (N_24597,N_15284,N_17890);
and U24598 (N_24598,N_18927,N_19430);
and U24599 (N_24599,N_18411,N_18919);
and U24600 (N_24600,N_17560,N_19525);
nor U24601 (N_24601,N_17395,N_16109);
and U24602 (N_24602,N_15776,N_19312);
xor U24603 (N_24603,N_18688,N_15000);
and U24604 (N_24604,N_19564,N_17495);
and U24605 (N_24605,N_15614,N_18910);
nand U24606 (N_24606,N_19841,N_16885);
or U24607 (N_24607,N_17185,N_16913);
and U24608 (N_24608,N_19304,N_15154);
or U24609 (N_24609,N_16960,N_17852);
nor U24610 (N_24610,N_17585,N_19473);
nor U24611 (N_24611,N_15165,N_15240);
nand U24612 (N_24612,N_16617,N_18334);
nor U24613 (N_24613,N_15882,N_18600);
nand U24614 (N_24614,N_19207,N_15519);
or U24615 (N_24615,N_16199,N_16551);
nand U24616 (N_24616,N_17285,N_19980);
nand U24617 (N_24617,N_16389,N_18847);
xnor U24618 (N_24618,N_16259,N_15622);
nand U24619 (N_24619,N_18142,N_16538);
nor U24620 (N_24620,N_16193,N_19132);
or U24621 (N_24621,N_19132,N_16696);
or U24622 (N_24622,N_15132,N_19249);
and U24623 (N_24623,N_15246,N_17179);
nor U24624 (N_24624,N_18476,N_18559);
nor U24625 (N_24625,N_15587,N_15811);
nand U24626 (N_24626,N_17886,N_18551);
or U24627 (N_24627,N_17853,N_15062);
nand U24628 (N_24628,N_19966,N_16528);
nand U24629 (N_24629,N_19506,N_19401);
nor U24630 (N_24630,N_16501,N_16921);
nor U24631 (N_24631,N_15259,N_15323);
xnor U24632 (N_24632,N_17451,N_19280);
and U24633 (N_24633,N_19458,N_17510);
and U24634 (N_24634,N_18143,N_17889);
and U24635 (N_24635,N_16790,N_15595);
nand U24636 (N_24636,N_19733,N_18829);
or U24637 (N_24637,N_19155,N_19842);
or U24638 (N_24638,N_17475,N_15966);
or U24639 (N_24639,N_18580,N_15128);
xnor U24640 (N_24640,N_17741,N_19733);
and U24641 (N_24641,N_16660,N_15485);
or U24642 (N_24642,N_16185,N_18333);
or U24643 (N_24643,N_15680,N_17476);
nand U24644 (N_24644,N_15229,N_19632);
nand U24645 (N_24645,N_18377,N_17785);
or U24646 (N_24646,N_15632,N_19373);
xnor U24647 (N_24647,N_17400,N_18512);
xnor U24648 (N_24648,N_15654,N_18177);
nand U24649 (N_24649,N_19116,N_15510);
nor U24650 (N_24650,N_16395,N_17287);
or U24651 (N_24651,N_18092,N_17345);
or U24652 (N_24652,N_19090,N_17588);
nor U24653 (N_24653,N_19905,N_16107);
nor U24654 (N_24654,N_15747,N_18251);
or U24655 (N_24655,N_19359,N_17612);
and U24656 (N_24656,N_17500,N_19990);
or U24657 (N_24657,N_16794,N_19163);
nor U24658 (N_24658,N_16857,N_16987);
nor U24659 (N_24659,N_17461,N_15570);
or U24660 (N_24660,N_15519,N_15617);
and U24661 (N_24661,N_16734,N_17325);
or U24662 (N_24662,N_19613,N_16678);
xor U24663 (N_24663,N_15358,N_17217);
nor U24664 (N_24664,N_18121,N_19049);
and U24665 (N_24665,N_19285,N_19348);
xor U24666 (N_24666,N_18872,N_19570);
or U24667 (N_24667,N_16574,N_18729);
nand U24668 (N_24668,N_18885,N_17031);
and U24669 (N_24669,N_17771,N_17881);
or U24670 (N_24670,N_19249,N_18139);
and U24671 (N_24671,N_17508,N_16967);
or U24672 (N_24672,N_17695,N_17535);
and U24673 (N_24673,N_15743,N_16916);
xor U24674 (N_24674,N_18253,N_18172);
nand U24675 (N_24675,N_17788,N_15783);
nand U24676 (N_24676,N_16014,N_19236);
nor U24677 (N_24677,N_18169,N_17476);
nand U24678 (N_24678,N_16710,N_17790);
nor U24679 (N_24679,N_15749,N_16907);
or U24680 (N_24680,N_19808,N_18382);
or U24681 (N_24681,N_16084,N_18516);
or U24682 (N_24682,N_16134,N_15668);
and U24683 (N_24683,N_17794,N_15262);
nand U24684 (N_24684,N_17606,N_15207);
or U24685 (N_24685,N_17399,N_16139);
and U24686 (N_24686,N_19624,N_17633);
or U24687 (N_24687,N_15024,N_15116);
and U24688 (N_24688,N_15393,N_16873);
and U24689 (N_24689,N_15391,N_17026);
nand U24690 (N_24690,N_19151,N_15954);
and U24691 (N_24691,N_17866,N_16804);
or U24692 (N_24692,N_16457,N_18812);
and U24693 (N_24693,N_17783,N_17496);
or U24694 (N_24694,N_15947,N_17037);
xnor U24695 (N_24695,N_16378,N_16795);
or U24696 (N_24696,N_19197,N_19847);
nor U24697 (N_24697,N_15695,N_15201);
nor U24698 (N_24698,N_16237,N_19766);
nand U24699 (N_24699,N_17642,N_18867);
nand U24700 (N_24700,N_16528,N_17443);
nor U24701 (N_24701,N_17899,N_18201);
or U24702 (N_24702,N_17753,N_19373);
and U24703 (N_24703,N_15619,N_18649);
or U24704 (N_24704,N_18940,N_17662);
and U24705 (N_24705,N_18902,N_16085);
or U24706 (N_24706,N_16794,N_15048);
xor U24707 (N_24707,N_18050,N_18931);
or U24708 (N_24708,N_19289,N_16777);
nor U24709 (N_24709,N_17362,N_16902);
or U24710 (N_24710,N_18399,N_18670);
nand U24711 (N_24711,N_18442,N_15037);
nor U24712 (N_24712,N_16683,N_18984);
nor U24713 (N_24713,N_17994,N_16064);
and U24714 (N_24714,N_16725,N_18376);
xor U24715 (N_24715,N_16825,N_19739);
nand U24716 (N_24716,N_18651,N_16054);
nor U24717 (N_24717,N_19103,N_19721);
or U24718 (N_24718,N_17082,N_16072);
xor U24719 (N_24719,N_15399,N_18423);
xnor U24720 (N_24720,N_16695,N_19667);
and U24721 (N_24721,N_15125,N_18045);
or U24722 (N_24722,N_18670,N_15941);
nor U24723 (N_24723,N_18632,N_15716);
nand U24724 (N_24724,N_15410,N_16103);
or U24725 (N_24725,N_19539,N_19746);
xor U24726 (N_24726,N_18831,N_18064);
nand U24727 (N_24727,N_17708,N_19330);
or U24728 (N_24728,N_17236,N_18710);
and U24729 (N_24729,N_17862,N_19062);
and U24730 (N_24730,N_15438,N_18307);
nor U24731 (N_24731,N_17775,N_16966);
or U24732 (N_24732,N_19208,N_15435);
nor U24733 (N_24733,N_19590,N_17003);
nor U24734 (N_24734,N_18828,N_19066);
or U24735 (N_24735,N_15407,N_17822);
and U24736 (N_24736,N_18649,N_15410);
nand U24737 (N_24737,N_17338,N_18782);
nor U24738 (N_24738,N_18850,N_18532);
or U24739 (N_24739,N_15361,N_19684);
and U24740 (N_24740,N_16509,N_15172);
and U24741 (N_24741,N_19846,N_15644);
and U24742 (N_24742,N_18324,N_18762);
nor U24743 (N_24743,N_18526,N_17169);
and U24744 (N_24744,N_16658,N_19734);
nand U24745 (N_24745,N_15212,N_17889);
nand U24746 (N_24746,N_16165,N_15066);
nand U24747 (N_24747,N_19091,N_15370);
or U24748 (N_24748,N_18040,N_19719);
or U24749 (N_24749,N_19315,N_17291);
nor U24750 (N_24750,N_17603,N_15064);
and U24751 (N_24751,N_18920,N_17198);
nor U24752 (N_24752,N_15468,N_19859);
and U24753 (N_24753,N_18193,N_17426);
nand U24754 (N_24754,N_17653,N_18062);
and U24755 (N_24755,N_18947,N_15078);
xor U24756 (N_24756,N_16001,N_18375);
or U24757 (N_24757,N_16656,N_19263);
xor U24758 (N_24758,N_16729,N_18778);
or U24759 (N_24759,N_19155,N_19848);
or U24760 (N_24760,N_19279,N_17078);
or U24761 (N_24761,N_15093,N_15441);
nor U24762 (N_24762,N_17830,N_15898);
or U24763 (N_24763,N_16523,N_18348);
or U24764 (N_24764,N_17970,N_19116);
or U24765 (N_24765,N_16218,N_19576);
nand U24766 (N_24766,N_17650,N_17484);
nand U24767 (N_24767,N_16234,N_15918);
or U24768 (N_24768,N_17637,N_17618);
or U24769 (N_24769,N_17288,N_18086);
or U24770 (N_24770,N_18909,N_17308);
nand U24771 (N_24771,N_16113,N_15616);
nor U24772 (N_24772,N_16725,N_18888);
and U24773 (N_24773,N_16758,N_15456);
or U24774 (N_24774,N_17899,N_16745);
and U24775 (N_24775,N_15753,N_15735);
nor U24776 (N_24776,N_15116,N_18881);
nor U24777 (N_24777,N_15489,N_15176);
nand U24778 (N_24778,N_15209,N_16401);
nand U24779 (N_24779,N_18263,N_18522);
nor U24780 (N_24780,N_15551,N_15539);
nand U24781 (N_24781,N_16369,N_18398);
and U24782 (N_24782,N_16381,N_16300);
nor U24783 (N_24783,N_17636,N_15458);
and U24784 (N_24784,N_15478,N_17201);
and U24785 (N_24785,N_17545,N_17764);
nor U24786 (N_24786,N_17622,N_17678);
or U24787 (N_24787,N_15523,N_16689);
nand U24788 (N_24788,N_19897,N_17592);
and U24789 (N_24789,N_16012,N_17699);
nand U24790 (N_24790,N_16987,N_16666);
and U24791 (N_24791,N_16598,N_17659);
or U24792 (N_24792,N_17458,N_19561);
and U24793 (N_24793,N_19309,N_18114);
or U24794 (N_24794,N_15380,N_18655);
nand U24795 (N_24795,N_16213,N_18766);
and U24796 (N_24796,N_18530,N_17726);
nand U24797 (N_24797,N_15197,N_15355);
or U24798 (N_24798,N_19556,N_17936);
or U24799 (N_24799,N_17558,N_16702);
nand U24800 (N_24800,N_18071,N_15588);
and U24801 (N_24801,N_17640,N_17658);
nand U24802 (N_24802,N_17747,N_18932);
and U24803 (N_24803,N_19124,N_17958);
nor U24804 (N_24804,N_18370,N_17647);
xor U24805 (N_24805,N_17754,N_16885);
nor U24806 (N_24806,N_15597,N_19061);
nor U24807 (N_24807,N_16365,N_18480);
nand U24808 (N_24808,N_19421,N_17178);
nor U24809 (N_24809,N_19393,N_18617);
nor U24810 (N_24810,N_16666,N_16735);
or U24811 (N_24811,N_17577,N_17129);
nand U24812 (N_24812,N_17869,N_15088);
nand U24813 (N_24813,N_17629,N_15778);
nand U24814 (N_24814,N_17318,N_18157);
and U24815 (N_24815,N_19523,N_16034);
nand U24816 (N_24816,N_19171,N_16307);
nor U24817 (N_24817,N_15542,N_15828);
nand U24818 (N_24818,N_17965,N_17910);
nand U24819 (N_24819,N_18366,N_15597);
nor U24820 (N_24820,N_18374,N_16771);
nor U24821 (N_24821,N_18406,N_19407);
and U24822 (N_24822,N_15220,N_16561);
or U24823 (N_24823,N_15074,N_16400);
and U24824 (N_24824,N_17512,N_17716);
and U24825 (N_24825,N_17760,N_19254);
nand U24826 (N_24826,N_17416,N_17217);
or U24827 (N_24827,N_17368,N_18853);
and U24828 (N_24828,N_17870,N_18078);
nand U24829 (N_24829,N_15262,N_18367);
nand U24830 (N_24830,N_15815,N_17833);
nand U24831 (N_24831,N_15105,N_16974);
nor U24832 (N_24832,N_17785,N_17006);
xnor U24833 (N_24833,N_16977,N_16748);
nor U24834 (N_24834,N_17075,N_15640);
and U24835 (N_24835,N_15635,N_15630);
or U24836 (N_24836,N_17190,N_18311);
nand U24837 (N_24837,N_16792,N_18538);
xor U24838 (N_24838,N_16770,N_19646);
or U24839 (N_24839,N_17200,N_16495);
and U24840 (N_24840,N_19117,N_17643);
and U24841 (N_24841,N_15236,N_17981);
or U24842 (N_24842,N_16975,N_18083);
nor U24843 (N_24843,N_19025,N_18640);
nand U24844 (N_24844,N_19037,N_15324);
and U24845 (N_24845,N_15458,N_19083);
or U24846 (N_24846,N_15244,N_17182);
xnor U24847 (N_24847,N_19806,N_18638);
and U24848 (N_24848,N_17865,N_16835);
nand U24849 (N_24849,N_19530,N_15269);
xnor U24850 (N_24850,N_17890,N_16033);
xnor U24851 (N_24851,N_16264,N_16518);
xor U24852 (N_24852,N_17861,N_18090);
nand U24853 (N_24853,N_19323,N_19856);
nand U24854 (N_24854,N_19856,N_16040);
nor U24855 (N_24855,N_18956,N_18478);
nor U24856 (N_24856,N_18240,N_19235);
or U24857 (N_24857,N_16358,N_18727);
or U24858 (N_24858,N_17032,N_19575);
nand U24859 (N_24859,N_17104,N_16849);
and U24860 (N_24860,N_15751,N_19922);
nor U24861 (N_24861,N_16977,N_19155);
nand U24862 (N_24862,N_19588,N_16704);
nand U24863 (N_24863,N_18023,N_16580);
nor U24864 (N_24864,N_15853,N_17226);
xor U24865 (N_24865,N_19835,N_17605);
nor U24866 (N_24866,N_16437,N_16549);
xor U24867 (N_24867,N_17186,N_19109);
nand U24868 (N_24868,N_19442,N_16957);
or U24869 (N_24869,N_19038,N_15132);
nor U24870 (N_24870,N_19553,N_18261);
nor U24871 (N_24871,N_19601,N_17077);
xor U24872 (N_24872,N_18203,N_15967);
nand U24873 (N_24873,N_15028,N_17579);
nor U24874 (N_24874,N_17737,N_19670);
xor U24875 (N_24875,N_16718,N_18634);
xor U24876 (N_24876,N_16355,N_16768);
nor U24877 (N_24877,N_15329,N_15214);
or U24878 (N_24878,N_17829,N_18008);
nor U24879 (N_24879,N_18104,N_15824);
and U24880 (N_24880,N_18882,N_17087);
or U24881 (N_24881,N_17696,N_16923);
and U24882 (N_24882,N_15257,N_16408);
and U24883 (N_24883,N_15341,N_17819);
nor U24884 (N_24884,N_17840,N_15856);
and U24885 (N_24885,N_17815,N_17252);
and U24886 (N_24886,N_19417,N_17460);
or U24887 (N_24887,N_17959,N_17743);
and U24888 (N_24888,N_15346,N_17350);
nand U24889 (N_24889,N_18345,N_16475);
nor U24890 (N_24890,N_17637,N_16588);
xor U24891 (N_24891,N_18054,N_17361);
nand U24892 (N_24892,N_19024,N_16854);
nand U24893 (N_24893,N_15693,N_17742);
or U24894 (N_24894,N_15678,N_15826);
and U24895 (N_24895,N_16479,N_19224);
nor U24896 (N_24896,N_18538,N_17152);
nor U24897 (N_24897,N_17070,N_17002);
and U24898 (N_24898,N_15266,N_18473);
nand U24899 (N_24899,N_18182,N_15081);
xnor U24900 (N_24900,N_15784,N_15924);
and U24901 (N_24901,N_15711,N_16739);
nor U24902 (N_24902,N_17177,N_17357);
nand U24903 (N_24903,N_16802,N_19748);
nor U24904 (N_24904,N_16381,N_18610);
nand U24905 (N_24905,N_18415,N_18110);
and U24906 (N_24906,N_17762,N_17164);
or U24907 (N_24907,N_19035,N_17302);
nand U24908 (N_24908,N_18949,N_16889);
nand U24909 (N_24909,N_17013,N_17399);
or U24910 (N_24910,N_17640,N_18371);
nand U24911 (N_24911,N_16347,N_19723);
or U24912 (N_24912,N_15722,N_17665);
or U24913 (N_24913,N_17497,N_19267);
nand U24914 (N_24914,N_18639,N_16852);
nand U24915 (N_24915,N_15394,N_17658);
or U24916 (N_24916,N_18278,N_19112);
or U24917 (N_24917,N_17517,N_15946);
xor U24918 (N_24918,N_18657,N_18656);
or U24919 (N_24919,N_16667,N_18026);
nand U24920 (N_24920,N_15214,N_19558);
and U24921 (N_24921,N_18516,N_16427);
nand U24922 (N_24922,N_16135,N_18193);
nand U24923 (N_24923,N_19613,N_15078);
and U24924 (N_24924,N_15631,N_17425);
nand U24925 (N_24925,N_19412,N_17500);
and U24926 (N_24926,N_19586,N_16170);
xnor U24927 (N_24927,N_15526,N_15838);
nand U24928 (N_24928,N_16301,N_17548);
xnor U24929 (N_24929,N_19167,N_16232);
nand U24930 (N_24930,N_16406,N_18649);
and U24931 (N_24931,N_19309,N_19469);
xnor U24932 (N_24932,N_19268,N_15905);
and U24933 (N_24933,N_17157,N_16777);
xor U24934 (N_24934,N_17264,N_18020);
nand U24935 (N_24935,N_15167,N_15718);
and U24936 (N_24936,N_19103,N_18437);
or U24937 (N_24937,N_18862,N_19874);
and U24938 (N_24938,N_18229,N_15268);
and U24939 (N_24939,N_16427,N_17636);
nor U24940 (N_24940,N_19964,N_15684);
nor U24941 (N_24941,N_16835,N_17344);
nor U24942 (N_24942,N_17819,N_17554);
and U24943 (N_24943,N_15736,N_15561);
or U24944 (N_24944,N_15521,N_17693);
and U24945 (N_24945,N_18635,N_17006);
nor U24946 (N_24946,N_18826,N_19106);
and U24947 (N_24947,N_16901,N_17901);
nor U24948 (N_24948,N_19533,N_16415);
nand U24949 (N_24949,N_18642,N_15205);
and U24950 (N_24950,N_18298,N_18737);
or U24951 (N_24951,N_16517,N_17772);
nand U24952 (N_24952,N_17975,N_16864);
nor U24953 (N_24953,N_17685,N_19997);
nand U24954 (N_24954,N_17640,N_18953);
nand U24955 (N_24955,N_16427,N_19306);
nor U24956 (N_24956,N_19729,N_18410);
nor U24957 (N_24957,N_16713,N_15159);
xnor U24958 (N_24958,N_16690,N_15134);
and U24959 (N_24959,N_16143,N_19342);
and U24960 (N_24960,N_17426,N_19823);
and U24961 (N_24961,N_19376,N_18725);
nand U24962 (N_24962,N_18144,N_16385);
xor U24963 (N_24963,N_16529,N_15990);
nor U24964 (N_24964,N_19901,N_19360);
nand U24965 (N_24965,N_16018,N_19248);
and U24966 (N_24966,N_16971,N_19260);
and U24967 (N_24967,N_17063,N_18504);
nand U24968 (N_24968,N_17648,N_19605);
xor U24969 (N_24969,N_18995,N_16095);
or U24970 (N_24970,N_15894,N_15697);
nand U24971 (N_24971,N_19827,N_17622);
nor U24972 (N_24972,N_15544,N_15022);
nand U24973 (N_24973,N_19789,N_19707);
nor U24974 (N_24974,N_18069,N_19094);
nor U24975 (N_24975,N_18006,N_19855);
nand U24976 (N_24976,N_15245,N_15963);
or U24977 (N_24977,N_18827,N_18847);
nand U24978 (N_24978,N_18614,N_15860);
and U24979 (N_24979,N_16261,N_19638);
nor U24980 (N_24980,N_19486,N_19002);
xor U24981 (N_24981,N_15477,N_15638);
and U24982 (N_24982,N_18629,N_19117);
nand U24983 (N_24983,N_16083,N_19156);
nand U24984 (N_24984,N_15209,N_18066);
nor U24985 (N_24985,N_16452,N_17080);
or U24986 (N_24986,N_18338,N_18675);
nor U24987 (N_24987,N_18490,N_16907);
nand U24988 (N_24988,N_17633,N_17453);
nor U24989 (N_24989,N_18180,N_16762);
and U24990 (N_24990,N_19717,N_17806);
nand U24991 (N_24991,N_15804,N_19513);
nor U24992 (N_24992,N_19107,N_19115);
nor U24993 (N_24993,N_19327,N_19154);
xnor U24994 (N_24994,N_16131,N_16103);
or U24995 (N_24995,N_17454,N_18213);
nor U24996 (N_24996,N_17251,N_19557);
and U24997 (N_24997,N_15604,N_16557);
nand U24998 (N_24998,N_18065,N_18206);
or U24999 (N_24999,N_19546,N_19261);
or U25000 (N_25000,N_20823,N_22140);
nor U25001 (N_25001,N_23810,N_24555);
nand U25002 (N_25002,N_23986,N_22908);
and U25003 (N_25003,N_23397,N_22191);
nor U25004 (N_25004,N_24976,N_20839);
nand U25005 (N_25005,N_22825,N_21092);
or U25006 (N_25006,N_21660,N_24291);
or U25007 (N_25007,N_20526,N_22528);
or U25008 (N_25008,N_24488,N_21135);
nand U25009 (N_25009,N_21507,N_21825);
and U25010 (N_25010,N_24372,N_20500);
nand U25011 (N_25011,N_21590,N_22621);
nand U25012 (N_25012,N_20595,N_23516);
nand U25013 (N_25013,N_20181,N_24609);
and U25014 (N_25014,N_24161,N_24296);
and U25015 (N_25015,N_20545,N_22796);
or U25016 (N_25016,N_20961,N_20536);
nor U25017 (N_25017,N_23559,N_23126);
or U25018 (N_25018,N_24029,N_20202);
nor U25019 (N_25019,N_24962,N_21969);
or U25020 (N_25020,N_24384,N_24589);
nand U25021 (N_25021,N_20194,N_21000);
or U25022 (N_25022,N_23094,N_22453);
or U25023 (N_25023,N_22917,N_23467);
or U25024 (N_25024,N_24688,N_21465);
nand U25025 (N_25025,N_23602,N_20227);
nand U25026 (N_25026,N_23763,N_23342);
nand U25027 (N_25027,N_24238,N_20184);
or U25028 (N_25028,N_24708,N_20251);
nor U25029 (N_25029,N_20681,N_23685);
or U25030 (N_25030,N_20862,N_22260);
or U25031 (N_25031,N_22185,N_21118);
or U25032 (N_25032,N_20178,N_24464);
xnor U25033 (N_25033,N_24395,N_21805);
xnor U25034 (N_25034,N_20702,N_24800);
nor U25035 (N_25035,N_24821,N_22276);
or U25036 (N_25036,N_23834,N_22334);
nand U25037 (N_25037,N_23452,N_22840);
and U25038 (N_25038,N_23201,N_21966);
or U25039 (N_25039,N_20639,N_22524);
nor U25040 (N_25040,N_24135,N_23881);
and U25041 (N_25041,N_20112,N_21180);
nor U25042 (N_25042,N_24943,N_24436);
nor U25043 (N_25043,N_23059,N_24846);
and U25044 (N_25044,N_21948,N_20241);
or U25045 (N_25045,N_24293,N_21619);
nor U25046 (N_25046,N_22118,N_23999);
nand U25047 (N_25047,N_23522,N_23012);
and U25048 (N_25048,N_20389,N_22707);
nand U25049 (N_25049,N_20344,N_22009);
and U25050 (N_25050,N_24583,N_23941);
xnor U25051 (N_25051,N_20569,N_22475);
nor U25052 (N_25052,N_23242,N_23387);
xor U25053 (N_25053,N_21566,N_22685);
nand U25054 (N_25054,N_23064,N_24379);
or U25055 (N_25055,N_22561,N_23952);
nor U25056 (N_25056,N_24777,N_21833);
and U25057 (N_25057,N_20663,N_23272);
nand U25058 (N_25058,N_22277,N_23130);
nor U25059 (N_25059,N_23486,N_21959);
and U25060 (N_25060,N_21239,N_21737);
nor U25061 (N_25061,N_24919,N_24932);
nor U25062 (N_25062,N_20816,N_24234);
or U25063 (N_25063,N_22947,N_20185);
and U25064 (N_25064,N_24328,N_21129);
nand U25065 (N_25065,N_21168,N_20798);
and U25066 (N_25066,N_24792,N_21922);
nor U25067 (N_25067,N_23389,N_21537);
nor U25068 (N_25068,N_23571,N_20568);
nand U25069 (N_25069,N_23707,N_22173);
nand U25070 (N_25070,N_22636,N_23463);
nand U25071 (N_25071,N_23944,N_22697);
and U25072 (N_25072,N_23636,N_23847);
or U25073 (N_25073,N_23800,N_21269);
nand U25074 (N_25074,N_21624,N_22097);
nand U25075 (N_25075,N_23494,N_24219);
nor U25076 (N_25076,N_20606,N_20266);
nor U25077 (N_25077,N_21491,N_23036);
or U25078 (N_25078,N_21081,N_20180);
nand U25079 (N_25079,N_23395,N_23438);
xor U25080 (N_25080,N_20844,N_23381);
nand U25081 (N_25081,N_24856,N_23578);
nor U25082 (N_25082,N_20063,N_20054);
or U25083 (N_25083,N_21440,N_24515);
and U25084 (N_25084,N_22807,N_24838);
xnor U25085 (N_25085,N_21207,N_24370);
nor U25086 (N_25086,N_23660,N_24718);
xnor U25087 (N_25087,N_22152,N_24368);
nand U25088 (N_25088,N_22294,N_24223);
nand U25089 (N_25089,N_21100,N_21525);
and U25090 (N_25090,N_21375,N_24433);
or U25091 (N_25091,N_23243,N_22049);
or U25092 (N_25092,N_24710,N_21576);
nor U25093 (N_25093,N_23882,N_21898);
and U25094 (N_25094,N_20600,N_23157);
nor U25095 (N_25095,N_22045,N_21606);
and U25096 (N_25096,N_23801,N_22133);
and U25097 (N_25097,N_20279,N_20323);
nor U25098 (N_25098,N_24017,N_23367);
xnor U25099 (N_25099,N_21094,N_21668);
xor U25100 (N_25100,N_23984,N_23319);
nand U25101 (N_25101,N_23219,N_20611);
or U25102 (N_25102,N_23436,N_24117);
xor U25103 (N_25103,N_23412,N_24252);
nor U25104 (N_25104,N_24648,N_21865);
or U25105 (N_25105,N_22497,N_24891);
and U25106 (N_25106,N_22808,N_23980);
nor U25107 (N_25107,N_22650,N_20701);
or U25108 (N_25108,N_24629,N_20775);
or U25109 (N_25109,N_22229,N_24620);
nand U25110 (N_25110,N_20292,N_21199);
nand U25111 (N_25111,N_23916,N_20086);
nand U25112 (N_25112,N_23727,N_23799);
and U25113 (N_25113,N_23089,N_23599);
or U25114 (N_25114,N_23354,N_23226);
and U25115 (N_25115,N_20693,N_23159);
nand U25116 (N_25116,N_23449,N_22035);
nand U25117 (N_25117,N_24011,N_22230);
nand U25118 (N_25118,N_24256,N_24386);
and U25119 (N_25119,N_23456,N_22777);
and U25120 (N_25120,N_23920,N_20091);
nand U25121 (N_25121,N_21071,N_20578);
nand U25122 (N_25122,N_21244,N_21846);
and U25123 (N_25123,N_23379,N_22871);
nor U25124 (N_25124,N_21643,N_22929);
nand U25125 (N_25125,N_24495,N_21413);
and U25126 (N_25126,N_24260,N_21336);
or U25127 (N_25127,N_23097,N_24142);
or U25128 (N_25128,N_20311,N_20274);
nand U25129 (N_25129,N_20803,N_21773);
and U25130 (N_25130,N_20215,N_22040);
xor U25131 (N_25131,N_23924,N_23241);
and U25132 (N_25132,N_20937,N_24640);
or U25133 (N_25133,N_20341,N_22199);
nand U25134 (N_25134,N_21400,N_21160);
nand U25135 (N_25135,N_24305,N_20940);
nor U25136 (N_25136,N_23079,N_20919);
nand U25137 (N_25137,N_23992,N_23435);
nand U25138 (N_25138,N_22417,N_21720);
or U25139 (N_25139,N_23408,N_22309);
and U25140 (N_25140,N_23674,N_20784);
and U25141 (N_25141,N_20127,N_24186);
nand U25142 (N_25142,N_24568,N_20947);
or U25143 (N_25143,N_24724,N_24155);
and U25144 (N_25144,N_23694,N_24143);
and U25145 (N_25145,N_20932,N_20361);
nand U25146 (N_25146,N_22301,N_20668);
nor U25147 (N_25147,N_22938,N_20665);
nand U25148 (N_25148,N_23929,N_20108);
or U25149 (N_25149,N_22200,N_23465);
nor U25150 (N_25150,N_21884,N_21623);
or U25151 (N_25151,N_22443,N_20087);
and U25152 (N_25152,N_23560,N_22131);
xor U25153 (N_25153,N_22243,N_21323);
xnor U25154 (N_25154,N_22498,N_23060);
nor U25155 (N_25155,N_20019,N_24054);
or U25156 (N_25156,N_22911,N_24764);
nor U25157 (N_25157,N_23006,N_24771);
nand U25158 (N_25158,N_20735,N_24803);
nor U25159 (N_25159,N_24320,N_20859);
nor U25160 (N_25160,N_21298,N_24828);
or U25161 (N_25161,N_20074,N_23355);
nor U25162 (N_25162,N_22375,N_20878);
nand U25163 (N_25163,N_24214,N_24335);
nor U25164 (N_25164,N_22029,N_20783);
nor U25165 (N_25165,N_23209,N_23528);
and U25166 (N_25166,N_23915,N_22404);
nor U25167 (N_25167,N_22771,N_24626);
or U25168 (N_25168,N_20676,N_24141);
nor U25169 (N_25169,N_20880,N_22635);
or U25170 (N_25170,N_21258,N_22177);
nand U25171 (N_25171,N_21049,N_24426);
or U25172 (N_25172,N_23294,N_20722);
nor U25173 (N_25173,N_21495,N_20166);
or U25174 (N_25174,N_21126,N_22366);
and U25175 (N_25175,N_22623,N_21883);
nor U25176 (N_25176,N_22566,N_24675);
or U25177 (N_25177,N_21591,N_23865);
and U25178 (N_25178,N_20220,N_21847);
xnor U25179 (N_25179,N_24535,N_20228);
xnor U25180 (N_25180,N_24663,N_20043);
nand U25181 (N_25181,N_24352,N_20540);
or U25182 (N_25182,N_23550,N_21514);
or U25183 (N_25183,N_21377,N_21220);
or U25184 (N_25184,N_23945,N_21320);
nand U25185 (N_25185,N_24714,N_22345);
nand U25186 (N_25186,N_22515,N_20280);
nor U25187 (N_25187,N_20532,N_24888);
nor U25188 (N_25188,N_20244,N_24804);
nor U25189 (N_25189,N_24922,N_24517);
nand U25190 (N_25190,N_21785,N_20260);
and U25191 (N_25191,N_23966,N_23190);
xor U25192 (N_25192,N_21947,N_23982);
or U25193 (N_25193,N_22665,N_21638);
nand U25194 (N_25194,N_23101,N_21649);
and U25195 (N_25195,N_20754,N_23298);
nor U25196 (N_25196,N_23940,N_23797);
and U25197 (N_25197,N_20337,N_23848);
or U25198 (N_25198,N_20000,N_23587);
nand U25199 (N_25199,N_21264,N_23121);
and U25200 (N_25200,N_24079,N_24067);
or U25201 (N_25201,N_21074,N_20865);
nor U25202 (N_25202,N_20449,N_20513);
or U25203 (N_25203,N_24231,N_20629);
nand U25204 (N_25204,N_21988,N_21146);
or U25205 (N_25205,N_24940,N_21840);
or U25206 (N_25206,N_22849,N_23661);
nor U25207 (N_25207,N_21257,N_23195);
or U25208 (N_25208,N_21289,N_20902);
or U25209 (N_25209,N_24659,N_22487);
nand U25210 (N_25210,N_22760,N_23268);
nor U25211 (N_25211,N_22711,N_23380);
nand U25212 (N_25212,N_21291,N_23365);
nor U25213 (N_25213,N_20135,N_23204);
and U25214 (N_25214,N_22226,N_21792);
xnor U25215 (N_25215,N_23814,N_23754);
or U25216 (N_25216,N_20814,N_22741);
nand U25217 (N_25217,N_23642,N_21829);
nor U25218 (N_25218,N_21231,N_20424);
and U25219 (N_25219,N_21625,N_23025);
or U25220 (N_25220,N_21822,N_21471);
nor U25221 (N_25221,N_20928,N_21504);
xnor U25222 (N_25222,N_21172,N_20841);
and U25223 (N_25223,N_24298,N_24654);
nor U25224 (N_25224,N_23886,N_21395);
and U25225 (N_25225,N_23816,N_21637);
nand U25226 (N_25226,N_24059,N_24516);
and U25227 (N_25227,N_22662,N_20088);
nand U25228 (N_25228,N_21962,N_20896);
or U25229 (N_25229,N_23584,N_24192);
nand U25230 (N_25230,N_20277,N_21232);
and U25231 (N_25231,N_21658,N_24383);
xnor U25232 (N_25232,N_24807,N_23464);
nor U25233 (N_25233,N_21084,N_20633);
nand U25234 (N_25234,N_23370,N_24413);
nand U25235 (N_25235,N_21263,N_20934);
and U25236 (N_25236,N_24778,N_22794);
or U25237 (N_25237,N_22306,N_21645);
nand U25238 (N_25238,N_23231,N_24531);
xor U25239 (N_25239,N_21589,N_21817);
nor U25240 (N_25240,N_21972,N_20486);
nor U25241 (N_25241,N_23472,N_21411);
nor U25242 (N_25242,N_21615,N_22939);
xnor U25243 (N_25243,N_22074,N_23705);
xor U25244 (N_25244,N_24990,N_20697);
nor U25245 (N_25245,N_24462,N_20522);
nand U25246 (N_25246,N_23739,N_22480);
and U25247 (N_25247,N_20307,N_21524);
or U25248 (N_25248,N_22601,N_23649);
or U25249 (N_25249,N_21787,N_20363);
nor U25250 (N_25250,N_20604,N_22019);
nor U25251 (N_25251,N_23679,N_20939);
or U25252 (N_25252,N_22872,N_24797);
nand U25253 (N_25253,N_21562,N_24162);
or U25254 (N_25254,N_24077,N_24184);
or U25255 (N_25255,N_22891,N_23021);
and U25256 (N_25256,N_20335,N_24088);
xnor U25257 (N_25257,N_23360,N_23755);
and U25258 (N_25258,N_21500,N_21321);
xnor U25259 (N_25259,N_20198,N_24506);
nand U25260 (N_25260,N_24596,N_23453);
and U25261 (N_25261,N_23738,N_22839);
xor U25262 (N_25262,N_20739,N_23548);
or U25263 (N_25263,N_23022,N_20590);
nor U25264 (N_25264,N_24884,N_24574);
or U25265 (N_25265,N_24805,N_20137);
xnor U25266 (N_25266,N_20142,N_22778);
and U25267 (N_25267,N_22383,N_21498);
nand U25268 (N_25268,N_21812,N_21794);
and U25269 (N_25269,N_21770,N_24720);
and U25270 (N_25270,N_22881,N_23524);
nand U25271 (N_25271,N_23840,N_21148);
nor U25272 (N_25272,N_22928,N_24968);
nand U25273 (N_25273,N_23115,N_21088);
and U25274 (N_25274,N_22408,N_21974);
or U25275 (N_25275,N_21598,N_21360);
nand U25276 (N_25276,N_21136,N_21497);
or U25277 (N_25277,N_20471,N_20485);
and U25278 (N_25278,N_21861,N_20774);
nor U25279 (N_25279,N_21515,N_20123);
xnor U25280 (N_25280,N_24348,N_23736);
nor U25281 (N_25281,N_20340,N_22661);
and U25282 (N_25282,N_21201,N_24530);
nor U25283 (N_25283,N_22394,N_24621);
nand U25284 (N_25284,N_23903,N_21695);
nand U25285 (N_25285,N_21076,N_24867);
nand U25286 (N_25286,N_20908,N_20695);
nand U25287 (N_25287,N_22395,N_23304);
or U25288 (N_25288,N_22257,N_23518);
and U25289 (N_25289,N_21016,N_22556);
nand U25290 (N_25290,N_23374,N_23414);
or U25291 (N_25291,N_23724,N_20929);
xor U25292 (N_25292,N_24965,N_24206);
nand U25293 (N_25293,N_22570,N_21985);
nor U25294 (N_25294,N_23122,N_20685);
nand U25295 (N_25295,N_21732,N_22682);
and U25296 (N_25296,N_21130,N_20012);
or U25297 (N_25297,N_24097,N_22368);
nand U25298 (N_25298,N_23895,N_23844);
and U25299 (N_25299,N_22392,N_20484);
or U25300 (N_25300,N_20560,N_23155);
nand U25301 (N_25301,N_24406,N_21225);
and U25302 (N_25302,N_21570,N_24679);
and U25303 (N_25303,N_21422,N_24443);
or U25304 (N_25304,N_22823,N_21245);
and U25305 (N_25305,N_21032,N_22735);
and U25306 (N_25306,N_22992,N_22514);
or U25307 (N_25307,N_23855,N_22533);
nand U25308 (N_25308,N_21679,N_24566);
or U25309 (N_25309,N_24120,N_24354);
or U25310 (N_25310,N_22400,N_22985);
or U25311 (N_25311,N_23504,N_23968);
or U25312 (N_25312,N_22637,N_22071);
nor U25313 (N_25313,N_23545,N_21909);
and U25314 (N_25314,N_21192,N_21858);
nor U25315 (N_25315,N_21534,N_24561);
xnor U25316 (N_25316,N_24716,N_24420);
nor U25317 (N_25317,N_22645,N_23106);
and U25318 (N_25318,N_20231,N_21956);
nor U25319 (N_25319,N_21064,N_22154);
and U25320 (N_25320,N_23215,N_23054);
and U25321 (N_25321,N_20730,N_20162);
xor U25322 (N_25322,N_24519,N_20339);
and U25323 (N_25323,N_21155,N_23282);
and U25324 (N_25324,N_21282,N_21359);
nor U25325 (N_25325,N_22100,N_21877);
or U25326 (N_25326,N_20188,N_22675);
and U25327 (N_25327,N_20981,N_24330);
or U25328 (N_25328,N_21421,N_24437);
nor U25329 (N_25329,N_23067,N_24432);
or U25330 (N_25330,N_23203,N_23643);
and U25331 (N_25331,N_22585,N_22885);
nand U25332 (N_25332,N_24133,N_23111);
or U25333 (N_25333,N_21450,N_21803);
and U25334 (N_25334,N_24246,N_21484);
nor U25335 (N_25335,N_23476,N_21611);
or U25336 (N_25336,N_22797,N_21675);
nor U25337 (N_25337,N_20238,N_20009);
nand U25338 (N_25338,N_23720,N_24020);
and U25339 (N_25339,N_21114,N_24830);
and U25340 (N_25340,N_23393,N_24118);
xnor U25341 (N_25341,N_24013,N_23768);
and U25342 (N_25342,N_22411,N_20772);
or U25343 (N_25343,N_24496,N_23893);
nor U25344 (N_25344,N_24979,N_23985);
nand U25345 (N_25345,N_21584,N_22716);
nand U25346 (N_25346,N_21296,N_22884);
or U25347 (N_25347,N_23260,N_24014);
nor U25348 (N_25348,N_24934,N_20157);
and U25349 (N_25349,N_24652,N_22804);
or U25350 (N_25350,N_21487,N_24085);
nand U25351 (N_25351,N_20799,N_21699);
nand U25352 (N_25352,N_23134,N_24910);
or U25353 (N_25353,N_22592,N_21086);
nand U25354 (N_25354,N_24964,N_24952);
nor U25355 (N_25355,N_23131,N_21188);
nand U25356 (N_25356,N_20375,N_22695);
and U25357 (N_25357,N_20331,N_22936);
nand U25358 (N_25358,N_21496,N_24373);
or U25359 (N_25359,N_21242,N_24887);
nand U25360 (N_25360,N_22657,N_23451);
nand U25361 (N_25361,N_23049,N_23652);
nand U25362 (N_25362,N_21236,N_22630);
xnor U25363 (N_25363,N_22237,N_23280);
nand U25364 (N_25364,N_20834,N_23008);
or U25365 (N_25365,N_23507,N_23444);
nor U25366 (N_25366,N_22416,N_23969);
and U25367 (N_25367,N_20926,N_22008);
and U25368 (N_25368,N_23618,N_20398);
nand U25369 (N_25369,N_20942,N_22166);
nor U25370 (N_25370,N_23626,N_23346);
nand U25371 (N_25371,N_20868,N_20721);
xnor U25372 (N_25372,N_24048,N_20423);
nand U25373 (N_25373,N_20014,N_21713);
xor U25374 (N_25374,N_23933,N_20421);
xnor U25375 (N_25375,N_22783,N_24216);
nand U25376 (N_25376,N_24410,N_20535);
or U25377 (N_25377,N_21018,N_22362);
nor U25378 (N_25378,N_22587,N_21511);
and U25379 (N_25379,N_21080,N_21597);
nor U25380 (N_25380,N_24545,N_22494);
or U25381 (N_25381,N_24146,N_20999);
or U25382 (N_25382,N_22412,N_23363);
nand U25383 (N_25383,N_23748,N_23867);
and U25384 (N_25384,N_22983,N_22349);
or U25385 (N_25385,N_24906,N_23311);
xnor U25386 (N_25386,N_22111,N_24448);
or U25387 (N_25387,N_20347,N_24992);
or U25388 (N_25388,N_21572,N_23430);
xnor U25389 (N_25389,N_23468,N_23339);
nand U25390 (N_25390,N_21857,N_24282);
and U25391 (N_25391,N_22397,N_23778);
nor U25392 (N_25392,N_21733,N_24752);
or U25393 (N_25393,N_21617,N_23492);
or U25394 (N_25394,N_20512,N_24265);
and U25395 (N_25395,N_24055,N_21738);
and U25396 (N_25396,N_24336,N_20516);
and U25397 (N_25397,N_24984,N_22844);
and U25398 (N_25398,N_23854,N_22244);
nand U25399 (N_25399,N_20904,N_23017);
nand U25400 (N_25400,N_23588,N_24969);
xor U25401 (N_25401,N_22754,N_21169);
xnor U25402 (N_25402,N_22128,N_23706);
nand U25403 (N_25403,N_24164,N_20313);
and U25404 (N_25404,N_24447,N_20534);
or U25405 (N_25405,N_24202,N_20410);
nand U25406 (N_25406,N_22119,N_24889);
and U25407 (N_25407,N_22041,N_24614);
or U25408 (N_25408,N_21548,N_20315);
and U25409 (N_25409,N_22036,N_21218);
or U25410 (N_25410,N_20236,N_23872);
nand U25411 (N_25411,N_23296,N_23330);
nand U25412 (N_25412,N_24485,N_24457);
nand U25413 (N_25413,N_20778,N_23841);
nor U25414 (N_25414,N_21430,N_20890);
nor U25415 (N_25415,N_22496,N_22543);
and U25416 (N_25416,N_23759,N_21328);
nand U25417 (N_25417,N_20317,N_23258);
or U25418 (N_25418,N_21585,N_23782);
nand U25419 (N_25419,N_24949,N_20973);
and U25420 (N_25420,N_24405,N_23827);
nand U25421 (N_25421,N_21299,N_22051);
and U25422 (N_25422,N_21594,N_24998);
nand U25423 (N_25423,N_24418,N_20698);
nor U25424 (N_25424,N_20687,N_23836);
or U25425 (N_25425,N_20713,N_23216);
and U25426 (N_25426,N_22452,N_24435);
nor U25427 (N_25427,N_20630,N_23005);
nand U25428 (N_25428,N_23349,N_20777);
nand U25429 (N_25429,N_20064,N_21826);
and U25430 (N_25430,N_23657,N_23352);
and U25431 (N_25431,N_24820,N_21272);
nand U25432 (N_25432,N_22761,N_24378);
and U25433 (N_25433,N_21653,N_21103);
and U25434 (N_25434,N_21120,N_23116);
and U25435 (N_25435,N_23956,N_22999);
xor U25436 (N_25436,N_24560,N_24149);
and U25437 (N_25437,N_23270,N_21429);
nor U25438 (N_25438,N_24624,N_21670);
nor U25439 (N_25439,N_23417,N_23338);
nor U25440 (N_25440,N_24997,N_24063);
nand U25441 (N_25441,N_24078,N_20933);
and U25442 (N_25442,N_20971,N_23611);
nor U25443 (N_25443,N_21486,N_22210);
nand U25444 (N_25444,N_23109,N_20505);
and U25445 (N_25445,N_22098,N_20978);
and U25446 (N_25446,N_24595,N_22755);
or U25447 (N_25447,N_22337,N_20243);
nor U25448 (N_25448,N_20051,N_24955);
nor U25449 (N_25449,N_22335,N_22278);
nand U25450 (N_25450,N_23150,N_20343);
and U25451 (N_25451,N_20916,N_21751);
or U25452 (N_25452,N_22921,N_21179);
xnor U25453 (N_25453,N_21930,N_20224);
nand U25454 (N_25454,N_20993,N_22263);
or U25455 (N_25455,N_24001,N_24070);
nor U25456 (N_25456,N_22591,N_23491);
nor U25457 (N_25457,N_23133,N_23870);
or U25458 (N_25458,N_24611,N_21804);
or U25459 (N_25459,N_22221,N_20822);
and U25460 (N_25460,N_21979,N_23108);
nand U25461 (N_25461,N_22284,N_22866);
xnor U25462 (N_25462,N_21655,N_20764);
nand U25463 (N_25463,N_23223,N_23563);
xnor U25464 (N_25464,N_24637,N_22510);
xnor U25465 (N_25465,N_22747,N_22973);
and U25466 (N_25466,N_24254,N_24774);
and U25467 (N_25467,N_23890,N_21467);
nor U25468 (N_25468,N_22135,N_23011);
or U25469 (N_25469,N_24908,N_24757);
and U25470 (N_25470,N_21676,N_20298);
xor U25471 (N_25471,N_23271,N_22932);
nor U25472 (N_25472,N_20710,N_24257);
or U25473 (N_25473,N_24333,N_20502);
nor U25474 (N_25474,N_24662,N_22781);
or U25475 (N_25475,N_22553,N_22901);
nor U25476 (N_25476,N_20818,N_21993);
or U25477 (N_25477,N_21480,N_20434);
and U25478 (N_25478,N_20474,N_22419);
and U25479 (N_25479,N_20567,N_22664);
nand U25480 (N_25480,N_23832,N_22252);
or U25481 (N_25481,N_21708,N_24314);
or U25482 (N_25482,N_24930,N_22205);
and U25483 (N_25483,N_20021,N_23628);
or U25484 (N_25484,N_24579,N_21006);
and U25485 (N_25485,N_24538,N_24036);
nand U25486 (N_25486,N_21905,N_22956);
and U25487 (N_25487,N_22421,N_20979);
nand U25488 (N_25488,N_20734,N_21902);
xor U25489 (N_25489,N_24490,N_23525);
nand U25490 (N_25490,N_21651,N_22508);
nor U25491 (N_25491,N_23697,N_23220);
nor U25492 (N_25492,N_23441,N_21193);
nand U25493 (N_25493,N_20518,N_20376);
xnor U25494 (N_25494,N_21116,N_24750);
nor U25495 (N_25495,N_23206,N_24492);
and U25496 (N_25496,N_23345,N_23478);
nor U25497 (N_25497,N_24107,N_24529);
nand U25498 (N_25498,N_22900,N_21780);
or U25499 (N_25499,N_21221,N_23781);
nand U25500 (N_25500,N_20571,N_21262);
nor U25501 (N_25501,N_21513,N_21381);
nor U25502 (N_25502,N_22355,N_22038);
nand U25503 (N_25503,N_21227,N_22204);
nand U25504 (N_25504,N_21364,N_22762);
nand U25505 (N_25505,N_21629,N_22527);
nand U25506 (N_25506,N_22841,N_22256);
nor U25507 (N_25507,N_20432,N_22668);
nand U25508 (N_25508,N_21012,N_22679);
nor U25509 (N_25509,N_23301,N_21752);
xnor U25510 (N_25510,N_23796,N_23600);
nand U25511 (N_25511,N_24670,N_23990);
nor U25512 (N_25512,N_23087,N_21712);
nor U25513 (N_25513,N_21784,N_24890);
nand U25514 (N_25514,N_24172,N_22271);
xnor U25515 (N_25515,N_22802,N_20742);
or U25516 (N_25516,N_20189,N_22867);
nor U25517 (N_25517,N_22085,N_20860);
nor U25518 (N_25518,N_22779,N_20580);
nand U25519 (N_25519,N_22300,N_24781);
or U25520 (N_25520,N_20334,N_23018);
xor U25521 (N_25521,N_21944,N_23068);
nand U25522 (N_25522,N_20027,N_20883);
and U25523 (N_25523,N_24267,N_20422);
xor U25524 (N_25524,N_22320,N_24102);
xor U25525 (N_25525,N_24513,N_21137);
and U25526 (N_25526,N_20373,N_24871);
nor U25527 (N_25527,N_23960,N_21771);
nor U25528 (N_25528,N_22731,N_23061);
and U25529 (N_25529,N_21442,N_23678);
or U25530 (N_25530,N_21078,N_23539);
or U25531 (N_25531,N_20163,N_24493);
or U25532 (N_25532,N_21023,N_21229);
nor U25533 (N_25533,N_23048,N_20179);
xnor U25534 (N_25534,N_23041,N_22367);
and U25535 (N_25535,N_21910,N_21407);
nor U25536 (N_25536,N_23020,N_22902);
nand U25537 (N_25537,N_23780,N_22095);
nor U25538 (N_25538,N_24879,N_21308);
or U25539 (N_25539,N_24342,N_20465);
xor U25540 (N_25540,N_22788,N_23230);
or U25541 (N_25541,N_24207,N_22325);
and U25542 (N_25542,N_22634,N_21709);
nand U25543 (N_25543,N_22445,N_24967);
nand U25544 (N_25544,N_20053,N_24737);
nor U25545 (N_25545,N_24111,N_22491);
nor U25546 (N_25546,N_23922,N_20404);
nand U25547 (N_25547,N_20128,N_23149);
nand U25548 (N_25548,N_20766,N_20662);
and U25549 (N_25549,N_24853,N_20254);
nor U25550 (N_25550,N_21459,N_20072);
xor U25551 (N_25551,N_21517,N_23750);
nand U25552 (N_25552,N_20538,N_22838);
nand U25553 (N_25553,N_21690,N_22120);
nand U25554 (N_25554,N_20106,N_20643);
or U25555 (N_25555,N_22162,N_24950);
nor U25556 (N_25556,N_20195,N_20609);
nor U25557 (N_25557,N_21678,N_21431);
nor U25558 (N_25558,N_23932,N_22670);
nor U25559 (N_25559,N_22604,N_22304);
nor U25560 (N_25560,N_20959,N_24822);
or U25561 (N_25561,N_20483,N_24527);
or U25562 (N_25562,N_23863,N_22490);
or U25563 (N_25563,N_23948,N_20007);
nor U25564 (N_25564,N_22544,N_23324);
xnor U25565 (N_25565,N_22422,N_23426);
nor U25566 (N_25566,N_21565,N_21319);
and U25567 (N_25567,N_24061,N_23098);
or U25568 (N_25568,N_24936,N_21276);
and U25569 (N_25569,N_21786,N_23634);
xnor U25570 (N_25570,N_24116,N_24458);
and U25571 (N_25571,N_20281,N_20969);
nor U25572 (N_25572,N_22582,N_23371);
or U25573 (N_25573,N_23889,N_21281);
or U25574 (N_25574,N_22050,N_20468);
xor U25575 (N_25575,N_22242,N_23176);
nand U25576 (N_25576,N_23798,N_21474);
and U25577 (N_25577,N_20488,N_23034);
and U25578 (N_25578,N_20924,N_24575);
nand U25579 (N_25579,N_24677,N_21604);
or U25580 (N_25580,N_20792,N_22080);
nand U25581 (N_25581,N_23987,N_22192);
nand U25582 (N_25582,N_22141,N_22217);
or U25583 (N_25583,N_21592,N_24726);
nand U25584 (N_25584,N_24809,N_24366);
or U25585 (N_25585,N_20183,N_24369);
nor U25586 (N_25586,N_22768,N_22603);
nand U25587 (N_25587,N_20305,N_23107);
nor U25588 (N_25588,N_22676,N_22843);
nor U25589 (N_25589,N_21582,N_21349);
nor U25590 (N_25590,N_20297,N_21931);
and U25591 (N_25591,N_20399,N_22212);
nand U25592 (N_25592,N_23536,N_21243);
or U25593 (N_25593,N_21749,N_24518);
nor U25594 (N_25594,N_20028,N_24428);
and U25595 (N_25595,N_22156,N_23862);
or U25596 (N_25596,N_20230,N_22894);
and U25597 (N_25597,N_23429,N_20820);
or U25598 (N_25598,N_23983,N_22190);
nand U25599 (N_25599,N_21482,N_21834);
nand U25600 (N_25600,N_23335,N_24126);
or U25601 (N_25601,N_24053,N_21772);
and U25602 (N_25602,N_23078,N_24041);
or U25603 (N_25603,N_23630,N_22672);
xnor U25604 (N_25604,N_22403,N_20673);
nor U25605 (N_25605,N_24152,N_24294);
nor U25606 (N_25606,N_22865,N_23719);
nor U25607 (N_25607,N_22158,N_20237);
nor U25608 (N_25608,N_21929,N_21519);
nor U25609 (N_25609,N_22898,N_22574);
nand U25610 (N_25610,N_20067,N_22203);
or U25611 (N_25611,N_22774,N_23459);
nor U25612 (N_25612,N_20977,N_21721);
or U25613 (N_25613,N_21705,N_20700);
xnor U25614 (N_25614,N_23624,N_20499);
and U25615 (N_25615,N_24885,N_20160);
nand U25616 (N_25616,N_20296,N_23158);
and U25617 (N_25617,N_20105,N_24883);
nand U25618 (N_25618,N_22361,N_22608);
or U25619 (N_25619,N_20118,N_22954);
nor U25620 (N_25620,N_23955,N_23809);
nor U25621 (N_25621,N_23266,N_21424);
nand U25622 (N_25622,N_22854,N_21579);
nand U25623 (N_25623,N_23103,N_21398);
nand U25624 (N_25624,N_24235,N_20650);
or U25625 (N_25625,N_23182,N_23306);
nor U25626 (N_25626,N_22642,N_21404);
nor U25627 (N_25627,N_23473,N_23237);
nand U25628 (N_25628,N_20174,N_22409);
nor U25629 (N_25629,N_22577,N_24074);
or U25630 (N_25630,N_23957,N_21195);
nand U25631 (N_25631,N_21880,N_22913);
nand U25632 (N_25632,N_23937,N_23648);
and U25633 (N_25633,N_20678,N_21370);
or U25634 (N_25634,N_24303,N_20035);
nor U25635 (N_25635,N_20061,N_21158);
nand U25636 (N_25636,N_24550,N_23723);
and U25637 (N_25637,N_23631,N_22742);
nor U25638 (N_25638,N_24281,N_21756);
or U25639 (N_25639,N_21631,N_21776);
xor U25640 (N_25640,N_22389,N_20656);
and U25641 (N_25641,N_20392,N_20390);
or U25642 (N_25642,N_24251,N_23047);
nor U25643 (N_25643,N_22460,N_24364);
xor U25644 (N_25644,N_21161,N_20728);
and U25645 (N_25645,N_23073,N_21964);
and U25646 (N_25646,N_24416,N_22449);
xnor U25647 (N_25647,N_23256,N_22018);
and U25648 (N_25648,N_21121,N_21415);
and U25649 (N_25649,N_21823,N_23805);
nor U25650 (N_25650,N_24080,N_22324);
xnor U25651 (N_25651,N_21314,N_20750);
and U25652 (N_25652,N_21197,N_24478);
or U25653 (N_25653,N_24732,N_24317);
nand U25654 (N_25654,N_22084,N_24907);
nor U25655 (N_25655,N_20819,N_22907);
or U25656 (N_25656,N_22398,N_22348);
nor U25657 (N_25657,N_22495,N_24586);
nor U25658 (N_25658,N_22889,N_24593);
or U25659 (N_25659,N_21790,N_24835);
and U25660 (N_25660,N_20885,N_21564);
nand U25661 (N_25661,N_23977,N_22091);
nor U25662 (N_25662,N_23919,N_22671);
nand U25663 (N_25663,N_22997,N_23289);
or U25664 (N_25664,N_24319,N_21134);
nand U25665 (N_25665,N_22336,N_20922);
xnor U25666 (N_25666,N_24359,N_21997);
and U25667 (N_25667,N_22569,N_22817);
nand U25668 (N_25668,N_21141,N_22236);
nand U25669 (N_25669,N_24963,N_22955);
nor U25670 (N_25670,N_21070,N_21607);
nand U25671 (N_25671,N_22931,N_21952);
or U25672 (N_25672,N_24877,N_21358);
xor U25673 (N_25673,N_24588,N_22145);
xor U25674 (N_25674,N_23586,N_21154);
or U25675 (N_25675,N_24403,N_23052);
nand U25676 (N_25676,N_21067,N_22425);
and U25677 (N_25677,N_22168,N_20167);
xor U25678 (N_25678,N_22127,N_20915);
or U25679 (N_25679,N_21710,N_21209);
nor U25680 (N_25680,N_20621,N_22328);
xnor U25681 (N_25681,N_20460,N_22589);
xnor U25682 (N_25682,N_24722,N_20594);
or U25683 (N_25683,N_23553,N_20077);
and U25684 (N_25684,N_24543,N_21991);
and U25685 (N_25685,N_23019,N_24743);
nand U25686 (N_25686,N_23787,N_24084);
nand U25687 (N_25687,N_22241,N_22012);
or U25688 (N_25688,N_23807,N_23625);
nand U25689 (N_25689,N_24604,N_22146);
and U25690 (N_25690,N_24179,N_22991);
or U25691 (N_25691,N_24340,N_21734);
or U25692 (N_25692,N_21935,N_22951);
nor U25693 (N_25693,N_21028,N_23030);
or U25694 (N_25694,N_20645,N_21108);
xor U25695 (N_25695,N_24845,N_21378);
or U25696 (N_25696,N_23415,N_20548);
nor U25697 (N_25697,N_24977,N_24449);
nand U25698 (N_25698,N_20737,N_20755);
and U25699 (N_25699,N_22883,N_24617);
or U25700 (N_25700,N_23316,N_20956);
or U25701 (N_25701,N_20125,N_24010);
xor U25702 (N_25702,N_23655,N_22385);
nand U25703 (N_25703,N_22208,N_23573);
and U25704 (N_25704,N_21026,N_24315);
and U25705 (N_25705,N_20328,N_24758);
or U25706 (N_25706,N_21925,N_22597);
nor U25707 (N_25707,N_20093,N_20152);
nor U25708 (N_25708,N_24258,N_22406);
nand U25709 (N_25709,N_21706,N_20554);
xnor U25710 (N_25710,N_21181,N_20425);
nand U25711 (N_25711,N_21975,N_24991);
nand U25712 (N_25712,N_22072,N_22869);
nor U25713 (N_25713,N_20131,N_23859);
nand U25714 (N_25714,N_22580,N_22732);
and U25715 (N_25715,N_22520,N_21949);
nand U25716 (N_25716,N_23619,N_21133);
nand U25717 (N_25717,N_20338,N_20610);
xor U25718 (N_25718,N_23007,N_22545);
or U25719 (N_25719,N_24183,N_20412);
xnor U25720 (N_25720,N_24066,N_22934);
xnor U25721 (N_25721,N_24701,N_22317);
or U25722 (N_25722,N_20843,N_23469);
nand U25723 (N_25723,N_22752,N_20849);
or U25724 (N_25724,N_20989,N_24880);
nor U25725 (N_25725,N_24297,N_24082);
nor U25726 (N_25726,N_23579,N_24279);
nor U25727 (N_25727,N_22612,N_20100);
xnor U25728 (N_25728,N_22506,N_21224);
and U25729 (N_25729,N_22622,N_20666);
and U25730 (N_25730,N_21249,N_21390);
and U25731 (N_25731,N_21351,N_21009);
nand U25732 (N_25732,N_24641,N_22522);
and U25733 (N_25733,N_21961,N_22151);
and U25734 (N_25734,N_23302,N_22681);
and U25735 (N_25735,N_21163,N_21444);
nand U25736 (N_25736,N_23564,N_21600);
and U25737 (N_25737,N_24801,N_23818);
or U25738 (N_25738,N_23285,N_23917);
nand U25739 (N_25739,N_20032,N_20634);
nor U25740 (N_25740,N_23547,N_20330);
or U25741 (N_25741,N_24032,N_22848);
or U25742 (N_25742,N_22851,N_24759);
nor U25743 (N_25743,N_22811,N_24230);
and U25744 (N_25744,N_24220,N_21342);
or U25745 (N_25745,N_20531,N_22459);
and U25746 (N_25746,N_21832,N_24338);
or U25747 (N_25747,N_24563,N_24477);
and U25748 (N_25748,N_22792,N_20738);
and U25749 (N_25749,N_21062,N_21639);
and U25750 (N_25750,N_22968,N_22196);
nor U25751 (N_25751,N_21315,N_20954);
nor U25752 (N_25752,N_24438,N_21950);
nand U25753 (N_25753,N_21543,N_22618);
and U25754 (N_25754,N_23811,N_21698);
xor U25755 (N_25755,N_21473,N_24430);
and U25756 (N_25756,N_22194,N_20262);
or U25757 (N_25757,N_24878,N_21819);
and U25758 (N_25758,N_24431,N_22766);
and U25759 (N_25759,N_20866,N_23138);
nor U25760 (N_25760,N_22734,N_24556);
xnor U25761 (N_25761,N_20041,N_20359);
nor U25762 (N_25762,N_20519,N_20636);
or U25763 (N_25763,N_20065,N_23320);
and U25764 (N_25764,N_22189,N_20173);
or U25765 (N_25765,N_24788,N_24239);
nand U25766 (N_25766,N_21233,N_20763);
nor U25767 (N_25767,N_23789,N_21657);
or U25768 (N_25768,N_21970,N_24236);
or U25769 (N_25769,N_24684,N_22673);
nor U25770 (N_25770,N_23099,N_20414);
or U25771 (N_25771,N_22677,N_24043);
nand U25772 (N_25772,N_23398,N_24429);
xnor U25773 (N_25773,N_20970,N_20658);
and U25774 (N_25774,N_22896,N_21438);
or U25775 (N_25775,N_21849,N_24866);
nor U25776 (N_25776,N_24746,N_21672);
nor U25777 (N_25777,N_24407,N_23341);
and U25778 (N_25778,N_21726,N_22926);
xor U25779 (N_25779,N_23257,N_24608);
or U25780 (N_25780,N_21287,N_21481);
and U25781 (N_25781,N_21273,N_24134);
nand U25782 (N_25782,N_21492,N_23267);
nand U25783 (N_25783,N_20440,N_23044);
nand U25784 (N_25784,N_23632,N_24795);
xor U25785 (N_25785,N_20056,N_24042);
and U25786 (N_25786,N_21106,N_21848);
nand U25787 (N_25787,N_20787,N_24334);
nor U25788 (N_25788,N_22255,N_23093);
nor U25789 (N_25789,N_24473,N_21642);
or U25790 (N_25790,N_20443,N_20632);
nor U25791 (N_25791,N_21361,N_21339);
nand U25792 (N_25792,N_24818,N_23621);
or U25793 (N_25793,N_23066,N_22530);
and U25794 (N_25794,N_20952,N_20913);
nor U25795 (N_25795,N_22503,N_23071);
or U25796 (N_25796,N_21477,N_23549);
and U25797 (N_25797,N_20680,N_22970);
nand U25798 (N_25798,N_22446,N_24549);
and U25799 (N_25799,N_20852,N_20256);
or U25800 (N_25800,N_24019,N_20062);
nor U25801 (N_25801,N_23262,N_20884);
nor U25802 (N_25802,N_24669,N_23928);
or U25803 (N_25803,N_23198,N_21455);
xnor U25804 (N_25804,N_23165,N_23425);
and U25805 (N_25805,N_23521,N_20893);
and U25806 (N_25806,N_24768,N_23383);
and U25807 (N_25807,N_21654,N_20172);
nand U25808 (N_25808,N_23498,N_21723);
or U25809 (N_25809,N_22104,N_22683);
or U25810 (N_25810,N_23480,N_21418);
nor U25811 (N_25811,N_21799,N_23028);
or U25812 (N_25812,N_22903,N_20097);
or U25813 (N_25813,N_24696,N_20217);
and U25814 (N_25814,N_20581,N_20771);
or U25815 (N_25815,N_23185,N_20807);
nand U25816 (N_25816,N_20039,N_23733);
nor U25817 (N_25817,N_23749,N_20439);
nor U25818 (N_25818,N_22596,N_24819);
xor U25819 (N_25819,N_24497,N_24502);
nand U25820 (N_25820,N_23213,N_23804);
and U25821 (N_25821,N_23416,N_24105);
xnor U25822 (N_25822,N_20158,N_20200);
nor U25823 (N_25823,N_20757,N_22980);
or U25824 (N_25824,N_20631,N_20825);
or U25825 (N_25825,N_20199,N_23869);
nor U25826 (N_25826,N_24189,N_23812);
and U25827 (N_25827,N_23765,N_24510);
nand U25828 (N_25828,N_23527,N_22853);
and U25829 (N_25829,N_20800,N_22897);
nand U25830 (N_25830,N_21104,N_20618);
nor U25831 (N_25831,N_21238,N_22784);
nor U25832 (N_25832,N_20442,N_22467);
or U25833 (N_25833,N_22831,N_23662);
or U25834 (N_25834,N_20306,N_21237);
or U25835 (N_25835,N_22481,N_24785);
and U25836 (N_25836,N_21754,N_23233);
nor U25837 (N_25837,N_23934,N_23609);
or U25838 (N_25838,N_24101,N_20603);
xor U25839 (N_25839,N_24259,N_24988);
nand U25840 (N_25840,N_20249,N_24355);
xnor U25841 (N_25841,N_20677,N_24633);
xor U25842 (N_25842,N_21926,N_23376);
nand U25843 (N_25843,N_20965,N_20229);
nand U25844 (N_25844,N_24049,N_23428);
and U25845 (N_25845,N_21346,N_23831);
nor U25846 (N_25846,N_20674,N_23063);
nor U25847 (N_25847,N_22060,N_20126);
nor U25848 (N_25848,N_22169,N_20848);
xor U25849 (N_25849,N_24138,N_23152);
nor U25850 (N_25850,N_20216,N_24918);
nor U25851 (N_25851,N_20070,N_24931);
xnor U25852 (N_25852,N_20891,N_20371);
or U25853 (N_25853,N_20177,N_20299);
and U25854 (N_25854,N_24250,N_20462);
xor U25855 (N_25855,N_22882,N_22377);
nand U25856 (N_25856,N_20809,N_21553);
or U25857 (N_25857,N_24182,N_21788);
xor U25858 (N_25858,N_20796,N_22715);
or U25859 (N_25859,N_23457,N_20095);
nor U25860 (N_25860,N_24773,N_24199);
and U25861 (N_25861,N_24012,N_23205);
nand U25862 (N_25862,N_23513,N_23568);
nor U25863 (N_25863,N_24747,N_24212);
nand U25864 (N_25864,N_20143,N_23144);
or U25865 (N_25865,N_23721,N_22423);
or U25866 (N_25866,N_20303,N_21419);
or U25867 (N_25867,N_21447,N_23731);
nor U25868 (N_25868,N_23647,N_23189);
and U25869 (N_25869,N_21664,N_24110);
and U25870 (N_25870,N_20503,N_20046);
nor U25871 (N_25871,N_22137,N_24958);
nor U25872 (N_25872,N_21938,N_23538);
nor U25873 (N_25873,N_23254,N_24625);
xor U25874 (N_25874,N_23331,N_21414);
or U25875 (N_25875,N_24397,N_21908);
nor U25876 (N_25876,N_22437,N_23835);
and U25877 (N_25877,N_22550,N_23830);
nor U25878 (N_25878,N_21596,N_23279);
nand U25879 (N_25879,N_22013,N_20293);
nand U25880 (N_25880,N_23500,N_21448);
xor U25881 (N_25881,N_23967,N_24736);
nand U25882 (N_25882,N_22032,N_21689);
or U25883 (N_25883,N_21707,N_20886);
nand U25884 (N_25884,N_21942,N_20426);
and U25885 (N_25885,N_22359,N_24542);
and U25886 (N_25886,N_22782,N_20467);
and U25887 (N_25887,N_24201,N_24094);
or U25888 (N_25888,N_21499,N_23766);
nand U25889 (N_25889,N_23169,N_22505);
nor U25890 (N_25890,N_23291,N_21716);
or U25891 (N_25891,N_24656,N_21363);
nand U25892 (N_25892,N_23259,N_24467);
and U25893 (N_25893,N_22314,N_22967);
xnor U25894 (N_25894,N_20549,N_23391);
or U25895 (N_25895,N_20129,N_21095);
xor U25896 (N_25896,N_23171,N_23989);
and U25897 (N_25897,N_22644,N_24249);
xnor U25898 (N_25898,N_24829,N_20972);
nor U25899 (N_25899,N_22113,N_23656);
nor U25900 (N_25900,N_23803,N_20030);
or U25901 (N_25901,N_21250,N_23070);
nand U25902 (N_25902,N_22178,N_24841);
nand U25903 (N_25903,N_23644,N_20116);
nand U25904 (N_25904,N_21920,N_22182);
nand U25905 (N_25905,N_21888,N_20557);
nand U25906 (N_25906,N_22435,N_24099);
nor U25907 (N_25907,N_23874,N_21873);
or U25908 (N_25908,N_24304,N_24713);
nor U25909 (N_25909,N_24240,N_24005);
nand U25910 (N_25910,N_21050,N_24361);
or U25911 (N_25911,N_21722,N_20583);
and U25912 (N_25912,N_20246,N_23042);
or U25913 (N_25913,N_20081,N_20983);
nand U25914 (N_25914,N_23758,N_23995);
and U25915 (N_25915,N_22039,N_22611);
nor U25916 (N_25916,N_22835,N_21982);
xor U25917 (N_25917,N_24044,N_22303);
nand U25918 (N_25918,N_23368,N_20923);
or U25919 (N_25919,N_22424,N_20209);
xor U25920 (N_25920,N_23462,N_21743);
and U25921 (N_25921,N_23015,N_22989);
nor U25922 (N_25922,N_23085,N_21051);
nor U25923 (N_25923,N_22919,N_23461);
nor U25924 (N_25924,N_20193,N_23240);
or U25925 (N_25925,N_20684,N_22380);
and U25926 (N_25926,N_24974,N_23308);
nand U25927 (N_25927,N_21563,N_22905);
or U25928 (N_25928,N_21850,N_23911);
or U25929 (N_25929,N_24711,N_20407);
nand U25930 (N_25930,N_22541,N_24564);
nand U25931 (N_25931,N_20769,N_22826);
or U25932 (N_25932,N_22620,N_23753);
nor U25933 (N_25933,N_21085,N_20707);
and U25934 (N_25934,N_23792,N_24664);
xor U25935 (N_25935,N_20864,N_20950);
nand U25936 (N_25936,N_21152,N_20588);
nand U25937 (N_25937,N_24008,N_20994);
or U25938 (N_25938,N_20478,N_21357);
or U25939 (N_25939,N_22870,N_20770);
and U25940 (N_25940,N_24093,N_23785);
xnor U25941 (N_25941,N_23475,N_22197);
nor U25942 (N_25942,N_24037,N_20605);
nor U25943 (N_25943,N_24494,N_24790);
nand U25944 (N_25944,N_22370,N_22474);
nand U25945 (N_25945,N_21310,N_23817);
or U25946 (N_25946,N_23434,N_23390);
xor U25947 (N_25947,N_20149,N_24444);
nand U25948 (N_25948,N_20316,N_24709);
or U25949 (N_25949,N_22861,N_21696);
nor U25950 (N_25950,N_24571,N_22486);
and U25951 (N_25951,N_21878,N_23535);
nand U25952 (N_25952,N_24039,N_21919);
nor U25953 (N_25953,N_24071,N_23726);
or U25954 (N_25954,N_21508,N_20463);
nand U25955 (N_25955,N_22836,N_20708);
nand U25956 (N_25956,N_21580,N_20627);
or U25957 (N_25957,N_23964,N_20614);
nor U25958 (N_25958,N_22770,N_23988);
nand U25959 (N_25959,N_20894,N_23160);
or U25960 (N_25960,N_21350,N_24414);
nand U25961 (N_25961,N_21386,N_22232);
nand U25962 (N_25962,N_20552,N_20638);
or U25963 (N_25963,N_24376,N_23377);
nand U25964 (N_25964,N_24948,N_20741);
xnor U25965 (N_25965,N_21586,N_23615);
and U25966 (N_25966,N_23653,N_23446);
nor U25967 (N_25967,N_22511,N_24533);
nand U25968 (N_25968,N_20948,N_22964);
or U25969 (N_25969,N_23269,N_21427);
xnor U25970 (N_25970,N_21240,N_22772);
xnor U25971 (N_25971,N_23821,N_21860);
nor U25972 (N_25972,N_20619,N_24453);
and U25973 (N_25973,N_21656,N_22720);
and U25974 (N_25974,N_22436,N_24668);
nand U25975 (N_25975,N_22687,N_20287);
and U25976 (N_25976,N_24087,N_21379);
nand U25977 (N_25977,N_23418,N_22824);
or U25978 (N_25978,N_21522,N_23406);
nand U25979 (N_25979,N_20250,N_24165);
nor U25980 (N_25980,N_21762,N_21216);
nor U25981 (N_25981,N_20596,N_23088);
or U25982 (N_25982,N_24623,N_21778);
or U25983 (N_25983,N_23004,N_21200);
and U25984 (N_25984,N_20378,N_24300);
nand U25985 (N_25985,N_23953,N_24526);
nand U25986 (N_25986,N_21228,N_23092);
and U25987 (N_25987,N_20551,N_22923);
or U25988 (N_25988,N_24893,N_24501);
nor U25989 (N_25989,N_22063,N_22942);
nand U25990 (N_25990,N_24959,N_22022);
nor U25991 (N_25991,N_21864,N_23253);
nand U25992 (N_25992,N_24802,N_23074);
or U25993 (N_25993,N_23357,N_24380);
nand U25994 (N_25994,N_23769,N_23313);
and U25995 (N_25995,N_24683,N_20746);
nor U25996 (N_25996,N_21933,N_22322);
or U25997 (N_25997,N_23359,N_23181);
nand U25998 (N_25998,N_24157,N_20055);
or U25999 (N_25999,N_23825,N_20473);
nor U26000 (N_26000,N_20564,N_22663);
or U26001 (N_26001,N_23883,N_20830);
or U26002 (N_26002,N_23575,N_24022);
nand U26003 (N_26003,N_24460,N_21853);
nor U26004 (N_26004,N_20804,N_24479);
or U26005 (N_26005,N_20955,N_22382);
nand U26006 (N_26006,N_24947,N_20308);
or U26007 (N_26007,N_24203,N_23483);
or U26008 (N_26008,N_24128,N_21571);
nor U26009 (N_26009,N_24487,N_23305);
nor U26010 (N_26010,N_22646,N_21729);
nand U26011 (N_26011,N_24409,N_22648);
and U26012 (N_26012,N_23080,N_20345);
nor U26013 (N_26013,N_22225,N_22180);
or U26014 (N_26014,N_23437,N_23445);
and U26015 (N_26015,N_20490,N_22105);
nand U26016 (N_26016,N_20197,N_20133);
or U26017 (N_26017,N_24901,N_24824);
xor U26018 (N_26018,N_24009,N_23764);
nand U26019 (N_26019,N_24026,N_22744);
and U26020 (N_26020,N_24942,N_21408);
and U26021 (N_26021,N_23845,N_20802);
and U26022 (N_26022,N_21567,N_21622);
and U26023 (N_26023,N_22567,N_20899);
or U26024 (N_26024,N_22987,N_20026);
or U26025 (N_26025,N_20089,N_21663);
and U26026 (N_26026,N_21963,N_23248);
nor U26027 (N_26027,N_21292,N_21391);
nor U26028 (N_26028,N_20290,N_20356);
nor U26029 (N_26029,N_22376,N_24742);
and U26030 (N_26030,N_23950,N_22061);
and U26031 (N_26031,N_22895,N_24981);
and U26032 (N_26032,N_20723,N_21494);
nor U26033 (N_26033,N_20539,N_24499);
nand U26034 (N_26034,N_20083,N_23689);
xor U26035 (N_26035,N_22202,N_22147);
nand U26036 (N_26036,N_20094,N_21166);
and U26037 (N_26037,N_22535,N_20541);
nor U26038 (N_26038,N_23312,N_21186);
and U26039 (N_26039,N_24247,N_21082);
or U26040 (N_26040,N_23167,N_20213);
or U26041 (N_26041,N_24914,N_22722);
nor U26042 (N_26042,N_23635,N_21774);
nor U26043 (N_26043,N_23582,N_24174);
nor U26044 (N_26044,N_20033,N_23404);
or U26045 (N_26045,N_24690,N_22058);
nand U26046 (N_26046,N_21052,N_24045);
nor U26047 (N_26047,N_22727,N_22456);
and U26048 (N_26048,N_24144,N_20909);
nand U26049 (N_26049,N_23014,N_20879);
or U26050 (N_26050,N_23364,N_23317);
nand U26051 (N_26051,N_24163,N_22607);
or U26052 (N_26052,N_24350,N_22950);
or U26053 (N_26053,N_20873,N_24817);
and U26054 (N_26054,N_23493,N_22099);
nand U26055 (N_26055,N_24970,N_21445);
and U26056 (N_26056,N_24038,N_20544);
nand U26057 (N_26057,N_24916,N_23829);
nand U26058 (N_26058,N_23671,N_23958);
nand U26059 (N_26059,N_23795,N_20507);
nand U26060 (N_26060,N_20099,N_23925);
or U26061 (N_26061,N_22605,N_22126);
or U26062 (N_26062,N_22856,N_23978);
or U26063 (N_26063,N_21601,N_22700);
nor U26064 (N_26064,N_22482,N_24125);
nor U26065 (N_26065,N_22439,N_21627);
nor U26066 (N_26066,N_24576,N_22155);
xnor U26067 (N_26067,N_24392,N_24076);
and U26068 (N_26068,N_20186,N_24307);
or U26069 (N_26069,N_24140,N_20747);
nand U26070 (N_26070,N_21010,N_21204);
nor U26071 (N_26071,N_20907,N_20372);
or U26072 (N_26072,N_22447,N_22201);
and U26073 (N_26073,N_21210,N_24616);
nor U26074 (N_26074,N_22026,N_20333);
or U26075 (N_26075,N_24408,N_23132);
or U26076 (N_26076,N_20966,N_23757);
or U26077 (N_26077,N_23629,N_20925);
nor U26078 (N_26078,N_22307,N_20648);
nand U26079 (N_26079,N_24951,N_24031);
or U26080 (N_26080,N_22046,N_22615);
and U26081 (N_26081,N_20835,N_22207);
or U26082 (N_26082,N_20458,N_21226);
and U26083 (N_26083,N_23487,N_24103);
nor U26084 (N_26084,N_23396,N_21433);
nor U26085 (N_26085,N_21035,N_20874);
nand U26086 (N_26086,N_21017,N_22927);
and U26087 (N_26087,N_21998,N_21392);
nor U26088 (N_26088,N_21464,N_21167);
nor U26089 (N_26089,N_23129,N_23222);
or U26090 (N_26090,N_23244,N_21483);
and U26091 (N_26091,N_23722,N_21174);
or U26092 (N_26092,N_22536,N_22492);
or U26093 (N_26093,N_20150,N_21014);
nand U26094 (N_26094,N_21863,N_24196);
nand U26095 (N_26095,N_24204,N_23399);
or U26096 (N_26096,N_20689,N_21388);
nor U26097 (N_26097,N_20640,N_20773);
xor U26098 (N_26098,N_21428,N_23936);
nand U26099 (N_26099,N_22786,N_21536);
nand U26100 (N_26100,N_23343,N_24213);
and U26101 (N_26101,N_21958,N_24591);
nor U26102 (N_26102,N_23403,N_23820);
or U26103 (N_26103,N_21801,N_24980);
and U26104 (N_26104,N_22288,N_24933);
and U26105 (N_26105,N_22594,N_24343);
xnor U26106 (N_26106,N_21446,N_21648);
nor U26107 (N_26107,N_24973,N_21117);
or U26108 (N_26108,N_23875,N_20352);
or U26109 (N_26109,N_21164,N_24909);
nand U26110 (N_26110,N_22690,N_23716);
or U26111 (N_26111,N_24456,N_24173);
or U26112 (N_26112,N_21520,N_21072);
or U26113 (N_26113,N_22982,N_20521);
nand U26114 (N_26114,N_22773,N_22287);
nor U26115 (N_26115,N_20696,N_21402);
nor U26116 (N_26116,N_23384,N_22791);
and U26117 (N_26117,N_24861,N_23147);
nor U26118 (N_26118,N_21882,N_24717);
or U26119 (N_26119,N_21449,N_24870);
nand U26120 (N_26120,N_20793,N_20078);
and U26121 (N_26121,N_20406,N_24693);
nor U26122 (N_26122,N_24131,N_24848);
nand U26123 (N_26123,N_23695,N_24188);
or U26124 (N_26124,N_20837,N_20011);
nand U26125 (N_26125,N_22647,N_22388);
or U26126 (N_26126,N_23191,N_23861);
nor U26127 (N_26127,N_22175,N_22052);
xor U26128 (N_26128,N_20882,N_23850);
and U26129 (N_26129,N_23114,N_22653);
xnor U26130 (N_26130,N_20466,N_22476);
and U26131 (N_26131,N_22946,N_22001);
and U26132 (N_26132,N_21340,N_21115);
and U26133 (N_26133,N_22116,N_24631);
nand U26134 (N_26134,N_21286,N_22552);
nor U26135 (N_26135,N_20672,N_23179);
xnor U26136 (N_26136,N_20653,N_22948);
nor U26137 (N_26137,N_21781,N_23616);
or U26138 (N_26138,N_23650,N_23708);
nand U26139 (N_26139,N_21951,N_22065);
nor U26140 (N_26140,N_24862,N_23569);
and U26141 (N_26141,N_24986,N_20608);
nor U26142 (N_26142,N_21182,N_21341);
nor U26143 (N_26143,N_24928,N_20489);
and U26144 (N_26144,N_24600,N_24358);
or U26145 (N_26145,N_24661,N_20943);
or U26146 (N_26146,N_22440,N_22290);
or U26147 (N_26147,N_24472,N_20642);
nand U26148 (N_26148,N_20895,N_21159);
and U26149 (N_26149,N_23424,N_21196);
or U26150 (N_26150,N_21303,N_23340);
or U26151 (N_26151,N_24051,N_21541);
nor U26152 (N_26152,N_20533,N_20472);
nand U26153 (N_26153,N_21587,N_21896);
and U26154 (N_26154,N_21149,N_20703);
or U26155 (N_26155,N_21140,N_23284);
nor U26156 (N_26156,N_24123,N_23939);
nand U26157 (N_26157,N_24401,N_20836);
or U26158 (N_26158,N_20918,N_22654);
nor U26159 (N_26159,N_20364,N_21841);
xnor U26160 (N_26160,N_21043,N_20761);
and U26161 (N_26161,N_23623,N_20740);
nand U26162 (N_26162,N_21322,N_24154);
or U26163 (N_26163,N_22102,N_24289);
and U26164 (N_26164,N_21110,N_23664);
xor U26165 (N_26165,N_22371,N_24783);
and U26166 (N_26166,N_22822,N_23485);
nand U26167 (N_26167,N_20867,N_23894);
nand U26168 (N_26168,N_21501,N_24365);
or U26169 (N_26169,N_21538,N_24832);
or U26170 (N_26170,N_23154,N_22886);
nand U26171 (N_26171,N_22321,N_22583);
nand U26172 (N_26172,N_23192,N_23681);
or U26173 (N_26173,N_21530,N_23902);
and U26174 (N_26174,N_23238,N_23214);
nand U26175 (N_26175,N_22659,N_23590);
xor U26176 (N_26176,N_24592,N_23849);
nand U26177 (N_26177,N_21252,N_20013);
or U26178 (N_26178,N_23505,N_22134);
nor U26179 (N_26179,N_20795,N_22736);
nand U26180 (N_26180,N_24960,N_20438);
nor U26181 (N_26181,N_22565,N_24917);
nor U26182 (N_26182,N_23229,N_22044);
nor U26183 (N_26183,N_24434,N_22924);
nor U26184 (N_26184,N_22420,N_23842);
nor U26185 (N_26185,N_21573,N_22251);
nor U26186 (N_26186,N_23954,N_23161);
and U26187 (N_26187,N_21759,N_24902);
nand U26188 (N_26188,N_20582,N_20525);
nor U26189 (N_26189,N_21362,N_22563);
nand U26190 (N_26190,N_23808,N_23970);
nand U26191 (N_26191,N_24655,N_23082);
nand U26192 (N_26192,N_24181,N_20445);
or U26193 (N_26193,N_21630,N_20022);
nor U26194 (N_26194,N_21183,N_24266);
or U26195 (N_26195,N_22979,N_21533);
nor U26196 (N_26196,N_20527,N_21973);
nand U26197 (N_26197,N_20420,N_23402);
nand U26198 (N_26198,N_24766,N_21652);
xor U26199 (N_26199,N_24095,N_20824);
nand U26200 (N_26200,N_20282,N_24491);
or U26201 (N_26201,N_21329,N_20524);
and U26202 (N_26202,N_20963,N_23714);
and U26203 (N_26203,N_20104,N_24876);
or U26204 (N_26204,N_20130,N_22092);
nand U26205 (N_26205,N_21892,N_21124);
or U26206 (N_26206,N_21045,N_23877);
or U26207 (N_26207,N_20808,N_21936);
or U26208 (N_26208,N_21704,N_24035);
nand U26209 (N_26209,N_20393,N_24514);
nor U26210 (N_26210,N_23696,N_21462);
or U26211 (N_26211,N_22333,N_20622);
nand U26212 (N_26212,N_21297,N_23194);
or U26213 (N_26213,N_23433,N_20649);
nor U26214 (N_26214,N_20354,N_22590);
nor U26215 (N_26215,N_20960,N_21529);
nand U26216 (N_26216,N_21409,N_21127);
nand U26217 (N_26217,N_23120,N_24331);
xor U26218 (N_26218,N_24839,N_20005);
nor U26219 (N_26219,N_20122,N_24073);
or U26220 (N_26220,N_22248,N_21410);
nor U26221 (N_26221,N_24971,N_21616);
nand U26222 (N_26222,N_24176,N_22415);
or U26223 (N_26223,N_24793,N_22087);
xnor U26224 (N_26224,N_21715,N_23348);
nand U26225 (N_26225,N_24347,N_24264);
xnor U26226 (N_26226,N_22238,N_21347);
or U26227 (N_26227,N_21122,N_24394);
nand U26228 (N_26228,N_20897,N_24357);
nor U26229 (N_26229,N_21856,N_22254);
nor U26230 (N_26230,N_23691,N_23593);
or U26231 (N_26231,N_23310,N_20208);
xnor U26232 (N_26232,N_21374,N_20261);
xnor U26233 (N_26233,N_23677,N_20577);
and U26234 (N_26234,N_23802,N_21518);
or U26235 (N_26235,N_21551,N_21128);
or U26236 (N_26236,N_20559,N_24327);
xor U26237 (N_26237,N_22558,N_22083);
and U26238 (N_26238,N_22925,N_23175);
nor U26239 (N_26239,N_23421,N_21396);
nor U26240 (N_26240,N_20921,N_23712);
nor U26241 (N_26241,N_22037,N_23118);
and U26242 (N_26242,N_23264,N_21602);
nor U26243 (N_26243,N_24869,N_23489);
nor U26244 (N_26244,N_23675,N_21561);
nand U26245 (N_26245,N_23551,N_21859);
and U26246 (N_26246,N_21091,N_21684);
xnor U26247 (N_26247,N_23183,N_21633);
nand U26248 (N_26248,N_23250,N_22223);
or U26249 (N_26249,N_22270,N_23273);
nor U26250 (N_26250,N_21844,N_23050);
nor U26251 (N_26251,N_24248,N_21916);
nor U26252 (N_26252,N_21345,N_23062);
and U26253 (N_26253,N_20858,N_20498);
or U26254 (N_26254,N_21102,N_24222);
or U26255 (N_26255,N_21545,N_23432);
or U26256 (N_26256,N_23502,N_20692);
nor U26257 (N_26257,N_20556,N_20655);
or U26258 (N_26258,N_22444,N_24894);
or U26259 (N_26259,N_24540,N_22624);
or U26260 (N_26260,N_22298,N_21147);
or U26261 (N_26261,N_20626,N_24552);
or U26262 (N_26262,N_23344,N_20815);
nor U26263 (N_26263,N_23742,N_24509);
and U26264 (N_26264,N_20029,N_22652);
nor U26265 (N_26265,N_20001,N_23297);
nor U26266 (N_26266,N_21694,N_21077);
nor U26267 (N_26267,N_20615,N_22575);
nand U26268 (N_26268,N_24057,N_20550);
or U26269 (N_26269,N_22743,N_23979);
nor U26270 (N_26270,N_24996,N_20427);
nor U26271 (N_26271,N_21206,N_23760);
and U26272 (N_26272,N_24927,N_21621);
nand U26273 (N_26273,N_22418,N_22125);
nor U26274 (N_26274,N_22179,N_21797);
or U26275 (N_26275,N_21033,N_22696);
nor U26276 (N_26276,N_24423,N_20917);
or U26277 (N_26277,N_24826,N_24613);
or U26278 (N_26278,N_20624,N_23744);
nand U26279 (N_26279,N_24666,N_20667);
nand U26280 (N_26280,N_23926,N_21003);
or U26281 (N_26281,N_21485,N_23824);
xnor U26282 (N_26282,N_22988,N_20975);
and U26283 (N_26283,N_22391,N_21306);
or U26284 (N_26284,N_22666,N_21089);
or U26285 (N_26285,N_22401,N_24698);
and U26286 (N_26286,N_20168,N_24261);
or U26287 (N_26287,N_23358,N_21505);
and U26288 (N_26288,N_20791,N_22340);
nor U26289 (N_26289,N_23963,N_22067);
or U26290 (N_26290,N_24705,N_22352);
xor U26291 (N_26291,N_23931,N_24895);
or U26292 (N_26292,N_23419,N_24345);
or U26293 (N_26293,N_23591,N_22466);
nor U26294 (N_26294,N_23255,N_23638);
xnor U26295 (N_26295,N_23239,N_23998);
and U26296 (N_26296,N_23127,N_21559);
and U26297 (N_26297,N_22477,N_22537);
or U26298 (N_26298,N_22240,N_21332);
nor U26299 (N_26299,N_21369,N_22433);
and U26300 (N_26300,N_21215,N_23580);
nor U26301 (N_26301,N_24868,N_24539);
xnor U26302 (N_26302,N_22164,N_20048);
or U26303 (N_26303,N_21075,N_21099);
nor U26304 (N_26304,N_24089,N_24411);
nand U26305 (N_26305,N_21523,N_22316);
nand U26306 (N_26306,N_24911,N_23822);
and U26307 (N_26307,N_23519,N_24421);
or U26308 (N_26308,N_22330,N_22998);
nand U26309 (N_26309,N_24995,N_24827);
nand U26310 (N_26310,N_23447,N_24603);
nand U26311 (N_26311,N_23897,N_24476);
and U26312 (N_26312,N_22910,N_21093);
nand U26313 (N_26313,N_20144,N_24178);
and U26314 (N_26314,N_24903,N_24627);
nand U26315 (N_26315,N_23823,N_20494);
nand U26316 (N_26316,N_23938,N_20419);
nor U26317 (N_26317,N_22629,N_22943);
nand U26318 (N_26318,N_22529,N_20255);
and U26319 (N_26319,N_21946,N_21554);
nor U26320 (N_26320,N_20134,N_23537);
or U26321 (N_26321,N_24280,N_20170);
or U26322 (N_26322,N_22501,N_20855);
nor U26323 (N_26323,N_21811,N_20998);
and U26324 (N_26324,N_20395,N_20437);
nand U26325 (N_26325,N_23139,N_23236);
xor U26326 (N_26326,N_24198,N_20821);
or U26327 (N_26327,N_21109,N_23973);
and U26328 (N_26328,N_21885,N_22724);
and U26329 (N_26329,N_24834,N_22821);
nand U26330 (N_26330,N_21697,N_20098);
nand U26331 (N_26331,N_24461,N_20312);
or U26332 (N_26332,N_22610,N_21994);
nand U26333 (N_26333,N_22273,N_21376);
or U26334 (N_26334,N_20042,N_21907);
and U26335 (N_26335,N_23856,N_24610);
nand U26336 (N_26336,N_22372,N_22430);
or U26337 (N_26337,N_20047,N_22365);
or U26338 (N_26338,N_20579,N_21309);
or U26339 (N_26339,N_23866,N_21924);
or U26340 (N_26340,N_21719,N_24961);
nor U26341 (N_26341,N_22613,N_22918);
and U26342 (N_26342,N_21394,N_22053);
or U26343 (N_26343,N_22094,N_22730);
nand U26344 (N_26344,N_20286,N_20905);
and U26345 (N_26345,N_20319,N_20140);
or U26346 (N_26346,N_20327,N_22030);
and U26347 (N_26347,N_21325,N_24811);
nor U26348 (N_26348,N_24700,N_21976);
nand U26349 (N_26349,N_24227,N_24702);
nand U26350 (N_26350,N_24287,N_22093);
and U26351 (N_26351,N_22628,N_22387);
nor U26352 (N_26352,N_24905,N_20670);
or U26353 (N_26353,N_22464,N_22705);
xor U26354 (N_26354,N_22562,N_21259);
or U26355 (N_26355,N_21766,N_23394);
and U26356 (N_26356,N_22709,N_20329);
and U26357 (N_26357,N_20976,N_20107);
nor U26358 (N_26358,N_24329,N_21333);
nor U26359 (N_26359,N_24425,N_20377);
or U26360 (N_26360,N_24644,N_21673);
and U26361 (N_26361,N_21044,N_23745);
nand U26362 (N_26362,N_22595,N_24404);
xor U26363 (N_26363,N_21700,N_22357);
and U26364 (N_26364,N_20415,N_20617);
or U26365 (N_26365,N_23482,N_23217);
xnor U26366 (N_26366,N_23168,N_20234);
and U26367 (N_26367,N_21725,N_20927);
or U26368 (N_26368,N_20487,N_22684);
and U26369 (N_26369,N_23879,N_20257);
and U26370 (N_26370,N_20931,N_22215);
nand U26371 (N_26371,N_24731,N_23177);
nand U26372 (N_26372,N_21217,N_22165);
nor U26373 (N_26373,N_21097,N_21512);
and U26374 (N_26374,N_22448,N_24982);
xor U26375 (N_26375,N_23032,N_23232);
nand U26376 (N_26376,N_20827,N_20946);
and U26377 (N_26377,N_22728,N_20068);
nor U26378 (N_26378,N_20071,N_23128);
nor U26379 (N_26379,N_20113,N_24957);
xnor U26380 (N_26380,N_23730,N_24630);
and U26381 (N_26381,N_24638,N_20232);
nor U26382 (N_26382,N_22834,N_23839);
xor U26383 (N_26383,N_23900,N_20218);
and U26384 (N_26384,N_24295,N_21890);
or U26385 (N_26385,N_21937,N_21190);
nor U26386 (N_26386,N_23333,N_20196);
xor U26387 (N_26387,N_20876,N_21317);
and U26388 (N_26388,N_22265,N_24313);
or U26389 (N_26389,N_24452,N_21662);
and U26390 (N_26390,N_21613,N_22703);
xor U26391 (N_26391,N_20247,N_22064);
xnor U26392 (N_26392,N_24782,N_21002);
and U26393 (N_26393,N_21443,N_23422);
xnor U26394 (N_26394,N_21187,N_22581);
nor U26395 (N_26395,N_24362,N_24780);
xor U26396 (N_26396,N_24326,N_22234);
nand U26397 (N_26397,N_20387,N_20391);
and U26398 (N_26398,N_24689,N_24730);
nor U26399 (N_26399,N_20017,N_23994);
or U26400 (N_26400,N_23554,N_21488);
and U26401 (N_26401,N_20694,N_24855);
nand U26402 (N_26402,N_23793,N_20138);
nand U26403 (N_26403,N_24288,N_23292);
nand U26404 (N_26404,N_23794,N_24686);
nand U26405 (N_26405,N_21365,N_22651);
nor U26406 (N_26406,N_22081,N_24694);
nand U26407 (N_26407,N_22691,N_21008);
or U26408 (N_26408,N_23885,N_22331);
nor U26409 (N_26409,N_24755,N_23752);
nor U26410 (N_26410,N_22517,N_21646);
and U26411 (N_26411,N_21380,N_23514);
nand U26412 (N_26412,N_21058,N_24441);
nor U26413 (N_26413,N_21560,N_24210);
nand U26414 (N_26414,N_22143,N_21437);
nand U26415 (N_26415,N_20749,N_20758);
and U26416 (N_26416,N_24541,N_21157);
nor U26417 (N_26417,N_24023,N_21255);
nor U26418 (N_26418,N_23037,N_24525);
xor U26419 (N_26419,N_22572,N_24537);
nand U26420 (N_26420,N_24745,N_20191);
or U26421 (N_26421,N_20493,N_22313);
xor U26422 (N_26422,N_23622,N_20853);
nor U26423 (N_26423,N_24439,N_22502);
nand U26424 (N_26424,N_23604,N_24283);
nor U26425 (N_26425,N_20452,N_20520);
or U26426 (N_26426,N_23113,N_21742);
nor U26427 (N_26427,N_23930,N_24033);
or U26428 (N_26428,N_23761,N_21830);
nand U26429 (N_26429,N_22969,N_22332);
nand U26430 (N_26430,N_23251,N_23164);
and U26431 (N_26431,N_24628,N_21691);
nand U26432 (N_26432,N_24385,N_24544);
xnor U26433 (N_26433,N_21041,N_23711);
nand U26434 (N_26434,N_24649,N_22451);
nand U26435 (N_26435,N_22386,N_22698);
and U26436 (N_26436,N_21912,N_21185);
nor U26437 (N_26437,N_24756,N_20448);
nand U26438 (N_26438,N_21162,N_24075);
nand U26439 (N_26439,N_21417,N_21671);
and U26440 (N_26440,N_21005,N_20647);
and U26441 (N_26441,N_23200,N_23667);
xor U26442 (N_26442,N_20073,N_20654);
and U26443 (N_26443,N_24685,N_24594);
and U26444 (N_26444,N_23775,N_23140);
nand U26445 (N_26445,N_20141,N_24171);
xor U26446 (N_26446,N_21644,N_20797);
nor U26447 (N_26447,N_21055,N_24302);
nor U26448 (N_26448,N_24137,N_21578);
or U26449 (N_26449,N_23687,N_20461);
or U26450 (N_26450,N_22228,N_21004);
and U26451 (N_26451,N_23735,N_20575);
or U26452 (N_26452,N_21641,N_22427);
or U26453 (N_26453,N_20732,N_24486);
nor U26454 (N_26454,N_24647,N_21125);
nand U26455 (N_26455,N_21510,N_22981);
nor U26456 (N_26456,N_20997,N_24622);
xor U26457 (N_26457,N_21490,N_23583);
and U26458 (N_26458,N_20203,N_23443);
or U26459 (N_26459,N_24024,N_23603);
xor U26460 (N_26460,N_24177,N_22560);
nand U26461 (N_26461,N_20563,N_23576);
nor U26462 (N_26462,N_21680,N_24489);
nor U26463 (N_26463,N_21040,N_24786);
and U26464 (N_26464,N_22748,N_20900);
and U26465 (N_26465,N_24898,N_24081);
xor U26466 (N_26466,N_21452,N_20457);
xnor U26467 (N_26467,N_22521,N_21416);
or U26468 (N_26468,N_24027,N_22806);
xnor U26469 (N_26469,N_22674,N_21852);
nand U26470 (N_26470,N_21870,N_22887);
and U26471 (N_26471,N_21191,N_22573);
and U26472 (N_26472,N_24915,N_22342);
or U26473 (N_26473,N_20669,N_24999);
nor U26474 (N_26474,N_20613,N_20854);
or U26475 (N_26475,N_22803,N_22000);
nand U26476 (N_26476,N_22272,N_20991);
xor U26477 (N_26477,N_23076,N_23283);
nand U26478 (N_26478,N_24578,N_20018);
xor U26479 (N_26479,N_24228,N_20936);
xnor U26480 (N_26480,N_20060,N_24812);
nor U26481 (N_26481,N_22879,N_22148);
xnor U26482 (N_26482,N_21087,N_23943);
nor U26483 (N_26483,N_20601,N_21921);
or U26484 (N_26484,N_24419,N_21502);
or U26485 (N_26485,N_21876,N_22547);
or U26486 (N_26486,N_21279,N_23334);
or U26487 (N_26487,N_24551,N_21546);
or U26488 (N_26488,N_20528,N_20620);
or U26489 (N_26489,N_23997,N_22513);
nor U26490 (N_26490,N_20084,N_22089);
nor U26491 (N_26491,N_23746,N_20768);
nor U26492 (N_26492,N_24226,N_21059);
and U26493 (N_26493,N_20147,N_23401);
and U26494 (N_26494,N_21113,N_20066);
and U26495 (N_26495,N_22719,N_24209);
nand U26496 (N_26496,N_21355,N_21143);
nor U26497 (N_26497,N_22216,N_20258);
nand U26498 (N_26498,N_23896,N_21891);
and U26499 (N_26499,N_23314,N_22075);
nand U26500 (N_26500,N_20374,N_22219);
or U26501 (N_26501,N_22112,N_22218);
xnor U26502 (N_26502,N_23207,N_23776);
and U26503 (N_26503,N_22940,N_23162);
nor U26504 (N_26504,N_20623,N_21061);
or U26505 (N_26505,N_20264,N_22374);
or U26506 (N_26506,N_22833,N_22130);
nor U26507 (N_26507,N_23375,N_23965);
or U26508 (N_26508,N_20417,N_22526);
xor U26509 (N_26509,N_21977,N_21798);
xnor U26510 (N_26510,N_21019,N_21953);
xor U26511 (N_26511,N_20811,N_24881);
nor U26512 (N_26512,N_24825,N_20846);
or U26513 (N_26513,N_24598,N_20477);
nand U26514 (N_26514,N_24692,N_23448);
nor U26515 (N_26515,N_22267,N_20987);
nand U26516 (N_26516,N_20192,N_21899);
and U26517 (N_26517,N_21441,N_20938);
nor U26518 (N_26518,N_24612,N_20565);
and U26519 (N_26519,N_24639,N_23806);
nand U26520 (N_26520,N_22546,N_22025);
and U26521 (N_26521,N_22222,N_22077);
and U26522 (N_26522,N_23332,N_20322);
nand U26523 (N_26523,N_24108,N_21039);
nor U26524 (N_26524,N_20146,N_22678);
nor U26525 (N_26525,N_21837,N_24978);
nand U26526 (N_26526,N_24815,N_22704);
nor U26527 (N_26527,N_22738,N_22123);
or U26528 (N_26528,N_21693,N_21618);
xor U26529 (N_26529,N_21903,N_22892);
nand U26530 (N_26530,N_20660,N_20139);
or U26531 (N_26531,N_23627,N_22571);
nand U26532 (N_26532,N_23670,N_21274);
xor U26533 (N_26533,N_22235,N_24636);
nand U26534 (N_26534,N_21893,N_22209);
or U26535 (N_26535,N_21054,N_23698);
and U26536 (N_26536,N_23224,N_24680);
and U26537 (N_26537,N_24699,N_21478);
or U26538 (N_26538,N_21918,N_20362);
or U26539 (N_26539,N_22739,N_23440);
nand U26540 (N_26540,N_22930,N_21165);
or U26541 (N_26541,N_21875,N_24929);
and U26542 (N_26542,N_21940,N_21034);
and U26543 (N_26543,N_22007,N_23503);
nand U26544 (N_26544,N_23567,N_21312);
or U26545 (N_26545,N_21468,N_23557);
and U26546 (N_26546,N_23826,N_21112);
nand U26547 (N_26547,N_24615,N_20454);
and U26548 (N_26548,N_21472,N_22429);
or U26549 (N_26549,N_22712,N_23193);
nand U26550 (N_26550,N_24512,N_21911);
and U26551 (N_26551,N_24813,N_23595);
nand U26552 (N_26552,N_20201,N_21605);
and U26553 (N_26553,N_20023,N_23442);
nand U26554 (N_26554,N_22878,N_22478);
nand U26555 (N_26555,N_21435,N_24553);
and U26556 (N_26556,N_23055,N_21986);
or U26557 (N_26557,N_20295,N_24374);
nand U26558 (N_26558,N_20543,N_21423);
and U26559 (N_26559,N_22935,N_21711);
and U26560 (N_26560,N_24484,N_22578);
nand U26561 (N_26561,N_24121,N_23901);
nor U26562 (N_26562,N_20888,N_22082);
and U26563 (N_26563,N_20394,N_20589);
nand U26564 (N_26564,N_22812,N_20240);
and U26565 (N_26565,N_22710,N_21222);
and U26566 (N_26566,N_22689,N_23974);
xor U26567 (N_26567,N_21318,N_21219);
nor U26568 (N_26568,N_23188,N_23075);
or U26569 (N_26569,N_22764,N_23790);
and U26570 (N_26570,N_21432,N_20004);
or U26571 (N_26571,N_22830,N_21775);
nor U26572 (N_26572,N_22442,N_24507);
or U26573 (N_26573,N_21304,N_22504);
nand U26574 (N_26574,N_23002,N_20671);
nor U26575 (N_26575,N_21782,N_24205);
nor U26576 (N_26576,N_23684,N_20537);
or U26577 (N_26577,N_23323,N_22559);
nor U26578 (N_26578,N_20992,N_24938);
nor U26579 (N_26579,N_20686,N_22899);
and U26580 (N_26580,N_22338,N_24584);
nand U26581 (N_26581,N_23427,N_24115);
xnor U26582 (N_26582,N_20509,N_21479);
or U26583 (N_26583,N_24375,N_21352);
nor U26584 (N_26584,N_24570,N_24925);
xor U26585 (N_26585,N_24941,N_21038);
nand U26586 (N_26586,N_24284,N_23734);
or U26587 (N_26587,N_24836,N_23592);
xor U26588 (N_26588,N_24065,N_22912);
nand U26589 (N_26589,N_22986,N_20857);
nor U26590 (N_26590,N_21107,N_22434);
and U26591 (N_26591,N_24450,N_23838);
and U26592 (N_26592,N_22702,N_21862);
nor U26593 (N_26593,N_21995,N_20418);
nand U26594 (N_26594,N_24136,N_20283);
nand U26595 (N_26595,N_21031,N_23423);
and U26596 (N_26596,N_21313,N_24166);
or U26597 (N_26597,N_24794,N_22602);
or U26598 (N_26598,N_21889,N_20762);
nor U26599 (N_26599,N_20402,N_21683);
or U26600 (N_26600,N_24469,N_22539);
and U26601 (N_26601,N_21368,N_23555);
nand U26602 (N_26602,N_20057,N_23009);
or U26603 (N_26603,N_22658,N_20455);
or U26604 (N_26604,N_23385,N_22283);
and U26605 (N_26605,N_20856,N_22107);
and U26606 (N_26606,N_21692,N_24442);
and U26607 (N_26607,N_24058,N_23142);
and U26608 (N_26608,N_23084,N_23470);
nand U26609 (N_26609,N_22318,N_22857);
or U26610 (N_26610,N_20990,N_21268);
and U26611 (N_26611,N_20788,N_22937);
or U26612 (N_26612,N_20988,N_22888);
and U26613 (N_26613,N_20661,N_21069);
nor U26614 (N_26614,N_24814,N_21338);
nand U26615 (N_26615,N_21682,N_24754);
nor U26616 (N_26616,N_20382,N_23846);
and U26617 (N_26617,N_20336,N_22548);
and U26618 (N_26618,N_21917,N_22101);
and U26619 (N_26619,N_20271,N_22787);
or U26620 (N_26620,N_24498,N_24844);
or U26621 (N_26621,N_20357,N_22186);
or U26622 (N_26622,N_23038,N_21779);
and U26623 (N_26623,N_24900,N_23153);
or U26624 (N_26624,N_22669,N_21677);
xnor U26625 (N_26625,N_20850,N_21636);
or U26626 (N_26626,N_23321,N_24466);
xnor U26627 (N_26627,N_21763,N_20092);
and U26628 (N_26628,N_21588,N_22299);
xnor U26629 (N_26629,N_22356,N_21401);
xnor U26630 (N_26630,N_23645,N_22028);
or U26631 (N_26631,N_21053,N_24072);
or U26632 (N_26632,N_22977,N_22027);
or U26633 (N_26633,N_23510,N_23659);
xor U26634 (N_26634,N_22863,N_21326);
nor U26635 (N_26635,N_22538,N_24025);
or U26636 (N_26636,N_24318,N_20429);
and U26637 (N_26637,N_22211,N_22233);
nor U26638 (N_26638,N_24272,N_20284);
or U26639 (N_26639,N_21271,N_22699);
or U26640 (N_26640,N_22680,N_20301);
xnor U26641 (N_26641,N_21090,N_23247);
and U26642 (N_26642,N_23946,N_20576);
and U26643 (N_26643,N_22132,N_20428);
xnor U26644 (N_26644,N_21205,N_24534);
or U26645 (N_26645,N_20044,N_20076);
or U26646 (N_26646,N_22996,N_23594);
and U26647 (N_26647,N_22319,N_20342);
nor U26648 (N_26648,N_24015,N_22994);
nand U26649 (N_26649,N_20637,N_23741);
nor U26650 (N_26650,N_21702,N_22245);
and U26651 (N_26651,N_23858,N_23001);
nor U26652 (N_26652,N_20059,N_23178);
nand U26653 (N_26653,N_23287,N_21527);
nor U26654 (N_26654,N_24482,N_23199);
and U26655 (N_26655,N_23013,N_21528);
nor U26656 (N_26656,N_21132,N_24323);
nor U26657 (N_26657,N_22606,N_22157);
or U26658 (N_26658,N_21175,N_20435);
nor U26659 (N_26659,N_24715,N_24651);
nand U26660 (N_26660,N_24602,N_24729);
and U26661 (N_26661,N_24122,N_20431);
nor U26662 (N_26662,N_20031,N_22280);
nand U26663 (N_26663,N_20515,N_24389);
nand U26664 (N_26664,N_20300,N_22890);
or U26665 (N_26665,N_20119,N_24520);
nor U26666 (N_26666,N_24402,N_21599);
and U26667 (N_26667,N_24218,N_24695);
and U26668 (N_26668,N_21810,N_20090);
xnor U26669 (N_26669,N_21879,N_20910);
xor U26670 (N_26670,N_24532,N_21261);
nor U26671 (N_26671,N_24273,N_22076);
and U26672 (N_26672,N_22465,N_21789);
and U26673 (N_26673,N_24471,N_21305);
or U26674 (N_26674,N_21119,N_20845);
nand U26675 (N_26675,N_22862,N_20517);
and U26676 (N_26676,N_24064,N_21549);
or U26677 (N_26677,N_24255,N_21184);
and U26678 (N_26678,N_22031,N_20470);
nand U26679 (N_26679,N_22315,N_21614);
nor U26680 (N_26680,N_20176,N_24167);
nand U26681 (N_26681,N_20405,N_24865);
or U26682 (N_26682,N_22827,N_21741);
xnor U26683 (N_26683,N_22945,N_22953);
nor U26684 (N_26684,N_21595,N_23413);
or U26685 (N_26685,N_23665,N_22339);
and U26686 (N_26686,N_21640,N_23574);
nor U26687 (N_26687,N_21550,N_20156);
nand U26688 (N_26688,N_21765,N_24159);
xor U26689 (N_26689,N_24440,N_23288);
or U26690 (N_26690,N_23913,N_20914);
nor U26691 (N_26691,N_23083,N_21913);
or U26692 (N_26692,N_20269,N_24728);
and U26693 (N_26693,N_24643,N_22011);
nand U26694 (N_26694,N_23170,N_22523);
and U26695 (N_26695,N_20996,N_24299);
or U26696 (N_26696,N_23040,N_24642);
or U26697 (N_26697,N_23353,N_22048);
and U26698 (N_26698,N_22852,N_20812);
or U26699 (N_26699,N_24356,N_21150);
or U26700 (N_26700,N_23673,N_23682);
xnor U26701 (N_26701,N_24193,N_22110);
nor U26702 (N_26702,N_23466,N_22828);
or U26703 (N_26703,N_23474,N_24899);
nor U26704 (N_26704,N_20153,N_21557);
and U26705 (N_26705,N_22115,N_21748);
or U26706 (N_26706,N_23410,N_24657);
nand U26707 (N_26707,N_23137,N_24091);
nor U26708 (N_26708,N_21198,N_21001);
nor U26709 (N_26709,N_21796,N_24483);
nand U26710 (N_26710,N_21915,N_22837);
nand U26711 (N_26711,N_21827,N_24840);
nand U26712 (N_26712,N_21020,N_22765);
nor U26713 (N_26713,N_22455,N_20383);
and U26714 (N_26714,N_22033,N_22941);
xor U26715 (N_26715,N_24100,N_24113);
and U26716 (N_26716,N_20058,N_23552);
and U26717 (N_26717,N_24306,N_22227);
xnor U26718 (N_26718,N_23740,N_22369);
nand U26719 (N_26719,N_24006,N_23293);
nor U26720 (N_26720,N_21583,N_21212);
and U26721 (N_26721,N_20616,N_23299);
xor U26722 (N_26722,N_24114,N_24850);
or U26723 (N_26723,N_23774,N_22142);
and U26724 (N_26724,N_24769,N_22819);
or U26725 (N_26725,N_20964,N_20024);
nand U26726 (N_26726,N_23912,N_22159);
and U26727 (N_26727,N_22144,N_22625);
or U26728 (N_26728,N_22262,N_21266);
nor U26729 (N_26729,N_22015,N_21176);
or U26730 (N_26730,N_21063,N_20949);
xnor U26731 (N_26731,N_21838,N_23851);
or U26732 (N_26732,N_22708,N_22274);
xnor U26733 (N_26733,N_22990,N_24187);
and U26734 (N_26734,N_23119,N_24559);
or U26735 (N_26735,N_23556,N_21632);
nor U26736 (N_26736,N_24092,N_22059);
and U26737 (N_26737,N_20935,N_23228);
and U26738 (N_26738,N_20325,N_21021);
nor U26739 (N_26739,N_23891,N_22096);
nand U26740 (N_26740,N_22640,N_21955);
nand U26741 (N_26741,N_21506,N_22874);
or U26742 (N_26742,N_23581,N_20318);
nand U26743 (N_26743,N_20210,N_20265);
or U26744 (N_26744,N_20204,N_21724);
and U26745 (N_26745,N_24132,N_20756);
nand U26746 (N_26746,N_23496,N_21750);
xor U26747 (N_26747,N_22193,N_21027);
or U26748 (N_26748,N_21385,N_22916);
nand U26749 (N_26749,N_22457,N_22350);
xnor U26750 (N_26750,N_24875,N_23163);
or U26751 (N_26751,N_20397,N_21828);
nor U26752 (N_26752,N_21739,N_21744);
and U26753 (N_26753,N_21981,N_20496);
and U26754 (N_26754,N_20476,N_24050);
or U26755 (N_26755,N_22701,N_20175);
nor U26756 (N_26756,N_24744,N_24872);
nand U26757 (N_26757,N_23315,N_22450);
nand U26758 (N_26758,N_24704,N_21894);
nor U26759 (N_26759,N_24480,N_21757);
nand U26760 (N_26760,N_23852,N_20291);
nor U26761 (N_26761,N_21300,N_22003);
nor U26762 (N_26762,N_20349,N_23234);
and U26763 (N_26763,N_24147,N_22181);
or U26764 (N_26764,N_20572,N_21516);
nand U26765 (N_26765,N_24301,N_21029);
nand U26766 (N_26766,N_20715,N_20982);
or U26767 (N_26767,N_23786,N_21793);
nand U26768 (N_26768,N_21509,N_21382);
or U26769 (N_26769,N_21932,N_21854);
or U26770 (N_26770,N_20159,N_21647);
nand U26771 (N_26771,N_23562,N_24393);
nor U26772 (N_26772,N_21371,N_21727);
nor U26773 (N_26773,N_24653,N_24873);
nand U26774 (N_26774,N_20690,N_24806);
and U26775 (N_26775,N_20324,N_24424);
and U26776 (N_26776,N_20765,N_24946);
or U26777 (N_26777,N_21470,N_21945);
xor U26778 (N_26778,N_22258,N_21753);
nor U26779 (N_26779,N_24935,N_20753);
nand U26780 (N_26780,N_22721,N_23045);
or U26781 (N_26781,N_22993,N_23942);
nand U26782 (N_26782,N_23325,N_24554);
xor U26783 (N_26783,N_23935,N_23654);
or U26784 (N_26784,N_24500,N_23771);
and U26785 (N_26785,N_20652,N_24068);
nor U26786 (N_26786,N_20302,N_24391);
nor U26787 (N_26787,N_21476,N_24672);
or U26788 (N_26788,N_21603,N_21904);
or U26789 (N_26789,N_21251,N_22499);
and U26790 (N_26790,N_23290,N_24854);
nor U26791 (N_26791,N_21897,N_22713);
nand U26792 (N_26792,N_20278,N_23700);
nor U26793 (N_26793,N_22588,N_24286);
and U26794 (N_26794,N_23490,N_21302);
nor U26795 (N_26795,N_23454,N_23187);
nand U26796 (N_26796,N_23729,N_20211);
nand U26797 (N_26797,N_22023,N_21267);
and U26798 (N_26798,N_20733,N_21189);
nor U26799 (N_26799,N_21769,N_21768);
and U26800 (N_26800,N_20906,N_21992);
or U26801 (N_26801,N_23221,N_20679);
and U26802 (N_26802,N_23029,N_22976);
or U26803 (N_26803,N_24707,N_23972);
and U26804 (N_26804,N_22042,N_23779);
and U26805 (N_26805,N_22213,N_20779);
nor U26806 (N_26806,N_22758,N_22286);
or U26807 (N_26807,N_24721,N_22692);
and U26808 (N_26808,N_21568,N_22617);
and U26809 (N_26809,N_23857,N_22471);
or U26810 (N_26810,N_21030,N_22470);
and U26811 (N_26811,N_20040,N_20599);
nand U26812 (N_26812,N_23788,N_21869);
or U26813 (N_26813,N_20872,N_21489);
nand U26814 (N_26814,N_21253,N_20711);
nor U26815 (N_26815,N_23725,N_22750);
xnor U26816 (N_26816,N_22557,N_23680);
or U26817 (N_26817,N_24665,N_21057);
nor U26818 (N_26818,N_20124,N_22292);
or U26819 (N_26819,N_23876,N_22749);
nand U26820 (N_26820,N_24200,N_24060);
nor U26821 (N_26821,N_22458,N_22832);
or U26822 (N_26822,N_24417,N_21728);
nor U26823 (N_26823,N_22483,N_24723);
nand U26824 (N_26824,N_23898,N_21542);
or U26825 (N_26825,N_22859,N_22846);
nor U26826 (N_26826,N_22047,N_23703);
nor U26827 (N_26827,N_24197,N_20504);
or U26828 (N_26828,N_24523,N_20782);
and U26829 (N_26829,N_21868,N_22694);
nor U26830 (N_26830,N_22776,N_24590);
or U26831 (N_26831,N_24158,N_22667);
and U26832 (N_26832,N_21806,N_22176);
nor U26833 (N_26833,N_21687,N_23439);
nor U26834 (N_26834,N_24145,N_24360);
or U26835 (N_26835,N_22995,N_23717);
or U26836 (N_26836,N_22161,N_21943);
or U26837 (N_26837,N_24597,N_20396);
and U26838 (N_26838,N_24119,N_24926);
nand U26839 (N_26839,N_21866,N_24681);
and U26840 (N_26840,N_20870,N_22078);
and U26841 (N_26841,N_20451,N_22540);
or U26842 (N_26842,N_21886,N_22876);
and U26843 (N_26843,N_23906,N_24733);
nand U26844 (N_26844,N_21079,N_23197);
and U26845 (N_26845,N_20584,N_22718);
or U26846 (N_26846,N_22297,N_20984);
and U26847 (N_26847,N_24508,N_23756);
and U26848 (N_26848,N_23031,N_22584);
nor U26849 (N_26849,N_20861,N_20944);
xor U26850 (N_26850,N_22136,N_22323);
nor U26851 (N_26851,N_24243,N_22842);
xnor U26852 (N_26852,N_24310,N_22246);
or U26853 (N_26853,N_20350,N_20433);
nor U26854 (N_26854,N_23318,N_21042);
xnor U26855 (N_26855,N_22214,N_23235);
nand U26856 (N_26856,N_22643,N_21714);
and U26857 (N_26857,N_20411,N_20120);
nor U26858 (N_26858,N_21650,N_23471);
nor U26859 (N_26859,N_22915,N_22963);
nor U26860 (N_26860,N_21060,N_23112);
xnor U26861 (N_26861,N_24339,N_20829);
or U26862 (N_26862,N_24459,N_24660);
nor U26863 (N_26863,N_23303,N_20320);
nand U26864 (N_26864,N_22799,N_21635);
xnor U26865 (N_26865,N_24697,N_20592);
or U26866 (N_26866,N_20683,N_21469);
and U26867 (N_26867,N_23058,N_21327);
or U26868 (N_26868,N_21170,N_21758);
and U26869 (N_26869,N_24148,N_22358);
or U26870 (N_26870,N_20602,N_21717);
or U26871 (N_26871,N_21316,N_24090);
or U26872 (N_26872,N_22893,N_23328);
nor U26873 (N_26873,N_23450,N_24727);
and U26874 (N_26874,N_22170,N_22829);
or U26875 (N_26875,N_21048,N_24843);
nor U26876 (N_26876,N_23690,N_24607);
xnor U26877 (N_26877,N_24558,N_23910);
or U26878 (N_26878,N_24185,N_24052);
and U26879 (N_26879,N_23274,N_20953);
nand U26880 (N_26880,N_23174,N_20887);
nand U26881 (N_26881,N_24667,N_24505);
nand U26882 (N_26882,N_23392,N_22438);
or U26883 (N_26883,N_22614,N_23326);
or U26884 (N_26884,N_20190,N_20263);
or U26885 (N_26885,N_22693,N_22960);
xor U26886 (N_26886,N_22626,N_22809);
or U26887 (N_26887,N_22965,N_23959);
nor U26888 (N_26888,N_20049,N_21022);
and U26889 (N_26889,N_22933,N_23541);
nand U26890 (N_26890,N_20358,N_23907);
and U26891 (N_26891,N_21466,N_24028);
nand U26892 (N_26892,N_22733,N_22469);
nand U26893 (N_26893,N_21839,N_21984);
and U26894 (N_26894,N_22978,N_20409);
nand U26895 (N_26895,N_20182,N_24632);
nor U26896 (N_26896,N_20360,N_23526);
or U26897 (N_26897,N_23123,N_20659);
nand U26898 (N_26898,N_22171,N_22068);
and U26899 (N_26899,N_21761,N_24463);
or U26900 (N_26900,N_24398,N_21577);
nand U26901 (N_26901,N_21457,N_23976);
xnor U26902 (N_26902,N_22518,N_21608);
nand U26903 (N_26903,N_24371,N_23908);
nor U26904 (N_26904,N_22746,N_22542);
nor U26905 (N_26905,N_20833,N_22198);
xor U26906 (N_26906,N_23713,N_20813);
nor U26907 (N_26907,N_20889,N_24784);
nand U26908 (N_26908,N_20877,N_20480);
nor U26909 (N_26909,N_20205,N_24211);
nor U26910 (N_26910,N_22549,N_21397);
xor U26911 (N_26911,N_24585,N_21816);
nand U26912 (N_26912,N_20207,N_23641);
or U26913 (N_26913,N_22302,N_22079);
nand U26914 (N_26914,N_23561,N_24311);
xnor U26915 (N_26915,N_23515,N_24725);
nand U26916 (N_26916,N_20546,N_22641);
nor U26917 (N_26917,N_22472,N_22780);
nand U26918 (N_26918,N_24016,N_24635);
nor U26919 (N_26919,N_22247,N_20242);
nand U26920 (N_26920,N_22407,N_21436);
nor U26921 (N_26921,N_20898,N_23046);
xor U26922 (N_26922,N_24776,N_21795);
and U26923 (N_26923,N_21971,N_20714);
nand U26924 (N_26924,N_23732,N_22275);
and U26925 (N_26925,N_24349,N_21842);
or U26926 (N_26926,N_20585,N_24377);
or U26927 (N_26927,N_23668,N_22961);
nand U26928 (N_26928,N_20368,N_20712);
nand U26929 (N_26929,N_21372,N_24671);
or U26930 (N_26930,N_24021,N_23156);
xor U26931 (N_26931,N_21755,N_20400);
nor U26932 (N_26932,N_23718,N_21138);
nor U26933 (N_26933,N_21453,N_24858);
xnor U26934 (N_26934,N_24276,N_20781);
nor U26935 (N_26935,N_20801,N_23709);
and U26936 (N_26936,N_24367,N_24153);
nand U26937 (N_26937,N_22974,N_24069);
or U26938 (N_26938,N_24422,N_22004);
xnor U26939 (N_26939,N_23669,N_22906);
or U26940 (N_26940,N_22639,N_23529);
and U26941 (N_26941,N_24739,N_24983);
or U26942 (N_26942,N_23495,N_24475);
xnor U26943 (N_26943,N_23813,N_22269);
and U26944 (N_26944,N_23373,N_23878);
and U26945 (N_26945,N_22160,N_22860);
and U26946 (N_26946,N_21836,N_24740);
nand U26947 (N_26947,N_21037,N_21526);
or U26948 (N_26948,N_20052,N_20748);
nand U26949 (N_26949,N_24789,N_24892);
and U26950 (N_26950,N_23904,N_21967);
nand U26951 (N_26951,N_23252,N_23184);
xor U26952 (N_26952,N_22249,N_23546);
or U26953 (N_26953,N_21777,N_21234);
and U26954 (N_26954,N_21927,N_20986);
nor U26955 (N_26955,N_20233,N_21575);
and U26956 (N_26956,N_24445,N_23520);
nand U26957 (N_26957,N_23143,N_22062);
nand U26958 (N_26958,N_21831,N_24913);
nor U26959 (N_26959,N_21901,N_22086);
or U26960 (N_26960,N_24953,N_23035);
nor U26961 (N_26961,N_24275,N_23105);
and U26962 (N_26962,N_22525,N_20718);
nand U26963 (N_26963,N_22405,N_21685);
or U26964 (N_26964,N_23975,N_22971);
and U26965 (N_26965,N_20321,N_22291);
or U26966 (N_26966,N_23613,N_23508);
nand U26967 (N_26967,N_24325,N_23077);
or U26968 (N_26968,N_22858,N_20214);
nor U26969 (N_26969,N_24129,N_23135);
xnor U26970 (N_26970,N_22984,N_20644);
and U26971 (N_26971,N_23091,N_20664);
xnor U26972 (N_26972,N_23186,N_20553);
nor U26973 (N_26973,N_20831,N_23828);
and U26974 (N_26974,N_24751,N_22493);
nor U26975 (N_26975,N_24290,N_23777);
xnor U26976 (N_26976,N_24388,N_23914);
or U26977 (N_26977,N_22489,N_21254);
or U26978 (N_26978,N_21353,N_20020);
xnor U26979 (N_26979,N_20109,N_24634);
and U26980 (N_26980,N_21047,N_24975);
nand U26981 (N_26981,N_22266,N_21983);
and U26982 (N_26982,N_23378,N_22959);
nand U26983 (N_26983,N_23873,N_21223);
nand U26984 (N_26984,N_22751,N_22798);
and U26985 (N_26985,N_21914,N_20111);
and U26986 (N_26986,N_20510,N_21343);
or U26987 (N_26987,N_20036,N_21144);
and U26988 (N_26988,N_21384,N_21458);
nand U26989 (N_26989,N_21990,N_22507);
or U26990 (N_26990,N_22441,N_24601);
nor U26991 (N_26991,N_20851,N_20453);
or U26992 (N_26992,N_23477,N_24047);
xnor U26993 (N_26993,N_23212,N_22914);
or U26994 (N_26994,N_23909,N_21978);
nor U26995 (N_26995,N_24779,N_22034);
or U26996 (N_26996,N_24124,N_24577);
nand U26997 (N_26997,N_22129,N_22564);
nand U26998 (N_26998,N_21256,N_20045);
and U26999 (N_26999,N_20719,N_21270);
nand U27000 (N_27000,N_20780,N_20481);
xor U27001 (N_27001,N_20817,N_23218);
nand U27002 (N_27002,N_20930,N_20309);
and U27003 (N_27003,N_24390,N_21581);
nand U27004 (N_27004,N_23351,N_24691);
nand U27005 (N_27005,N_20367,N_21211);
nor U27006 (N_27006,N_20165,N_24468);
nand U27007 (N_27007,N_21493,N_22054);
or U27008 (N_27008,N_21399,N_20842);
or U27009 (N_27009,N_23095,N_24191);
and U27010 (N_27010,N_20038,N_24130);
and U27011 (N_27011,N_23728,N_22329);
nor U27012 (N_27012,N_24524,N_21011);
xor U27013 (N_27013,N_24221,N_24562);
nand U27014 (N_27014,N_20151,N_22958);
or U27015 (N_27015,N_24270,N_24034);
and U27016 (N_27016,N_20252,N_23499);
nand U27017 (N_27017,N_20682,N_23737);
nor U27018 (N_27018,N_21461,N_20506);
or U27019 (N_27019,N_24451,N_24569);
nand U27020 (N_27020,N_21747,N_20273);
and U27021 (N_27021,N_20239,N_23601);
nor U27022 (N_27022,N_24194,N_22163);
and U27023 (N_27023,N_21278,N_20727);
xnor U27024 (N_27024,N_22753,N_22949);
nor U27025 (N_27025,N_23460,N_24658);
nand U27026 (N_27026,N_23565,N_23024);
or U27027 (N_27027,N_21293,N_20558);
and U27028 (N_27028,N_24096,N_20456);
or U27029 (N_27029,N_24170,N_24772);
or U27030 (N_27030,N_20752,N_23276);
nor U27031 (N_27031,N_20598,N_24673);
nor U27032 (N_27032,N_21558,N_24896);
nand U27033 (N_27033,N_24269,N_23971);
nand U27034 (N_27034,N_20482,N_22121);
or U27035 (N_27035,N_20716,N_23307);
nand U27036 (N_27036,N_22253,N_21098);
xor U27037 (N_27037,N_22402,N_20871);
nor U27038 (N_27038,N_22073,N_20459);
nor U27039 (N_27039,N_22183,N_24678);
nand U27040 (N_27040,N_22512,N_24573);
nor U27041 (N_27041,N_21802,N_20646);
and U27042 (N_27042,N_22172,N_21764);
or U27043 (N_27043,N_21821,N_20008);
xor U27044 (N_27044,N_24312,N_22184);
and U27045 (N_27045,N_20838,N_21307);
nor U27046 (N_27046,N_20767,N_20464);
nor U27047 (N_27047,N_22231,N_20187);
nand U27048 (N_27048,N_23598,N_24341);
nor U27049 (N_27049,N_22066,N_22598);
xor U27050 (N_27050,N_23202,N_20348);
or U27051 (N_27051,N_20212,N_23027);
nor U27052 (N_27052,N_23686,N_23610);
nand U27053 (N_27053,N_23166,N_23277);
xor U27054 (N_27054,N_24749,N_24920);
nand U27055 (N_27055,N_22756,N_21324);
and U27056 (N_27056,N_20495,N_20691);
nor U27057 (N_27057,N_20355,N_23261);
nand U27058 (N_27058,N_23263,N_20332);
or U27059 (N_27059,N_23658,N_23388);
xnor U27060 (N_27060,N_21145,N_24381);
nor U27061 (N_27061,N_21987,N_22002);
and U27062 (N_27062,N_24674,N_24241);
nor U27063 (N_27063,N_24816,N_20154);
or U27064 (N_27064,N_20751,N_21277);
and U27065 (N_27065,N_20760,N_21740);
xnor U27066 (N_27066,N_23227,N_22364);
nor U27067 (N_27067,N_20523,N_22790);
nor U27068 (N_27068,N_22814,N_21999);
nor U27069 (N_27069,N_21330,N_21383);
nor U27070 (N_27070,N_23455,N_22726);
nor U27071 (N_27071,N_24939,N_21767);
nand U27072 (N_27072,N_22920,N_21610);
or U27073 (N_27073,N_20096,N_23372);
nand U27074 (N_27074,N_24646,N_22795);
or U27075 (N_27075,N_23819,N_20826);
nand U27076 (N_27076,N_21434,N_22327);
xnor U27077 (N_27077,N_23110,N_23386);
nor U27078 (N_27078,N_23211,N_22463);
and U27079 (N_27079,N_23589,N_21412);
nor U27080 (N_27080,N_24581,N_23382);
xnor U27081 (N_27081,N_24337,N_24582);
or U27082 (N_27082,N_22810,N_21111);
and U27083 (N_27083,N_22972,N_23329);
nor U27084 (N_27084,N_23637,N_24002);
nor U27085 (N_27085,N_24277,N_20003);
and U27086 (N_27086,N_20901,N_23000);
or U27087 (N_27087,N_24787,N_22619);
and U27088 (N_27088,N_24454,N_22922);
and U27089 (N_27089,N_22426,N_22576);
or U27090 (N_27090,N_20447,N_23543);
and U27091 (N_27091,N_24703,N_21275);
nor U27092 (N_27092,N_22800,N_21661);
or U27093 (N_27093,N_22688,N_24353);
nor U27094 (N_27094,N_23540,N_22484);
xnor U27095 (N_27095,N_22088,N_22785);
and U27096 (N_27096,N_21337,N_23871);
and U27097 (N_27097,N_22815,N_22379);
or U27098 (N_27098,N_21096,N_22725);
nand U27099 (N_27099,N_22532,N_20492);
nor U27100 (N_27100,N_20786,N_22554);
nand U27101 (N_27101,N_23651,N_24104);
and U27102 (N_27102,N_20962,N_20235);
nor U27103 (N_27103,N_23784,N_20155);
nor U27104 (N_27104,N_20508,N_20903);
nor U27105 (N_27105,N_21230,N_21389);
or U27106 (N_27106,N_23918,N_21503);
nor U27107 (N_27107,N_20974,N_24321);
nor U27108 (N_27108,N_24831,N_21535);
nor U27109 (N_27109,N_24278,N_23053);
nand U27110 (N_27110,N_21845,N_24987);
or U27111 (N_27111,N_24446,N_22873);
or U27112 (N_27112,N_23286,N_23899);
or U27113 (N_27113,N_21173,N_24007);
and U27114 (N_27114,N_24481,N_24217);
and U27115 (N_27115,N_22106,N_21612);
xor U27116 (N_27116,N_21957,N_22043);
nand U27117 (N_27117,N_21989,N_22310);
nand U27118 (N_27118,N_23511,N_23125);
and U27119 (N_27119,N_24567,N_23702);
or U27120 (N_27120,N_20219,N_23884);
and U27121 (N_27121,N_21235,N_20366);
nor U27122 (N_27122,N_22757,N_21900);
nor U27123 (N_27123,N_21311,N_23993);
nand U27124 (N_27124,N_23146,N_23065);
nor U27125 (N_27125,N_20010,N_24382);
and U27126 (N_27126,N_24735,N_20436);
nor U27127 (N_27127,N_21887,N_24863);
or U27128 (N_27128,N_22962,N_20408);
and U27129 (N_27129,N_21718,N_22384);
nand U27130 (N_27130,N_21941,N_22057);
nand U27131 (N_27131,N_22729,N_20289);
and U27132 (N_27132,N_21285,N_23927);
or U27133 (N_27133,N_23843,N_22109);
xor U27134 (N_27134,N_21813,N_23003);
or U27135 (N_27135,N_21387,N_23136);
nand U27136 (N_27136,N_20416,N_20912);
nor U27137 (N_27137,N_23947,N_21214);
xor U27138 (N_27138,N_24232,N_22855);
and U27139 (N_27139,N_23023,N_23405);
nor U27140 (N_27140,N_24775,N_21960);
or U27141 (N_27141,N_23039,N_23747);
or U27142 (N_27142,N_22150,N_21131);
and U27143 (N_27143,N_21367,N_24344);
or U27144 (N_27144,N_20657,N_24676);
or U27145 (N_27145,N_21818,N_24547);
nor U27146 (N_27146,N_23148,N_22769);
nor U27147 (N_27147,N_20968,N_23853);
nand U27148 (N_27148,N_23639,N_24851);
and U27149 (N_27149,N_24229,N_20717);
or U27150 (N_27150,N_22805,N_21290);
nand U27151 (N_27151,N_20832,N_20840);
nand U27152 (N_27152,N_22904,N_20491);
nand U27153 (N_27153,N_20171,N_21425);
or U27154 (N_27154,N_22239,N_20079);
nor U27155 (N_27155,N_23517,N_23633);
nor U27156 (N_27156,N_24000,N_22282);
nand U27157 (N_27157,N_23542,N_21294);
nand U27158 (N_27158,N_24521,N_24030);
nor U27159 (N_27159,N_20365,N_21348);
nand U27160 (N_27160,N_20353,N_20709);
and U27161 (N_27161,N_20980,N_21665);
nand U27162 (N_27162,N_20828,N_20386);
or U27163 (N_27163,N_22957,N_22759);
or U27164 (N_27164,N_23249,N_20805);
or U27165 (N_27165,N_20941,N_24760);
and U27166 (N_27166,N_20294,N_22351);
nor U27167 (N_27167,N_20381,N_20869);
and U27168 (N_27168,N_24263,N_20607);
nor U27169 (N_27169,N_21815,N_22414);
and U27170 (N_27170,N_24242,N_24897);
nand U27171 (N_27171,N_22341,N_20222);
or U27172 (N_27172,N_22410,N_21065);
nor U27173 (N_27173,N_22308,N_23923);
and U27174 (N_27174,N_20276,N_21835);
xor U27175 (N_27175,N_20164,N_22305);
or U27176 (N_27176,N_22393,N_20025);
xnor U27177 (N_27177,N_22016,N_20145);
nor U27178 (N_27178,N_24536,N_21015);
nand U27179 (N_27179,N_20450,N_24599);
or U27180 (N_27180,N_21555,N_23791);
nor U27181 (N_27181,N_23322,N_21393);
and U27182 (N_27182,N_24156,N_20511);
and U27183 (N_27183,N_20248,N_22373);
or U27184 (N_27184,N_22296,N_23362);
or U27185 (N_27185,N_20401,N_24109);
or U27186 (N_27186,N_23265,N_21284);
and U27187 (N_27187,N_24308,N_22289);
or U27188 (N_27188,N_20110,N_22259);
and U27189 (N_27189,N_20892,N_20326);
nor U27190 (N_27190,N_24285,N_20736);
or U27191 (N_27191,N_20847,N_22818);
and U27192 (N_27192,N_24504,N_20380);
and U27193 (N_27193,N_23366,N_22473);
or U27194 (N_27194,N_24945,N_23361);
nor U27195 (N_27195,N_23605,N_22122);
nor U27196 (N_27196,N_20759,N_24056);
nor U27197 (N_27197,N_24004,N_23278);
and U27198 (N_27198,N_24712,N_22789);
nor U27199 (N_27199,N_23141,N_22326);
or U27200 (N_27200,N_20542,N_21335);
and U27201 (N_27201,N_24580,N_24292);
nand U27202 (N_27202,N_24618,N_24985);
or U27203 (N_27203,N_21843,N_23676);
nor U27204 (N_27204,N_22220,N_21426);
and U27205 (N_27205,N_20441,N_22813);
or U27206 (N_27206,N_20806,N_23743);
nand U27207 (N_27207,N_24018,N_21544);
nand U27208 (N_27208,N_21807,N_21439);
and U27209 (N_27209,N_23585,N_24098);
nor U27210 (N_27210,N_24546,N_23860);
and U27211 (N_27211,N_24706,N_23892);
or U27212 (N_27212,N_24767,N_22462);
xor U27213 (N_27213,N_22660,N_23701);
xnor U27214 (N_27214,N_23704,N_21046);
xnor U27215 (N_27215,N_21906,N_20115);
nor U27216 (N_27216,N_23275,N_22737);
nand U27217 (N_27217,N_22479,N_24399);
nor U27218 (N_27218,N_20745,N_22250);
or U27219 (N_27219,N_22793,N_24151);
or U27220 (N_27220,N_23666,N_23300);
nand U27221 (N_27221,N_22531,N_20863);
or U27222 (N_27222,N_23833,N_23086);
nand U27223 (N_27223,N_23762,N_20161);
and U27224 (N_27224,N_23090,N_22017);
or U27225 (N_27225,N_22850,N_20267);
nand U27226 (N_27226,N_24040,N_20688);
nand U27227 (N_27227,N_22006,N_21013);
nand U27228 (N_27228,N_23411,N_24994);
or U27229 (N_27229,N_22343,N_22432);
and U27230 (N_27230,N_23533,N_23072);
and U27231 (N_27231,N_20413,N_21667);
nor U27232 (N_27232,N_24847,N_22845);
nand U27233 (N_27233,N_24921,N_24619);
nor U27234 (N_27234,N_22311,N_24470);
or U27235 (N_27235,N_23327,N_21808);
and U27236 (N_27236,N_23096,N_22485);
and U27237 (N_27237,N_21965,N_22103);
nor U27238 (N_27238,N_22399,N_23996);
and U27239 (N_27239,N_20789,N_21373);
or U27240 (N_27240,N_22293,N_23409);
nand U27241 (N_27241,N_20785,N_22024);
nand U27242 (N_27242,N_21334,N_22609);
and U27243 (N_27243,N_22346,N_23350);
or U27244 (N_27244,N_22378,N_23614);
nand U27245 (N_27245,N_20911,N_22021);
or U27246 (N_27246,N_21101,N_24833);
nand U27247 (N_27247,N_22312,N_22740);
and U27248 (N_27248,N_24412,N_20114);
xor U27249 (N_27249,N_21331,N_23145);
xnor U27250 (N_27250,N_23693,N_22413);
nor U27251 (N_27251,N_21105,N_21791);
xor U27252 (N_27252,N_20530,N_20379);
or U27253 (N_27253,N_22390,N_21809);
or U27254 (N_27254,N_21083,N_23172);
and U27255 (N_27255,N_21456,N_21928);
nor U27256 (N_27256,N_24511,N_22010);
nand U27257 (N_27257,N_21241,N_21593);
xor U27258 (N_27258,N_22114,N_21354);
and U27259 (N_27259,N_20006,N_20069);
xor U27260 (N_27260,N_21142,N_23699);
nor U27261 (N_27261,N_22966,N_22281);
nand U27262 (N_27262,N_21366,N_23431);
or U27263 (N_27263,N_22593,N_24160);
and U27264 (N_27264,N_21139,N_23772);
or U27265 (N_27265,N_20085,N_20794);
and U27266 (N_27266,N_22816,N_24741);
and U27267 (N_27267,N_23523,N_24823);
nand U27268 (N_27268,N_21783,N_24734);
nand U27269 (N_27269,N_22285,N_21177);
nand U27270 (N_27270,N_24874,N_22655);
nor U27271 (N_27271,N_21295,N_24753);
xnor U27272 (N_27272,N_21521,N_20304);
or U27273 (N_27273,N_20810,N_22363);
or U27274 (N_27274,N_22519,N_21703);
and U27275 (N_27275,N_22090,N_23458);
or U27276 (N_27276,N_20479,N_23991);
or U27277 (N_27277,N_24606,N_24857);
and U27278 (N_27278,N_22579,N_21686);
xnor U27279 (N_27279,N_21451,N_20206);
nand U27280 (N_27280,N_24139,N_24427);
and U27281 (N_27281,N_24244,N_23497);
xor U27282 (N_27282,N_24474,N_24195);
or U27283 (N_27283,N_20675,N_24346);
nor U27284 (N_27284,N_24309,N_24522);
and U27285 (N_27285,N_24796,N_22551);
nor U27286 (N_27286,N_24253,N_23640);
and U27287 (N_27287,N_20388,N_24168);
nand U27288 (N_27288,N_21881,N_20726);
or U27289 (N_27289,N_23210,N_21540);
and U27290 (N_27290,N_21246,N_21872);
nand U27291 (N_27291,N_20957,N_22656);
nor U27292 (N_27292,N_24886,N_24859);
and U27293 (N_27293,N_20385,N_22020);
or U27294 (N_27294,N_22706,N_23100);
or U27295 (N_27295,N_24799,N_22261);
nand U27296 (N_27296,N_23104,N_21800);
nor U27297 (N_27297,N_24770,N_20699);
nor U27298 (N_27298,N_20705,N_21556);
and U27299 (N_27299,N_23281,N_23509);
nand U27300 (N_27300,N_22195,N_24415);
nor U27301 (N_27301,N_21171,N_20082);
nand U27302 (N_27302,N_22224,N_24324);
or U27303 (N_27303,N_20034,N_21288);
and U27304 (N_27304,N_23225,N_22627);
nor U27305 (N_27305,N_23606,N_24062);
nor U27306 (N_27306,N_20724,N_20587);
and U27307 (N_27307,N_20514,N_21735);
and U27308 (N_27308,N_23488,N_21280);
and U27309 (N_27309,N_23479,N_23033);
nor U27310 (N_27310,N_24904,N_22599);
or U27311 (N_27311,N_21569,N_20570);
or U27312 (N_27312,N_20102,N_21123);
nand U27313 (N_27313,N_23921,N_23888);
nor U27314 (N_27314,N_21855,N_21609);
nand U27315 (N_27315,N_24937,N_21824);
and U27316 (N_27316,N_24682,N_24808);
nand U27317 (N_27317,N_24262,N_22014);
and U27318 (N_27318,N_21736,N_24455);
nor U27319 (N_27319,N_21475,N_21669);
nor U27320 (N_27320,N_20016,N_21760);
and U27321 (N_27321,N_21626,N_20628);
or U27322 (N_27322,N_24316,N_22056);
nand U27323 (N_27323,N_24748,N_24798);
and U27324 (N_27324,N_23336,N_21247);
and U27325 (N_27325,N_22264,N_20706);
nor U27326 (N_27326,N_20430,N_24190);
nor U27327 (N_27327,N_21968,N_23544);
nor U27328 (N_27328,N_21178,N_21260);
and U27329 (N_27329,N_22468,N_23512);
nand U27330 (N_27330,N_24083,N_23057);
nor U27331 (N_27331,N_24923,N_22454);
or U27332 (N_27332,N_24842,N_23597);
nand U27333 (N_27333,N_21073,N_23773);
nand U27334 (N_27334,N_21153,N_23180);
xnor U27335 (N_27335,N_20226,N_20591);
nor U27336 (N_27336,N_20597,N_20015);
and U27337 (N_27337,N_21701,N_24322);
nor U27338 (N_27338,N_20050,N_24882);
and U27339 (N_27339,N_23016,N_20725);
xor U27340 (N_27340,N_20148,N_23566);
nand U27341 (N_27341,N_21460,N_21874);
or U27342 (N_27342,N_21547,N_24645);
nand U27343 (N_27343,N_20497,N_21996);
or U27344 (N_27344,N_20310,N_22347);
or U27345 (N_27345,N_20881,N_21356);
and U27346 (N_27346,N_23951,N_24274);
nand U27347 (N_27347,N_23558,N_22516);
xor U27348 (N_27348,N_23420,N_24738);
nor U27349 (N_27349,N_23051,N_23962);
and U27350 (N_27350,N_24849,N_22360);
and U27351 (N_27351,N_22649,N_21895);
nand U27352 (N_27352,N_22206,N_22354);
nand U27353 (N_27353,N_24112,N_23069);
nand U27354 (N_27354,N_21745,N_20635);
and U27355 (N_27355,N_22509,N_20225);
and U27356 (N_27356,N_20245,N_21194);
nor U27357 (N_27357,N_22820,N_21151);
nand U27358 (N_27358,N_20561,N_22952);
xnor U27359 (N_27359,N_23646,N_23043);
xnor U27360 (N_27360,N_21820,N_24587);
nor U27361 (N_27361,N_24912,N_20985);
nand U27362 (N_27362,N_23245,N_23617);
and U27363 (N_27363,N_20103,N_22767);
nor U27364 (N_27364,N_23608,N_24966);
xnor U27365 (N_27365,N_22638,N_24763);
or U27366 (N_27366,N_20555,N_23570);
xor U27367 (N_27367,N_24224,N_24989);
and U27368 (N_27368,N_22174,N_20469);
or U27369 (N_27369,N_22488,N_24396);
nand U27370 (N_27370,N_22139,N_23484);
xnor U27371 (N_27371,N_23124,N_20275);
xor U27372 (N_27372,N_24993,N_24400);
or U27373 (N_27373,N_22880,N_23356);
or U27374 (N_27374,N_21024,N_22149);
or U27375 (N_27375,N_21666,N_23864);
nor U27376 (N_27376,N_21851,N_24810);
nor U27377 (N_27377,N_22847,N_22396);
and U27378 (N_27378,N_24924,N_23751);
and U27379 (N_27379,N_23102,N_21454);
nor U27380 (N_27380,N_23710,N_23531);
nor U27381 (N_27381,N_20169,N_23407);
xor U27382 (N_27382,N_21574,N_23612);
or U27383 (N_27383,N_22631,N_21531);
nor U27384 (N_27384,N_22431,N_22117);
or U27385 (N_27385,N_21552,N_22801);
nand U27386 (N_27386,N_23337,N_21688);
or U27387 (N_27387,N_22909,N_20574);
or U27388 (N_27388,N_23905,N_24956);
or U27389 (N_27389,N_21056,N_24565);
and U27390 (N_27390,N_23501,N_24548);
nand U27391 (N_27391,N_23056,N_23295);
nor U27392 (N_27392,N_22500,N_20501);
nand U27393 (N_27393,N_20731,N_20920);
and U27394 (N_27394,N_23770,N_22763);
and U27395 (N_27395,N_24351,N_23208);
nor U27396 (N_27396,N_23596,N_24046);
xor U27397 (N_27397,N_20221,N_22295);
xnor U27398 (N_27398,N_21248,N_21025);
nand U27399 (N_27399,N_21939,N_23887);
or U27400 (N_27400,N_24762,N_20080);
xor U27401 (N_27401,N_23880,N_23767);
and U27402 (N_27402,N_24150,N_24972);
or U27403 (N_27403,N_20945,N_21634);
nand U27404 (N_27404,N_20729,N_24106);
nand U27405 (N_27405,N_22461,N_23530);
nor U27406 (N_27406,N_20995,N_21036);
and U27407 (N_27407,N_21156,N_22188);
and U27408 (N_27408,N_24127,N_24791);
or U27409 (N_27409,N_20586,N_22868);
xnor U27410 (N_27410,N_22381,N_23837);
and U27411 (N_27411,N_22344,N_22723);
xor U27412 (N_27412,N_24180,N_20593);
xnor U27413 (N_27413,N_20272,N_24271);
xor U27414 (N_27414,N_20403,N_22555);
and U27415 (N_27415,N_24944,N_21203);
or U27416 (N_27416,N_21420,N_20259);
and U27417 (N_27417,N_24852,N_21403);
nor U27418 (N_27418,N_20037,N_21659);
and U27419 (N_27419,N_23196,N_22775);
nor U27420 (N_27420,N_21867,N_23532);
nor U27421 (N_27421,N_24086,N_22268);
nor U27422 (N_27422,N_22568,N_20625);
xor U27423 (N_27423,N_22055,N_20370);
nor U27424 (N_27424,N_22944,N_22586);
or U27425 (N_27425,N_23663,N_20744);
nor U27426 (N_27426,N_20253,N_24528);
and U27427 (N_27427,N_20958,N_24225);
or U27428 (N_27428,N_21620,N_24215);
nand U27429 (N_27429,N_23961,N_24765);
or U27430 (N_27430,N_23949,N_21068);
or U27431 (N_27431,N_23783,N_21954);
nor U27432 (N_27432,N_24761,N_23010);
nor U27433 (N_27433,N_24268,N_22632);
or U27434 (N_27434,N_24687,N_20612);
nor U27435 (N_27435,N_20136,N_24169);
and U27436 (N_27436,N_21746,N_21934);
xor U27437 (N_27437,N_22877,N_23369);
xor U27438 (N_27438,N_20475,N_20223);
nor U27439 (N_27439,N_21532,N_23683);
and U27440 (N_27440,N_24237,N_23981);
nand U27441 (N_27441,N_21463,N_20446);
or U27442 (N_27442,N_23868,N_21301);
nor U27443 (N_27443,N_24363,N_20951);
or U27444 (N_27444,N_23173,N_20075);
and U27445 (N_27445,N_21674,N_24233);
nand U27446 (N_27446,N_22279,N_21980);
or U27447 (N_27447,N_20720,N_22975);
or U27448 (N_27448,N_23577,N_23151);
nand U27449 (N_27449,N_24837,N_22717);
nor U27450 (N_27450,N_23400,N_21731);
or U27451 (N_27451,N_21208,N_24557);
and U27452 (N_27452,N_20369,N_20547);
nand U27453 (N_27453,N_22686,N_24605);
nand U27454 (N_27454,N_22124,N_20875);
nor U27455 (N_27455,N_21871,N_20121);
nand U27456 (N_27456,N_21265,N_22600);
or U27457 (N_27457,N_22070,N_21344);
nand U27458 (N_27458,N_23607,N_23506);
and U27459 (N_27459,N_23026,N_23688);
and U27460 (N_27460,N_20384,N_20270);
nand U27461 (N_27461,N_24650,N_23081);
nor U27462 (N_27462,N_22745,N_22875);
nand U27463 (N_27463,N_22138,N_24572);
or U27464 (N_27464,N_23309,N_20562);
and U27465 (N_27465,N_24245,N_22616);
nand U27466 (N_27466,N_22534,N_21405);
or U27467 (N_27467,N_21202,N_20132);
nor U27468 (N_27468,N_21406,N_20351);
or U27469 (N_27469,N_24860,N_21681);
or U27470 (N_27470,N_20444,N_20268);
nor U27471 (N_27471,N_20651,N_24719);
xor U27472 (N_27472,N_21628,N_23117);
or U27473 (N_27473,N_23347,N_23572);
or U27474 (N_27474,N_21007,N_22108);
nand U27475 (N_27475,N_22153,N_22633);
or U27476 (N_27476,N_22069,N_24175);
nand U27477 (N_27477,N_23620,N_20288);
or U27478 (N_27478,N_23672,N_21066);
xnor U27479 (N_27479,N_24387,N_23481);
nand U27480 (N_27480,N_24208,N_21814);
and U27481 (N_27481,N_20101,N_20117);
nor U27482 (N_27482,N_20314,N_23715);
nand U27483 (N_27483,N_20566,N_22005);
and U27484 (N_27484,N_20641,N_22714);
nor U27485 (N_27485,N_20743,N_24954);
and U27486 (N_27486,N_24332,N_20967);
nand U27487 (N_27487,N_20573,N_23692);
xnor U27488 (N_27488,N_24864,N_22167);
nor U27489 (N_27489,N_23815,N_20002);
nand U27490 (N_27490,N_22428,N_21283);
and U27491 (N_27491,N_24465,N_24003);
nand U27492 (N_27492,N_23534,N_21730);
nand U27493 (N_27493,N_20529,N_21213);
nand U27494 (N_27494,N_20790,N_21923);
nand U27495 (N_27495,N_22187,N_22353);
xor U27496 (N_27496,N_20704,N_20776);
nor U27497 (N_27497,N_22864,N_24503);
xnor U27498 (N_27498,N_21539,N_20346);
or U27499 (N_27499,N_20285,N_23246);
or U27500 (N_27500,N_23564,N_23106);
and U27501 (N_27501,N_22706,N_21523);
and U27502 (N_27502,N_20647,N_24666);
nand U27503 (N_27503,N_20744,N_22649);
and U27504 (N_27504,N_22946,N_23809);
or U27505 (N_27505,N_22571,N_22529);
nand U27506 (N_27506,N_20924,N_24620);
nor U27507 (N_27507,N_20497,N_21242);
xor U27508 (N_27508,N_20223,N_20935);
nor U27509 (N_27509,N_24654,N_22291);
nand U27510 (N_27510,N_23786,N_24238);
nand U27511 (N_27511,N_24844,N_23701);
and U27512 (N_27512,N_23078,N_23502);
nand U27513 (N_27513,N_21215,N_21398);
and U27514 (N_27514,N_22139,N_23252);
or U27515 (N_27515,N_23674,N_24879);
nor U27516 (N_27516,N_22593,N_20466);
nor U27517 (N_27517,N_21238,N_21123);
nand U27518 (N_27518,N_24378,N_23707);
nor U27519 (N_27519,N_24667,N_22123);
nor U27520 (N_27520,N_24288,N_22404);
xor U27521 (N_27521,N_24863,N_23803);
nand U27522 (N_27522,N_22412,N_20796);
or U27523 (N_27523,N_21843,N_20542);
or U27524 (N_27524,N_20609,N_22122);
xnor U27525 (N_27525,N_20607,N_24043);
or U27526 (N_27526,N_21857,N_20588);
or U27527 (N_27527,N_24856,N_24172);
or U27528 (N_27528,N_22943,N_24954);
nand U27529 (N_27529,N_23514,N_21357);
or U27530 (N_27530,N_24618,N_22605);
nor U27531 (N_27531,N_20121,N_24673);
and U27532 (N_27532,N_24184,N_24469);
and U27533 (N_27533,N_22609,N_20651);
nor U27534 (N_27534,N_21864,N_22417);
xnor U27535 (N_27535,N_21170,N_24483);
and U27536 (N_27536,N_21017,N_20232);
nor U27537 (N_27537,N_22941,N_21354);
nand U27538 (N_27538,N_21917,N_22973);
and U27539 (N_27539,N_24777,N_21848);
nand U27540 (N_27540,N_23039,N_21202);
nand U27541 (N_27541,N_23020,N_21191);
nand U27542 (N_27542,N_20105,N_24834);
nor U27543 (N_27543,N_23164,N_24317);
xor U27544 (N_27544,N_23412,N_21129);
nor U27545 (N_27545,N_21903,N_20014);
nor U27546 (N_27546,N_24036,N_24151);
nor U27547 (N_27547,N_22511,N_23413);
and U27548 (N_27548,N_21667,N_24306);
and U27549 (N_27549,N_24785,N_22292);
or U27550 (N_27550,N_22880,N_22417);
or U27551 (N_27551,N_24810,N_21085);
and U27552 (N_27552,N_20758,N_23775);
or U27553 (N_27553,N_22123,N_23440);
and U27554 (N_27554,N_23445,N_24626);
nor U27555 (N_27555,N_22547,N_20737);
xnor U27556 (N_27556,N_23876,N_23549);
and U27557 (N_27557,N_20105,N_23255);
nor U27558 (N_27558,N_20738,N_20407);
and U27559 (N_27559,N_23691,N_22581);
nor U27560 (N_27560,N_23272,N_24148);
nand U27561 (N_27561,N_22752,N_21007);
and U27562 (N_27562,N_23432,N_24968);
or U27563 (N_27563,N_24056,N_24845);
and U27564 (N_27564,N_23628,N_24112);
and U27565 (N_27565,N_23956,N_22582);
nand U27566 (N_27566,N_22259,N_23228);
and U27567 (N_27567,N_22963,N_20345);
nor U27568 (N_27568,N_23596,N_22926);
or U27569 (N_27569,N_24245,N_20311);
nand U27570 (N_27570,N_21384,N_23078);
xor U27571 (N_27571,N_24695,N_21858);
or U27572 (N_27572,N_24606,N_23300);
nand U27573 (N_27573,N_21978,N_20427);
nor U27574 (N_27574,N_22566,N_23889);
and U27575 (N_27575,N_23050,N_23210);
and U27576 (N_27576,N_24326,N_24579);
nand U27577 (N_27577,N_21297,N_22889);
or U27578 (N_27578,N_22609,N_20370);
nand U27579 (N_27579,N_23168,N_21675);
and U27580 (N_27580,N_20117,N_22139);
nand U27581 (N_27581,N_21290,N_23177);
xnor U27582 (N_27582,N_24913,N_21168);
or U27583 (N_27583,N_24894,N_23134);
nand U27584 (N_27584,N_24520,N_20089);
and U27585 (N_27585,N_21523,N_20728);
or U27586 (N_27586,N_22556,N_24514);
nand U27587 (N_27587,N_22879,N_23408);
nor U27588 (N_27588,N_23287,N_22157);
xnor U27589 (N_27589,N_22138,N_20734);
nor U27590 (N_27590,N_24617,N_23082);
nand U27591 (N_27591,N_24669,N_20824);
nand U27592 (N_27592,N_24718,N_24314);
and U27593 (N_27593,N_24537,N_20111);
nor U27594 (N_27594,N_24492,N_22293);
and U27595 (N_27595,N_24606,N_23469);
xnor U27596 (N_27596,N_23371,N_22906);
nor U27597 (N_27597,N_21172,N_24799);
or U27598 (N_27598,N_22226,N_24739);
xor U27599 (N_27599,N_22575,N_20657);
and U27600 (N_27600,N_24260,N_20668);
and U27601 (N_27601,N_23218,N_20693);
nand U27602 (N_27602,N_21759,N_20979);
nand U27603 (N_27603,N_20794,N_23430);
or U27604 (N_27604,N_21946,N_20164);
and U27605 (N_27605,N_20107,N_24192);
nand U27606 (N_27606,N_20727,N_24932);
or U27607 (N_27607,N_23442,N_23007);
nor U27608 (N_27608,N_23997,N_22000);
nand U27609 (N_27609,N_21133,N_24831);
nor U27610 (N_27610,N_24435,N_22369);
nor U27611 (N_27611,N_20287,N_24334);
nand U27612 (N_27612,N_23438,N_23766);
and U27613 (N_27613,N_21012,N_21752);
and U27614 (N_27614,N_23721,N_24953);
or U27615 (N_27615,N_23847,N_22068);
nand U27616 (N_27616,N_23347,N_20032);
nand U27617 (N_27617,N_23166,N_22008);
xnor U27618 (N_27618,N_23298,N_23448);
nor U27619 (N_27619,N_24179,N_24927);
xnor U27620 (N_27620,N_23543,N_21213);
or U27621 (N_27621,N_24021,N_20618);
nor U27622 (N_27622,N_24863,N_23418);
nor U27623 (N_27623,N_20151,N_22334);
nand U27624 (N_27624,N_23220,N_23859);
nand U27625 (N_27625,N_20404,N_20250);
and U27626 (N_27626,N_23622,N_21638);
nand U27627 (N_27627,N_24493,N_21143);
or U27628 (N_27628,N_23830,N_23477);
or U27629 (N_27629,N_22877,N_21614);
xor U27630 (N_27630,N_24986,N_22429);
nand U27631 (N_27631,N_21874,N_20509);
xnor U27632 (N_27632,N_23029,N_21040);
or U27633 (N_27633,N_23164,N_23720);
nor U27634 (N_27634,N_21141,N_20573);
nand U27635 (N_27635,N_21423,N_21752);
nor U27636 (N_27636,N_24766,N_24145);
or U27637 (N_27637,N_24644,N_24468);
or U27638 (N_27638,N_20332,N_23648);
nor U27639 (N_27639,N_22813,N_24917);
nand U27640 (N_27640,N_23307,N_22171);
nand U27641 (N_27641,N_20775,N_22150);
nor U27642 (N_27642,N_24117,N_22991);
nand U27643 (N_27643,N_24721,N_21744);
or U27644 (N_27644,N_20848,N_24127);
and U27645 (N_27645,N_24587,N_23959);
nand U27646 (N_27646,N_20489,N_23042);
or U27647 (N_27647,N_24652,N_22035);
nand U27648 (N_27648,N_23058,N_24387);
nor U27649 (N_27649,N_21128,N_21020);
xnor U27650 (N_27650,N_20756,N_23018);
and U27651 (N_27651,N_23170,N_21360);
or U27652 (N_27652,N_20312,N_23023);
xnor U27653 (N_27653,N_24283,N_21399);
and U27654 (N_27654,N_20116,N_23456);
and U27655 (N_27655,N_24321,N_23549);
nand U27656 (N_27656,N_20949,N_23724);
or U27657 (N_27657,N_24592,N_24333);
or U27658 (N_27658,N_22081,N_22700);
nor U27659 (N_27659,N_22760,N_22511);
and U27660 (N_27660,N_24262,N_22069);
nand U27661 (N_27661,N_23394,N_24026);
nand U27662 (N_27662,N_22754,N_23817);
nor U27663 (N_27663,N_22773,N_20366);
nand U27664 (N_27664,N_24406,N_24785);
nor U27665 (N_27665,N_24361,N_24870);
or U27666 (N_27666,N_21988,N_20519);
xor U27667 (N_27667,N_21936,N_20394);
nand U27668 (N_27668,N_23094,N_21943);
nor U27669 (N_27669,N_20239,N_21424);
and U27670 (N_27670,N_20142,N_24322);
nor U27671 (N_27671,N_20448,N_21325);
nor U27672 (N_27672,N_24433,N_22632);
nand U27673 (N_27673,N_20013,N_20461);
and U27674 (N_27674,N_23740,N_22667);
nand U27675 (N_27675,N_20759,N_21227);
nand U27676 (N_27676,N_22315,N_23446);
or U27677 (N_27677,N_24518,N_23051);
nor U27678 (N_27678,N_21307,N_24663);
nand U27679 (N_27679,N_21573,N_23851);
nor U27680 (N_27680,N_23402,N_23180);
nor U27681 (N_27681,N_20696,N_23983);
or U27682 (N_27682,N_22347,N_24609);
or U27683 (N_27683,N_24172,N_22031);
nor U27684 (N_27684,N_24927,N_20617);
nor U27685 (N_27685,N_24136,N_20551);
xor U27686 (N_27686,N_20615,N_20997);
and U27687 (N_27687,N_22539,N_24827);
xor U27688 (N_27688,N_21202,N_21892);
nand U27689 (N_27689,N_22907,N_23468);
nand U27690 (N_27690,N_20714,N_24630);
nand U27691 (N_27691,N_23414,N_24563);
or U27692 (N_27692,N_22197,N_21927);
nor U27693 (N_27693,N_24734,N_21348);
nand U27694 (N_27694,N_21291,N_22192);
nand U27695 (N_27695,N_23557,N_21037);
or U27696 (N_27696,N_21820,N_24005);
nand U27697 (N_27697,N_23343,N_20064);
or U27698 (N_27698,N_23181,N_23412);
nor U27699 (N_27699,N_21842,N_22736);
and U27700 (N_27700,N_24868,N_21834);
and U27701 (N_27701,N_22851,N_21807);
nand U27702 (N_27702,N_22960,N_21627);
nand U27703 (N_27703,N_20058,N_20087);
xor U27704 (N_27704,N_20995,N_21291);
nand U27705 (N_27705,N_23142,N_24888);
nor U27706 (N_27706,N_22962,N_21067);
nand U27707 (N_27707,N_24614,N_23218);
and U27708 (N_27708,N_24717,N_22009);
and U27709 (N_27709,N_23050,N_23735);
and U27710 (N_27710,N_24107,N_23758);
or U27711 (N_27711,N_21965,N_22031);
or U27712 (N_27712,N_20500,N_20633);
nand U27713 (N_27713,N_20260,N_20463);
and U27714 (N_27714,N_23447,N_21292);
nand U27715 (N_27715,N_21262,N_21079);
or U27716 (N_27716,N_21363,N_20853);
nand U27717 (N_27717,N_21693,N_23122);
xor U27718 (N_27718,N_24727,N_22952);
and U27719 (N_27719,N_24181,N_21823);
nand U27720 (N_27720,N_21350,N_23417);
or U27721 (N_27721,N_20224,N_21230);
nand U27722 (N_27722,N_22708,N_23880);
or U27723 (N_27723,N_21182,N_21769);
nand U27724 (N_27724,N_23041,N_24077);
or U27725 (N_27725,N_22166,N_23926);
nor U27726 (N_27726,N_20366,N_21023);
nor U27727 (N_27727,N_22783,N_20778);
nand U27728 (N_27728,N_21477,N_23481);
nand U27729 (N_27729,N_20059,N_21594);
or U27730 (N_27730,N_24036,N_21165);
nand U27731 (N_27731,N_20844,N_20870);
xor U27732 (N_27732,N_20854,N_24002);
or U27733 (N_27733,N_23780,N_22691);
xor U27734 (N_27734,N_24937,N_21505);
xnor U27735 (N_27735,N_20829,N_23234);
nor U27736 (N_27736,N_23893,N_22585);
nand U27737 (N_27737,N_23141,N_23322);
and U27738 (N_27738,N_24750,N_21224);
nand U27739 (N_27739,N_22911,N_21205);
nand U27740 (N_27740,N_20038,N_23902);
nor U27741 (N_27741,N_24305,N_22110);
nor U27742 (N_27742,N_23227,N_24630);
or U27743 (N_27743,N_20333,N_24076);
and U27744 (N_27744,N_24166,N_21932);
nand U27745 (N_27745,N_24569,N_23904);
nand U27746 (N_27746,N_22905,N_20467);
nor U27747 (N_27747,N_22524,N_20905);
and U27748 (N_27748,N_22124,N_23834);
xor U27749 (N_27749,N_24574,N_23090);
and U27750 (N_27750,N_20879,N_20916);
nor U27751 (N_27751,N_22107,N_21609);
and U27752 (N_27752,N_23701,N_24245);
nand U27753 (N_27753,N_24073,N_21320);
or U27754 (N_27754,N_22025,N_24495);
or U27755 (N_27755,N_24771,N_21781);
nand U27756 (N_27756,N_21214,N_22184);
nand U27757 (N_27757,N_21554,N_24048);
and U27758 (N_27758,N_23282,N_21206);
and U27759 (N_27759,N_24088,N_24624);
nor U27760 (N_27760,N_24835,N_20845);
nor U27761 (N_27761,N_23569,N_21515);
and U27762 (N_27762,N_22614,N_22431);
and U27763 (N_27763,N_21137,N_23295);
nand U27764 (N_27764,N_21664,N_20176);
or U27765 (N_27765,N_21389,N_24152);
nand U27766 (N_27766,N_22940,N_20966);
xnor U27767 (N_27767,N_23702,N_22184);
or U27768 (N_27768,N_22813,N_23764);
nor U27769 (N_27769,N_21049,N_24495);
and U27770 (N_27770,N_24017,N_20723);
or U27771 (N_27771,N_22406,N_23123);
nor U27772 (N_27772,N_21979,N_22262);
xor U27773 (N_27773,N_20673,N_22985);
nor U27774 (N_27774,N_24892,N_21500);
nand U27775 (N_27775,N_24980,N_23598);
or U27776 (N_27776,N_21814,N_23652);
or U27777 (N_27777,N_21176,N_20224);
and U27778 (N_27778,N_23054,N_20789);
nand U27779 (N_27779,N_20146,N_20502);
nor U27780 (N_27780,N_23765,N_22754);
or U27781 (N_27781,N_22564,N_21172);
or U27782 (N_27782,N_20505,N_20951);
nor U27783 (N_27783,N_21327,N_21111);
nor U27784 (N_27784,N_21135,N_22559);
nor U27785 (N_27785,N_22460,N_20490);
nor U27786 (N_27786,N_23055,N_20667);
nand U27787 (N_27787,N_23529,N_22331);
and U27788 (N_27788,N_22977,N_20669);
or U27789 (N_27789,N_23737,N_22107);
nand U27790 (N_27790,N_20387,N_23510);
xnor U27791 (N_27791,N_20784,N_20478);
or U27792 (N_27792,N_24614,N_21234);
or U27793 (N_27793,N_21401,N_23164);
and U27794 (N_27794,N_23445,N_23618);
or U27795 (N_27795,N_23906,N_23298);
nand U27796 (N_27796,N_23886,N_23126);
and U27797 (N_27797,N_22070,N_24931);
nor U27798 (N_27798,N_21365,N_22096);
nand U27799 (N_27799,N_23632,N_24711);
or U27800 (N_27800,N_21026,N_20494);
nor U27801 (N_27801,N_23331,N_20676);
nor U27802 (N_27802,N_23267,N_24202);
nor U27803 (N_27803,N_20993,N_22362);
and U27804 (N_27804,N_22384,N_21052);
nand U27805 (N_27805,N_20602,N_22861);
nand U27806 (N_27806,N_21171,N_24652);
and U27807 (N_27807,N_22534,N_22033);
nor U27808 (N_27808,N_23479,N_24419);
and U27809 (N_27809,N_22274,N_21629);
nor U27810 (N_27810,N_21340,N_23801);
or U27811 (N_27811,N_24929,N_24166);
nand U27812 (N_27812,N_20567,N_24652);
nand U27813 (N_27813,N_20268,N_23316);
nor U27814 (N_27814,N_20221,N_23863);
and U27815 (N_27815,N_22211,N_20855);
nand U27816 (N_27816,N_22977,N_21798);
nor U27817 (N_27817,N_21406,N_20579);
nor U27818 (N_27818,N_22864,N_21171);
or U27819 (N_27819,N_23376,N_20054);
nor U27820 (N_27820,N_22326,N_22405);
and U27821 (N_27821,N_21504,N_23479);
or U27822 (N_27822,N_22599,N_20771);
nor U27823 (N_27823,N_20523,N_22722);
nor U27824 (N_27824,N_23566,N_20891);
or U27825 (N_27825,N_22023,N_20425);
nor U27826 (N_27826,N_24759,N_24219);
or U27827 (N_27827,N_20357,N_24249);
and U27828 (N_27828,N_21459,N_22459);
xor U27829 (N_27829,N_24599,N_24485);
xnor U27830 (N_27830,N_22662,N_22509);
xnor U27831 (N_27831,N_21552,N_23269);
or U27832 (N_27832,N_20148,N_22302);
nor U27833 (N_27833,N_22484,N_24821);
and U27834 (N_27834,N_24408,N_24200);
or U27835 (N_27835,N_22540,N_23788);
nand U27836 (N_27836,N_24066,N_21225);
nand U27837 (N_27837,N_24987,N_24815);
nor U27838 (N_27838,N_24552,N_22546);
nor U27839 (N_27839,N_22018,N_20674);
nor U27840 (N_27840,N_22344,N_20865);
nor U27841 (N_27841,N_22944,N_24340);
or U27842 (N_27842,N_24071,N_21066);
or U27843 (N_27843,N_22589,N_24816);
and U27844 (N_27844,N_24450,N_20440);
and U27845 (N_27845,N_22823,N_24603);
or U27846 (N_27846,N_23046,N_22100);
or U27847 (N_27847,N_20621,N_20149);
and U27848 (N_27848,N_23424,N_23131);
nor U27849 (N_27849,N_23123,N_22811);
nand U27850 (N_27850,N_20824,N_24763);
nand U27851 (N_27851,N_20012,N_20156);
or U27852 (N_27852,N_24933,N_24187);
nor U27853 (N_27853,N_23222,N_23459);
nand U27854 (N_27854,N_22183,N_20527);
xnor U27855 (N_27855,N_23597,N_24537);
xnor U27856 (N_27856,N_22386,N_24003);
nand U27857 (N_27857,N_20513,N_21646);
nor U27858 (N_27858,N_24706,N_22651);
nor U27859 (N_27859,N_21003,N_20361);
or U27860 (N_27860,N_20913,N_20831);
and U27861 (N_27861,N_20087,N_23866);
xnor U27862 (N_27862,N_24439,N_23001);
and U27863 (N_27863,N_21429,N_22503);
xnor U27864 (N_27864,N_20359,N_24337);
nand U27865 (N_27865,N_23851,N_21602);
xor U27866 (N_27866,N_23539,N_24745);
and U27867 (N_27867,N_22006,N_21371);
xor U27868 (N_27868,N_22439,N_23299);
nor U27869 (N_27869,N_22662,N_22325);
and U27870 (N_27870,N_21791,N_23347);
or U27871 (N_27871,N_23068,N_24661);
nand U27872 (N_27872,N_24572,N_24698);
nor U27873 (N_27873,N_21798,N_21822);
nor U27874 (N_27874,N_24665,N_21399);
and U27875 (N_27875,N_21322,N_21046);
nand U27876 (N_27876,N_23375,N_24797);
nor U27877 (N_27877,N_20243,N_21382);
or U27878 (N_27878,N_23681,N_21471);
nor U27879 (N_27879,N_23464,N_21879);
nor U27880 (N_27880,N_21917,N_24772);
and U27881 (N_27881,N_22011,N_23558);
nor U27882 (N_27882,N_20983,N_24357);
nor U27883 (N_27883,N_20749,N_24498);
xnor U27884 (N_27884,N_21833,N_21507);
nor U27885 (N_27885,N_23248,N_23500);
nand U27886 (N_27886,N_23086,N_21649);
nor U27887 (N_27887,N_20623,N_21449);
or U27888 (N_27888,N_24710,N_23586);
or U27889 (N_27889,N_23128,N_22883);
and U27890 (N_27890,N_23459,N_21966);
xor U27891 (N_27891,N_21644,N_23322);
or U27892 (N_27892,N_24894,N_24672);
and U27893 (N_27893,N_21837,N_24493);
or U27894 (N_27894,N_21229,N_23848);
nor U27895 (N_27895,N_22612,N_23728);
nand U27896 (N_27896,N_20050,N_22141);
nor U27897 (N_27897,N_21319,N_20576);
nand U27898 (N_27898,N_24876,N_21961);
and U27899 (N_27899,N_21767,N_21367);
nor U27900 (N_27900,N_22031,N_21360);
nand U27901 (N_27901,N_21557,N_24318);
and U27902 (N_27902,N_23572,N_23505);
nand U27903 (N_27903,N_24780,N_20123);
or U27904 (N_27904,N_24169,N_21604);
nand U27905 (N_27905,N_23836,N_21770);
or U27906 (N_27906,N_20075,N_22997);
and U27907 (N_27907,N_22053,N_22146);
nand U27908 (N_27908,N_23015,N_20589);
and U27909 (N_27909,N_21098,N_21152);
or U27910 (N_27910,N_22145,N_20974);
and U27911 (N_27911,N_23571,N_22231);
nor U27912 (N_27912,N_21056,N_24728);
xor U27913 (N_27913,N_23504,N_23883);
or U27914 (N_27914,N_21436,N_21758);
or U27915 (N_27915,N_21088,N_23340);
nand U27916 (N_27916,N_20718,N_23432);
nand U27917 (N_27917,N_23572,N_20324);
or U27918 (N_27918,N_22636,N_24095);
nor U27919 (N_27919,N_20132,N_21527);
or U27920 (N_27920,N_24290,N_22628);
xnor U27921 (N_27921,N_20938,N_22497);
nand U27922 (N_27922,N_23599,N_20677);
nand U27923 (N_27923,N_22174,N_24704);
nand U27924 (N_27924,N_24165,N_20917);
or U27925 (N_27925,N_20193,N_22878);
or U27926 (N_27926,N_24422,N_22595);
xor U27927 (N_27927,N_24007,N_20789);
and U27928 (N_27928,N_24912,N_20880);
nor U27929 (N_27929,N_23548,N_20008);
xnor U27930 (N_27930,N_22504,N_21499);
or U27931 (N_27931,N_20951,N_23670);
nand U27932 (N_27932,N_24353,N_20429);
nor U27933 (N_27933,N_23443,N_24987);
nand U27934 (N_27934,N_24035,N_24771);
xor U27935 (N_27935,N_21463,N_20366);
or U27936 (N_27936,N_22418,N_24163);
and U27937 (N_27937,N_20686,N_21154);
nor U27938 (N_27938,N_23118,N_21375);
or U27939 (N_27939,N_22073,N_23213);
xor U27940 (N_27940,N_23763,N_23789);
and U27941 (N_27941,N_23574,N_24162);
nor U27942 (N_27942,N_20989,N_20053);
or U27943 (N_27943,N_22224,N_22798);
or U27944 (N_27944,N_20340,N_24449);
nand U27945 (N_27945,N_23588,N_21474);
nand U27946 (N_27946,N_22876,N_20137);
and U27947 (N_27947,N_24168,N_21377);
nor U27948 (N_27948,N_21345,N_24111);
xnor U27949 (N_27949,N_23494,N_23454);
nor U27950 (N_27950,N_23794,N_23920);
or U27951 (N_27951,N_21138,N_22253);
xnor U27952 (N_27952,N_22817,N_24366);
or U27953 (N_27953,N_24709,N_22046);
xor U27954 (N_27954,N_22753,N_21050);
and U27955 (N_27955,N_20856,N_21062);
nand U27956 (N_27956,N_20767,N_21250);
nor U27957 (N_27957,N_24069,N_20740);
nor U27958 (N_27958,N_24792,N_20262);
and U27959 (N_27959,N_20782,N_23369);
and U27960 (N_27960,N_20943,N_21785);
nand U27961 (N_27961,N_20232,N_21967);
nand U27962 (N_27962,N_23629,N_22421);
xnor U27963 (N_27963,N_24892,N_21675);
nand U27964 (N_27964,N_21054,N_20470);
xor U27965 (N_27965,N_20460,N_22348);
xnor U27966 (N_27966,N_23883,N_21221);
nand U27967 (N_27967,N_21050,N_21754);
nor U27968 (N_27968,N_23378,N_21201);
nor U27969 (N_27969,N_24552,N_24901);
and U27970 (N_27970,N_22033,N_20050);
xor U27971 (N_27971,N_22799,N_22912);
or U27972 (N_27972,N_23697,N_23309);
nand U27973 (N_27973,N_20971,N_22850);
and U27974 (N_27974,N_22180,N_24760);
nand U27975 (N_27975,N_22378,N_22414);
and U27976 (N_27976,N_23184,N_23084);
and U27977 (N_27977,N_21099,N_21691);
xnor U27978 (N_27978,N_21182,N_23252);
or U27979 (N_27979,N_22086,N_24503);
nand U27980 (N_27980,N_23863,N_22021);
and U27981 (N_27981,N_20453,N_22840);
and U27982 (N_27982,N_22671,N_21330);
or U27983 (N_27983,N_22625,N_21853);
nand U27984 (N_27984,N_23510,N_22003);
or U27985 (N_27985,N_20489,N_20029);
or U27986 (N_27986,N_23849,N_20410);
nor U27987 (N_27987,N_21597,N_21620);
nor U27988 (N_27988,N_20220,N_21725);
nand U27989 (N_27989,N_22764,N_23020);
nand U27990 (N_27990,N_20379,N_20846);
nor U27991 (N_27991,N_20095,N_21021);
nand U27992 (N_27992,N_21075,N_22368);
and U27993 (N_27993,N_21533,N_20728);
and U27994 (N_27994,N_21210,N_23104);
nand U27995 (N_27995,N_24397,N_20722);
xnor U27996 (N_27996,N_22591,N_24789);
nor U27997 (N_27997,N_23410,N_24300);
xnor U27998 (N_27998,N_22871,N_22068);
nand U27999 (N_27999,N_23691,N_20189);
nand U28000 (N_28000,N_20573,N_23953);
nor U28001 (N_28001,N_24582,N_21448);
nand U28002 (N_28002,N_24272,N_23045);
or U28003 (N_28003,N_24618,N_21555);
nor U28004 (N_28004,N_20989,N_20360);
and U28005 (N_28005,N_20220,N_20494);
nand U28006 (N_28006,N_21303,N_20195);
nand U28007 (N_28007,N_24489,N_23552);
nand U28008 (N_28008,N_24807,N_22621);
or U28009 (N_28009,N_21557,N_23239);
nor U28010 (N_28010,N_20844,N_23260);
or U28011 (N_28011,N_23665,N_24841);
and U28012 (N_28012,N_21697,N_23015);
nor U28013 (N_28013,N_22145,N_20641);
and U28014 (N_28014,N_21616,N_20552);
nand U28015 (N_28015,N_21427,N_22759);
or U28016 (N_28016,N_24039,N_20109);
and U28017 (N_28017,N_23728,N_21027);
nand U28018 (N_28018,N_22758,N_21659);
or U28019 (N_28019,N_23196,N_22342);
and U28020 (N_28020,N_24000,N_24102);
nand U28021 (N_28021,N_24242,N_20057);
and U28022 (N_28022,N_23826,N_23791);
nand U28023 (N_28023,N_22311,N_20235);
nand U28024 (N_28024,N_23869,N_23861);
and U28025 (N_28025,N_21931,N_24911);
and U28026 (N_28026,N_24588,N_22258);
nand U28027 (N_28027,N_21561,N_22395);
and U28028 (N_28028,N_23125,N_22833);
nand U28029 (N_28029,N_23403,N_22550);
nor U28030 (N_28030,N_21800,N_23717);
nand U28031 (N_28031,N_23062,N_20269);
or U28032 (N_28032,N_23058,N_24126);
and U28033 (N_28033,N_23946,N_22081);
nand U28034 (N_28034,N_24518,N_22114);
xnor U28035 (N_28035,N_24863,N_24207);
nand U28036 (N_28036,N_24696,N_21802);
or U28037 (N_28037,N_20136,N_21427);
nand U28038 (N_28038,N_21694,N_23946);
nand U28039 (N_28039,N_20475,N_23991);
nor U28040 (N_28040,N_23817,N_20312);
or U28041 (N_28041,N_20373,N_22311);
or U28042 (N_28042,N_23176,N_21391);
nand U28043 (N_28043,N_24963,N_22809);
nand U28044 (N_28044,N_24314,N_23006);
and U28045 (N_28045,N_21150,N_22847);
or U28046 (N_28046,N_21394,N_20169);
nand U28047 (N_28047,N_20338,N_23129);
nor U28048 (N_28048,N_24280,N_20785);
nand U28049 (N_28049,N_20736,N_21211);
or U28050 (N_28050,N_23244,N_24994);
and U28051 (N_28051,N_22153,N_20520);
xor U28052 (N_28052,N_22934,N_24045);
nand U28053 (N_28053,N_24777,N_23357);
and U28054 (N_28054,N_24954,N_23839);
and U28055 (N_28055,N_23618,N_22805);
or U28056 (N_28056,N_22198,N_22671);
nor U28057 (N_28057,N_20946,N_21236);
nand U28058 (N_28058,N_21210,N_22481);
nor U28059 (N_28059,N_21793,N_22366);
and U28060 (N_28060,N_23550,N_24986);
or U28061 (N_28061,N_20937,N_24422);
and U28062 (N_28062,N_21065,N_22517);
nor U28063 (N_28063,N_22542,N_23746);
or U28064 (N_28064,N_23183,N_22589);
nor U28065 (N_28065,N_24189,N_23729);
nor U28066 (N_28066,N_21128,N_23724);
xnor U28067 (N_28067,N_21182,N_24580);
nand U28068 (N_28068,N_23887,N_21960);
and U28069 (N_28069,N_22687,N_24370);
nor U28070 (N_28070,N_20923,N_22843);
and U28071 (N_28071,N_21770,N_23392);
or U28072 (N_28072,N_20611,N_21447);
and U28073 (N_28073,N_21219,N_21852);
and U28074 (N_28074,N_21626,N_23508);
xor U28075 (N_28075,N_22985,N_22298);
nand U28076 (N_28076,N_23865,N_22588);
or U28077 (N_28077,N_20616,N_21878);
xnor U28078 (N_28078,N_24503,N_24645);
or U28079 (N_28079,N_22233,N_21080);
and U28080 (N_28080,N_24905,N_21848);
xor U28081 (N_28081,N_22866,N_22903);
and U28082 (N_28082,N_20706,N_22218);
nand U28083 (N_28083,N_23559,N_22215);
nor U28084 (N_28084,N_22024,N_21272);
nand U28085 (N_28085,N_22870,N_21847);
or U28086 (N_28086,N_20130,N_21206);
nor U28087 (N_28087,N_21087,N_24254);
and U28088 (N_28088,N_23112,N_24380);
xor U28089 (N_28089,N_21237,N_20322);
or U28090 (N_28090,N_24964,N_23272);
xor U28091 (N_28091,N_20687,N_24458);
xnor U28092 (N_28092,N_24070,N_20902);
and U28093 (N_28093,N_23220,N_22969);
nor U28094 (N_28094,N_22444,N_21993);
nor U28095 (N_28095,N_22391,N_21105);
xor U28096 (N_28096,N_20189,N_20673);
nand U28097 (N_28097,N_24624,N_23701);
and U28098 (N_28098,N_20848,N_23993);
xnor U28099 (N_28099,N_20586,N_22048);
xnor U28100 (N_28100,N_21452,N_20041);
nor U28101 (N_28101,N_20454,N_22950);
and U28102 (N_28102,N_22156,N_22874);
nor U28103 (N_28103,N_20705,N_24480);
xor U28104 (N_28104,N_22514,N_22131);
nand U28105 (N_28105,N_24257,N_20120);
or U28106 (N_28106,N_21836,N_23740);
xor U28107 (N_28107,N_20838,N_21274);
nor U28108 (N_28108,N_24243,N_22441);
nor U28109 (N_28109,N_21923,N_22406);
or U28110 (N_28110,N_20779,N_21827);
or U28111 (N_28111,N_24204,N_22087);
or U28112 (N_28112,N_21155,N_23662);
nand U28113 (N_28113,N_24413,N_23241);
nor U28114 (N_28114,N_22051,N_20089);
or U28115 (N_28115,N_21575,N_20933);
xnor U28116 (N_28116,N_23775,N_21602);
and U28117 (N_28117,N_21628,N_20670);
nor U28118 (N_28118,N_23429,N_23778);
nor U28119 (N_28119,N_23823,N_20654);
and U28120 (N_28120,N_24166,N_24699);
nand U28121 (N_28121,N_23680,N_23545);
and U28122 (N_28122,N_23367,N_23021);
and U28123 (N_28123,N_20815,N_23186);
and U28124 (N_28124,N_22691,N_20985);
nor U28125 (N_28125,N_23624,N_22927);
or U28126 (N_28126,N_24743,N_24299);
and U28127 (N_28127,N_20199,N_22330);
nand U28128 (N_28128,N_20877,N_23812);
nand U28129 (N_28129,N_21618,N_22173);
and U28130 (N_28130,N_20329,N_20711);
or U28131 (N_28131,N_22252,N_24560);
nand U28132 (N_28132,N_23429,N_21926);
nor U28133 (N_28133,N_21395,N_23761);
or U28134 (N_28134,N_24029,N_21983);
nor U28135 (N_28135,N_22422,N_21494);
nand U28136 (N_28136,N_20615,N_20713);
nor U28137 (N_28137,N_23445,N_24927);
nand U28138 (N_28138,N_22008,N_21725);
xnor U28139 (N_28139,N_23058,N_22667);
nand U28140 (N_28140,N_23773,N_23948);
and U28141 (N_28141,N_20669,N_23062);
nand U28142 (N_28142,N_20333,N_24806);
and U28143 (N_28143,N_23759,N_21206);
or U28144 (N_28144,N_24036,N_24267);
nor U28145 (N_28145,N_22401,N_23801);
xnor U28146 (N_28146,N_22760,N_21278);
or U28147 (N_28147,N_24730,N_23427);
nand U28148 (N_28148,N_20531,N_22711);
or U28149 (N_28149,N_24269,N_21994);
and U28150 (N_28150,N_21517,N_23564);
nor U28151 (N_28151,N_20571,N_24545);
xor U28152 (N_28152,N_20154,N_20398);
nand U28153 (N_28153,N_22786,N_24234);
nand U28154 (N_28154,N_23214,N_24806);
and U28155 (N_28155,N_21389,N_23934);
nand U28156 (N_28156,N_20889,N_20475);
or U28157 (N_28157,N_21785,N_20072);
nand U28158 (N_28158,N_22502,N_22274);
and U28159 (N_28159,N_24322,N_21853);
nor U28160 (N_28160,N_20637,N_20099);
and U28161 (N_28161,N_23917,N_21530);
xor U28162 (N_28162,N_22914,N_21855);
nand U28163 (N_28163,N_21564,N_21154);
and U28164 (N_28164,N_20403,N_22295);
nand U28165 (N_28165,N_22317,N_21303);
nor U28166 (N_28166,N_24090,N_24453);
nor U28167 (N_28167,N_20812,N_21725);
xor U28168 (N_28168,N_23066,N_20089);
xor U28169 (N_28169,N_22271,N_22021);
nand U28170 (N_28170,N_21950,N_24817);
and U28171 (N_28171,N_24784,N_24365);
nand U28172 (N_28172,N_21095,N_22078);
nand U28173 (N_28173,N_21856,N_22216);
nand U28174 (N_28174,N_22677,N_21105);
or U28175 (N_28175,N_22653,N_23460);
and U28176 (N_28176,N_20281,N_22281);
and U28177 (N_28177,N_22388,N_21710);
nor U28178 (N_28178,N_24288,N_20447);
nor U28179 (N_28179,N_24301,N_23696);
or U28180 (N_28180,N_22897,N_21700);
nor U28181 (N_28181,N_20206,N_22432);
or U28182 (N_28182,N_24098,N_21055);
nand U28183 (N_28183,N_20013,N_21584);
xnor U28184 (N_28184,N_20311,N_21819);
or U28185 (N_28185,N_24651,N_23746);
nand U28186 (N_28186,N_24348,N_20780);
xor U28187 (N_28187,N_21252,N_23498);
or U28188 (N_28188,N_22306,N_24196);
xor U28189 (N_28189,N_20233,N_24823);
or U28190 (N_28190,N_24854,N_21573);
or U28191 (N_28191,N_22613,N_21225);
nand U28192 (N_28192,N_21770,N_22982);
and U28193 (N_28193,N_20122,N_22639);
and U28194 (N_28194,N_24654,N_24025);
nand U28195 (N_28195,N_23212,N_20649);
and U28196 (N_28196,N_24892,N_24004);
or U28197 (N_28197,N_22496,N_21772);
nand U28198 (N_28198,N_23089,N_20768);
nand U28199 (N_28199,N_22149,N_21942);
or U28200 (N_28200,N_20145,N_22983);
nand U28201 (N_28201,N_24691,N_22565);
or U28202 (N_28202,N_20252,N_21929);
nor U28203 (N_28203,N_22236,N_21865);
nand U28204 (N_28204,N_24519,N_21097);
and U28205 (N_28205,N_23575,N_24433);
nand U28206 (N_28206,N_21552,N_24223);
or U28207 (N_28207,N_22899,N_23965);
nand U28208 (N_28208,N_24815,N_24681);
or U28209 (N_28209,N_21333,N_24906);
and U28210 (N_28210,N_22763,N_20603);
xor U28211 (N_28211,N_23273,N_21381);
or U28212 (N_28212,N_24190,N_24263);
or U28213 (N_28213,N_21611,N_23030);
nor U28214 (N_28214,N_24481,N_24048);
nand U28215 (N_28215,N_23336,N_22132);
nor U28216 (N_28216,N_23408,N_22800);
xnor U28217 (N_28217,N_21483,N_20124);
nor U28218 (N_28218,N_20115,N_21252);
or U28219 (N_28219,N_21172,N_23995);
nor U28220 (N_28220,N_24929,N_21917);
xor U28221 (N_28221,N_23045,N_20802);
and U28222 (N_28222,N_23331,N_24075);
nand U28223 (N_28223,N_20365,N_21811);
or U28224 (N_28224,N_21145,N_20157);
xnor U28225 (N_28225,N_21169,N_20016);
or U28226 (N_28226,N_20388,N_23279);
nand U28227 (N_28227,N_21978,N_20211);
nor U28228 (N_28228,N_23820,N_22092);
nor U28229 (N_28229,N_23526,N_22435);
and U28230 (N_28230,N_21674,N_24931);
or U28231 (N_28231,N_20350,N_22070);
nor U28232 (N_28232,N_21195,N_23656);
nor U28233 (N_28233,N_23924,N_24850);
or U28234 (N_28234,N_20696,N_22376);
and U28235 (N_28235,N_20486,N_21981);
or U28236 (N_28236,N_24493,N_22198);
or U28237 (N_28237,N_20172,N_24436);
and U28238 (N_28238,N_22594,N_23296);
nand U28239 (N_28239,N_21145,N_23710);
or U28240 (N_28240,N_24210,N_20646);
xor U28241 (N_28241,N_20861,N_22092);
or U28242 (N_28242,N_22795,N_24168);
nand U28243 (N_28243,N_20457,N_23577);
xor U28244 (N_28244,N_23589,N_24618);
and U28245 (N_28245,N_23552,N_23208);
nand U28246 (N_28246,N_23628,N_24968);
xnor U28247 (N_28247,N_24944,N_21831);
nor U28248 (N_28248,N_23732,N_22353);
nand U28249 (N_28249,N_21714,N_21845);
and U28250 (N_28250,N_20578,N_21015);
nand U28251 (N_28251,N_22222,N_22604);
or U28252 (N_28252,N_21825,N_21738);
and U28253 (N_28253,N_23924,N_23691);
nand U28254 (N_28254,N_22077,N_23264);
nand U28255 (N_28255,N_22370,N_23443);
or U28256 (N_28256,N_23427,N_22929);
nor U28257 (N_28257,N_21090,N_20857);
or U28258 (N_28258,N_20381,N_21707);
nor U28259 (N_28259,N_20321,N_21771);
nand U28260 (N_28260,N_22166,N_21769);
nor U28261 (N_28261,N_21404,N_20819);
or U28262 (N_28262,N_22360,N_20067);
nand U28263 (N_28263,N_23706,N_21187);
and U28264 (N_28264,N_22302,N_20497);
nor U28265 (N_28265,N_24351,N_23338);
nand U28266 (N_28266,N_22636,N_20289);
or U28267 (N_28267,N_23773,N_24672);
nor U28268 (N_28268,N_20515,N_20715);
nor U28269 (N_28269,N_24312,N_23024);
nand U28270 (N_28270,N_24136,N_21601);
or U28271 (N_28271,N_21031,N_20930);
or U28272 (N_28272,N_21925,N_22150);
nand U28273 (N_28273,N_21934,N_24600);
nand U28274 (N_28274,N_22225,N_21925);
and U28275 (N_28275,N_23619,N_22389);
nand U28276 (N_28276,N_22772,N_22788);
nor U28277 (N_28277,N_23103,N_22787);
or U28278 (N_28278,N_20419,N_21395);
xor U28279 (N_28279,N_20128,N_22139);
and U28280 (N_28280,N_23529,N_20966);
or U28281 (N_28281,N_23648,N_24684);
nand U28282 (N_28282,N_22373,N_23097);
nor U28283 (N_28283,N_21133,N_22908);
nand U28284 (N_28284,N_21486,N_23927);
nand U28285 (N_28285,N_20387,N_22100);
nand U28286 (N_28286,N_23373,N_22029);
and U28287 (N_28287,N_22128,N_23291);
or U28288 (N_28288,N_23536,N_20272);
and U28289 (N_28289,N_22613,N_20800);
or U28290 (N_28290,N_20863,N_23371);
nand U28291 (N_28291,N_20214,N_23686);
nand U28292 (N_28292,N_23977,N_22716);
or U28293 (N_28293,N_23119,N_23232);
nor U28294 (N_28294,N_23551,N_21547);
nor U28295 (N_28295,N_23423,N_23753);
xnor U28296 (N_28296,N_23614,N_21340);
or U28297 (N_28297,N_22069,N_24759);
nand U28298 (N_28298,N_21578,N_24499);
and U28299 (N_28299,N_24958,N_22364);
nor U28300 (N_28300,N_20894,N_24781);
or U28301 (N_28301,N_21221,N_22608);
nor U28302 (N_28302,N_24014,N_21557);
or U28303 (N_28303,N_23729,N_24514);
or U28304 (N_28304,N_24800,N_22631);
nor U28305 (N_28305,N_23841,N_20987);
nand U28306 (N_28306,N_20457,N_21207);
nand U28307 (N_28307,N_20678,N_23433);
nor U28308 (N_28308,N_20663,N_20322);
and U28309 (N_28309,N_22980,N_21408);
nor U28310 (N_28310,N_22789,N_24218);
or U28311 (N_28311,N_22985,N_23117);
nor U28312 (N_28312,N_23594,N_22030);
or U28313 (N_28313,N_21893,N_24010);
xnor U28314 (N_28314,N_20242,N_23928);
nand U28315 (N_28315,N_21102,N_21144);
or U28316 (N_28316,N_23274,N_23306);
nand U28317 (N_28317,N_23518,N_21451);
nand U28318 (N_28318,N_24009,N_21597);
and U28319 (N_28319,N_21508,N_21651);
nand U28320 (N_28320,N_20994,N_21955);
or U28321 (N_28321,N_21523,N_21061);
nand U28322 (N_28322,N_23996,N_24856);
nand U28323 (N_28323,N_23018,N_24795);
nor U28324 (N_28324,N_21546,N_20445);
nor U28325 (N_28325,N_23171,N_20645);
xor U28326 (N_28326,N_20527,N_20749);
xnor U28327 (N_28327,N_23374,N_22433);
or U28328 (N_28328,N_24101,N_24564);
and U28329 (N_28329,N_22408,N_20517);
and U28330 (N_28330,N_24864,N_24227);
and U28331 (N_28331,N_22341,N_20467);
nor U28332 (N_28332,N_22085,N_21185);
xor U28333 (N_28333,N_23844,N_20608);
nor U28334 (N_28334,N_22363,N_20120);
nor U28335 (N_28335,N_21208,N_22641);
or U28336 (N_28336,N_24281,N_21148);
or U28337 (N_28337,N_24187,N_20447);
xnor U28338 (N_28338,N_23811,N_24393);
and U28339 (N_28339,N_21798,N_24152);
xnor U28340 (N_28340,N_24140,N_24311);
nor U28341 (N_28341,N_24790,N_21834);
nor U28342 (N_28342,N_21050,N_24149);
nor U28343 (N_28343,N_23957,N_24046);
nand U28344 (N_28344,N_21735,N_22543);
or U28345 (N_28345,N_24152,N_21714);
or U28346 (N_28346,N_24866,N_22530);
nand U28347 (N_28347,N_24584,N_20383);
xor U28348 (N_28348,N_24767,N_20493);
nor U28349 (N_28349,N_21853,N_20739);
nand U28350 (N_28350,N_20837,N_24180);
xnor U28351 (N_28351,N_23014,N_22778);
nand U28352 (N_28352,N_22204,N_23905);
or U28353 (N_28353,N_22437,N_23846);
xor U28354 (N_28354,N_21600,N_23812);
nor U28355 (N_28355,N_22056,N_22932);
nor U28356 (N_28356,N_22959,N_23669);
xor U28357 (N_28357,N_22035,N_24974);
nand U28358 (N_28358,N_21338,N_20210);
nor U28359 (N_28359,N_21613,N_22548);
nor U28360 (N_28360,N_21563,N_24909);
nor U28361 (N_28361,N_24877,N_23042);
or U28362 (N_28362,N_22349,N_23408);
and U28363 (N_28363,N_24354,N_22104);
nor U28364 (N_28364,N_24183,N_21884);
and U28365 (N_28365,N_23072,N_20833);
nand U28366 (N_28366,N_21054,N_22559);
nor U28367 (N_28367,N_24482,N_20389);
nand U28368 (N_28368,N_20157,N_24720);
or U28369 (N_28369,N_20878,N_21342);
nor U28370 (N_28370,N_21709,N_21361);
nor U28371 (N_28371,N_20260,N_23273);
and U28372 (N_28372,N_21482,N_22278);
and U28373 (N_28373,N_20958,N_22851);
nand U28374 (N_28374,N_24858,N_23719);
or U28375 (N_28375,N_21693,N_24878);
and U28376 (N_28376,N_20227,N_24035);
nor U28377 (N_28377,N_24082,N_22132);
and U28378 (N_28378,N_22945,N_23104);
or U28379 (N_28379,N_22531,N_21974);
or U28380 (N_28380,N_23318,N_20526);
or U28381 (N_28381,N_20625,N_20411);
nand U28382 (N_28382,N_21506,N_20973);
and U28383 (N_28383,N_24444,N_23595);
xor U28384 (N_28384,N_23838,N_23844);
and U28385 (N_28385,N_22870,N_22230);
or U28386 (N_28386,N_21814,N_20737);
nand U28387 (N_28387,N_24545,N_23639);
nand U28388 (N_28388,N_23544,N_20322);
nor U28389 (N_28389,N_24966,N_23399);
nand U28390 (N_28390,N_23130,N_20943);
nor U28391 (N_28391,N_23917,N_21230);
and U28392 (N_28392,N_23798,N_23355);
or U28393 (N_28393,N_24113,N_24155);
and U28394 (N_28394,N_20032,N_24485);
nor U28395 (N_28395,N_22056,N_20179);
nand U28396 (N_28396,N_24126,N_21726);
and U28397 (N_28397,N_23469,N_24130);
or U28398 (N_28398,N_21768,N_22076);
nand U28399 (N_28399,N_22060,N_24657);
or U28400 (N_28400,N_23979,N_23028);
or U28401 (N_28401,N_24337,N_22134);
and U28402 (N_28402,N_22103,N_21919);
nor U28403 (N_28403,N_22344,N_21825);
and U28404 (N_28404,N_20593,N_24041);
or U28405 (N_28405,N_20376,N_21846);
nand U28406 (N_28406,N_20935,N_24411);
nor U28407 (N_28407,N_24769,N_22454);
or U28408 (N_28408,N_22486,N_21045);
xnor U28409 (N_28409,N_24666,N_22898);
or U28410 (N_28410,N_21613,N_20589);
or U28411 (N_28411,N_20623,N_22943);
nor U28412 (N_28412,N_22521,N_23755);
nand U28413 (N_28413,N_23213,N_22741);
and U28414 (N_28414,N_24243,N_21739);
xnor U28415 (N_28415,N_22232,N_20355);
and U28416 (N_28416,N_23161,N_23617);
and U28417 (N_28417,N_21881,N_22809);
nor U28418 (N_28418,N_20858,N_22505);
xor U28419 (N_28419,N_24082,N_24456);
or U28420 (N_28420,N_22162,N_24504);
nand U28421 (N_28421,N_24746,N_22314);
nor U28422 (N_28422,N_22227,N_23678);
or U28423 (N_28423,N_20184,N_22204);
xor U28424 (N_28424,N_20513,N_23468);
xnor U28425 (N_28425,N_23149,N_22314);
or U28426 (N_28426,N_23492,N_22586);
nor U28427 (N_28427,N_20490,N_24706);
xnor U28428 (N_28428,N_20600,N_23158);
or U28429 (N_28429,N_21851,N_22018);
or U28430 (N_28430,N_24842,N_22870);
nand U28431 (N_28431,N_23347,N_21075);
xnor U28432 (N_28432,N_22887,N_21957);
or U28433 (N_28433,N_22413,N_24511);
nor U28434 (N_28434,N_20687,N_22405);
nor U28435 (N_28435,N_24522,N_21256);
nand U28436 (N_28436,N_21072,N_20705);
nor U28437 (N_28437,N_20871,N_24111);
or U28438 (N_28438,N_22334,N_20924);
nand U28439 (N_28439,N_20448,N_22719);
or U28440 (N_28440,N_21293,N_20800);
or U28441 (N_28441,N_23155,N_22341);
nand U28442 (N_28442,N_24555,N_21826);
xor U28443 (N_28443,N_24396,N_21713);
and U28444 (N_28444,N_24669,N_22263);
nand U28445 (N_28445,N_24993,N_20233);
nor U28446 (N_28446,N_22293,N_23750);
and U28447 (N_28447,N_24661,N_20873);
nand U28448 (N_28448,N_21800,N_23298);
xor U28449 (N_28449,N_21233,N_23667);
or U28450 (N_28450,N_23647,N_22869);
nor U28451 (N_28451,N_22895,N_21508);
xor U28452 (N_28452,N_24263,N_24311);
xor U28453 (N_28453,N_23135,N_21112);
and U28454 (N_28454,N_20451,N_24918);
nand U28455 (N_28455,N_23149,N_22477);
or U28456 (N_28456,N_20256,N_21347);
nand U28457 (N_28457,N_21634,N_23479);
nor U28458 (N_28458,N_22545,N_22872);
or U28459 (N_28459,N_24903,N_21073);
nand U28460 (N_28460,N_20420,N_22738);
xor U28461 (N_28461,N_23584,N_24266);
nor U28462 (N_28462,N_21070,N_22279);
xor U28463 (N_28463,N_23078,N_24872);
nor U28464 (N_28464,N_20179,N_21805);
nand U28465 (N_28465,N_23935,N_23232);
and U28466 (N_28466,N_24672,N_23914);
nor U28467 (N_28467,N_23034,N_23484);
nand U28468 (N_28468,N_24358,N_22715);
or U28469 (N_28469,N_22009,N_21776);
or U28470 (N_28470,N_21326,N_20931);
or U28471 (N_28471,N_23765,N_23829);
nand U28472 (N_28472,N_20259,N_24852);
and U28473 (N_28473,N_24658,N_23710);
or U28474 (N_28474,N_21137,N_24182);
xnor U28475 (N_28475,N_20301,N_23781);
nand U28476 (N_28476,N_24756,N_24146);
and U28477 (N_28477,N_23806,N_21286);
nor U28478 (N_28478,N_24340,N_22628);
and U28479 (N_28479,N_20886,N_24118);
and U28480 (N_28480,N_23405,N_23436);
nor U28481 (N_28481,N_24029,N_24397);
xnor U28482 (N_28482,N_24225,N_23103);
nand U28483 (N_28483,N_20946,N_20596);
or U28484 (N_28484,N_22893,N_21990);
nand U28485 (N_28485,N_20735,N_24130);
and U28486 (N_28486,N_24454,N_21831);
nor U28487 (N_28487,N_23957,N_22348);
nand U28488 (N_28488,N_20481,N_23005);
nand U28489 (N_28489,N_20023,N_20928);
and U28490 (N_28490,N_24368,N_20272);
and U28491 (N_28491,N_22106,N_24135);
and U28492 (N_28492,N_20950,N_23404);
and U28493 (N_28493,N_20238,N_23984);
nand U28494 (N_28494,N_21538,N_23727);
xnor U28495 (N_28495,N_23860,N_21462);
or U28496 (N_28496,N_23313,N_24824);
nor U28497 (N_28497,N_22201,N_21752);
nand U28498 (N_28498,N_21591,N_23543);
nor U28499 (N_28499,N_20984,N_21627);
nor U28500 (N_28500,N_20701,N_22908);
or U28501 (N_28501,N_22986,N_20993);
nand U28502 (N_28502,N_24884,N_20581);
xnor U28503 (N_28503,N_21409,N_23904);
and U28504 (N_28504,N_23639,N_24499);
or U28505 (N_28505,N_24882,N_24994);
nand U28506 (N_28506,N_24851,N_21533);
nor U28507 (N_28507,N_24971,N_24615);
nor U28508 (N_28508,N_20115,N_24999);
or U28509 (N_28509,N_22901,N_21294);
nand U28510 (N_28510,N_24959,N_21516);
or U28511 (N_28511,N_24490,N_20181);
or U28512 (N_28512,N_21055,N_21773);
or U28513 (N_28513,N_24810,N_22724);
and U28514 (N_28514,N_21239,N_22780);
and U28515 (N_28515,N_22492,N_24574);
nand U28516 (N_28516,N_23197,N_23075);
nor U28517 (N_28517,N_22204,N_23129);
and U28518 (N_28518,N_23540,N_24373);
and U28519 (N_28519,N_20845,N_20251);
and U28520 (N_28520,N_21847,N_23966);
nor U28521 (N_28521,N_23845,N_23337);
or U28522 (N_28522,N_21621,N_20340);
or U28523 (N_28523,N_23880,N_23989);
or U28524 (N_28524,N_22743,N_20547);
or U28525 (N_28525,N_21263,N_20344);
and U28526 (N_28526,N_20470,N_21201);
nand U28527 (N_28527,N_22914,N_21183);
or U28528 (N_28528,N_21472,N_21720);
and U28529 (N_28529,N_24898,N_24094);
or U28530 (N_28530,N_24891,N_22174);
nor U28531 (N_28531,N_22162,N_23347);
or U28532 (N_28532,N_21724,N_22336);
or U28533 (N_28533,N_24029,N_20244);
nand U28534 (N_28534,N_23872,N_22283);
and U28535 (N_28535,N_23935,N_23007);
xor U28536 (N_28536,N_21178,N_21383);
or U28537 (N_28537,N_22907,N_24171);
nor U28538 (N_28538,N_22549,N_24555);
nand U28539 (N_28539,N_23882,N_22998);
nand U28540 (N_28540,N_21483,N_22733);
and U28541 (N_28541,N_24320,N_22259);
and U28542 (N_28542,N_21953,N_20658);
nor U28543 (N_28543,N_20299,N_23829);
nand U28544 (N_28544,N_20504,N_20714);
or U28545 (N_28545,N_22105,N_21641);
nor U28546 (N_28546,N_24092,N_21781);
or U28547 (N_28547,N_22860,N_24911);
nand U28548 (N_28548,N_23303,N_23598);
xor U28549 (N_28549,N_23612,N_22066);
nor U28550 (N_28550,N_24774,N_21994);
xnor U28551 (N_28551,N_20515,N_22100);
nand U28552 (N_28552,N_22892,N_21781);
and U28553 (N_28553,N_21855,N_21245);
or U28554 (N_28554,N_23210,N_22429);
and U28555 (N_28555,N_24953,N_23518);
nand U28556 (N_28556,N_20251,N_23605);
nor U28557 (N_28557,N_21130,N_23188);
nand U28558 (N_28558,N_23000,N_24678);
nand U28559 (N_28559,N_23950,N_21964);
nor U28560 (N_28560,N_23021,N_22196);
nand U28561 (N_28561,N_20201,N_24594);
nand U28562 (N_28562,N_23550,N_24845);
and U28563 (N_28563,N_23602,N_22502);
nand U28564 (N_28564,N_21864,N_23825);
or U28565 (N_28565,N_20838,N_24398);
and U28566 (N_28566,N_24000,N_22160);
nand U28567 (N_28567,N_22193,N_22063);
nor U28568 (N_28568,N_23767,N_23047);
xor U28569 (N_28569,N_24233,N_22478);
nor U28570 (N_28570,N_23519,N_23172);
xnor U28571 (N_28571,N_24237,N_24146);
and U28572 (N_28572,N_22222,N_23202);
and U28573 (N_28573,N_21714,N_21226);
and U28574 (N_28574,N_22380,N_20213);
or U28575 (N_28575,N_21319,N_20640);
nor U28576 (N_28576,N_23515,N_23918);
and U28577 (N_28577,N_20373,N_23862);
nor U28578 (N_28578,N_20623,N_24868);
or U28579 (N_28579,N_22609,N_21257);
or U28580 (N_28580,N_20255,N_23994);
or U28581 (N_28581,N_23809,N_23238);
or U28582 (N_28582,N_21545,N_20483);
and U28583 (N_28583,N_20781,N_23136);
nand U28584 (N_28584,N_21242,N_21283);
nand U28585 (N_28585,N_24094,N_24537);
and U28586 (N_28586,N_22928,N_21272);
and U28587 (N_28587,N_24346,N_23724);
nand U28588 (N_28588,N_24874,N_20037);
and U28589 (N_28589,N_23544,N_23582);
xnor U28590 (N_28590,N_20652,N_23575);
nor U28591 (N_28591,N_23050,N_21090);
nor U28592 (N_28592,N_21394,N_23864);
nor U28593 (N_28593,N_22219,N_20801);
or U28594 (N_28594,N_22351,N_24554);
xnor U28595 (N_28595,N_22386,N_22985);
and U28596 (N_28596,N_24323,N_23994);
and U28597 (N_28597,N_24679,N_21569);
or U28598 (N_28598,N_21804,N_24279);
xor U28599 (N_28599,N_23213,N_22600);
or U28600 (N_28600,N_21376,N_20269);
xnor U28601 (N_28601,N_22656,N_24325);
or U28602 (N_28602,N_21910,N_23499);
xnor U28603 (N_28603,N_20284,N_24727);
nor U28604 (N_28604,N_20864,N_21114);
nor U28605 (N_28605,N_20667,N_20465);
nand U28606 (N_28606,N_21524,N_20402);
and U28607 (N_28607,N_23849,N_20716);
xor U28608 (N_28608,N_23858,N_22877);
nor U28609 (N_28609,N_20151,N_21499);
and U28610 (N_28610,N_20230,N_20192);
and U28611 (N_28611,N_23451,N_21684);
or U28612 (N_28612,N_20169,N_21989);
or U28613 (N_28613,N_21234,N_24423);
or U28614 (N_28614,N_21922,N_20282);
and U28615 (N_28615,N_24676,N_23352);
and U28616 (N_28616,N_21821,N_23745);
nor U28617 (N_28617,N_21518,N_21380);
and U28618 (N_28618,N_21110,N_20826);
nor U28619 (N_28619,N_23139,N_24848);
xnor U28620 (N_28620,N_24346,N_24900);
or U28621 (N_28621,N_21872,N_21906);
or U28622 (N_28622,N_21549,N_23479);
nor U28623 (N_28623,N_22799,N_20080);
and U28624 (N_28624,N_24714,N_21822);
and U28625 (N_28625,N_23867,N_22433);
and U28626 (N_28626,N_22554,N_22199);
or U28627 (N_28627,N_23703,N_23699);
nand U28628 (N_28628,N_24573,N_23417);
nor U28629 (N_28629,N_23697,N_20581);
nand U28630 (N_28630,N_21374,N_20529);
xnor U28631 (N_28631,N_23972,N_23949);
or U28632 (N_28632,N_22427,N_22714);
and U28633 (N_28633,N_23221,N_22116);
nor U28634 (N_28634,N_22749,N_23508);
xnor U28635 (N_28635,N_22662,N_23121);
and U28636 (N_28636,N_21308,N_21620);
and U28637 (N_28637,N_20235,N_22096);
or U28638 (N_28638,N_22438,N_22150);
nor U28639 (N_28639,N_22941,N_22992);
xor U28640 (N_28640,N_24603,N_20478);
or U28641 (N_28641,N_24083,N_23120);
or U28642 (N_28642,N_20907,N_21417);
and U28643 (N_28643,N_22378,N_21268);
or U28644 (N_28644,N_21790,N_21377);
nand U28645 (N_28645,N_22037,N_20635);
nand U28646 (N_28646,N_20359,N_22193);
nand U28647 (N_28647,N_21979,N_23397);
and U28648 (N_28648,N_24741,N_21897);
and U28649 (N_28649,N_22114,N_21008);
nand U28650 (N_28650,N_20611,N_24329);
or U28651 (N_28651,N_22092,N_21475);
nor U28652 (N_28652,N_20531,N_24056);
nor U28653 (N_28653,N_21916,N_21579);
and U28654 (N_28654,N_24670,N_22467);
and U28655 (N_28655,N_23557,N_20222);
nor U28656 (N_28656,N_24341,N_23060);
xor U28657 (N_28657,N_20178,N_22695);
xor U28658 (N_28658,N_23027,N_23606);
or U28659 (N_28659,N_20352,N_21872);
and U28660 (N_28660,N_20607,N_21575);
or U28661 (N_28661,N_20174,N_21930);
and U28662 (N_28662,N_22300,N_21568);
or U28663 (N_28663,N_24367,N_22779);
and U28664 (N_28664,N_21099,N_20924);
and U28665 (N_28665,N_24720,N_22553);
xnor U28666 (N_28666,N_24560,N_20804);
nor U28667 (N_28667,N_20213,N_23418);
nand U28668 (N_28668,N_20605,N_21421);
and U28669 (N_28669,N_20274,N_20211);
nand U28670 (N_28670,N_23887,N_21448);
xnor U28671 (N_28671,N_23697,N_22688);
or U28672 (N_28672,N_23279,N_21023);
and U28673 (N_28673,N_22393,N_21749);
and U28674 (N_28674,N_23346,N_23356);
nand U28675 (N_28675,N_20506,N_23235);
and U28676 (N_28676,N_21386,N_20092);
or U28677 (N_28677,N_22388,N_24631);
xor U28678 (N_28678,N_21456,N_21097);
or U28679 (N_28679,N_23518,N_20119);
nor U28680 (N_28680,N_20391,N_24116);
and U28681 (N_28681,N_22393,N_21397);
or U28682 (N_28682,N_20732,N_24949);
or U28683 (N_28683,N_20191,N_21849);
xnor U28684 (N_28684,N_21664,N_22481);
xnor U28685 (N_28685,N_21304,N_22248);
xnor U28686 (N_28686,N_20388,N_24489);
nand U28687 (N_28687,N_21520,N_22342);
and U28688 (N_28688,N_21724,N_23972);
nand U28689 (N_28689,N_23177,N_23256);
nor U28690 (N_28690,N_24674,N_22400);
and U28691 (N_28691,N_20445,N_23926);
and U28692 (N_28692,N_24135,N_24764);
nor U28693 (N_28693,N_21178,N_21353);
xor U28694 (N_28694,N_23075,N_23563);
nand U28695 (N_28695,N_23995,N_23903);
or U28696 (N_28696,N_22189,N_23687);
and U28697 (N_28697,N_23945,N_21385);
nor U28698 (N_28698,N_20000,N_24878);
nand U28699 (N_28699,N_23439,N_22531);
or U28700 (N_28700,N_20154,N_24242);
or U28701 (N_28701,N_21351,N_24508);
nand U28702 (N_28702,N_23367,N_24146);
xor U28703 (N_28703,N_21380,N_22669);
nor U28704 (N_28704,N_21082,N_23427);
or U28705 (N_28705,N_24174,N_24526);
nand U28706 (N_28706,N_23089,N_23684);
and U28707 (N_28707,N_24709,N_22633);
or U28708 (N_28708,N_24092,N_24039);
or U28709 (N_28709,N_23145,N_23372);
nand U28710 (N_28710,N_23600,N_22899);
and U28711 (N_28711,N_23292,N_23096);
nand U28712 (N_28712,N_24882,N_21372);
nor U28713 (N_28713,N_24223,N_23884);
xnor U28714 (N_28714,N_22381,N_23145);
nand U28715 (N_28715,N_21198,N_24484);
xor U28716 (N_28716,N_24398,N_22947);
or U28717 (N_28717,N_22984,N_20116);
and U28718 (N_28718,N_21184,N_22680);
or U28719 (N_28719,N_22467,N_20139);
nor U28720 (N_28720,N_24195,N_22804);
or U28721 (N_28721,N_22382,N_20091);
and U28722 (N_28722,N_21666,N_20876);
nand U28723 (N_28723,N_21600,N_21856);
nand U28724 (N_28724,N_24596,N_24364);
or U28725 (N_28725,N_20336,N_21272);
nor U28726 (N_28726,N_20521,N_22346);
or U28727 (N_28727,N_24657,N_20675);
and U28728 (N_28728,N_21719,N_20902);
and U28729 (N_28729,N_22286,N_24726);
or U28730 (N_28730,N_20498,N_20118);
nand U28731 (N_28731,N_22185,N_20658);
or U28732 (N_28732,N_23550,N_20531);
nand U28733 (N_28733,N_21903,N_23322);
or U28734 (N_28734,N_20659,N_24292);
nor U28735 (N_28735,N_20310,N_20726);
or U28736 (N_28736,N_23296,N_22786);
and U28737 (N_28737,N_20618,N_20596);
nand U28738 (N_28738,N_23788,N_20184);
and U28739 (N_28739,N_20786,N_20354);
or U28740 (N_28740,N_24462,N_23814);
nor U28741 (N_28741,N_21744,N_21498);
xnor U28742 (N_28742,N_22460,N_22469);
and U28743 (N_28743,N_21382,N_24078);
nand U28744 (N_28744,N_21249,N_23457);
nor U28745 (N_28745,N_23590,N_22239);
nand U28746 (N_28746,N_21041,N_21562);
nor U28747 (N_28747,N_24562,N_20907);
xor U28748 (N_28748,N_23447,N_21940);
nor U28749 (N_28749,N_23282,N_21905);
nand U28750 (N_28750,N_24783,N_21591);
or U28751 (N_28751,N_24543,N_22487);
nand U28752 (N_28752,N_23893,N_21292);
or U28753 (N_28753,N_23503,N_21334);
nor U28754 (N_28754,N_21740,N_22230);
nand U28755 (N_28755,N_22306,N_21613);
and U28756 (N_28756,N_23650,N_23063);
nor U28757 (N_28757,N_21550,N_22458);
and U28758 (N_28758,N_23885,N_24650);
and U28759 (N_28759,N_21356,N_23329);
nand U28760 (N_28760,N_24919,N_21273);
or U28761 (N_28761,N_24379,N_23029);
or U28762 (N_28762,N_24206,N_23062);
nand U28763 (N_28763,N_20115,N_23625);
and U28764 (N_28764,N_24373,N_20126);
and U28765 (N_28765,N_21623,N_24354);
and U28766 (N_28766,N_24375,N_23537);
and U28767 (N_28767,N_22957,N_24281);
nand U28768 (N_28768,N_23127,N_23122);
nor U28769 (N_28769,N_22192,N_22628);
nand U28770 (N_28770,N_22219,N_23630);
nand U28771 (N_28771,N_23653,N_24885);
nor U28772 (N_28772,N_20920,N_22384);
and U28773 (N_28773,N_21441,N_23138);
nor U28774 (N_28774,N_24282,N_24813);
nor U28775 (N_28775,N_20873,N_23937);
nor U28776 (N_28776,N_21759,N_23976);
and U28777 (N_28777,N_24372,N_21318);
and U28778 (N_28778,N_23065,N_24166);
and U28779 (N_28779,N_21912,N_24872);
or U28780 (N_28780,N_20185,N_20541);
xnor U28781 (N_28781,N_22281,N_22522);
or U28782 (N_28782,N_22684,N_20717);
nand U28783 (N_28783,N_20007,N_23565);
or U28784 (N_28784,N_23898,N_23089);
nor U28785 (N_28785,N_21350,N_23480);
or U28786 (N_28786,N_23269,N_20121);
or U28787 (N_28787,N_20256,N_20198);
and U28788 (N_28788,N_21926,N_20795);
nor U28789 (N_28789,N_23835,N_23507);
or U28790 (N_28790,N_22623,N_21252);
nor U28791 (N_28791,N_20587,N_24051);
nand U28792 (N_28792,N_23969,N_20974);
nand U28793 (N_28793,N_23192,N_24630);
and U28794 (N_28794,N_24741,N_22726);
or U28795 (N_28795,N_22856,N_24201);
xor U28796 (N_28796,N_22756,N_23524);
nand U28797 (N_28797,N_21664,N_22904);
nor U28798 (N_28798,N_24188,N_21479);
or U28799 (N_28799,N_22179,N_24303);
nand U28800 (N_28800,N_21823,N_22204);
nand U28801 (N_28801,N_21133,N_20168);
and U28802 (N_28802,N_23165,N_22417);
nor U28803 (N_28803,N_23783,N_24229);
and U28804 (N_28804,N_23017,N_21728);
and U28805 (N_28805,N_24973,N_24006);
xor U28806 (N_28806,N_20016,N_20497);
nand U28807 (N_28807,N_21564,N_24443);
and U28808 (N_28808,N_23857,N_20161);
nand U28809 (N_28809,N_24270,N_20298);
nor U28810 (N_28810,N_21139,N_21531);
nor U28811 (N_28811,N_22761,N_21642);
xor U28812 (N_28812,N_20028,N_24236);
or U28813 (N_28813,N_22089,N_20230);
and U28814 (N_28814,N_20644,N_23820);
or U28815 (N_28815,N_23861,N_20959);
nor U28816 (N_28816,N_21971,N_23440);
or U28817 (N_28817,N_23057,N_24903);
and U28818 (N_28818,N_22089,N_20619);
xnor U28819 (N_28819,N_22490,N_20321);
and U28820 (N_28820,N_22113,N_24602);
xnor U28821 (N_28821,N_21708,N_23950);
or U28822 (N_28822,N_20368,N_21051);
nand U28823 (N_28823,N_21489,N_22819);
nand U28824 (N_28824,N_23277,N_23759);
and U28825 (N_28825,N_22816,N_21914);
nor U28826 (N_28826,N_24533,N_22646);
or U28827 (N_28827,N_20252,N_20598);
nor U28828 (N_28828,N_24018,N_20908);
nand U28829 (N_28829,N_24322,N_20388);
or U28830 (N_28830,N_24185,N_20253);
or U28831 (N_28831,N_22533,N_22917);
xor U28832 (N_28832,N_24287,N_21341);
and U28833 (N_28833,N_20305,N_21125);
nor U28834 (N_28834,N_24763,N_22305);
nor U28835 (N_28835,N_20977,N_22387);
or U28836 (N_28836,N_24525,N_20074);
or U28837 (N_28837,N_23069,N_22280);
or U28838 (N_28838,N_24073,N_24588);
nor U28839 (N_28839,N_23796,N_20344);
and U28840 (N_28840,N_24111,N_23854);
and U28841 (N_28841,N_24912,N_22101);
nor U28842 (N_28842,N_24722,N_21923);
and U28843 (N_28843,N_22475,N_23091);
xor U28844 (N_28844,N_20630,N_20749);
and U28845 (N_28845,N_21426,N_22471);
nor U28846 (N_28846,N_22643,N_24599);
nand U28847 (N_28847,N_22179,N_24181);
or U28848 (N_28848,N_20348,N_24430);
xnor U28849 (N_28849,N_24906,N_23931);
nand U28850 (N_28850,N_20841,N_24640);
nand U28851 (N_28851,N_24580,N_22326);
or U28852 (N_28852,N_22883,N_22327);
nor U28853 (N_28853,N_22381,N_20336);
or U28854 (N_28854,N_21199,N_21153);
nand U28855 (N_28855,N_21210,N_24476);
or U28856 (N_28856,N_20911,N_20850);
nand U28857 (N_28857,N_20425,N_20295);
nand U28858 (N_28858,N_24480,N_20173);
nor U28859 (N_28859,N_23077,N_21636);
nor U28860 (N_28860,N_24985,N_24859);
nor U28861 (N_28861,N_22725,N_24761);
and U28862 (N_28862,N_22065,N_21040);
nand U28863 (N_28863,N_24343,N_24264);
and U28864 (N_28864,N_20690,N_24182);
nand U28865 (N_28865,N_22698,N_23334);
nand U28866 (N_28866,N_20923,N_23559);
nand U28867 (N_28867,N_23270,N_21744);
and U28868 (N_28868,N_21358,N_24382);
nand U28869 (N_28869,N_20570,N_24582);
or U28870 (N_28870,N_23665,N_22133);
nand U28871 (N_28871,N_20156,N_20124);
and U28872 (N_28872,N_23793,N_20072);
nor U28873 (N_28873,N_21148,N_22187);
nor U28874 (N_28874,N_22851,N_24295);
or U28875 (N_28875,N_21854,N_20950);
nor U28876 (N_28876,N_23878,N_23064);
or U28877 (N_28877,N_21684,N_22653);
nand U28878 (N_28878,N_20720,N_24092);
nand U28879 (N_28879,N_24808,N_20971);
or U28880 (N_28880,N_22164,N_24487);
and U28881 (N_28881,N_21400,N_20478);
nor U28882 (N_28882,N_24399,N_21398);
and U28883 (N_28883,N_22077,N_22631);
and U28884 (N_28884,N_22234,N_20943);
xor U28885 (N_28885,N_20420,N_22187);
nor U28886 (N_28886,N_22001,N_24908);
xnor U28887 (N_28887,N_21401,N_23712);
nand U28888 (N_28888,N_22884,N_23431);
or U28889 (N_28889,N_21701,N_20570);
and U28890 (N_28890,N_24704,N_23251);
nor U28891 (N_28891,N_22728,N_24877);
and U28892 (N_28892,N_21198,N_24460);
xnor U28893 (N_28893,N_24447,N_21427);
and U28894 (N_28894,N_22625,N_20484);
nor U28895 (N_28895,N_23847,N_21046);
and U28896 (N_28896,N_23611,N_22706);
nor U28897 (N_28897,N_23006,N_21857);
or U28898 (N_28898,N_23828,N_20135);
and U28899 (N_28899,N_23753,N_24081);
nand U28900 (N_28900,N_22206,N_23896);
nor U28901 (N_28901,N_23918,N_24636);
or U28902 (N_28902,N_21221,N_23058);
or U28903 (N_28903,N_22832,N_20351);
nor U28904 (N_28904,N_20856,N_24659);
nor U28905 (N_28905,N_21674,N_21772);
and U28906 (N_28906,N_22353,N_23574);
nand U28907 (N_28907,N_24273,N_24284);
nand U28908 (N_28908,N_22573,N_21085);
or U28909 (N_28909,N_22509,N_23017);
or U28910 (N_28910,N_23064,N_24022);
or U28911 (N_28911,N_20483,N_22331);
nor U28912 (N_28912,N_24136,N_21742);
nor U28913 (N_28913,N_24812,N_22439);
and U28914 (N_28914,N_20523,N_20051);
nor U28915 (N_28915,N_20937,N_24835);
xnor U28916 (N_28916,N_23036,N_22081);
nand U28917 (N_28917,N_21666,N_23860);
nand U28918 (N_28918,N_22028,N_21901);
or U28919 (N_28919,N_24859,N_20495);
and U28920 (N_28920,N_23993,N_22057);
and U28921 (N_28921,N_22129,N_24252);
and U28922 (N_28922,N_23369,N_21095);
and U28923 (N_28923,N_20942,N_23472);
and U28924 (N_28924,N_21072,N_22352);
nand U28925 (N_28925,N_24278,N_22714);
nand U28926 (N_28926,N_22016,N_22836);
nand U28927 (N_28927,N_24237,N_20910);
xor U28928 (N_28928,N_21052,N_21021);
or U28929 (N_28929,N_22762,N_23483);
nor U28930 (N_28930,N_23748,N_22934);
and U28931 (N_28931,N_22771,N_22681);
or U28932 (N_28932,N_22343,N_20303);
or U28933 (N_28933,N_24467,N_23983);
xor U28934 (N_28934,N_20639,N_22795);
nor U28935 (N_28935,N_20894,N_23917);
and U28936 (N_28936,N_20692,N_24642);
nand U28937 (N_28937,N_21675,N_21012);
nand U28938 (N_28938,N_23116,N_24832);
nand U28939 (N_28939,N_21758,N_20568);
or U28940 (N_28940,N_22609,N_20905);
nor U28941 (N_28941,N_20433,N_20769);
and U28942 (N_28942,N_21722,N_24526);
xor U28943 (N_28943,N_22064,N_24649);
and U28944 (N_28944,N_24366,N_24964);
or U28945 (N_28945,N_24746,N_21846);
xor U28946 (N_28946,N_22442,N_23358);
nor U28947 (N_28947,N_23282,N_23739);
nor U28948 (N_28948,N_24581,N_22736);
or U28949 (N_28949,N_20177,N_23262);
nand U28950 (N_28950,N_22830,N_24920);
nor U28951 (N_28951,N_22607,N_20602);
nand U28952 (N_28952,N_21514,N_23895);
or U28953 (N_28953,N_22397,N_23287);
and U28954 (N_28954,N_24228,N_24189);
xnor U28955 (N_28955,N_20349,N_24305);
and U28956 (N_28956,N_21488,N_20412);
nor U28957 (N_28957,N_24493,N_23499);
nand U28958 (N_28958,N_23014,N_20907);
nand U28959 (N_28959,N_24363,N_24650);
or U28960 (N_28960,N_24077,N_24277);
and U28961 (N_28961,N_20250,N_21099);
nor U28962 (N_28962,N_22170,N_24708);
or U28963 (N_28963,N_23839,N_22062);
nand U28964 (N_28964,N_21198,N_21275);
or U28965 (N_28965,N_24142,N_23994);
or U28966 (N_28966,N_21784,N_23864);
or U28967 (N_28967,N_22798,N_20698);
nand U28968 (N_28968,N_24034,N_21883);
nand U28969 (N_28969,N_23826,N_23589);
nor U28970 (N_28970,N_24421,N_21720);
nand U28971 (N_28971,N_24283,N_20795);
or U28972 (N_28972,N_20733,N_23005);
nor U28973 (N_28973,N_21450,N_22745);
or U28974 (N_28974,N_21959,N_21073);
and U28975 (N_28975,N_20723,N_20554);
nor U28976 (N_28976,N_22914,N_22910);
or U28977 (N_28977,N_21914,N_24867);
nor U28978 (N_28978,N_21470,N_20744);
xnor U28979 (N_28979,N_20328,N_22412);
xnor U28980 (N_28980,N_22458,N_23671);
nor U28981 (N_28981,N_22896,N_24166);
and U28982 (N_28982,N_24170,N_24790);
and U28983 (N_28983,N_22741,N_23159);
nor U28984 (N_28984,N_23470,N_21299);
or U28985 (N_28985,N_20595,N_24872);
and U28986 (N_28986,N_22170,N_23236);
nor U28987 (N_28987,N_24178,N_21116);
nand U28988 (N_28988,N_20900,N_24181);
nor U28989 (N_28989,N_22587,N_20620);
nor U28990 (N_28990,N_23877,N_22542);
nand U28991 (N_28991,N_22025,N_21837);
or U28992 (N_28992,N_21382,N_23371);
xnor U28993 (N_28993,N_20526,N_23454);
nand U28994 (N_28994,N_20734,N_24144);
and U28995 (N_28995,N_20606,N_21736);
and U28996 (N_28996,N_24996,N_23113);
or U28997 (N_28997,N_24003,N_20851);
nand U28998 (N_28998,N_22028,N_21135);
and U28999 (N_28999,N_23573,N_24403);
and U29000 (N_29000,N_22047,N_24888);
xor U29001 (N_29001,N_24605,N_24850);
or U29002 (N_29002,N_21378,N_24150);
or U29003 (N_29003,N_20536,N_22294);
and U29004 (N_29004,N_20506,N_21691);
xnor U29005 (N_29005,N_23520,N_21842);
or U29006 (N_29006,N_21783,N_24663);
or U29007 (N_29007,N_22534,N_21194);
and U29008 (N_29008,N_24004,N_23699);
nor U29009 (N_29009,N_20323,N_22041);
and U29010 (N_29010,N_23490,N_24824);
nor U29011 (N_29011,N_23732,N_24225);
nor U29012 (N_29012,N_24266,N_20311);
or U29013 (N_29013,N_21771,N_21469);
or U29014 (N_29014,N_23261,N_21402);
or U29015 (N_29015,N_20360,N_22286);
or U29016 (N_29016,N_23901,N_22866);
or U29017 (N_29017,N_24070,N_23085);
nand U29018 (N_29018,N_23532,N_20353);
or U29019 (N_29019,N_23726,N_21868);
nand U29020 (N_29020,N_23402,N_21076);
or U29021 (N_29021,N_22378,N_23015);
nor U29022 (N_29022,N_24093,N_20514);
or U29023 (N_29023,N_22074,N_22614);
nand U29024 (N_29024,N_23104,N_23885);
nand U29025 (N_29025,N_22097,N_24440);
or U29026 (N_29026,N_21384,N_21719);
nand U29027 (N_29027,N_20887,N_20466);
or U29028 (N_29028,N_22861,N_24220);
xnor U29029 (N_29029,N_20116,N_22385);
nand U29030 (N_29030,N_20870,N_23708);
and U29031 (N_29031,N_20499,N_20373);
nand U29032 (N_29032,N_21579,N_20930);
nor U29033 (N_29033,N_23461,N_22905);
nor U29034 (N_29034,N_20688,N_20957);
and U29035 (N_29035,N_22294,N_24124);
nor U29036 (N_29036,N_24919,N_24828);
and U29037 (N_29037,N_20115,N_22650);
or U29038 (N_29038,N_20434,N_20143);
or U29039 (N_29039,N_20626,N_21346);
or U29040 (N_29040,N_20713,N_24735);
nand U29041 (N_29041,N_20143,N_21730);
nand U29042 (N_29042,N_20060,N_20135);
nand U29043 (N_29043,N_21765,N_22930);
nor U29044 (N_29044,N_21270,N_23302);
or U29045 (N_29045,N_20237,N_22215);
or U29046 (N_29046,N_20468,N_24639);
or U29047 (N_29047,N_21901,N_24958);
or U29048 (N_29048,N_23296,N_23534);
and U29049 (N_29049,N_23243,N_24066);
nor U29050 (N_29050,N_24012,N_22364);
nor U29051 (N_29051,N_20458,N_24108);
nand U29052 (N_29052,N_24521,N_24528);
nor U29053 (N_29053,N_21674,N_21912);
nand U29054 (N_29054,N_24627,N_21918);
nand U29055 (N_29055,N_21333,N_24790);
nand U29056 (N_29056,N_22826,N_23982);
nor U29057 (N_29057,N_22029,N_22426);
and U29058 (N_29058,N_21161,N_23059);
or U29059 (N_29059,N_21137,N_22578);
nand U29060 (N_29060,N_24437,N_21776);
nor U29061 (N_29061,N_24556,N_21305);
nor U29062 (N_29062,N_24365,N_21368);
nand U29063 (N_29063,N_21765,N_21788);
xnor U29064 (N_29064,N_22260,N_23747);
and U29065 (N_29065,N_21382,N_20198);
and U29066 (N_29066,N_24730,N_22566);
and U29067 (N_29067,N_20907,N_24111);
and U29068 (N_29068,N_23719,N_22876);
xor U29069 (N_29069,N_22600,N_21173);
nand U29070 (N_29070,N_23361,N_21158);
nor U29071 (N_29071,N_24123,N_21553);
and U29072 (N_29072,N_24099,N_20097);
or U29073 (N_29073,N_24411,N_23767);
or U29074 (N_29074,N_21168,N_22409);
or U29075 (N_29075,N_24247,N_23231);
xnor U29076 (N_29076,N_23990,N_20133);
nor U29077 (N_29077,N_20204,N_22328);
nor U29078 (N_29078,N_23756,N_24959);
or U29079 (N_29079,N_24975,N_20845);
xor U29080 (N_29080,N_23570,N_23342);
or U29081 (N_29081,N_21279,N_24803);
and U29082 (N_29082,N_21548,N_22511);
or U29083 (N_29083,N_20727,N_20158);
or U29084 (N_29084,N_21814,N_24109);
xor U29085 (N_29085,N_22768,N_20589);
nor U29086 (N_29086,N_21655,N_20607);
or U29087 (N_29087,N_24225,N_20629);
and U29088 (N_29088,N_23752,N_22879);
and U29089 (N_29089,N_21691,N_24450);
nand U29090 (N_29090,N_22650,N_23418);
nand U29091 (N_29091,N_24993,N_22180);
nor U29092 (N_29092,N_24995,N_22421);
xnor U29093 (N_29093,N_21886,N_20089);
nand U29094 (N_29094,N_22816,N_21832);
xor U29095 (N_29095,N_24095,N_22137);
xor U29096 (N_29096,N_23948,N_20225);
or U29097 (N_29097,N_24639,N_24508);
xnor U29098 (N_29098,N_20774,N_21651);
nand U29099 (N_29099,N_20600,N_20085);
nor U29100 (N_29100,N_22571,N_21939);
nor U29101 (N_29101,N_21158,N_23184);
nor U29102 (N_29102,N_21344,N_22747);
nor U29103 (N_29103,N_23054,N_20182);
nor U29104 (N_29104,N_23790,N_20445);
nor U29105 (N_29105,N_23725,N_23354);
or U29106 (N_29106,N_23904,N_24244);
nor U29107 (N_29107,N_24399,N_24944);
or U29108 (N_29108,N_21008,N_23751);
nand U29109 (N_29109,N_23126,N_23929);
nand U29110 (N_29110,N_21027,N_21261);
and U29111 (N_29111,N_20322,N_22211);
xor U29112 (N_29112,N_22165,N_22861);
xor U29113 (N_29113,N_20784,N_20299);
nor U29114 (N_29114,N_20604,N_21259);
and U29115 (N_29115,N_24453,N_22702);
nor U29116 (N_29116,N_21899,N_24532);
nand U29117 (N_29117,N_20818,N_24220);
xor U29118 (N_29118,N_20317,N_20696);
nor U29119 (N_29119,N_21901,N_21524);
nor U29120 (N_29120,N_21930,N_20754);
nand U29121 (N_29121,N_20628,N_24185);
nor U29122 (N_29122,N_21507,N_20370);
or U29123 (N_29123,N_21517,N_21163);
nor U29124 (N_29124,N_21668,N_24678);
and U29125 (N_29125,N_21852,N_22536);
xor U29126 (N_29126,N_21590,N_22325);
xnor U29127 (N_29127,N_22122,N_24521);
nand U29128 (N_29128,N_22700,N_22598);
nand U29129 (N_29129,N_22982,N_20804);
and U29130 (N_29130,N_23507,N_23330);
nor U29131 (N_29131,N_20459,N_23734);
nor U29132 (N_29132,N_24200,N_20142);
xnor U29133 (N_29133,N_24976,N_24688);
nor U29134 (N_29134,N_23732,N_23193);
xnor U29135 (N_29135,N_20953,N_22568);
nor U29136 (N_29136,N_21803,N_21204);
or U29137 (N_29137,N_21170,N_24811);
or U29138 (N_29138,N_23617,N_23503);
nor U29139 (N_29139,N_22931,N_23260);
nand U29140 (N_29140,N_22350,N_24704);
and U29141 (N_29141,N_21822,N_20080);
and U29142 (N_29142,N_22044,N_22540);
nand U29143 (N_29143,N_23723,N_23737);
xor U29144 (N_29144,N_22871,N_20919);
xor U29145 (N_29145,N_22547,N_20940);
or U29146 (N_29146,N_24997,N_24625);
nand U29147 (N_29147,N_22289,N_20020);
or U29148 (N_29148,N_21538,N_23547);
nor U29149 (N_29149,N_21693,N_21463);
xnor U29150 (N_29150,N_20814,N_20597);
nand U29151 (N_29151,N_23528,N_22070);
and U29152 (N_29152,N_23433,N_24515);
or U29153 (N_29153,N_23993,N_24226);
and U29154 (N_29154,N_22171,N_23501);
nor U29155 (N_29155,N_24877,N_22809);
and U29156 (N_29156,N_21322,N_22566);
nand U29157 (N_29157,N_24602,N_20270);
and U29158 (N_29158,N_23766,N_21936);
or U29159 (N_29159,N_23630,N_20014);
nor U29160 (N_29160,N_20123,N_20715);
nand U29161 (N_29161,N_23771,N_24892);
nor U29162 (N_29162,N_22542,N_20402);
and U29163 (N_29163,N_21583,N_24326);
nand U29164 (N_29164,N_24759,N_21554);
and U29165 (N_29165,N_24767,N_24188);
nor U29166 (N_29166,N_20003,N_22382);
and U29167 (N_29167,N_20172,N_23041);
nand U29168 (N_29168,N_22365,N_23479);
and U29169 (N_29169,N_24763,N_22535);
or U29170 (N_29170,N_21246,N_24529);
xnor U29171 (N_29171,N_22309,N_22262);
and U29172 (N_29172,N_24308,N_24943);
xor U29173 (N_29173,N_20460,N_24474);
or U29174 (N_29174,N_21737,N_22776);
nand U29175 (N_29175,N_20806,N_24705);
nand U29176 (N_29176,N_21484,N_21246);
xnor U29177 (N_29177,N_23892,N_23870);
nor U29178 (N_29178,N_23366,N_24696);
nand U29179 (N_29179,N_24368,N_20088);
nand U29180 (N_29180,N_23889,N_20150);
nor U29181 (N_29181,N_20155,N_23463);
or U29182 (N_29182,N_24496,N_23218);
or U29183 (N_29183,N_21130,N_23687);
nor U29184 (N_29184,N_23189,N_21365);
and U29185 (N_29185,N_22312,N_24788);
nor U29186 (N_29186,N_23257,N_20039);
and U29187 (N_29187,N_22294,N_24908);
nor U29188 (N_29188,N_24581,N_23487);
or U29189 (N_29189,N_21065,N_24483);
nor U29190 (N_29190,N_20014,N_20707);
nor U29191 (N_29191,N_23448,N_21755);
and U29192 (N_29192,N_23218,N_23952);
and U29193 (N_29193,N_21501,N_23236);
xor U29194 (N_29194,N_20093,N_23159);
xnor U29195 (N_29195,N_22108,N_24426);
xor U29196 (N_29196,N_23889,N_23735);
or U29197 (N_29197,N_21270,N_21508);
nand U29198 (N_29198,N_23641,N_20097);
nor U29199 (N_29199,N_24611,N_24732);
and U29200 (N_29200,N_24787,N_20444);
xor U29201 (N_29201,N_20690,N_21416);
or U29202 (N_29202,N_20025,N_22594);
or U29203 (N_29203,N_21475,N_21392);
nor U29204 (N_29204,N_24509,N_21077);
nand U29205 (N_29205,N_20481,N_21151);
nor U29206 (N_29206,N_20223,N_20205);
nor U29207 (N_29207,N_23851,N_23984);
nand U29208 (N_29208,N_24404,N_23725);
and U29209 (N_29209,N_20783,N_24130);
or U29210 (N_29210,N_20511,N_20465);
nand U29211 (N_29211,N_21974,N_21179);
nor U29212 (N_29212,N_21921,N_23304);
nor U29213 (N_29213,N_24370,N_23883);
nor U29214 (N_29214,N_20761,N_20039);
nand U29215 (N_29215,N_24642,N_24628);
or U29216 (N_29216,N_21407,N_23995);
xor U29217 (N_29217,N_23095,N_23530);
and U29218 (N_29218,N_21594,N_23967);
nand U29219 (N_29219,N_20205,N_23991);
or U29220 (N_29220,N_21729,N_21191);
nand U29221 (N_29221,N_23972,N_22787);
nand U29222 (N_29222,N_24379,N_23730);
xnor U29223 (N_29223,N_24704,N_21026);
nor U29224 (N_29224,N_23857,N_23797);
nor U29225 (N_29225,N_20234,N_23044);
nand U29226 (N_29226,N_22055,N_21874);
nor U29227 (N_29227,N_20910,N_21727);
or U29228 (N_29228,N_22157,N_23464);
and U29229 (N_29229,N_20310,N_23718);
nor U29230 (N_29230,N_21490,N_20912);
nor U29231 (N_29231,N_23560,N_20481);
xor U29232 (N_29232,N_21030,N_20010);
xnor U29233 (N_29233,N_24816,N_20059);
nand U29234 (N_29234,N_21796,N_22916);
and U29235 (N_29235,N_23234,N_24446);
or U29236 (N_29236,N_24599,N_24085);
and U29237 (N_29237,N_22572,N_24573);
nor U29238 (N_29238,N_20758,N_21091);
or U29239 (N_29239,N_20344,N_21428);
nand U29240 (N_29240,N_20057,N_22288);
nor U29241 (N_29241,N_24941,N_22856);
or U29242 (N_29242,N_22994,N_23173);
nor U29243 (N_29243,N_24839,N_23404);
or U29244 (N_29244,N_24875,N_24236);
nand U29245 (N_29245,N_22574,N_20311);
and U29246 (N_29246,N_21961,N_21789);
or U29247 (N_29247,N_24984,N_21960);
nor U29248 (N_29248,N_22357,N_24310);
nand U29249 (N_29249,N_23776,N_24143);
and U29250 (N_29250,N_24447,N_23903);
nand U29251 (N_29251,N_24978,N_21048);
and U29252 (N_29252,N_23707,N_23898);
xnor U29253 (N_29253,N_20273,N_23533);
nand U29254 (N_29254,N_23996,N_24824);
nor U29255 (N_29255,N_22960,N_22844);
nand U29256 (N_29256,N_21244,N_24032);
nand U29257 (N_29257,N_20861,N_24975);
or U29258 (N_29258,N_23809,N_21942);
xor U29259 (N_29259,N_20734,N_23289);
nand U29260 (N_29260,N_24049,N_24489);
nand U29261 (N_29261,N_23306,N_22272);
nand U29262 (N_29262,N_23345,N_21472);
and U29263 (N_29263,N_22259,N_23928);
or U29264 (N_29264,N_20824,N_24110);
and U29265 (N_29265,N_21379,N_23529);
or U29266 (N_29266,N_22465,N_24427);
nand U29267 (N_29267,N_20324,N_22537);
nor U29268 (N_29268,N_23828,N_20746);
and U29269 (N_29269,N_21303,N_20972);
nor U29270 (N_29270,N_22599,N_23921);
and U29271 (N_29271,N_21777,N_24633);
nor U29272 (N_29272,N_20829,N_20299);
nand U29273 (N_29273,N_24133,N_20425);
or U29274 (N_29274,N_24902,N_21213);
nand U29275 (N_29275,N_22020,N_22633);
nor U29276 (N_29276,N_20518,N_23233);
xnor U29277 (N_29277,N_21710,N_20560);
nor U29278 (N_29278,N_21387,N_23982);
or U29279 (N_29279,N_24291,N_21231);
nor U29280 (N_29280,N_21891,N_21416);
nor U29281 (N_29281,N_24661,N_21529);
and U29282 (N_29282,N_22244,N_22962);
xnor U29283 (N_29283,N_24641,N_22155);
nand U29284 (N_29284,N_22202,N_20181);
and U29285 (N_29285,N_24501,N_21960);
or U29286 (N_29286,N_21793,N_23597);
xor U29287 (N_29287,N_24537,N_22837);
or U29288 (N_29288,N_21633,N_23509);
nand U29289 (N_29289,N_20052,N_24704);
xnor U29290 (N_29290,N_24618,N_23592);
nor U29291 (N_29291,N_23706,N_24961);
nand U29292 (N_29292,N_21217,N_20227);
and U29293 (N_29293,N_22697,N_24267);
nand U29294 (N_29294,N_22204,N_23651);
xor U29295 (N_29295,N_23452,N_20630);
nor U29296 (N_29296,N_22247,N_24242);
nand U29297 (N_29297,N_20124,N_22545);
or U29298 (N_29298,N_23214,N_21783);
and U29299 (N_29299,N_23195,N_24413);
nand U29300 (N_29300,N_23063,N_23660);
and U29301 (N_29301,N_22601,N_21675);
nand U29302 (N_29302,N_20395,N_23160);
and U29303 (N_29303,N_23647,N_21499);
and U29304 (N_29304,N_23935,N_21360);
or U29305 (N_29305,N_23500,N_23202);
nor U29306 (N_29306,N_22052,N_20985);
nand U29307 (N_29307,N_21407,N_23547);
or U29308 (N_29308,N_20466,N_22713);
nand U29309 (N_29309,N_20532,N_22683);
nor U29310 (N_29310,N_22500,N_20636);
or U29311 (N_29311,N_20186,N_20437);
and U29312 (N_29312,N_22619,N_21312);
and U29313 (N_29313,N_20777,N_20239);
and U29314 (N_29314,N_21776,N_23513);
nand U29315 (N_29315,N_23126,N_22102);
or U29316 (N_29316,N_23585,N_20915);
and U29317 (N_29317,N_24850,N_21582);
nand U29318 (N_29318,N_20065,N_20995);
nor U29319 (N_29319,N_23088,N_22651);
nand U29320 (N_29320,N_20182,N_22287);
nand U29321 (N_29321,N_23984,N_21246);
nand U29322 (N_29322,N_20083,N_20909);
nand U29323 (N_29323,N_20404,N_21152);
and U29324 (N_29324,N_23384,N_20414);
and U29325 (N_29325,N_23682,N_20646);
nor U29326 (N_29326,N_24061,N_20379);
nor U29327 (N_29327,N_23600,N_21693);
or U29328 (N_29328,N_24586,N_22544);
or U29329 (N_29329,N_24990,N_23283);
and U29330 (N_29330,N_20318,N_21088);
xor U29331 (N_29331,N_21441,N_20553);
nand U29332 (N_29332,N_24896,N_21772);
nand U29333 (N_29333,N_23700,N_21564);
nand U29334 (N_29334,N_23359,N_22760);
nor U29335 (N_29335,N_22236,N_21615);
nor U29336 (N_29336,N_23846,N_22864);
or U29337 (N_29337,N_21744,N_24599);
nand U29338 (N_29338,N_21861,N_21536);
nor U29339 (N_29339,N_22344,N_23930);
nand U29340 (N_29340,N_24277,N_22144);
nand U29341 (N_29341,N_22019,N_23709);
nand U29342 (N_29342,N_20468,N_21949);
or U29343 (N_29343,N_23933,N_24242);
or U29344 (N_29344,N_21485,N_24081);
nor U29345 (N_29345,N_20159,N_24665);
and U29346 (N_29346,N_22474,N_22780);
xnor U29347 (N_29347,N_24254,N_20330);
and U29348 (N_29348,N_23730,N_21849);
and U29349 (N_29349,N_20320,N_24569);
or U29350 (N_29350,N_24539,N_21699);
and U29351 (N_29351,N_23458,N_20214);
or U29352 (N_29352,N_20065,N_23666);
and U29353 (N_29353,N_23105,N_23318);
or U29354 (N_29354,N_22316,N_20208);
and U29355 (N_29355,N_24349,N_21669);
xor U29356 (N_29356,N_24739,N_24020);
nor U29357 (N_29357,N_23889,N_21421);
or U29358 (N_29358,N_24366,N_21530);
and U29359 (N_29359,N_22590,N_20406);
or U29360 (N_29360,N_21341,N_24193);
nand U29361 (N_29361,N_24009,N_24030);
or U29362 (N_29362,N_20025,N_23118);
nand U29363 (N_29363,N_21907,N_22113);
and U29364 (N_29364,N_24896,N_20726);
nor U29365 (N_29365,N_24796,N_21329);
nor U29366 (N_29366,N_23855,N_24591);
and U29367 (N_29367,N_22509,N_24139);
nor U29368 (N_29368,N_21047,N_24673);
nor U29369 (N_29369,N_23330,N_20658);
nand U29370 (N_29370,N_21537,N_23868);
and U29371 (N_29371,N_24217,N_21532);
nand U29372 (N_29372,N_21711,N_22500);
nand U29373 (N_29373,N_21238,N_23920);
or U29374 (N_29374,N_24379,N_20404);
or U29375 (N_29375,N_21273,N_20635);
nand U29376 (N_29376,N_20553,N_21985);
nor U29377 (N_29377,N_20489,N_23286);
xnor U29378 (N_29378,N_20598,N_22340);
nor U29379 (N_29379,N_23606,N_23963);
and U29380 (N_29380,N_24148,N_24270);
nor U29381 (N_29381,N_24460,N_24353);
nand U29382 (N_29382,N_21036,N_23840);
nor U29383 (N_29383,N_24354,N_21083);
and U29384 (N_29384,N_23308,N_24567);
and U29385 (N_29385,N_24256,N_23633);
nand U29386 (N_29386,N_20975,N_22549);
nand U29387 (N_29387,N_21473,N_24510);
nor U29388 (N_29388,N_22978,N_20992);
or U29389 (N_29389,N_24427,N_24658);
and U29390 (N_29390,N_22036,N_24183);
or U29391 (N_29391,N_24076,N_22545);
nand U29392 (N_29392,N_20817,N_22985);
or U29393 (N_29393,N_24459,N_22048);
and U29394 (N_29394,N_24356,N_23338);
nor U29395 (N_29395,N_21574,N_22125);
xnor U29396 (N_29396,N_20242,N_21305);
nor U29397 (N_29397,N_22479,N_22939);
or U29398 (N_29398,N_23751,N_23044);
and U29399 (N_29399,N_21382,N_23992);
xor U29400 (N_29400,N_21907,N_20698);
nand U29401 (N_29401,N_21414,N_21945);
nor U29402 (N_29402,N_20644,N_22235);
nand U29403 (N_29403,N_20173,N_24455);
xor U29404 (N_29404,N_21060,N_21717);
nand U29405 (N_29405,N_20822,N_21607);
nor U29406 (N_29406,N_24036,N_21878);
nand U29407 (N_29407,N_23794,N_24107);
and U29408 (N_29408,N_24993,N_20168);
nor U29409 (N_29409,N_20813,N_22168);
nand U29410 (N_29410,N_24190,N_23260);
xnor U29411 (N_29411,N_24106,N_23943);
xor U29412 (N_29412,N_23284,N_23233);
and U29413 (N_29413,N_24931,N_24387);
nand U29414 (N_29414,N_22356,N_23871);
nor U29415 (N_29415,N_24180,N_24230);
nand U29416 (N_29416,N_21105,N_20778);
or U29417 (N_29417,N_24194,N_23546);
nor U29418 (N_29418,N_21165,N_23676);
and U29419 (N_29419,N_22071,N_22259);
or U29420 (N_29420,N_24290,N_20528);
and U29421 (N_29421,N_22918,N_21206);
and U29422 (N_29422,N_23136,N_23328);
and U29423 (N_29423,N_22649,N_21615);
and U29424 (N_29424,N_21433,N_20395);
or U29425 (N_29425,N_21588,N_23160);
and U29426 (N_29426,N_22907,N_21410);
xnor U29427 (N_29427,N_20181,N_22259);
or U29428 (N_29428,N_24633,N_23779);
nand U29429 (N_29429,N_24288,N_22550);
nand U29430 (N_29430,N_22745,N_22533);
and U29431 (N_29431,N_23889,N_24085);
or U29432 (N_29432,N_24853,N_20471);
and U29433 (N_29433,N_20927,N_21369);
and U29434 (N_29434,N_20373,N_24760);
nor U29435 (N_29435,N_21525,N_24414);
nand U29436 (N_29436,N_24748,N_21220);
nand U29437 (N_29437,N_20763,N_20501);
or U29438 (N_29438,N_20345,N_20250);
nor U29439 (N_29439,N_20533,N_21682);
xor U29440 (N_29440,N_20302,N_22096);
xnor U29441 (N_29441,N_24519,N_24434);
xor U29442 (N_29442,N_20058,N_23316);
nand U29443 (N_29443,N_20078,N_21136);
nand U29444 (N_29444,N_20383,N_23301);
and U29445 (N_29445,N_23497,N_23369);
nand U29446 (N_29446,N_21340,N_22635);
and U29447 (N_29447,N_20491,N_21741);
or U29448 (N_29448,N_20011,N_22551);
or U29449 (N_29449,N_21732,N_23904);
nand U29450 (N_29450,N_21450,N_24790);
nor U29451 (N_29451,N_24089,N_20002);
and U29452 (N_29452,N_23841,N_23027);
nor U29453 (N_29453,N_23482,N_21860);
or U29454 (N_29454,N_23733,N_21648);
or U29455 (N_29455,N_21992,N_24823);
and U29456 (N_29456,N_22679,N_22296);
or U29457 (N_29457,N_24692,N_24010);
and U29458 (N_29458,N_21023,N_22448);
nand U29459 (N_29459,N_21862,N_21131);
nand U29460 (N_29460,N_20133,N_24144);
and U29461 (N_29461,N_21321,N_22496);
and U29462 (N_29462,N_23892,N_24307);
and U29463 (N_29463,N_22349,N_24273);
nor U29464 (N_29464,N_20799,N_23461);
nand U29465 (N_29465,N_22055,N_21733);
nor U29466 (N_29466,N_23037,N_22200);
and U29467 (N_29467,N_21148,N_21509);
nor U29468 (N_29468,N_21364,N_20150);
or U29469 (N_29469,N_22513,N_22999);
and U29470 (N_29470,N_22580,N_23890);
nor U29471 (N_29471,N_22306,N_24815);
and U29472 (N_29472,N_22864,N_21053);
nor U29473 (N_29473,N_21331,N_21199);
nor U29474 (N_29474,N_24879,N_21039);
nand U29475 (N_29475,N_21532,N_22756);
or U29476 (N_29476,N_24772,N_22558);
nand U29477 (N_29477,N_21995,N_24214);
nor U29478 (N_29478,N_22039,N_23084);
or U29479 (N_29479,N_24038,N_22218);
or U29480 (N_29480,N_20545,N_24138);
nor U29481 (N_29481,N_20156,N_20439);
and U29482 (N_29482,N_22474,N_20947);
nor U29483 (N_29483,N_20253,N_21638);
nor U29484 (N_29484,N_23230,N_22309);
and U29485 (N_29485,N_22180,N_21552);
and U29486 (N_29486,N_21728,N_23564);
or U29487 (N_29487,N_24828,N_20374);
and U29488 (N_29488,N_24337,N_24895);
nand U29489 (N_29489,N_20342,N_20239);
and U29490 (N_29490,N_21973,N_23371);
or U29491 (N_29491,N_23487,N_21000);
nor U29492 (N_29492,N_20002,N_20537);
nor U29493 (N_29493,N_23472,N_23371);
or U29494 (N_29494,N_21754,N_20679);
or U29495 (N_29495,N_23841,N_21608);
nor U29496 (N_29496,N_23645,N_23028);
xnor U29497 (N_29497,N_24648,N_20440);
nor U29498 (N_29498,N_24192,N_23622);
and U29499 (N_29499,N_23782,N_20982);
and U29500 (N_29500,N_22806,N_21480);
xor U29501 (N_29501,N_23523,N_22597);
or U29502 (N_29502,N_23656,N_21310);
nor U29503 (N_29503,N_23189,N_24627);
nand U29504 (N_29504,N_23429,N_22036);
or U29505 (N_29505,N_20726,N_24916);
nand U29506 (N_29506,N_23580,N_22084);
nor U29507 (N_29507,N_23049,N_24426);
nand U29508 (N_29508,N_23502,N_22424);
xor U29509 (N_29509,N_21260,N_22979);
or U29510 (N_29510,N_20697,N_24127);
or U29511 (N_29511,N_21236,N_24325);
xor U29512 (N_29512,N_24268,N_22887);
nor U29513 (N_29513,N_24263,N_20219);
nand U29514 (N_29514,N_21998,N_22584);
nor U29515 (N_29515,N_24991,N_21203);
xor U29516 (N_29516,N_22079,N_21882);
or U29517 (N_29517,N_21711,N_20916);
nand U29518 (N_29518,N_22961,N_22335);
xnor U29519 (N_29519,N_24613,N_23721);
and U29520 (N_29520,N_24248,N_22678);
nand U29521 (N_29521,N_22904,N_23370);
or U29522 (N_29522,N_20781,N_24097);
nor U29523 (N_29523,N_21076,N_21406);
or U29524 (N_29524,N_23227,N_20825);
nor U29525 (N_29525,N_20321,N_24338);
nor U29526 (N_29526,N_23680,N_24069);
nand U29527 (N_29527,N_24122,N_24716);
or U29528 (N_29528,N_20126,N_20007);
or U29529 (N_29529,N_24745,N_21060);
and U29530 (N_29530,N_24660,N_23942);
nor U29531 (N_29531,N_22898,N_23749);
xnor U29532 (N_29532,N_21635,N_23584);
nand U29533 (N_29533,N_22340,N_23961);
nand U29534 (N_29534,N_20665,N_22546);
or U29535 (N_29535,N_24345,N_24282);
xnor U29536 (N_29536,N_21000,N_24788);
or U29537 (N_29537,N_23379,N_20236);
xor U29538 (N_29538,N_23343,N_21888);
nand U29539 (N_29539,N_22229,N_20487);
nand U29540 (N_29540,N_22577,N_24361);
and U29541 (N_29541,N_22069,N_23075);
xor U29542 (N_29542,N_22607,N_23464);
and U29543 (N_29543,N_24811,N_20303);
nor U29544 (N_29544,N_22429,N_21870);
and U29545 (N_29545,N_24715,N_23070);
nor U29546 (N_29546,N_24462,N_20465);
or U29547 (N_29547,N_20278,N_21633);
nor U29548 (N_29548,N_23001,N_22214);
nand U29549 (N_29549,N_24534,N_22714);
nand U29550 (N_29550,N_24330,N_21160);
and U29551 (N_29551,N_23655,N_22712);
nor U29552 (N_29552,N_23569,N_21795);
and U29553 (N_29553,N_20977,N_21447);
nand U29554 (N_29554,N_24900,N_23091);
nor U29555 (N_29555,N_23813,N_23639);
nand U29556 (N_29556,N_24104,N_24654);
xnor U29557 (N_29557,N_24302,N_24963);
or U29558 (N_29558,N_23563,N_20199);
nor U29559 (N_29559,N_21589,N_20410);
nand U29560 (N_29560,N_22478,N_20112);
nand U29561 (N_29561,N_20060,N_21690);
xnor U29562 (N_29562,N_24023,N_21922);
nand U29563 (N_29563,N_20840,N_23504);
nand U29564 (N_29564,N_20167,N_24533);
or U29565 (N_29565,N_20489,N_21260);
and U29566 (N_29566,N_22756,N_21859);
or U29567 (N_29567,N_24561,N_22874);
xor U29568 (N_29568,N_21791,N_22856);
nor U29569 (N_29569,N_23797,N_21326);
xor U29570 (N_29570,N_24301,N_20914);
or U29571 (N_29571,N_23175,N_23261);
xnor U29572 (N_29572,N_24849,N_21960);
and U29573 (N_29573,N_23747,N_23012);
or U29574 (N_29574,N_21520,N_24406);
nand U29575 (N_29575,N_22804,N_22049);
nor U29576 (N_29576,N_23510,N_23040);
nand U29577 (N_29577,N_23083,N_20383);
or U29578 (N_29578,N_24089,N_20873);
nand U29579 (N_29579,N_21075,N_23914);
nand U29580 (N_29580,N_23160,N_24494);
nand U29581 (N_29581,N_22610,N_24647);
or U29582 (N_29582,N_21686,N_20476);
or U29583 (N_29583,N_21551,N_20229);
nand U29584 (N_29584,N_24358,N_23900);
nor U29585 (N_29585,N_22799,N_21879);
nand U29586 (N_29586,N_20185,N_20537);
or U29587 (N_29587,N_22376,N_24487);
or U29588 (N_29588,N_23349,N_21176);
nor U29589 (N_29589,N_20584,N_20119);
nor U29590 (N_29590,N_24077,N_21878);
nand U29591 (N_29591,N_21352,N_22904);
nor U29592 (N_29592,N_22713,N_21347);
nor U29593 (N_29593,N_20564,N_20482);
nand U29594 (N_29594,N_24421,N_23285);
or U29595 (N_29595,N_21475,N_23258);
xor U29596 (N_29596,N_22486,N_22835);
nor U29597 (N_29597,N_23756,N_22845);
nand U29598 (N_29598,N_24217,N_24542);
or U29599 (N_29599,N_20901,N_20805);
and U29600 (N_29600,N_20021,N_24784);
xnor U29601 (N_29601,N_24535,N_23805);
or U29602 (N_29602,N_21336,N_21792);
and U29603 (N_29603,N_23852,N_23422);
or U29604 (N_29604,N_20817,N_23623);
and U29605 (N_29605,N_22557,N_21267);
nand U29606 (N_29606,N_22032,N_24745);
nand U29607 (N_29607,N_24712,N_21083);
and U29608 (N_29608,N_23046,N_23988);
nand U29609 (N_29609,N_24617,N_22297);
and U29610 (N_29610,N_24830,N_21635);
and U29611 (N_29611,N_21775,N_20817);
nor U29612 (N_29612,N_22304,N_20999);
or U29613 (N_29613,N_22002,N_20358);
nand U29614 (N_29614,N_20616,N_20805);
nor U29615 (N_29615,N_24135,N_22470);
nor U29616 (N_29616,N_20808,N_22802);
xor U29617 (N_29617,N_21881,N_21739);
or U29618 (N_29618,N_24567,N_23727);
nor U29619 (N_29619,N_23083,N_24125);
or U29620 (N_29620,N_24371,N_20657);
nand U29621 (N_29621,N_21686,N_24251);
and U29622 (N_29622,N_24938,N_22657);
and U29623 (N_29623,N_22889,N_24626);
xnor U29624 (N_29624,N_20886,N_22327);
nor U29625 (N_29625,N_24872,N_20147);
or U29626 (N_29626,N_20265,N_20659);
or U29627 (N_29627,N_21784,N_23840);
xor U29628 (N_29628,N_21180,N_23680);
nor U29629 (N_29629,N_24697,N_24235);
or U29630 (N_29630,N_22408,N_23360);
and U29631 (N_29631,N_20880,N_21932);
nand U29632 (N_29632,N_23587,N_23653);
nand U29633 (N_29633,N_20579,N_21750);
or U29634 (N_29634,N_20730,N_20471);
nand U29635 (N_29635,N_22420,N_20182);
or U29636 (N_29636,N_22842,N_23588);
nand U29637 (N_29637,N_23058,N_24262);
xor U29638 (N_29638,N_21950,N_20668);
and U29639 (N_29639,N_24450,N_23485);
nor U29640 (N_29640,N_23033,N_21164);
and U29641 (N_29641,N_20393,N_23621);
or U29642 (N_29642,N_24580,N_20002);
nand U29643 (N_29643,N_20302,N_21020);
nand U29644 (N_29644,N_20575,N_24678);
xor U29645 (N_29645,N_22176,N_22834);
and U29646 (N_29646,N_24662,N_24800);
or U29647 (N_29647,N_20427,N_21259);
nor U29648 (N_29648,N_22654,N_21904);
nand U29649 (N_29649,N_22312,N_22658);
nand U29650 (N_29650,N_24693,N_23400);
nand U29651 (N_29651,N_23531,N_22606);
and U29652 (N_29652,N_20246,N_22053);
or U29653 (N_29653,N_20460,N_21068);
nand U29654 (N_29654,N_23314,N_22113);
and U29655 (N_29655,N_22123,N_23650);
or U29656 (N_29656,N_24180,N_23701);
and U29657 (N_29657,N_21744,N_24301);
nor U29658 (N_29658,N_21806,N_23614);
or U29659 (N_29659,N_24035,N_22167);
and U29660 (N_29660,N_20816,N_20586);
nor U29661 (N_29661,N_22965,N_21562);
and U29662 (N_29662,N_20912,N_20580);
nor U29663 (N_29663,N_21760,N_21990);
or U29664 (N_29664,N_24347,N_21376);
and U29665 (N_29665,N_21421,N_23954);
nand U29666 (N_29666,N_24607,N_23476);
nor U29667 (N_29667,N_22418,N_24337);
and U29668 (N_29668,N_23291,N_24567);
xor U29669 (N_29669,N_22503,N_23804);
xnor U29670 (N_29670,N_23186,N_24531);
xor U29671 (N_29671,N_21009,N_24725);
and U29672 (N_29672,N_21313,N_20204);
nor U29673 (N_29673,N_20032,N_22870);
nand U29674 (N_29674,N_22849,N_24517);
and U29675 (N_29675,N_23209,N_22352);
nor U29676 (N_29676,N_23934,N_23102);
and U29677 (N_29677,N_23443,N_22601);
xor U29678 (N_29678,N_23423,N_24807);
and U29679 (N_29679,N_20081,N_23104);
xnor U29680 (N_29680,N_22910,N_22644);
and U29681 (N_29681,N_20367,N_24761);
or U29682 (N_29682,N_24716,N_24642);
nand U29683 (N_29683,N_20209,N_20355);
or U29684 (N_29684,N_24933,N_21680);
and U29685 (N_29685,N_24979,N_23053);
xor U29686 (N_29686,N_23183,N_24311);
and U29687 (N_29687,N_21211,N_21779);
or U29688 (N_29688,N_22082,N_21480);
and U29689 (N_29689,N_23238,N_22718);
or U29690 (N_29690,N_21641,N_22350);
nand U29691 (N_29691,N_23169,N_20511);
and U29692 (N_29692,N_22470,N_24081);
nand U29693 (N_29693,N_23685,N_22089);
nand U29694 (N_29694,N_23669,N_24075);
xor U29695 (N_29695,N_24083,N_21791);
or U29696 (N_29696,N_23359,N_23513);
and U29697 (N_29697,N_23748,N_21124);
or U29698 (N_29698,N_22777,N_23024);
nor U29699 (N_29699,N_22096,N_24927);
nor U29700 (N_29700,N_24734,N_20066);
nand U29701 (N_29701,N_20770,N_21386);
nor U29702 (N_29702,N_24855,N_20460);
nor U29703 (N_29703,N_24129,N_21346);
nand U29704 (N_29704,N_24725,N_20661);
nand U29705 (N_29705,N_20319,N_22679);
nor U29706 (N_29706,N_24310,N_22536);
nand U29707 (N_29707,N_22001,N_23288);
nor U29708 (N_29708,N_24133,N_20600);
or U29709 (N_29709,N_20939,N_23742);
and U29710 (N_29710,N_24381,N_24980);
xnor U29711 (N_29711,N_23750,N_23347);
nor U29712 (N_29712,N_23546,N_23807);
nand U29713 (N_29713,N_23531,N_22016);
nor U29714 (N_29714,N_21105,N_22327);
and U29715 (N_29715,N_24374,N_23496);
or U29716 (N_29716,N_22004,N_21102);
or U29717 (N_29717,N_20029,N_23433);
nand U29718 (N_29718,N_20372,N_24321);
and U29719 (N_29719,N_20470,N_21689);
or U29720 (N_29720,N_24563,N_23406);
nor U29721 (N_29721,N_22345,N_20762);
nor U29722 (N_29722,N_24847,N_20886);
and U29723 (N_29723,N_24708,N_21867);
and U29724 (N_29724,N_20535,N_23352);
nand U29725 (N_29725,N_20264,N_22062);
nand U29726 (N_29726,N_23305,N_22074);
nand U29727 (N_29727,N_21979,N_20273);
nand U29728 (N_29728,N_24182,N_22604);
and U29729 (N_29729,N_23822,N_20024);
nor U29730 (N_29730,N_21635,N_20354);
or U29731 (N_29731,N_22108,N_21638);
nand U29732 (N_29732,N_24753,N_22018);
nand U29733 (N_29733,N_24296,N_22370);
nand U29734 (N_29734,N_23136,N_24814);
xor U29735 (N_29735,N_23306,N_20664);
nor U29736 (N_29736,N_21415,N_20092);
nor U29737 (N_29737,N_24225,N_23854);
and U29738 (N_29738,N_21711,N_20457);
nand U29739 (N_29739,N_21267,N_23406);
nor U29740 (N_29740,N_24250,N_21809);
and U29741 (N_29741,N_22377,N_21997);
xor U29742 (N_29742,N_23924,N_24623);
nor U29743 (N_29743,N_24648,N_22363);
and U29744 (N_29744,N_21924,N_21758);
nand U29745 (N_29745,N_20657,N_20718);
nor U29746 (N_29746,N_22635,N_21049);
xor U29747 (N_29747,N_21666,N_22643);
and U29748 (N_29748,N_21532,N_21876);
and U29749 (N_29749,N_22002,N_24886);
or U29750 (N_29750,N_21406,N_20725);
or U29751 (N_29751,N_20274,N_24578);
nand U29752 (N_29752,N_21341,N_24900);
or U29753 (N_29753,N_23683,N_23905);
and U29754 (N_29754,N_20479,N_21275);
nand U29755 (N_29755,N_22813,N_23721);
or U29756 (N_29756,N_20578,N_21735);
nor U29757 (N_29757,N_23379,N_21513);
and U29758 (N_29758,N_20763,N_22891);
or U29759 (N_29759,N_24911,N_21762);
nand U29760 (N_29760,N_23964,N_22653);
and U29761 (N_29761,N_20316,N_22685);
and U29762 (N_29762,N_20899,N_22617);
and U29763 (N_29763,N_24472,N_22101);
and U29764 (N_29764,N_24378,N_24803);
nand U29765 (N_29765,N_20446,N_22206);
or U29766 (N_29766,N_24551,N_23823);
nor U29767 (N_29767,N_22420,N_23927);
nor U29768 (N_29768,N_22387,N_23042);
and U29769 (N_29769,N_20758,N_23693);
nor U29770 (N_29770,N_22467,N_21535);
and U29771 (N_29771,N_23414,N_24307);
nor U29772 (N_29772,N_22407,N_20925);
nand U29773 (N_29773,N_20206,N_20269);
or U29774 (N_29774,N_21691,N_24569);
nor U29775 (N_29775,N_23909,N_23401);
nor U29776 (N_29776,N_24851,N_20747);
nand U29777 (N_29777,N_20113,N_20304);
and U29778 (N_29778,N_23227,N_22748);
nor U29779 (N_29779,N_24087,N_22927);
and U29780 (N_29780,N_23867,N_21316);
nand U29781 (N_29781,N_24591,N_23328);
or U29782 (N_29782,N_22345,N_20618);
or U29783 (N_29783,N_24076,N_22232);
or U29784 (N_29784,N_22934,N_23173);
or U29785 (N_29785,N_23061,N_22204);
nand U29786 (N_29786,N_21009,N_21028);
nor U29787 (N_29787,N_20825,N_23969);
or U29788 (N_29788,N_20182,N_23126);
nor U29789 (N_29789,N_24514,N_21226);
or U29790 (N_29790,N_21985,N_20927);
and U29791 (N_29791,N_23478,N_22528);
and U29792 (N_29792,N_24132,N_21754);
xor U29793 (N_29793,N_24735,N_22947);
xnor U29794 (N_29794,N_20206,N_24629);
nand U29795 (N_29795,N_20568,N_23394);
and U29796 (N_29796,N_24186,N_20436);
and U29797 (N_29797,N_21415,N_22116);
nand U29798 (N_29798,N_20911,N_24629);
or U29799 (N_29799,N_22930,N_22338);
nand U29800 (N_29800,N_23842,N_24181);
and U29801 (N_29801,N_20782,N_22586);
nor U29802 (N_29802,N_23061,N_22801);
or U29803 (N_29803,N_22677,N_22308);
nor U29804 (N_29804,N_21112,N_22110);
and U29805 (N_29805,N_22340,N_20299);
nand U29806 (N_29806,N_23747,N_22030);
and U29807 (N_29807,N_24958,N_22314);
or U29808 (N_29808,N_20296,N_23155);
nor U29809 (N_29809,N_23760,N_22144);
nand U29810 (N_29810,N_23107,N_21876);
xnor U29811 (N_29811,N_24023,N_22840);
or U29812 (N_29812,N_23971,N_23558);
or U29813 (N_29813,N_24903,N_24629);
and U29814 (N_29814,N_20391,N_23303);
and U29815 (N_29815,N_21687,N_21078);
nor U29816 (N_29816,N_21888,N_21350);
or U29817 (N_29817,N_20448,N_24585);
or U29818 (N_29818,N_22897,N_22108);
nor U29819 (N_29819,N_24367,N_22989);
or U29820 (N_29820,N_21091,N_23974);
nor U29821 (N_29821,N_24623,N_21543);
or U29822 (N_29822,N_24179,N_21774);
and U29823 (N_29823,N_22878,N_20131);
nand U29824 (N_29824,N_24654,N_20396);
nor U29825 (N_29825,N_22843,N_22217);
and U29826 (N_29826,N_24519,N_23530);
or U29827 (N_29827,N_23704,N_24447);
and U29828 (N_29828,N_21652,N_21559);
nand U29829 (N_29829,N_21502,N_22739);
nor U29830 (N_29830,N_22767,N_23216);
and U29831 (N_29831,N_23263,N_22014);
nor U29832 (N_29832,N_21007,N_21343);
and U29833 (N_29833,N_20551,N_21769);
or U29834 (N_29834,N_21238,N_20481);
nor U29835 (N_29835,N_23538,N_24488);
nand U29836 (N_29836,N_21456,N_24267);
xor U29837 (N_29837,N_22113,N_20275);
nor U29838 (N_29838,N_21672,N_21238);
nand U29839 (N_29839,N_23411,N_20482);
nand U29840 (N_29840,N_24601,N_24296);
and U29841 (N_29841,N_23593,N_24563);
nand U29842 (N_29842,N_23582,N_21398);
xnor U29843 (N_29843,N_23885,N_23372);
and U29844 (N_29844,N_22728,N_24227);
and U29845 (N_29845,N_22268,N_23861);
and U29846 (N_29846,N_21148,N_22104);
nand U29847 (N_29847,N_24990,N_23622);
nor U29848 (N_29848,N_20327,N_20817);
and U29849 (N_29849,N_24168,N_23827);
nor U29850 (N_29850,N_20253,N_21482);
and U29851 (N_29851,N_21955,N_22649);
nor U29852 (N_29852,N_20416,N_20091);
nand U29853 (N_29853,N_23601,N_22787);
nand U29854 (N_29854,N_23781,N_22858);
nor U29855 (N_29855,N_20398,N_23494);
nand U29856 (N_29856,N_20066,N_22149);
nand U29857 (N_29857,N_24918,N_23034);
or U29858 (N_29858,N_20215,N_24717);
nor U29859 (N_29859,N_20172,N_23382);
and U29860 (N_29860,N_21171,N_20404);
and U29861 (N_29861,N_24639,N_21222);
nand U29862 (N_29862,N_20722,N_24474);
or U29863 (N_29863,N_24487,N_23922);
nor U29864 (N_29864,N_23294,N_20002);
and U29865 (N_29865,N_24442,N_22076);
xor U29866 (N_29866,N_23774,N_24464);
nor U29867 (N_29867,N_22234,N_22150);
nand U29868 (N_29868,N_21898,N_24359);
or U29869 (N_29869,N_24262,N_24182);
nor U29870 (N_29870,N_24292,N_23040);
nor U29871 (N_29871,N_24300,N_20657);
and U29872 (N_29872,N_21774,N_22924);
nand U29873 (N_29873,N_23925,N_21200);
or U29874 (N_29874,N_22722,N_22734);
nand U29875 (N_29875,N_21933,N_20600);
and U29876 (N_29876,N_22403,N_20014);
and U29877 (N_29877,N_22985,N_24051);
xor U29878 (N_29878,N_24976,N_22934);
nand U29879 (N_29879,N_24904,N_22315);
or U29880 (N_29880,N_20824,N_24192);
nand U29881 (N_29881,N_22992,N_23715);
xnor U29882 (N_29882,N_23797,N_23002);
nand U29883 (N_29883,N_24999,N_21891);
nand U29884 (N_29884,N_24633,N_22711);
nand U29885 (N_29885,N_21361,N_20553);
nand U29886 (N_29886,N_22441,N_24019);
nand U29887 (N_29887,N_20565,N_22639);
or U29888 (N_29888,N_21358,N_21573);
and U29889 (N_29889,N_20980,N_22189);
nor U29890 (N_29890,N_23694,N_24776);
and U29891 (N_29891,N_21384,N_22083);
or U29892 (N_29892,N_21541,N_22345);
or U29893 (N_29893,N_23872,N_23983);
or U29894 (N_29894,N_24129,N_22498);
nand U29895 (N_29895,N_22781,N_20045);
or U29896 (N_29896,N_21428,N_23294);
or U29897 (N_29897,N_20043,N_24158);
nor U29898 (N_29898,N_23737,N_21111);
and U29899 (N_29899,N_20095,N_21072);
nand U29900 (N_29900,N_20508,N_24483);
or U29901 (N_29901,N_22369,N_20178);
nand U29902 (N_29902,N_22557,N_20578);
nor U29903 (N_29903,N_24299,N_24162);
and U29904 (N_29904,N_23964,N_24939);
xor U29905 (N_29905,N_21502,N_20640);
nor U29906 (N_29906,N_20361,N_20601);
or U29907 (N_29907,N_21378,N_20831);
and U29908 (N_29908,N_21627,N_23496);
nor U29909 (N_29909,N_24364,N_22001);
nor U29910 (N_29910,N_20740,N_23030);
xnor U29911 (N_29911,N_24479,N_20087);
nand U29912 (N_29912,N_22318,N_23211);
nor U29913 (N_29913,N_20956,N_20551);
xor U29914 (N_29914,N_23410,N_20119);
nor U29915 (N_29915,N_22130,N_22481);
or U29916 (N_29916,N_22398,N_20049);
or U29917 (N_29917,N_24537,N_20579);
and U29918 (N_29918,N_20267,N_24217);
xor U29919 (N_29919,N_24405,N_20114);
or U29920 (N_29920,N_21367,N_20247);
nor U29921 (N_29921,N_22688,N_24661);
or U29922 (N_29922,N_24363,N_22233);
and U29923 (N_29923,N_24752,N_21981);
nand U29924 (N_29924,N_20976,N_21992);
nand U29925 (N_29925,N_21167,N_20105);
and U29926 (N_29926,N_22076,N_23580);
nand U29927 (N_29927,N_20558,N_23849);
or U29928 (N_29928,N_23167,N_22078);
and U29929 (N_29929,N_20911,N_22870);
nor U29930 (N_29930,N_21850,N_24031);
or U29931 (N_29931,N_22894,N_22153);
nand U29932 (N_29932,N_23108,N_21062);
nor U29933 (N_29933,N_20154,N_22113);
and U29934 (N_29934,N_23768,N_23388);
or U29935 (N_29935,N_23848,N_21150);
nand U29936 (N_29936,N_21099,N_23546);
xor U29937 (N_29937,N_22361,N_20836);
or U29938 (N_29938,N_24491,N_22939);
or U29939 (N_29939,N_21260,N_23995);
nand U29940 (N_29940,N_23945,N_21468);
and U29941 (N_29941,N_21010,N_21692);
or U29942 (N_29942,N_21426,N_22526);
nand U29943 (N_29943,N_21059,N_20988);
or U29944 (N_29944,N_22253,N_23549);
nor U29945 (N_29945,N_24078,N_22091);
or U29946 (N_29946,N_23199,N_21311);
and U29947 (N_29947,N_24355,N_24426);
nand U29948 (N_29948,N_23974,N_24547);
or U29949 (N_29949,N_22140,N_23689);
nand U29950 (N_29950,N_20574,N_20111);
or U29951 (N_29951,N_23508,N_20066);
xor U29952 (N_29952,N_22992,N_23282);
nor U29953 (N_29953,N_22863,N_23633);
nand U29954 (N_29954,N_21346,N_22968);
xor U29955 (N_29955,N_20152,N_24307);
or U29956 (N_29956,N_23499,N_23021);
or U29957 (N_29957,N_22117,N_22035);
or U29958 (N_29958,N_24511,N_22829);
nor U29959 (N_29959,N_23961,N_20889);
nor U29960 (N_29960,N_23510,N_21604);
nand U29961 (N_29961,N_23627,N_22941);
and U29962 (N_29962,N_23216,N_22053);
nor U29963 (N_29963,N_20655,N_22130);
or U29964 (N_29964,N_22544,N_21283);
nand U29965 (N_29965,N_20751,N_21066);
and U29966 (N_29966,N_20689,N_22777);
nand U29967 (N_29967,N_20059,N_21312);
nand U29968 (N_29968,N_23248,N_21100);
nand U29969 (N_29969,N_20545,N_21350);
and U29970 (N_29970,N_22842,N_20137);
xor U29971 (N_29971,N_21030,N_21397);
and U29972 (N_29972,N_20494,N_21764);
xnor U29973 (N_29973,N_23465,N_20555);
and U29974 (N_29974,N_21538,N_21466);
or U29975 (N_29975,N_24479,N_21215);
nand U29976 (N_29976,N_20712,N_20287);
and U29977 (N_29977,N_23260,N_22615);
nor U29978 (N_29978,N_24536,N_23746);
nor U29979 (N_29979,N_22174,N_21577);
and U29980 (N_29980,N_23091,N_24345);
xor U29981 (N_29981,N_24307,N_23536);
or U29982 (N_29982,N_20036,N_23728);
or U29983 (N_29983,N_24067,N_23781);
nor U29984 (N_29984,N_22899,N_22716);
and U29985 (N_29985,N_22903,N_22435);
nor U29986 (N_29986,N_21378,N_21767);
or U29987 (N_29987,N_24178,N_23854);
or U29988 (N_29988,N_22106,N_22707);
xnor U29989 (N_29989,N_21765,N_21483);
nand U29990 (N_29990,N_20526,N_20238);
nand U29991 (N_29991,N_24286,N_20894);
and U29992 (N_29992,N_21146,N_23256);
or U29993 (N_29993,N_20284,N_22572);
or U29994 (N_29994,N_20764,N_20950);
or U29995 (N_29995,N_20318,N_20129);
and U29996 (N_29996,N_23216,N_22376);
nand U29997 (N_29997,N_20605,N_21298);
or U29998 (N_29998,N_20747,N_24997);
xnor U29999 (N_29999,N_24707,N_24257);
nor U30000 (N_30000,N_26632,N_26729);
nor U30001 (N_30001,N_25040,N_25719);
xnor U30002 (N_30002,N_27574,N_25486);
nor U30003 (N_30003,N_28300,N_26268);
xor U30004 (N_30004,N_27486,N_29041);
nor U30005 (N_30005,N_26830,N_26566);
xnor U30006 (N_30006,N_25720,N_26071);
nand U30007 (N_30007,N_25726,N_25877);
nand U30008 (N_30008,N_25105,N_26090);
or U30009 (N_30009,N_27637,N_29957);
and U30010 (N_30010,N_27862,N_26937);
nand U30011 (N_30011,N_28655,N_26685);
and U30012 (N_30012,N_29239,N_25947);
xnor U30013 (N_30013,N_29656,N_27300);
and U30014 (N_30014,N_26537,N_26372);
nand U30015 (N_30015,N_29737,N_25513);
nor U30016 (N_30016,N_29860,N_27547);
nor U30017 (N_30017,N_25721,N_28801);
or U30018 (N_30018,N_26654,N_27457);
nand U30019 (N_30019,N_27554,N_29241);
or U30020 (N_30020,N_27046,N_28844);
or U30021 (N_30021,N_26263,N_26210);
or U30022 (N_30022,N_28348,N_29251);
nor U30023 (N_30023,N_28529,N_29775);
and U30024 (N_30024,N_25598,N_28284);
or U30025 (N_30025,N_26317,N_28140);
nand U30026 (N_30026,N_28755,N_29166);
nand U30027 (N_30027,N_26167,N_27111);
and U30028 (N_30028,N_28314,N_27347);
or U30029 (N_30029,N_27353,N_27285);
nor U30030 (N_30030,N_25966,N_28857);
nand U30031 (N_30031,N_25714,N_26986);
nand U30032 (N_30032,N_29893,N_28063);
and U30033 (N_30033,N_28675,N_28738);
nor U30034 (N_30034,N_28530,N_28347);
nand U30035 (N_30035,N_25799,N_25081);
nand U30036 (N_30036,N_28405,N_28029);
nand U30037 (N_30037,N_27061,N_26631);
xor U30038 (N_30038,N_26875,N_28250);
nor U30039 (N_30039,N_26097,N_29335);
nor U30040 (N_30040,N_25389,N_27215);
or U30041 (N_30041,N_27688,N_28240);
and U30042 (N_30042,N_25977,N_25065);
or U30043 (N_30043,N_28929,N_26351);
xor U30044 (N_30044,N_25694,N_25018);
and U30045 (N_30045,N_26383,N_26367);
xnor U30046 (N_30046,N_26754,N_27770);
nand U30047 (N_30047,N_25242,N_29324);
or U30048 (N_30048,N_29009,N_27963);
nor U30049 (N_30049,N_26034,N_28193);
xnor U30050 (N_30050,N_28587,N_25152);
nor U30051 (N_30051,N_29887,N_27582);
nand U30052 (N_30052,N_28433,N_25371);
nor U30053 (N_30053,N_26811,N_27911);
or U30054 (N_30054,N_27157,N_29851);
and U30055 (N_30055,N_28438,N_27489);
nor U30056 (N_30056,N_26294,N_25588);
nor U30057 (N_30057,N_29849,N_25507);
and U30058 (N_30058,N_25473,N_27145);
nand U30059 (N_30059,N_27287,N_25928);
xor U30060 (N_30060,N_26267,N_28797);
or U30061 (N_30061,N_27456,N_28377);
and U30062 (N_30062,N_29913,N_26256);
and U30063 (N_30063,N_29058,N_26499);
or U30064 (N_30064,N_27063,N_28648);
nor U30065 (N_30065,N_25829,N_25216);
and U30066 (N_30066,N_25149,N_26823);
xnor U30067 (N_30067,N_25963,N_26241);
and U30068 (N_30068,N_27234,N_29633);
and U30069 (N_30069,N_27533,N_28730);
and U30070 (N_30070,N_26431,N_28480);
nand U30071 (N_30071,N_26790,N_27081);
or U30072 (N_30072,N_28039,N_29279);
and U30073 (N_30073,N_25000,N_27584);
or U30074 (N_30074,N_26198,N_27222);
nand U30075 (N_30075,N_25992,N_29881);
nand U30076 (N_30076,N_29606,N_25739);
or U30077 (N_30077,N_29475,N_29210);
and U30078 (N_30078,N_29404,N_26743);
and U30079 (N_30079,N_28399,N_27834);
or U30080 (N_30080,N_28065,N_27967);
or U30081 (N_30081,N_29135,N_29966);
or U30082 (N_30082,N_26932,N_26737);
or U30083 (N_30083,N_26669,N_29052);
and U30084 (N_30084,N_26543,N_27108);
nor U30085 (N_30085,N_29092,N_25136);
and U30086 (N_30086,N_27957,N_28912);
xnor U30087 (N_30087,N_29638,N_28069);
or U30088 (N_30088,N_29502,N_29422);
nand U30089 (N_30089,N_25421,N_27600);
nor U30090 (N_30090,N_26358,N_28682);
nor U30091 (N_30091,N_26032,N_25047);
or U30092 (N_30092,N_29038,N_29529);
and U30093 (N_30093,N_29131,N_29163);
nor U30094 (N_30094,N_26377,N_27049);
nand U30095 (N_30095,N_28249,N_28926);
and U30096 (N_30096,N_28391,N_28335);
nand U30097 (N_30097,N_29112,N_25482);
or U30098 (N_30098,N_26553,N_29193);
nor U30099 (N_30099,N_28280,N_25681);
nand U30100 (N_30100,N_25887,N_27281);
xnor U30101 (N_30101,N_25317,N_29876);
nor U30102 (N_30102,N_27331,N_26187);
and U30103 (N_30103,N_27781,N_25344);
and U30104 (N_30104,N_27601,N_25703);
xor U30105 (N_30105,N_26460,N_26018);
nand U30106 (N_30106,N_28763,N_25478);
and U30107 (N_30107,N_29442,N_28518);
and U30108 (N_30108,N_25207,N_26174);
and U30109 (N_30109,N_28515,N_29890);
nor U30110 (N_30110,N_29740,N_27943);
xor U30111 (N_30111,N_27738,N_25821);
nand U30112 (N_30112,N_27598,N_26336);
nor U30113 (N_30113,N_28051,N_27727);
or U30114 (N_30114,N_29892,N_28867);
nor U30115 (N_30115,N_28878,N_26013);
and U30116 (N_30116,N_25087,N_28232);
nor U30117 (N_30117,N_29297,N_26374);
nand U30118 (N_30118,N_25808,N_28877);
nor U30119 (N_30119,N_27659,N_25810);
nor U30120 (N_30120,N_27627,N_25903);
and U30121 (N_30121,N_27101,N_27759);
nand U30122 (N_30122,N_25015,N_26946);
or U30123 (N_30123,N_28308,N_25825);
nor U30124 (N_30124,N_27602,N_27459);
nand U30125 (N_30125,N_27882,N_26767);
nor U30126 (N_30126,N_28323,N_27211);
and U30127 (N_30127,N_27761,N_27237);
and U30128 (N_30128,N_25575,N_28044);
nand U30129 (N_30129,N_28264,N_25777);
or U30130 (N_30130,N_26794,N_26453);
or U30131 (N_30131,N_27744,N_29726);
xor U30132 (N_30132,N_27613,N_27571);
nor U30133 (N_30133,N_27067,N_25611);
and U30134 (N_30134,N_25819,N_25595);
nand U30135 (N_30135,N_29445,N_29456);
or U30136 (N_30136,N_27359,N_25673);
and U30137 (N_30137,N_26853,N_25809);
xnor U30138 (N_30138,N_28026,N_29412);
nand U30139 (N_30139,N_25290,N_27426);
nor U30140 (N_30140,N_29671,N_26515);
nand U30141 (N_30141,N_25100,N_26793);
and U30142 (N_30142,N_27815,N_27380);
nand U30143 (N_30143,N_25875,N_25376);
xor U30144 (N_30144,N_26678,N_25935);
and U30145 (N_30145,N_27888,N_25048);
and U30146 (N_30146,N_26834,N_26440);
nor U30147 (N_30147,N_29353,N_25060);
and U30148 (N_30148,N_26176,N_28533);
or U30149 (N_30149,N_25988,N_25792);
or U30150 (N_30150,N_29730,N_29394);
nand U30151 (N_30151,N_29078,N_28141);
and U30152 (N_30152,N_27516,N_26520);
nand U30153 (N_30153,N_28916,N_26973);
xnor U30154 (N_30154,N_27989,N_26974);
nand U30155 (N_30155,N_29944,N_27166);
and U30156 (N_30156,N_25471,N_28829);
xor U30157 (N_30157,N_29548,N_25349);
and U30158 (N_30158,N_28237,N_29348);
xor U30159 (N_30159,N_28610,N_25836);
nand U30160 (N_30160,N_28118,N_27649);
nand U30161 (N_30161,N_25646,N_26542);
and U30162 (N_30162,N_29197,N_29342);
nand U30163 (N_30163,N_29296,N_26378);
nand U30164 (N_30164,N_27055,N_27236);
and U30165 (N_30165,N_28368,N_25049);
and U30166 (N_30166,N_27549,N_27025);
nor U30167 (N_30167,N_25323,N_25658);
and U30168 (N_30168,N_27464,N_25549);
nor U30169 (N_30169,N_27408,N_28503);
nand U30170 (N_30170,N_27762,N_27003);
or U30171 (N_30171,N_29660,N_28490);
and U30172 (N_30172,N_27253,N_29792);
nand U30173 (N_30173,N_26745,N_27954);
xor U30174 (N_30174,N_27853,N_28189);
nor U30175 (N_30175,N_28167,N_25700);
or U30176 (N_30176,N_27608,N_29341);
and U30177 (N_30177,N_27151,N_29327);
nand U30178 (N_30178,N_26252,N_29861);
xor U30179 (N_30179,N_27133,N_29395);
nand U30180 (N_30180,N_25094,N_25969);
and U30181 (N_30181,N_27488,N_27418);
nand U30182 (N_30182,N_28547,N_29277);
nand U30183 (N_30183,N_29469,N_25517);
and U30184 (N_30184,N_25820,N_27315);
and U30185 (N_30185,N_28413,N_25350);
nor U30186 (N_30186,N_28718,N_28680);
or U30187 (N_30187,N_28639,N_25390);
nor U30188 (N_30188,N_25538,N_25175);
nor U30189 (N_30189,N_25064,N_25251);
nor U30190 (N_30190,N_25042,N_25248);
and U30191 (N_30191,N_28524,N_26370);
nand U30192 (N_30192,N_25727,N_28743);
and U30193 (N_30193,N_27280,N_25837);
and U30194 (N_30194,N_25543,N_25164);
or U30195 (N_30195,N_29350,N_28714);
nor U30196 (N_30196,N_27631,N_26056);
and U30197 (N_30197,N_25539,N_28853);
xnor U30198 (N_30198,N_29776,N_25070);
or U30199 (N_30199,N_27956,N_27412);
xnor U30200 (N_30200,N_25982,N_29698);
nand U30201 (N_30201,N_25174,N_29495);
nand U30202 (N_30202,N_28922,N_27527);
nor U30203 (N_30203,N_28288,N_27844);
or U30204 (N_30204,N_27490,N_25102);
nand U30205 (N_30205,N_29199,N_29274);
nand U30206 (N_30206,N_25937,N_29271);
nand U30207 (N_30207,N_27142,N_25456);
nand U30208 (N_30208,N_26560,N_28905);
nand U30209 (N_30209,N_28523,N_25041);
or U30210 (N_30210,N_26569,N_25879);
or U30211 (N_30211,N_28061,N_29732);
and U30212 (N_30212,N_28998,N_27594);
or U30213 (N_30213,N_25217,N_25795);
and U30214 (N_30214,N_25537,N_28387);
nand U30215 (N_30215,N_28016,N_26825);
and U30216 (N_30216,N_25274,N_28373);
xor U30217 (N_30217,N_25560,N_27886);
and U30218 (N_30218,N_29108,N_28759);
and U30219 (N_30219,N_26180,N_26108);
and U30220 (N_30220,N_29276,N_26707);
or U30221 (N_30221,N_27419,N_26861);
or U30222 (N_30222,N_28129,N_27648);
or U30223 (N_30223,N_28823,N_28709);
nor U30224 (N_30224,N_28132,N_29380);
nand U30225 (N_30225,N_29285,N_25632);
or U30226 (N_30226,N_29448,N_25710);
or U30227 (N_30227,N_29617,N_25083);
and U30228 (N_30228,N_27047,N_27842);
nor U30229 (N_30229,N_26143,N_27243);
and U30230 (N_30230,N_29855,N_29922);
nor U30231 (N_30231,N_28213,N_25626);
nor U30232 (N_30232,N_25874,N_25062);
nor U30233 (N_30233,N_26417,N_27019);
nand U30234 (N_30234,N_26872,N_28400);
and U30235 (N_30235,N_26259,N_25336);
and U30236 (N_30236,N_28021,N_28705);
nand U30237 (N_30237,N_26410,N_25522);
nor U30238 (N_30238,N_26068,N_27891);
nand U30239 (N_30239,N_25990,N_29713);
and U30240 (N_30240,N_29240,N_26592);
and U30241 (N_30241,N_27104,N_29772);
or U30242 (N_30242,N_29269,N_29461);
and U30243 (N_30243,N_29684,N_27766);
or U30244 (N_30244,N_29289,N_25145);
nor U30245 (N_30245,N_25692,N_25247);
and U30246 (N_30246,N_27736,N_29185);
and U30247 (N_30247,N_26369,N_26082);
or U30248 (N_30248,N_29584,N_28012);
nor U30249 (N_30249,N_25017,N_28441);
or U30250 (N_30250,N_26916,N_25748);
nand U30251 (N_30251,N_29852,N_27093);
xor U30252 (N_30252,N_26432,N_29111);
and U30253 (N_30253,N_26910,N_26833);
or U30254 (N_30254,N_29653,N_25245);
nand U30255 (N_30255,N_28505,N_26302);
or U30256 (N_30256,N_25728,N_29019);
and U30257 (N_30257,N_28054,N_27346);
and U30258 (N_30258,N_26433,N_29280);
and U30259 (N_30259,N_28080,N_26730);
nor U30260 (N_30260,N_29843,N_27473);
or U30261 (N_30261,N_27259,N_26172);
nand U30262 (N_30262,N_25150,N_26675);
nand U30263 (N_30263,N_27128,N_25036);
or U30264 (N_30264,N_29723,N_26679);
xnor U30265 (N_30265,N_28430,N_29015);
nand U30266 (N_30266,N_29367,N_28301);
and U30267 (N_30267,N_25555,N_26297);
nand U30268 (N_30268,N_29156,N_25212);
nor U30269 (N_30269,N_25976,N_27877);
nand U30270 (N_30270,N_26043,N_28402);
xnor U30271 (N_30271,N_27849,N_25892);
or U30272 (N_30272,N_28047,N_25378);
nor U30273 (N_30273,N_29013,N_27854);
nor U30274 (N_30274,N_29321,N_27779);
nand U30275 (N_30275,N_29867,N_27981);
and U30276 (N_30276,N_29786,N_28669);
xor U30277 (N_30277,N_29609,N_25080);
and U30278 (N_30278,N_26792,N_25237);
nand U30279 (N_30279,N_26398,N_29414);
and U30280 (N_30280,N_29362,N_26663);
nand U30281 (N_30281,N_28398,N_26442);
and U30282 (N_30282,N_25832,N_29034);
nor U30283 (N_30283,N_26044,N_25587);
nand U30284 (N_30284,N_29573,N_27732);
or U30285 (N_30285,N_25337,N_26371);
and U30286 (N_30286,N_28152,N_29508);
and U30287 (N_30287,N_25238,N_26009);
or U30288 (N_30288,N_29071,N_26286);
and U30289 (N_30289,N_26444,N_25960);
or U30290 (N_30290,N_29856,N_26429);
or U30291 (N_30291,N_26870,N_26321);
nor U30292 (N_30292,N_28657,N_29416);
or U30293 (N_30293,N_27553,N_29267);
and U30294 (N_30294,N_29547,N_25604);
nand U30295 (N_30295,N_28270,N_26506);
xnor U30296 (N_30296,N_26243,N_28153);
or U30297 (N_30297,N_25715,N_28765);
nand U30298 (N_30298,N_26512,N_28479);
nor U30299 (N_30299,N_27544,N_29478);
or U30300 (N_30300,N_25627,N_28628);
nor U30301 (N_30301,N_27062,N_26047);
nand U30302 (N_30302,N_26615,N_26538);
xor U30303 (N_30303,N_29134,N_25847);
xnor U30304 (N_30304,N_29787,N_27368);
and U30305 (N_30305,N_28170,N_26918);
or U30306 (N_30306,N_27207,N_29374);
or U30307 (N_30307,N_28125,N_25030);
xnor U30308 (N_30308,N_29190,N_27424);
nor U30309 (N_30309,N_25278,N_27343);
nand U30310 (N_30310,N_25252,N_28581);
xor U30311 (N_30311,N_27113,N_27268);
xor U30312 (N_30312,N_26805,N_28356);
nor U30313 (N_30313,N_27860,N_28919);
or U30314 (N_30314,N_26558,N_29702);
and U30315 (N_30315,N_28297,N_25031);
or U30316 (N_30316,N_28785,N_25026);
nor U30317 (N_30317,N_29433,N_27054);
xnor U30318 (N_30318,N_28334,N_28494);
nand U30319 (N_30319,N_26462,N_27221);
xnor U30320 (N_30320,N_26171,N_27152);
xnor U30321 (N_30321,N_26762,N_29945);
and U30322 (N_30322,N_28043,N_25128);
and U30323 (N_30323,N_28835,N_26579);
nor U30324 (N_30324,N_25452,N_25126);
nor U30325 (N_30325,N_27375,N_26924);
and U30326 (N_30326,N_27909,N_29074);
nand U30327 (N_30327,N_26150,N_26272);
or U30328 (N_30328,N_29001,N_29100);
nand U30329 (N_30329,N_28493,N_28219);
nor U30330 (N_30330,N_29828,N_29819);
and U30331 (N_30331,N_25725,N_29971);
nor U30332 (N_30332,N_26839,N_28848);
or U30333 (N_30333,N_25383,N_27689);
or U30334 (N_30334,N_26474,N_28290);
or U30335 (N_30335,N_25226,N_26261);
nor U30336 (N_30336,N_25756,N_28559);
nand U30337 (N_30337,N_25521,N_29593);
nor U30338 (N_30338,N_28071,N_29153);
or U30339 (N_30339,N_28800,N_27823);
nor U30340 (N_30340,N_28573,N_25256);
nor U30341 (N_30341,N_29915,N_25896);
or U30342 (N_30342,N_25599,N_27393);
nor U30343 (N_30343,N_29696,N_25730);
and U30344 (N_30344,N_28833,N_27563);
or U30345 (N_30345,N_25824,N_25610);
or U30346 (N_30346,N_29333,N_29232);
nand U30347 (N_30347,N_25529,N_25477);
or U30348 (N_30348,N_25057,N_26151);
nand U30349 (N_30349,N_29727,N_26340);
and U30350 (N_30350,N_26595,N_27141);
nand U30351 (N_30351,N_26091,N_27057);
and U30352 (N_30352,N_25330,N_29755);
and U30353 (N_30353,N_27785,N_29579);
and U30354 (N_30354,N_25377,N_29005);
and U30355 (N_30355,N_27468,N_29816);
nand U30356 (N_30356,N_28576,N_27182);
nor U30357 (N_30357,N_26397,N_28428);
or U30358 (N_30358,N_28178,N_28603);
nor U30359 (N_30359,N_29051,N_25639);
xnor U30360 (N_30360,N_28066,N_27454);
and U30361 (N_30361,N_28013,N_26731);
xnor U30362 (N_30362,N_29494,N_29368);
nor U30363 (N_30363,N_25165,N_26234);
nor U30364 (N_30364,N_28318,N_28339);
nand U30365 (N_30365,N_29118,N_25420);
and U30366 (N_30366,N_28673,N_26664);
nor U30367 (N_30367,N_25939,N_27297);
and U30368 (N_30368,N_25436,N_26925);
nand U30369 (N_30369,N_29569,N_26457);
nand U30370 (N_30370,N_28049,N_26426);
or U30371 (N_30371,N_29972,N_26724);
nor U30372 (N_30372,N_29568,N_29284);
and U30373 (N_30373,N_26634,N_28647);
nor U30374 (N_30374,N_28475,N_28983);
and U30375 (N_30375,N_27518,N_27514);
or U30376 (N_30376,N_26332,N_28027);
nand U30377 (N_30377,N_29325,N_28298);
or U30378 (N_30378,N_29227,N_29809);
nor U30379 (N_30379,N_26469,N_27639);
and U30380 (N_30380,N_28561,N_27576);
nor U30381 (N_30381,N_27256,N_28435);
nor U30382 (N_30382,N_25270,N_26969);
and U30383 (N_30383,N_27745,N_27229);
nand U30384 (N_30384,N_29756,N_27317);
nand U30385 (N_30385,N_28964,N_27638);
nor U30386 (N_30386,N_27387,N_25932);
nand U30387 (N_30387,N_29378,N_26118);
nor U30388 (N_30388,N_25911,N_29449);
xnor U30389 (N_30389,N_28491,N_28052);
nor U30390 (N_30390,N_27717,N_28584);
nor U30391 (N_30391,N_26001,N_28594);
and U30392 (N_30392,N_28932,N_29686);
nand U30393 (N_30393,N_28664,N_26053);
nand U30394 (N_30394,N_26721,N_28397);
and U30395 (N_30395,N_28773,N_27710);
and U30396 (N_30396,N_27614,N_28355);
xor U30397 (N_30397,N_26025,N_25173);
nor U30398 (N_30398,N_25803,N_25373);
or U30399 (N_30399,N_28499,N_28843);
and U30400 (N_30400,N_25455,N_29479);
nor U30401 (N_30401,N_29334,N_25745);
nor U30402 (N_30402,N_27445,N_28936);
nand U30403 (N_30403,N_29583,N_29645);
or U30404 (N_30404,N_28163,N_28987);
nand U30405 (N_30405,N_28821,N_25056);
or U30406 (N_30406,N_26221,N_28073);
nor U30407 (N_30407,N_29516,N_27903);
nor U30408 (N_30408,N_29859,N_26067);
and U30409 (N_30409,N_29793,N_26593);
and U30410 (N_30410,N_26997,N_27086);
and U30411 (N_30411,N_28651,N_27254);
nor U30412 (N_30412,N_25052,N_29160);
and U30413 (N_30413,N_26352,N_25641);
and U30414 (N_30414,N_27333,N_26461);
nor U30415 (N_30415,N_26368,N_28366);
nand U30416 (N_30416,N_28942,N_26062);
and U30417 (N_30417,N_27180,N_28754);
and U30418 (N_30418,N_25086,N_25978);
and U30419 (N_30419,N_26092,N_26016);
nand U30420 (N_30420,N_25067,N_26695);
xnor U30421 (N_30421,N_25919,N_27365);
nor U30422 (N_30422,N_27120,N_28789);
or U30423 (N_30423,N_27179,N_25108);
xnor U30424 (N_30424,N_26657,N_26653);
and U30425 (N_30425,N_29714,N_29505);
nor U30426 (N_30426,N_28378,N_29965);
and U30427 (N_30427,N_28920,N_26339);
nor U30428 (N_30428,N_26482,N_25495);
nand U30429 (N_30429,N_29435,N_29635);
xnor U30430 (N_30430,N_26435,N_28341);
nand U30431 (N_30431,N_25503,N_25922);
xor U30432 (N_30432,N_29999,N_25561);
or U30433 (N_30433,N_25013,N_29132);
or U30434 (N_30434,N_26246,N_26753);
xnor U30435 (N_30435,N_28904,N_28960);
nor U30436 (N_30436,N_25335,N_28331);
xor U30437 (N_30437,N_27843,N_29098);
xnor U30438 (N_30438,N_26718,N_25084);
or U30439 (N_30439,N_29091,N_25872);
xnor U30440 (N_30440,N_28512,N_27805);
nor U30441 (N_30441,N_26552,N_27356);
and U30442 (N_30442,N_28064,N_28426);
nor U30443 (N_30443,N_26778,N_26237);
nand U30444 (N_30444,N_29758,N_25151);
nand U30445 (N_30445,N_25510,N_27984);
nor U30446 (N_30446,N_28181,N_27804);
or U30447 (N_30447,N_29365,N_28642);
or U30448 (N_30448,N_27425,N_28019);
or U30449 (N_30449,N_26005,N_27033);
nand U30450 (N_30450,N_25573,N_29674);
nand U30451 (N_30451,N_27325,N_28406);
and U30452 (N_30452,N_29719,N_25074);
nand U30453 (N_30453,N_25857,N_25442);
or U30454 (N_30454,N_26085,N_27103);
or U30455 (N_30455,N_28752,N_29838);
and U30456 (N_30456,N_28386,N_25112);
and U30457 (N_30457,N_27465,N_28006);
nand U30458 (N_30458,N_28943,N_29498);
nand U30459 (N_30459,N_26274,N_29905);
or U30460 (N_30460,N_27299,N_27806);
and U30461 (N_30461,N_26407,N_25124);
nor U30462 (N_30462,N_28191,N_29912);
nor U30463 (N_30463,N_29891,N_28055);
nor U30464 (N_30464,N_26803,N_26105);
nand U30465 (N_30465,N_29400,N_29451);
and U30466 (N_30466,N_29235,N_25007);
or U30467 (N_30467,N_27487,N_27716);
or U30468 (N_30468,N_28448,N_27754);
nand U30469 (N_30469,N_28900,N_29888);
or U30470 (N_30470,N_29387,N_25880);
or U30471 (N_30471,N_25757,N_27344);
nor U30472 (N_30472,N_29063,N_26464);
nand U30473 (N_30473,N_28045,N_25717);
and U30474 (N_30474,N_28194,N_25945);
or U30475 (N_30475,N_27700,N_28078);
or U30476 (N_30476,N_28575,N_27266);
nand U30477 (N_30477,N_28892,N_26990);
nand U30478 (N_30478,N_26546,N_28591);
nand U30479 (N_30479,N_26498,N_28018);
or U30480 (N_30480,N_25740,N_26994);
nand U30481 (N_30481,N_28910,N_25137);
nor U30482 (N_30482,N_29465,N_28199);
and U30483 (N_30483,N_25016,N_26361);
xor U30484 (N_30484,N_29658,N_27091);
nor U30485 (N_30485,N_26574,N_25179);
and U30486 (N_30486,N_26083,N_27453);
and U30487 (N_30487,N_27548,N_27379);
nor U30488 (N_30488,N_25733,N_26810);
nand U30489 (N_30489,N_25754,N_25622);
or U30490 (N_30490,N_26212,N_27220);
and U30491 (N_30491,N_26691,N_25097);
nor U30492 (N_30492,N_28053,N_29814);
nand U30493 (N_30493,N_27908,N_29429);
nand U30494 (N_30494,N_26114,N_28927);
or U30495 (N_30495,N_26158,N_27367);
or U30496 (N_30496,N_26270,N_27027);
xor U30497 (N_30497,N_28498,N_25569);
nor U30498 (N_30498,N_28982,N_27219);
and U30499 (N_30499,N_28084,N_28706);
nor U30500 (N_30500,N_26868,N_25944);
nand U30501 (N_30501,N_27959,N_28889);
and U30502 (N_30502,N_25422,N_26638);
and U30503 (N_30503,N_26519,N_29918);
nor U30504 (N_30504,N_27289,N_25955);
nand U30505 (N_30505,N_25002,N_29248);
or U30506 (N_30506,N_28296,N_26625);
nor U30507 (N_30507,N_28760,N_28941);
or U30508 (N_30508,N_28917,N_28562);
nor U30509 (N_30509,N_26882,N_27624);
nor U30510 (N_30510,N_26341,N_26201);
nand U30511 (N_30511,N_28003,N_25120);
and U30512 (N_30512,N_28796,N_27587);
and U30513 (N_30513,N_29426,N_28077);
and U30514 (N_30514,N_26907,N_27728);
and U30515 (N_30515,N_29874,N_25055);
and U30516 (N_30516,N_27520,N_29906);
nor U30517 (N_30517,N_28116,N_26285);
nand U30518 (N_30518,N_27201,N_29510);
xor U30519 (N_30519,N_26051,N_28635);
nor U30520 (N_30520,N_27997,N_27993);
and U30521 (N_30521,N_27181,N_27833);
nand U30522 (N_30522,N_27148,N_28209);
xor U30523 (N_30523,N_26766,N_28091);
and U30524 (N_30524,N_29612,N_28990);
or U30525 (N_30525,N_28149,N_25643);
and U30526 (N_30526,N_25855,N_28721);
nand U30527 (N_30527,N_29815,N_29557);
nor U30528 (N_30528,N_26576,N_25953);
or U30529 (N_30529,N_27200,N_28032);
nor U30530 (N_30530,N_28417,N_29268);
and U30531 (N_30531,N_29452,N_26800);
or U30532 (N_30532,N_28502,N_25333);
or U30533 (N_30533,N_28888,N_29546);
or U30534 (N_30534,N_27171,N_26389);
xor U30535 (N_30535,N_26318,N_25296);
nor U30536 (N_30536,N_27352,N_29916);
xnor U30537 (N_30537,N_26661,N_28715);
and U30538 (N_30538,N_26315,N_27175);
xor U30539 (N_30539,N_25468,N_27296);
nor U30540 (N_30540,N_27278,N_27397);
and U30541 (N_30541,N_27525,N_29018);
nand U30542 (N_30542,N_25523,N_25684);
xor U30543 (N_30543,N_28558,N_28712);
and U30544 (N_30544,N_25365,N_28344);
nor U30545 (N_30545,N_28906,N_26900);
xnor U30546 (N_30546,N_26817,N_28599);
nand U30547 (N_30547,N_26194,N_27556);
nand U30548 (N_30548,N_27270,N_27283);
xnor U30549 (N_30549,N_28452,N_28903);
or U30550 (N_30550,N_29164,N_28745);
or U30551 (N_30551,N_26603,N_27610);
nand U30552 (N_30552,N_29923,N_27098);
xor U30553 (N_30553,N_25965,N_29685);
nand U30554 (N_30554,N_29586,N_27513);
and U30555 (N_30555,N_25940,N_28202);
nand U30556 (N_30556,N_26905,N_25967);
and U30557 (N_30557,N_26760,N_28546);
nor U30558 (N_30558,N_26271,N_26776);
and U30559 (N_30559,N_27965,N_28251);
and U30560 (N_30560,N_28542,N_27483);
nor U30561 (N_30561,N_26602,N_26610);
nor U30562 (N_30562,N_28262,N_26393);
nand U30563 (N_30563,N_26844,N_29848);
nor U30564 (N_30564,N_26042,N_28117);
and U30565 (N_30565,N_28746,N_27966);
and U30566 (N_30566,N_26496,N_28396);
and U30567 (N_30567,N_25210,N_27307);
and U30568 (N_30568,N_28938,N_29613);
nand U30569 (N_30569,N_27497,N_28768);
nand U30570 (N_30570,N_29396,N_25178);
xnor U30571 (N_30571,N_25530,N_25861);
and U30572 (N_30572,N_27481,N_26459);
xnor U30573 (N_30573,N_28000,N_28067);
or U30574 (N_30574,N_25841,N_29234);
nor U30575 (N_30575,N_25366,N_26572);
nand U30576 (N_30576,N_26066,N_27752);
nor U30577 (N_30577,N_29564,N_26225);
and U30578 (N_30578,N_29046,N_25770);
xnor U30579 (N_30579,N_26236,N_29827);
and U30580 (N_30580,N_26054,N_26855);
nor U30581 (N_30581,N_28702,N_28271);
and U30582 (N_30582,N_25427,N_27264);
or U30583 (N_30583,N_25659,N_28028);
nor U30584 (N_30584,N_28269,N_28838);
and U30585 (N_30585,N_27354,N_28371);
nor U30586 (N_30586,N_26401,N_28733);
and U30587 (N_30587,N_27077,N_25869);
or U30588 (N_30588,N_26831,N_26550);
nand U30589 (N_30589,N_26616,N_29314);
nor U30590 (N_30590,N_26326,N_28307);
or U30591 (N_30591,N_29563,N_29937);
nor U30592 (N_30592,N_27392,N_27204);
nor U30593 (N_30593,N_29047,N_27557);
and U30594 (N_30594,N_27725,N_28588);
nor U30595 (N_30595,N_28585,N_28393);
and U30596 (N_30596,N_28999,N_28557);
nor U30597 (N_30597,N_29149,N_25329);
nand U30598 (N_30598,N_28617,N_28808);
nor U30599 (N_30599,N_29219,N_27656);
xor U30600 (N_30600,N_28470,N_25141);
and U30601 (N_30601,N_27743,N_28699);
nand U30602 (N_30602,N_27480,N_29604);
and U30603 (N_30603,N_29488,N_26149);
nand U30604 (N_30604,N_25493,N_25582);
and U30605 (N_30605,N_29694,N_27078);
xor U30606 (N_30606,N_27442,N_26979);
nand U30607 (N_30607,N_25211,N_29624);
and U30608 (N_30608,N_25785,N_29305);
nor U30609 (N_30609,N_28668,N_25813);
nor U30610 (N_30610,N_28762,N_25320);
and U30611 (N_30611,N_28360,N_29229);
nand U30612 (N_30612,N_26554,N_26406);
or U30613 (N_30613,N_26452,N_27786);
nand U30614 (N_30614,N_29590,N_25340);
or U30615 (N_30615,N_28563,N_26886);
nor U30616 (N_30616,N_29138,N_26972);
xnor U30617 (N_30617,N_25750,N_27472);
nor U30618 (N_30618,N_25104,N_25461);
or U30619 (N_30619,N_26684,N_29833);
and U30620 (N_30620,N_29477,N_26175);
nand U30621 (N_30621,N_25926,N_29585);
and U30622 (N_30622,N_29250,N_27110);
nand U30623 (N_30623,N_29120,N_27674);
nand U30624 (N_30624,N_28676,N_26074);
nand U30625 (N_30625,N_28662,N_29294);
nor U30626 (N_30626,N_27129,N_25962);
or U30627 (N_30627,N_25638,N_26298);
and U30628 (N_30628,N_29954,N_26156);
nand U30629 (N_30629,N_26945,N_29935);
and U30630 (N_30630,N_28818,N_25225);
nand U30631 (N_30631,N_25434,N_28370);
xnor U30632 (N_30632,N_29803,N_26484);
and U30633 (N_30633,N_26881,N_27642);
nand U30634 (N_30634,N_29857,N_27791);
nor U30635 (N_30635,N_29777,N_26555);
nor U30636 (N_30636,N_26284,N_27318);
or U30637 (N_30637,N_28868,N_29213);
nor U30638 (N_30638,N_29627,N_25751);
nor U30639 (N_30639,N_25884,N_28549);
nand U30640 (N_30640,N_29391,N_29863);
xor U30641 (N_30641,N_27644,N_25419);
or U30642 (N_30642,N_25213,N_25931);
nor U30643 (N_30643,N_28075,N_29877);
or U30644 (N_30644,N_26726,N_28579);
nor U30645 (N_30645,N_29802,N_28445);
nor U30646 (N_30646,N_29535,N_27947);
or U30647 (N_30647,N_25764,N_28590);
xor U30648 (N_30648,N_27377,N_27012);
and U30649 (N_30649,N_27240,N_25850);
xor U30650 (N_30650,N_26311,N_26599);
and U30651 (N_30651,N_27719,N_26942);
xnor U30652 (N_30652,N_29907,N_27138);
or U30653 (N_30653,N_27446,N_27802);
nand U30654 (N_30654,N_29467,N_28685);
nor U30655 (N_30655,N_26621,N_28875);
nand U30656 (N_30656,N_26020,N_28257);
xnor U30657 (N_30657,N_28120,N_28770);
nor U30658 (N_30658,N_25166,N_26015);
nor U30659 (N_30659,N_27664,N_28188);
or U30660 (N_30660,N_29531,N_25051);
nand U30661 (N_30661,N_29764,N_26828);
nand U30662 (N_30662,N_26671,N_25467);
nand U30663 (N_30663,N_28772,N_26033);
or U30664 (N_30664,N_25416,N_28226);
nand U30665 (N_30665,N_29716,N_26214);
and U30666 (N_30666,N_27482,N_27705);
or U30667 (N_30667,N_29979,N_25010);
and U30668 (N_30668,N_25737,N_25858);
and U30669 (N_30669,N_28036,N_27185);
nand U30670 (N_30670,N_29175,N_29329);
nand U30671 (N_30671,N_28312,N_27671);
or U30672 (N_30672,N_28211,N_27147);
or U30673 (N_30673,N_27796,N_27357);
nand U30674 (N_30674,N_27100,N_28521);
nand U30675 (N_30675,N_29552,N_29530);
and U30676 (N_30676,N_26022,N_25291);
xnor U30677 (N_30677,N_28467,N_25883);
nand U30678 (N_30678,N_25533,N_27540);
and U30679 (N_30679,N_27008,N_27939);
nor U30680 (N_30680,N_29963,N_27774);
and U30681 (N_30681,N_25612,N_28897);
nor U30682 (N_30682,N_27227,N_25499);
nor U30683 (N_30683,N_29733,N_29360);
nor U30684 (N_30684,N_25593,N_28830);
or U30685 (N_30685,N_26842,N_29553);
nor U30686 (N_30686,N_25601,N_25325);
xnor U30687 (N_30687,N_25313,N_25873);
nand U30688 (N_30688,N_26878,N_28485);
nor U30689 (N_30689,N_26379,N_25012);
nand U30690 (N_30690,N_25310,N_26470);
or U30691 (N_30691,N_28126,N_27376);
nor U30692 (N_30692,N_27373,N_25445);
or U30693 (N_30693,N_29050,N_27400);
nand U30694 (N_30694,N_28974,N_26136);
nor U30695 (N_30695,N_25395,N_27742);
nand U30696 (N_30696,N_26854,N_25146);
xnor U30697 (N_30697,N_26992,N_29223);
nand U30698 (N_30698,N_25272,N_28672);
and U30699 (N_30699,N_25901,N_25357);
and U30700 (N_30700,N_29381,N_26320);
nor U30701 (N_30701,N_28483,N_27696);
nor U30702 (N_30702,N_26301,N_28749);
or U30703 (N_30703,N_28074,N_27314);
nand U30704 (N_30704,N_27960,N_25121);
nand U30705 (N_30705,N_25849,N_25439);
or U30706 (N_30706,N_28114,N_26622);
nor U30707 (N_30707,N_29919,N_27210);
or U30708 (N_30708,N_25635,N_25624);
nand U30709 (N_30709,N_26568,N_29582);
nand U30710 (N_30710,N_25050,N_27428);
and U30711 (N_30711,N_28795,N_25838);
and U30712 (N_30712,N_28967,N_29027);
or U30713 (N_30713,N_29326,N_26570);
and U30714 (N_30714,N_27708,N_27050);
xor U30715 (N_30715,N_29821,N_28993);
and U30716 (N_30716,N_29008,N_27684);
or U30717 (N_30717,N_26075,N_26809);
nor U30718 (N_30718,N_28766,N_27431);
nand U30719 (N_30719,N_29114,N_29804);
and U30720 (N_30720,N_27566,N_27304);
nand U30721 (N_30721,N_28701,N_29541);
or U30722 (N_30722,N_26303,N_28783);
and U30723 (N_30723,N_29317,N_25775);
nand U30724 (N_30724,N_29113,N_27623);
nor U30725 (N_30725,N_27383,N_28429);
nand U30726 (N_30726,N_25667,N_28656);
xnor U30727 (N_30727,N_27884,N_28015);
nand U30728 (N_30728,N_27150,N_28414);
nand U30729 (N_30729,N_29345,N_25209);
or U30730 (N_30730,N_27187,N_29763);
or U30731 (N_30731,N_27542,N_29526);
nor U30732 (N_30732,N_26540,N_25630);
and U30733 (N_30733,N_29061,N_26098);
and U30734 (N_30734,N_27313,N_25182);
nand U30735 (N_30735,N_25028,N_26215);
nand U30736 (N_30736,N_28222,N_29415);
or U30737 (N_30737,N_29288,N_25765);
nor U30738 (N_30738,N_28729,N_26629);
or U30739 (N_30739,N_29688,N_27326);
and U30740 (N_30740,N_26646,N_27810);
and U30741 (N_30741,N_25072,N_26380);
nor U30742 (N_30742,N_26427,N_26993);
or U30743 (N_30743,N_25882,N_25675);
nor U30744 (N_30744,N_26796,N_29760);
and U30745 (N_30745,N_29509,N_28683);
nand U30746 (N_30746,N_27703,N_26505);
or U30747 (N_30747,N_25532,N_29187);
nand U30748 (N_30748,N_27134,N_29236);
or U30749 (N_30749,N_26985,N_28166);
and U30750 (N_30750,N_27937,N_25941);
nor U30751 (N_30751,N_29914,N_25243);
or U30752 (N_30752,N_28565,N_29955);
xnor U30753 (N_30753,N_25132,N_27874);
nand U30754 (N_30754,N_25581,N_28023);
nor U30755 (N_30755,N_27389,N_28395);
nand U30756 (N_30756,N_25563,N_26670);
and U30757 (N_30757,N_29921,N_28740);
nand U30758 (N_30758,N_29659,N_25413);
nor U30759 (N_30759,N_26240,N_28109);
nand U30760 (N_30760,N_29938,N_25699);
nor U30761 (N_30761,N_25197,N_29690);
or U30762 (N_30762,N_26052,N_29678);
or U30763 (N_30763,N_25856,N_28605);
nor U30764 (N_30764,N_25712,N_26395);
or U30765 (N_30765,N_29570,N_26818);
or U30766 (N_30766,N_29295,N_27709);
and U30767 (N_30767,N_28996,N_29930);
xor U30768 (N_30768,N_27076,N_26667);
nor U30769 (N_30769,N_29708,N_27813);
and U30770 (N_30770,N_29883,N_29290);
nand U30771 (N_30771,N_26903,N_28484);
nor U30772 (N_30772,N_27329,N_26473);
nand U30773 (N_30773,N_28372,N_29057);
or U30774 (N_30774,N_28309,N_25597);
or U30775 (N_30775,N_27149,N_26912);
or U30776 (N_30776,N_29810,N_28592);
or U30777 (N_30777,N_26103,N_28764);
xor U30778 (N_30778,N_25674,N_26017);
xor U30779 (N_30779,N_25600,N_26659);
nor U30780 (N_30780,N_26740,N_27724);
nand U30781 (N_30781,N_26182,N_26966);
xnor U30782 (N_30782,N_29226,N_29622);
or U30783 (N_30783,N_28157,N_29669);
nand U30784 (N_30784,N_25842,N_28583);
nor U30785 (N_30785,N_25053,N_27415);
nand U30786 (N_30786,N_27378,N_27809);
or U30787 (N_30787,N_28278,N_28690);
or U30788 (N_30788,N_29103,N_26471);
nand U30789 (N_30789,N_29712,N_25220);
xor U30790 (N_30790,N_27159,N_27360);
nor U30791 (N_30791,N_27538,N_25475);
nor U30792 (N_30792,N_26222,N_29094);
or U30793 (N_30793,N_25224,N_27746);
nand U30794 (N_30794,N_27827,N_28513);
xnor U30795 (N_30795,N_27016,N_27069);
or U30796 (N_30796,N_28361,N_28359);
or U30797 (N_30797,N_25304,N_28207);
and U30798 (N_30798,N_28455,N_29640);
nand U30799 (N_30799,N_27591,N_26962);
nand U30800 (N_30800,N_28338,N_26528);
nand U30801 (N_30801,N_29124,N_29666);
nand U30802 (N_30802,N_25705,N_27920);
xor U30803 (N_30803,N_25027,N_28185);
nand U30804 (N_30804,N_29007,N_26416);
nor U30805 (N_30805,N_26815,N_26698);
nand U30806 (N_30806,N_26446,N_28852);
nand U30807 (N_30807,N_29511,N_27124);
nor U30808 (N_30808,N_28358,N_28532);
or U30809 (N_30809,N_27214,N_25088);
or U30810 (N_30810,N_26772,N_27764);
nor U30811 (N_30811,N_26273,N_29667);
or U30812 (N_30812,N_26381,N_27662);
and U30813 (N_30813,N_25119,N_26660);
nand U30814 (N_30814,N_27982,N_25987);
or U30815 (N_30815,N_28062,N_29956);
nor U30816 (N_30816,N_28921,N_27213);
or U30817 (N_30817,N_28516,N_29879);
and U30818 (N_30818,N_25912,N_25647);
xnor U30819 (N_30819,N_29908,N_25285);
or U30820 (N_30820,N_25254,N_28879);
and U30821 (N_30821,N_26521,N_29483);
nor U30822 (N_30822,N_25263,N_28813);
or U30823 (N_30823,N_27485,N_25235);
nor U30824 (N_30824,N_27924,N_28953);
nand U30825 (N_30825,N_25942,N_27342);
and U30826 (N_30826,N_26683,N_26758);
xor U30827 (N_30827,N_27361,N_28177);
nand U30828 (N_30828,N_28088,N_28679);
nand U30829 (N_30829,N_28113,N_26163);
nand U30830 (N_30830,N_27763,N_29950);
or U30831 (N_30831,N_26587,N_25342);
nor U30832 (N_30832,N_27820,N_28861);
nand U30833 (N_30833,N_29369,N_29409);
nand U30834 (N_30834,N_27232,N_26089);
nor U30835 (N_30835,N_27978,N_27176);
or U30836 (N_30836,N_28162,N_29000);
and U30837 (N_30837,N_27094,N_29927);
and U30838 (N_30838,N_26642,N_28030);
nand U30839 (N_30839,N_29070,N_26293);
and U30840 (N_30840,N_28544,N_27616);
nor U30841 (N_30841,N_27948,N_29996);
nand U30842 (N_30842,N_25353,N_27570);
nand U30843 (N_30843,N_25822,N_26126);
nor U30844 (N_30844,N_26637,N_26862);
nand U30845 (N_30845,N_27801,N_27448);
nand U30846 (N_30846,N_29430,N_27889);
nand U30847 (N_30847,N_26424,N_28311);
or U30848 (N_30848,N_26892,N_25959);
or U30849 (N_30849,N_26475,N_26357);
or U30850 (N_30850,N_26674,N_28289);
nor U30851 (N_30851,N_28160,N_26816);
or U30852 (N_30852,N_26959,N_25685);
nand U30853 (N_30853,N_27037,N_26883);
nand U30854 (N_30854,N_28161,N_29097);
nand U30855 (N_30855,N_29661,N_28496);
xnor U30856 (N_30856,N_25479,N_27878);
nor U30857 (N_30857,N_26232,N_26257);
xor U30858 (N_30858,N_29003,N_26353);
nand U30859 (N_30859,N_25474,N_28991);
xor U30860 (N_30860,N_29835,N_28798);
nor U30861 (N_30861,N_27500,N_25447);
or U30862 (N_30862,N_25515,N_29011);
nor U30863 (N_30863,N_27756,N_29767);
or U30864 (N_30864,N_28914,N_25287);
or U30865 (N_30865,N_28951,N_26607);
nor U30866 (N_30866,N_27194,N_25921);
and U30867 (N_30867,N_26478,N_29785);
or U30868 (N_30868,N_26950,N_26347);
nor U30869 (N_30869,N_25854,N_25608);
and U30870 (N_30870,N_27881,N_26769);
and U30871 (N_30871,N_29252,N_27593);
nor U30872 (N_30872,N_28570,N_26779);
and U30873 (N_30873,N_27697,N_27177);
xnor U30874 (N_30874,N_28115,N_28627);
xnor U30875 (N_30875,N_29707,N_25642);
nand U30876 (N_30876,N_28267,N_28328);
nor U30877 (N_30877,N_28107,N_28658);
and U30878 (N_30878,N_26879,N_25222);
nor U30879 (N_30879,N_25781,N_27462);
xnor U30880 (N_30880,N_27399,N_29171);
nor U30881 (N_30881,N_25093,N_28275);
nand U30882 (N_30882,N_27840,N_27116);
nand U30883 (N_30883,N_26955,N_26179);
xnor U30884 (N_30884,N_25519,N_28569);
nand U30885 (N_30885,N_25045,N_28849);
and U30886 (N_30886,N_27421,N_28986);
nor U30887 (N_30887,N_25043,N_25246);
or U30888 (N_30888,N_28836,N_28303);
and U30889 (N_30889,N_25113,N_29493);
or U30890 (N_30890,N_27657,N_25407);
or U30891 (N_30891,N_28384,N_26438);
xor U30892 (N_30892,N_25347,N_27755);
xor U30893 (N_30893,N_28247,N_29941);
and U30894 (N_30894,N_25487,N_28719);
or U30895 (N_30895,N_29626,N_26617);
and U30896 (N_30896,N_26468,N_26229);
nor U30897 (N_30897,N_26915,N_27654);
or U30898 (N_30898,N_25432,N_28722);
nor U30899 (N_30899,N_27291,N_26938);
and U30900 (N_30900,N_25678,N_29718);
or U30901 (N_30901,N_25957,N_26975);
xnor U30902 (N_30902,N_27186,N_26901);
nand U30903 (N_30903,N_27469,N_27038);
nand U30904 (N_30904,N_29575,N_28948);
nand U30905 (N_30905,N_27866,N_28150);
nand U30906 (N_30906,N_26128,N_29144);
and U30907 (N_30907,N_26594,N_27043);
and U30908 (N_30908,N_27302,N_28828);
xnor U30909 (N_30909,N_26727,N_26354);
nor U30910 (N_30910,N_27381,N_29137);
or U30911 (N_30911,N_27267,N_25410);
nand U30912 (N_30912,N_25746,N_25267);
and U30913 (N_30913,N_27384,N_28460);
and U30914 (N_30914,N_27789,N_27350);
and U30915 (N_30915,N_27250,N_29233);
xor U30916 (N_30916,N_26633,N_29779);
nor U30917 (N_30917,N_26635,N_28629);
nor U30918 (N_30918,N_27336,N_27311);
xor U30919 (N_30919,N_25682,N_26590);
or U30920 (N_30920,N_26147,N_29581);
and U30921 (N_30921,N_29506,N_28094);
or U30922 (N_30922,N_28616,N_25186);
and U30923 (N_30923,N_26689,N_25443);
or U30924 (N_30924,N_29146,N_27726);
and U30925 (N_30925,N_26619,N_29757);
or U30926 (N_30926,N_29194,N_28870);
nand U30927 (N_30927,N_26951,N_27864);
nand U30928 (N_30928,N_26820,N_29749);
and U30929 (N_30929,N_28510,N_25654);
or U30930 (N_30930,N_29088,N_26690);
or U30931 (N_30931,N_27723,N_29419);
and U30932 (N_30932,N_29211,N_27053);
and U30933 (N_30933,N_28316,N_25878);
or U30934 (N_30934,N_25709,N_28192);
or U30935 (N_30935,N_27403,N_27084);
nor U30936 (N_30936,N_29168,N_26906);
nor U30937 (N_30937,N_29651,N_26451);
and U30938 (N_30938,N_29087,N_29262);
nor U30939 (N_30939,N_27846,N_28083);
nor U30940 (N_30940,N_26329,N_26913);
and U30941 (N_30941,N_29346,N_26880);
nand U30942 (N_30942,N_29520,N_29203);
or U30943 (N_30943,N_29245,N_27986);
nor U30944 (N_30944,N_29998,N_26195);
and U30945 (N_30945,N_29988,N_27112);
and U30946 (N_30946,N_26448,N_27863);
and U30947 (N_30947,N_29484,N_26423);
xor U30948 (N_30948,N_26144,N_25868);
xnor U30949 (N_30949,N_29964,N_26079);
nand U30950 (N_30950,N_29064,N_25092);
nand U30951 (N_30951,N_27665,N_28555);
and U30952 (N_30952,N_28434,N_29200);
or U30953 (N_30953,N_28761,N_28614);
nor U30954 (N_30954,N_27156,N_25005);
nor U30955 (N_30955,N_28206,N_25526);
and U30956 (N_30956,N_27366,N_28956);
nand U30957 (N_30957,N_27679,N_28265);
or U30958 (N_30958,N_25791,N_28945);
or U30959 (N_30959,N_29432,N_26449);
or U30960 (N_30960,N_28408,N_26491);
nor U30961 (N_30961,N_28686,N_28776);
or U30962 (N_30962,N_26988,N_25231);
nand U30963 (N_30963,N_27760,N_28971);
nand U30964 (N_30964,N_28564,N_27238);
nand U30965 (N_30965,N_28128,N_25788);
nor U30966 (N_30966,N_25952,N_26292);
xnor U30967 (N_30967,N_25818,N_25672);
nor U30968 (N_30968,N_26489,N_28858);
nand U30969 (N_30969,N_27995,N_28791);
or U30970 (N_30970,N_29650,N_26430);
nand U30971 (N_30971,N_28415,N_26527);
nor U30972 (N_30972,N_25865,N_28214);
nand U30973 (N_30973,N_28790,N_25852);
nor U30974 (N_30974,N_26159,N_29032);
or U30975 (N_30975,N_25956,N_28606);
or U30976 (N_30976,N_29540,N_27511);
nor U30977 (N_30977,N_25160,N_26363);
and U30978 (N_30978,N_27792,N_29215);
xnor U30979 (N_30979,N_27635,N_27775);
nand U30980 (N_30980,N_29172,N_29161);
nand U30981 (N_30981,N_28550,N_28787);
or U30982 (N_30982,N_25706,N_26238);
nor U30983 (N_30983,N_27951,N_28947);
nand U30984 (N_30984,N_27471,N_25095);
xor U30985 (N_30985,N_26153,N_28571);
nor U30986 (N_30986,N_29263,N_26647);
nand U30987 (N_30987,N_27174,N_26682);
nand U30988 (N_30988,N_25170,N_26641);
and U30989 (N_30989,N_25806,N_26283);
or U30990 (N_30990,N_28831,N_27030);
nand U30991 (N_30991,N_25747,N_26996);
nand U30992 (N_30992,N_28221,N_26911);
nand U30993 (N_30993,N_26456,N_26652);
xnor U30994 (N_30994,N_27865,N_28689);
nand U30995 (N_30995,N_26884,N_25172);
or U30996 (N_30996,N_26132,N_27298);
nand U30997 (N_30997,N_26687,N_26327);
nand U30998 (N_30998,N_28528,N_27672);
or U30999 (N_30999,N_29154,N_27417);
nand U31000 (N_31000,N_29292,N_29524);
xnor U31001 (N_31001,N_27409,N_29571);
or U31002 (N_31002,N_26312,N_27819);
nor U31003 (N_31003,N_25244,N_27869);
nand U31004 (N_31004,N_26838,N_27001);
nand U31005 (N_31005,N_29298,N_26387);
and U31006 (N_31006,N_27106,N_29191);
nor U31007 (N_31007,N_27004,N_26418);
nand U31008 (N_31008,N_28381,N_29774);
nand U31009 (N_31009,N_25387,N_29769);
nor U31010 (N_31010,N_27443,N_27011);
nand U31011 (N_31011,N_29853,N_27687);
nor U31012 (N_31012,N_27718,N_29151);
nand U31013 (N_31013,N_26503,N_26930);
nor U31014 (N_31014,N_27917,N_26786);
nor U31015 (N_31015,N_25762,N_27198);
nor U31016 (N_31016,N_29902,N_28713);
and U31017 (N_31017,N_25326,N_27083);
nand U31018 (N_31018,N_27855,N_29812);
nor U31019 (N_31019,N_28093,N_25392);
or U31020 (N_31020,N_25767,N_25797);
nand U31021 (N_31021,N_25793,N_26487);
nand U31022 (N_31022,N_26808,N_27747);
or U31023 (N_31023,N_26202,N_29082);
or U31024 (N_31024,N_28653,N_25232);
xnor U31025 (N_31025,N_28337,N_28527);
and U31026 (N_31026,N_29180,N_27539);
nor U31027 (N_31027,N_26676,N_26902);
nand U31028 (N_31028,N_29903,N_27546);
xnor U31029 (N_31029,N_29554,N_28165);
xor U31030 (N_31030,N_26024,N_25834);
and U31031 (N_31031,N_25891,N_29231);
xor U31032 (N_31032,N_28104,N_26516);
nor U31033 (N_31033,N_28287,N_28079);
and U31034 (N_31034,N_25665,N_26549);
or U31035 (N_31035,N_25397,N_27825);
and U31036 (N_31036,N_29778,N_27938);
and U31037 (N_31037,N_29320,N_26771);
nand U31038 (N_31038,N_27088,N_25729);
or U31039 (N_31039,N_28444,N_29826);
nand U31040 (N_31040,N_28876,N_29664);
nor U31041 (N_31041,N_27848,N_25249);
nor U31042 (N_31042,N_27452,N_26768);
or U31043 (N_31043,N_28645,N_26640);
nor U31044 (N_31044,N_26783,N_28595);
and U31045 (N_31045,N_28035,N_25438);
xor U31046 (N_31046,N_27114,N_26253);
nand U31047 (N_31047,N_29347,N_28637);
or U31048 (N_31048,N_25240,N_25621);
and U31049 (N_31049,N_27092,N_27233);
nor U31050 (N_31050,N_25316,N_25469);
and U31051 (N_31051,N_29352,N_29079);
nand U31052 (N_31052,N_27681,N_27737);
and U31053 (N_31053,N_28401,N_29446);
nand U31054 (N_31054,N_25840,N_29099);
and U31055 (N_31055,N_29044,N_25361);
and U31056 (N_31056,N_29746,N_29523);
and U31057 (N_31057,N_28908,N_28136);
and U31058 (N_31058,N_26738,N_25279);
nor U31059 (N_31059,N_25218,N_27821);
nand U31060 (N_31060,N_29599,N_28619);
xnor U31061 (N_31061,N_28034,N_27822);
xnor U31062 (N_31062,N_25743,N_28551);
nand U31063 (N_31063,N_29256,N_26782);
and U31064 (N_31064,N_26165,N_28171);
nor U31065 (N_31065,N_26821,N_25405);
nor U31066 (N_31066,N_27286,N_26342);
xnor U31067 (N_31067,N_26826,N_27776);
nand U31068 (N_31068,N_25860,N_26290);
or U31069 (N_31069,N_27632,N_28369);
or U31070 (N_31070,N_28175,N_29470);
and U31071 (N_31071,N_27479,N_25184);
nor U31072 (N_31072,N_28693,N_29619);
xor U31073 (N_31073,N_26706,N_29910);
nor U31074 (N_31074,N_29616,N_26208);
nand U31075 (N_31075,N_29150,N_25547);
or U31076 (N_31076,N_29423,N_28952);
or U31077 (N_31077,N_28596,N_27042);
nand U31078 (N_31078,N_27858,N_28096);
nor U31079 (N_31079,N_27615,N_28631);
nor U31080 (N_31080,N_29174,N_28268);
xor U31081 (N_31081,N_27940,N_28215);
and U31082 (N_31082,N_28234,N_25133);
nor U31083 (N_31083,N_26138,N_27934);
and U31084 (N_31084,N_26665,N_25307);
nor U31085 (N_31085,N_28081,N_27521);
and U31086 (N_31086,N_25071,N_26931);
or U31087 (N_31087,N_29865,N_25457);
or U31088 (N_31088,N_28601,N_28716);
or U31089 (N_31089,N_27009,N_29065);
nand U31090 (N_31090,N_26694,N_26941);
or U31091 (N_31091,N_28158,N_29377);
nand U31092 (N_31092,N_26967,N_25223);
nor U31093 (N_31093,N_25835,N_28017);
nor U31094 (N_31094,N_27080,N_25318);
nand U31095 (N_31095,N_26129,N_28135);
and U31096 (N_31096,N_25180,N_27455);
xnor U31097 (N_31097,N_25188,N_29832);
nand U31098 (N_31098,N_27926,N_26705);
or U31099 (N_31099,N_28164,N_26703);
nand U31100 (N_31100,N_29281,N_26192);
or U31101 (N_31101,N_27592,N_28970);
nand U31102 (N_31102,N_29076,N_25760);
or U31103 (N_31103,N_27125,N_28625);
and U31104 (N_31104,N_29143,N_27203);
xor U31105 (N_31105,N_25716,N_25215);
nor U31106 (N_31106,N_28577,N_27205);
or U31107 (N_31107,N_25023,N_28866);
and U31108 (N_31108,N_26281,N_29675);
nand U31109 (N_31109,N_25893,N_29911);
xor U31110 (N_31110,N_25609,N_26076);
nand U31111 (N_31111,N_27828,N_26465);
nor U31112 (N_31112,N_29405,N_26871);
nand U31113 (N_31113,N_29472,N_28097);
nand U31114 (N_31114,N_27701,N_27206);
nand U31115 (N_31115,N_29401,N_28477);
and U31116 (N_31116,N_26953,N_25637);
and U31117 (N_31117,N_26648,N_25035);
nand U31118 (N_31118,N_26713,N_28933);
nor U31119 (N_31119,N_28299,N_26249);
nor U31120 (N_31120,N_27578,N_27451);
nand U31121 (N_31121,N_25401,N_26623);
nand U31122 (N_31122,N_27589,N_25801);
and U31123 (N_31123,N_25541,N_28850);
nand U31124 (N_31124,N_29106,N_28735);
nand U31125 (N_31125,N_25738,N_27633);
and U31126 (N_31126,N_28883,N_28169);
nor U31127 (N_31127,N_28306,N_25628);
xor U31128 (N_31128,N_27330,N_26850);
or U31129 (N_31129,N_26073,N_27749);
nand U31130 (N_31130,N_25260,N_26987);
or U31131 (N_31131,N_28110,N_27603);
nand U31132 (N_31132,N_28352,N_29434);
and U31133 (N_31133,N_26710,N_28893);
or U31134 (N_31134,N_25280,N_29073);
and U31135 (N_31135,N_27395,N_27309);
xor U31136 (N_31136,N_29397,N_29982);
xnor U31137 (N_31137,N_27999,N_29042);
or U31138 (N_31138,N_29577,N_26494);
nand U31139 (N_31139,N_29476,N_25356);
and U31140 (N_31140,N_28235,N_27942);
and U31141 (N_31141,N_28345,N_26454);
xor U31142 (N_31142,N_25078,N_29066);
or U31143 (N_31143,N_28771,N_27118);
nor U31144 (N_31144,N_26041,N_26276);
and U31145 (N_31145,N_29343,N_29743);
or U31146 (N_31146,N_28266,N_28640);
and U31147 (N_31147,N_29754,N_25266);
nor U31148 (N_31148,N_27432,N_27517);
nor U31149 (N_31149,N_29004,N_25683);
nor U31150 (N_31150,N_28501,N_25525);
or U31151 (N_31151,N_29720,N_26154);
nor U31152 (N_31152,N_28436,N_27663);
nor U31153 (N_31153,N_27241,N_27099);
nor U31154 (N_31154,N_29873,N_25971);
nand U31155 (N_31155,N_27040,N_27675);
and U31156 (N_31156,N_27306,N_28108);
xor U31157 (N_31157,N_26244,N_27265);
or U31158 (N_31158,N_27961,N_25671);
and U31159 (N_31159,N_28238,N_25082);
nand U31160 (N_31160,N_27255,N_29544);
and U31161 (N_31161,N_29980,N_27340);
nor U31162 (N_31162,N_29499,N_25888);
xor U31163 (N_31163,N_29663,N_26420);
xnor U31164 (N_31164,N_27505,N_29705);
nand U31165 (N_31165,N_26876,N_27411);
or U31166 (N_31166,N_29457,N_26308);
and U31167 (N_31167,N_27429,N_26437);
and U31168 (N_31168,N_29983,N_29272);
xnor U31169 (N_31169,N_25201,N_28741);
or U31170 (N_31170,N_28684,N_26169);
or U31171 (N_31171,N_26757,N_27564);
xnor U31172 (N_31172,N_27652,N_26230);
nand U31173 (N_31173,N_25689,N_27900);
or U31174 (N_31174,N_26514,N_27039);
or U31175 (N_31175,N_29022,N_25107);
or U31176 (N_31176,N_27879,N_26701);
nand U31177 (N_31177,N_25129,N_27402);
and U31178 (N_31178,N_29676,N_28750);
nor U31179 (N_31179,N_29657,N_29771);
nor U31180 (N_31180,N_25037,N_26948);
nor U31181 (N_31181,N_26847,N_27165);
nand U31182 (N_31182,N_26548,N_29006);
and U31183 (N_31183,N_28634,N_28127);
nand U31184 (N_31184,N_26571,N_29115);
nand U31185 (N_31185,N_25589,N_25451);
or U31186 (N_31186,N_27867,N_29691);
nor U31187 (N_31187,N_25115,N_29654);
nor U31188 (N_31188,N_26226,N_27427);
or U31189 (N_31189,N_28968,N_28898);
nor U31190 (N_31190,N_25492,N_29313);
xor U31191 (N_31191,N_25343,N_25374);
or U31192 (N_31192,N_28090,N_26612);
nor U31193 (N_31193,N_28531,N_27085);
xor U31194 (N_31194,N_28807,N_29866);
or U31195 (N_31195,N_26213,N_26219);
xor U31196 (N_31196,N_29904,N_25920);
xnor U31197 (N_31197,N_29228,N_28786);
and U31198 (N_31198,N_25384,N_29961);
or U31199 (N_31199,N_29549,N_25915);
nand U31200 (N_31200,N_28748,N_28566);
nor U31201 (N_31201,N_29868,N_27524);
and U31202 (N_31202,N_26534,N_28954);
and U31203 (N_31203,N_26917,N_27915);
xor U31204 (N_31204,N_26428,N_29328);
or U31205 (N_31205,N_28362,N_25616);
xor U31206 (N_31206,N_25409,N_25505);
or U31207 (N_31207,N_25651,N_28058);
nand U31208 (N_31208,N_25360,N_28179);
or U31209 (N_31209,N_28696,N_25902);
nand U31210 (N_31210,N_27910,N_28934);
nor U31211 (N_31211,N_29373,N_28507);
nand U31212 (N_31212,N_25312,N_25143);
nand U31213 (N_31213,N_29315,N_28392);
nor U31214 (N_31214,N_28322,N_27051);
or U31215 (N_31215,N_25253,N_28780);
nand U31216 (N_31216,N_27183,N_25250);
and U31217 (N_31217,N_29782,N_29002);
nor U31218 (N_31218,N_28142,N_28310);
or U31219 (N_31219,N_26864,N_27284);
or U31220 (N_31220,N_29596,N_25289);
and U31221 (N_31221,N_26890,N_25660);
and U31222 (N_31222,N_29984,N_26561);
and U31223 (N_31223,N_26337,N_27163);
or U31224 (N_31224,N_26282,N_26189);
nand U31225 (N_31225,N_25500,N_27439);
xor U31226 (N_31226,N_28174,N_28805);
nand U31227 (N_31227,N_27492,N_26952);
nand U31228 (N_31228,N_26784,N_26197);
nand U31229 (N_31229,N_26030,N_26799);
nand U31230 (N_31230,N_25553,N_28451);
and U31231 (N_31231,N_25428,N_29030);
and U31232 (N_31232,N_26218,N_27733);
nand U31233 (N_31233,N_27780,N_28205);
or U31234 (N_31234,N_27625,N_26535);
nand U31235 (N_31235,N_26719,N_27288);
nand U31236 (N_31236,N_29791,N_29408);
nand U31237 (N_31237,N_28468,N_28567);
and U31238 (N_31238,N_28782,N_25578);
and U31239 (N_31239,N_28418,N_28525);
nor U31240 (N_31240,N_28248,N_29084);
or U31241 (N_31241,N_27420,N_26181);
nand U31242 (N_31242,N_29358,N_29450);
or U31243 (N_31243,N_26763,N_29628);
xor U31244 (N_31244,N_28383,N_25704);
nand U31245 (N_31245,N_25293,N_26806);
nor U31246 (N_31246,N_29040,N_25679);
nor U31247 (N_31247,N_25204,N_28665);
and U31248 (N_31248,N_28024,N_28085);
and U31249 (N_31249,N_25980,N_29119);
or U31250 (N_31250,N_26600,N_29817);
or U31251 (N_31251,N_25352,N_25096);
nand U31252 (N_31252,N_27137,N_27161);
xnor U31253 (N_31253,N_25214,N_29533);
or U31254 (N_31254,N_26099,N_28979);
and U31255 (N_31255,N_25568,N_29224);
or U31256 (N_31256,N_26045,N_27573);
nand U31257 (N_31257,N_25193,N_29023);
nor U31258 (N_31258,N_29580,N_25625);
nor U31259 (N_31259,N_25355,N_26046);
and U31260 (N_31260,N_25135,N_28880);
nand U31261 (N_31261,N_25906,N_26168);
nor U31262 (N_31262,N_26575,N_25288);
or U31263 (N_31263,N_29894,N_26000);
or U31264 (N_31264,N_29318,N_29932);
or U31265 (N_31265,N_29102,N_28364);
nand U31266 (N_31266,N_26686,N_25910);
or U31267 (N_31267,N_25815,N_29750);
nor U31268 (N_31268,N_25194,N_27226);
nand U31269 (N_31269,N_29121,N_27262);
or U31270 (N_31270,N_26998,N_29960);
or U31271 (N_31271,N_29993,N_27401);
nand U31272 (N_31272,N_28037,N_25736);
and U31273 (N_31273,N_27551,N_28082);
nor U31274 (N_31274,N_25590,N_25399);
and U31275 (N_31275,N_28447,N_25484);
and U31276 (N_31276,N_25008,N_29207);
nor U31277 (N_31277,N_25191,N_28208);
nand U31278 (N_31278,N_27936,N_28681);
nand U31279 (N_31279,N_29739,N_29538);
or U31280 (N_31280,N_29216,N_25779);
and U31281 (N_31281,N_27470,N_29225);
nor U31282 (N_31282,N_28884,N_26627);
nor U31283 (N_31283,N_28259,N_27355);
or U31284 (N_31284,N_27682,N_27838);
and U31285 (N_31285,N_29253,N_29039);
and U31286 (N_31286,N_29641,N_27034);
or U31287 (N_31287,N_28422,N_27933);
nand U31288 (N_31288,N_27875,N_28881);
nand U31289 (N_31289,N_27797,N_27994);
or U31290 (N_31290,N_29797,N_28825);
or U31291 (N_31291,N_29142,N_25454);
or U31292 (N_31292,N_26750,N_25722);
nor U31293 (N_31293,N_29620,N_25811);
or U31294 (N_31294,N_27117,N_26458);
or U31295 (N_31295,N_28196,N_28218);
and U31296 (N_31296,N_27944,N_29709);
and U31297 (N_31297,N_25098,N_28046);
and U31298 (N_31298,N_25558,N_27565);
and U31299 (N_31299,N_29839,N_29731);
xor U31300 (N_31300,N_28641,N_29319);
nor U31301 (N_31301,N_28148,N_26199);
and U31302 (N_31302,N_26173,N_28351);
or U31303 (N_31303,N_29811,N_28466);
nor U31304 (N_31304,N_28002,N_28442);
and U31305 (N_31305,N_28847,N_27153);
or U31306 (N_31306,N_25431,N_25933);
and U31307 (N_31307,N_29049,N_27799);
and U31308 (N_31308,N_29410,N_27730);
nand U31309 (N_31309,N_27385,N_29170);
nand U31310 (N_31310,N_27930,N_28031);
or U31311 (N_31311,N_29989,N_27461);
nor U31312 (N_31312,N_25759,N_25968);
or U31313 (N_31313,N_28139,N_27476);
and U31314 (N_31314,N_27146,N_28076);
or U31315 (N_31315,N_25506,N_25973);
or U31316 (N_31316,N_25206,N_26662);
nor U31317 (N_31317,N_28817,N_25406);
or U31318 (N_31318,N_29081,N_25192);
nand U31319 (N_31319,N_28688,N_25338);
and U31320 (N_31320,N_27410,N_27777);
and U31321 (N_31321,N_27508,N_29059);
nor U31322 (N_31322,N_29247,N_27247);
nor U31323 (N_31323,N_28902,N_25695);
nand U31324 (N_31324,N_29985,N_27335);
xnor U31325 (N_31325,N_28229,N_26961);
and U31326 (N_31326,N_25234,N_28459);
nor U31327 (N_31327,N_25025,N_27006);
and U31328 (N_31328,N_29901,N_25904);
and U31329 (N_31329,N_29220,N_25219);
nor U31330 (N_31330,N_28727,N_28508);
nor U31331 (N_31331,N_27577,N_28862);
nor U31332 (N_31332,N_28615,N_26480);
xnor U31333 (N_31333,N_29729,N_29266);
nor U31334 (N_31334,N_25900,N_26856);
and U31335 (N_31335,N_26078,N_25895);
nor U31336 (N_31336,N_27528,N_25196);
or U31337 (N_31337,N_26832,N_27349);
nand U31338 (N_31338,N_28279,N_25724);
nor U31339 (N_31339,N_26027,N_28354);
nor U31340 (N_31340,N_25789,N_28172);
and U31341 (N_31341,N_26928,N_26186);
nor U31342 (N_31342,N_29128,N_27068);
and U31343 (N_31343,N_28842,N_26531);
nor U31344 (N_31344,N_28841,N_27246);
and U31345 (N_31345,N_25019,N_25954);
nor U31346 (N_31346,N_26059,N_25766);
or U31347 (N_31347,N_27164,N_26316);
and U31348 (N_31348,N_26869,N_29715);
and U31349 (N_31349,N_25430,N_28295);
or U31350 (N_31350,N_28060,N_29455);
xnor U31351 (N_31351,N_28102,N_29075);
xor U31352 (N_31352,N_28201,N_29784);
nor U31353 (N_31353,N_26404,N_29196);
or U31354 (N_31354,N_26314,N_29594);
nand U31355 (N_31355,N_25412,N_28896);
and U31356 (N_31356,N_29936,N_27945);
and U31357 (N_31357,N_25607,N_27102);
xnor U31358 (N_31358,N_27987,N_26204);
and U31359 (N_31359,N_26012,N_27199);
nor U31360 (N_31360,N_27850,N_26227);
nand U31361 (N_31361,N_26562,N_29987);
xnor U31362 (N_31362,N_26680,N_28609);
nand U31363 (N_31363,N_26785,N_27818);
nor U31364 (N_31364,N_28050,N_29798);
and U31365 (N_31365,N_27983,N_29123);
and U31366 (N_31366,N_29307,N_29824);
xor U31367 (N_31367,N_27503,N_29195);
or U31368 (N_31368,N_28659,N_25372);
nor U31369 (N_31369,N_28865,N_29273);
nor U31370 (N_31370,N_29799,N_26639);
nand U31371 (N_31371,N_27139,N_29417);
or U31372 (N_31372,N_27595,N_29836);
nand U31373 (N_31373,N_25943,N_25698);
and U31374 (N_31374,N_27567,N_25633);
and U31375 (N_31375,N_27338,N_26206);
or U31376 (N_31376,N_28159,N_25131);
xor U31377 (N_31377,N_27115,N_29486);
nor U31378 (N_31378,N_25551,N_27765);
nand U31379 (N_31379,N_25314,N_29354);
xor U31380 (N_31380,N_26220,N_27498);
or U31381 (N_31381,N_27251,N_26224);
or U31382 (N_31382,N_26133,N_27169);
and U31383 (N_31383,N_26040,N_26233);
nor U31384 (N_31384,N_27041,N_29425);
or U31385 (N_31385,N_26626,N_27433);
or U31386 (N_31386,N_27316,N_25354);
and U31387 (N_31387,N_29371,N_27263);
or U31388 (N_31388,N_27661,N_27640);
nand U31389 (N_31389,N_25205,N_29818);
or U31390 (N_31390,N_26356,N_26196);
nor U31391 (N_31391,N_27036,N_25021);
or U31392 (N_31392,N_26405,N_28210);
and U31393 (N_31393,N_27704,N_27680);
and U31394 (N_31394,N_28963,N_25208);
or U31395 (N_31395,N_25494,N_26485);
nand U31396 (N_31396,N_26949,N_27467);
or U31397 (N_31397,N_27985,N_28173);
nand U31398 (N_31398,N_29634,N_25527);
and U31399 (N_31399,N_28225,N_28394);
nor U31400 (N_31400,N_28774,N_28572);
nand U31401 (N_31401,N_25394,N_27572);
nand U31402 (N_31402,N_27870,N_27323);
xor U31403 (N_31403,N_29801,N_27394);
and U31404 (N_31404,N_26824,N_27773);
or U31405 (N_31405,N_25491,N_26216);
nand U31406 (N_31406,N_26289,N_28407);
and U31407 (N_31407,N_26343,N_28263);
or U31408 (N_31408,N_29198,N_29162);
or U31409 (N_31409,N_25629,N_29576);
nor U31410 (N_31410,N_28190,N_28724);
nor U31411 (N_31411,N_27647,N_26260);
nand U31412 (N_31412,N_25460,N_26335);
xnor U31413 (N_31413,N_27890,N_29212);
nor U31414 (N_31414,N_27388,N_27293);
or U31415 (N_31415,N_28644,N_28156);
or U31416 (N_31416,N_28336,N_26483);
and U31417 (N_31417,N_29717,N_29035);
or U31418 (N_31418,N_26157,N_26620);
xnor U31419 (N_31419,N_26277,N_29202);
nand U31420 (N_31420,N_27167,N_26102);
and U31421 (N_31421,N_28985,N_26852);
nand U31422 (N_31422,N_26899,N_29109);
and U31423 (N_31423,N_25147,N_26893);
nand U31424 (N_31424,N_28464,N_25542);
and U31425 (N_31425,N_29302,N_25761);
nor U31426 (N_31426,N_27190,N_28495);
nand U31427 (N_31427,N_27173,N_27931);
xnor U31428 (N_31428,N_27494,N_27758);
or U31429 (N_31429,N_27276,N_28966);
nor U31430 (N_31430,N_27109,N_29356);
nor U31431 (N_31431,N_25268,N_29807);
and U31432 (N_31432,N_26529,N_26348);
nand U31433 (N_31433,N_26774,N_25668);
and U31434 (N_31434,N_29054,N_26840);
or U31435 (N_31435,N_28182,N_29080);
xnor U31436 (N_31436,N_27543,N_26296);
and U31437 (N_31437,N_29872,N_29411);
nor U31438 (N_31438,N_28155,N_25535);
or U31439 (N_31439,N_28453,N_26324);
nor U31440 (N_31440,N_29572,N_29644);
and U31441 (N_31441,N_27144,N_29805);
nor U31442 (N_31442,N_29973,N_27430);
nor U31443 (N_31443,N_25828,N_28255);
and U31444 (N_31444,N_29464,N_27729);
and U31445 (N_31445,N_25423,N_29463);
and U31446 (N_31446,N_26557,N_26614);
nand U31447 (N_31447,N_27628,N_27007);
or U31448 (N_31448,N_28005,N_27750);
nand U31449 (N_31449,N_26835,N_25844);
or U31450 (N_31450,N_26513,N_25584);
nand U31451 (N_31451,N_28340,N_26258);
nor U31452 (N_31452,N_28241,N_29337);
or U31453 (N_31453,N_26060,N_28553);
nor U31454 (N_31454,N_28258,N_27817);
nor U31455 (N_31455,N_25236,N_27899);
nand U31456 (N_31456,N_26742,N_27677);
and U31457 (N_31457,N_29943,N_27000);
and U31458 (N_31458,N_28374,N_26601);
nor U31459 (N_31459,N_29105,N_28846);
nor U31460 (N_31460,N_27605,N_28602);
nand U31461 (N_31461,N_25114,N_25570);
nand U31462 (N_31462,N_28636,N_28432);
xor U31463 (N_31463,N_28678,N_26688);
nor U31464 (N_31464,N_29221,N_28506);
and U31465 (N_31465,N_29167,N_26021);
nor U31466 (N_31466,N_27962,N_27976);
or U31467 (N_31467,N_25014,N_28410);
nor U31468 (N_31468,N_29864,N_26203);
nor U31469 (N_31469,N_25996,N_28887);
and U31470 (N_31470,N_29237,N_25054);
xor U31471 (N_31471,N_25550,N_27440);
nor U31472 (N_31472,N_29703,N_26095);
or U31473 (N_31473,N_29728,N_28469);
and U31474 (N_31474,N_27074,N_25981);
xnor U31475 (N_31475,N_26152,N_29460);
nor U31476 (N_31476,N_29773,N_27894);
nand U31477 (N_31477,N_27876,N_26242);
and U31478 (N_31478,N_25531,N_28792);
or U31479 (N_31479,N_27529,N_27170);
nand U31480 (N_31480,N_29722,N_27658);
or U31481 (N_31481,N_27499,N_28272);
xor U31482 (N_31482,N_27230,N_26069);
or U31483 (N_31483,N_29140,N_26547);
or U31484 (N_31484,N_27277,N_29402);
nor U31485 (N_31485,N_25923,N_29209);
nand U31486 (N_31486,N_25393,N_26845);
and U31487 (N_31487,N_29611,N_29385);
nand U31488 (N_31488,N_27535,N_26891);
nor U31489 (N_31489,N_26874,N_26131);
nand U31490 (N_31490,N_28568,N_26467);
or U31491 (N_31491,N_29261,N_28803);
nor U31492 (N_31492,N_29497,N_25862);
or U31493 (N_31493,N_26781,N_26309);
nand U31494 (N_31494,N_25402,N_26588);
or U31495 (N_31495,N_27090,N_26166);
xor U31496 (N_31496,N_29736,N_26338);
nand U31497 (N_31497,N_27072,N_25273);
xor U31498 (N_31498,N_29107,N_27988);
nand U31499 (N_31499,N_25690,N_29665);
nand U31500 (N_31500,N_28103,N_28143);
and U31501 (N_31501,N_27831,N_28180);
nor U31502 (N_31502,N_28137,N_25029);
nand U31503 (N_31503,N_29643,N_26476);
nand U31504 (N_31504,N_28224,N_27073);
or U31505 (N_31505,N_28598,N_28809);
or U31506 (N_31506,N_27969,N_25400);
or U31507 (N_31507,N_26331,N_28994);
and U31508 (N_31508,N_29850,N_29556);
and U31509 (N_31509,N_29967,N_25774);
and U31510 (N_31510,N_29699,N_28851);
nor U31511 (N_31511,N_27618,N_28624);
or U31512 (N_31512,N_26795,N_25557);
nand U31513 (N_31513,N_26307,N_27282);
nor U31514 (N_31514,N_27541,N_26700);
nor U31515 (N_31515,N_28376,N_26960);
or U31516 (N_31516,N_25708,N_27534);
nor U31517 (N_31517,N_28586,N_28895);
and U31518 (N_31518,N_29673,N_28885);
and U31519 (N_31519,N_25221,N_27382);
or U31520 (N_31520,N_28589,N_27303);
and U31521 (N_31521,N_26096,N_25264);
and U31522 (N_31522,N_28478,N_25640);
nor U31523 (N_31523,N_29629,N_27020);
and U31524 (N_31524,N_26065,N_27803);
nor U31525 (N_31525,N_27753,N_28471);
nor U31526 (N_31526,N_26366,N_25958);
and U31527 (N_31527,N_27685,N_25063);
xor U31528 (N_31528,N_26735,N_27504);
nor U31529 (N_31529,N_29104,N_28233);
nor U31530 (N_31530,N_29453,N_26447);
nor U31531 (N_31531,N_26813,N_28778);
nor U31532 (N_31532,N_26450,N_27328);
nand U31533 (N_31533,N_27807,N_29312);
and U31534 (N_31534,N_28660,N_25424);
or U31535 (N_31535,N_29390,N_27859);
nand U31536 (N_31536,N_28972,N_28704);
nand U31537 (N_31537,N_27127,N_28040);
xnor U31538 (N_31538,N_27414,N_26402);
nor U31539 (N_31539,N_28321,N_28260);
nand U31540 (N_31540,N_25183,N_29822);
and U31541 (N_31541,N_25148,N_29869);
nor U31542 (N_31542,N_29036,N_28138);
nor U31543 (N_31543,N_29532,N_27619);
and U31544 (N_31544,N_27014,N_28411);
and U31545 (N_31545,N_29693,N_27450);
and U31546 (N_31546,N_27673,N_25758);
nor U31547 (N_31547,N_27741,N_28486);
nand U31548 (N_31548,N_27404,N_29566);
xor U31549 (N_31549,N_25661,N_26522);
xor U31550 (N_31550,N_28649,N_28691);
or U31551 (N_31551,N_27245,N_26927);
nand U31552 (N_31552,N_26708,N_29968);
and U31553 (N_31553,N_28476,N_25572);
and U31554 (N_31554,N_26504,N_29436);
nor U31555 (N_31555,N_26211,N_29680);
or U31556 (N_31556,N_28784,N_27396);
nor U31557 (N_31557,N_25776,N_25929);
or U31558 (N_31558,N_28742,N_28068);
or U31559 (N_31559,N_27391,N_26773);
nand U31560 (N_31560,N_29847,N_27695);
or U31561 (N_31561,N_26007,N_26885);
or U31562 (N_31562,N_26291,N_25111);
nor U31563 (N_31563,N_29608,N_25362);
or U31564 (N_31564,N_25501,N_26981);
or U31565 (N_31565,N_28243,N_25229);
or U31566 (N_31566,N_25605,N_28072);
or U31567 (N_31567,N_27560,N_27327);
and U31568 (N_31568,N_29489,N_25999);
nand U31569 (N_31569,N_25851,N_28236);
or U31570 (N_31570,N_28554,N_27320);
nor U31571 (N_31571,N_27216,N_29555);
nand U31572 (N_31572,N_27438,N_28674);
nor U31573 (N_31573,N_26164,N_27946);
and U31574 (N_31574,N_29545,N_27002);
and U31575 (N_31575,N_29301,N_27022);
nor U31576 (N_31576,N_28981,N_25816);
and U31577 (N_31577,N_27784,N_27905);
xor U31578 (N_31578,N_26756,N_25162);
or U31579 (N_31579,N_26863,N_29093);
nand U31580 (N_31580,N_27189,N_26577);
and U31581 (N_31581,N_28890,N_29308);
or U31582 (N_31582,N_26466,N_29842);
nor U31583 (N_31583,N_28959,N_25463);
nand U31584 (N_31584,N_26807,N_27537);
and U31585 (N_31585,N_25465,N_25381);
nand U31586 (N_31586,N_29952,N_28481);
and U31587 (N_31587,N_28350,N_28461);
or U31588 (N_31588,N_29515,N_26170);
and U31589 (N_31589,N_25485,N_27324);
nand U31590 (N_31590,N_29522,N_29238);
or U31591 (N_31591,N_25831,N_27475);
nand U31592 (N_31592,N_25796,N_26551);
nand U31593 (N_31593,N_25742,N_25284);
xor U31594 (N_31594,N_26036,N_27122);
xor U31595 (N_31595,N_25497,N_27599);
nand U31596 (N_31596,N_26425,N_27029);
nor U31597 (N_31597,N_26741,N_26565);
and U31598 (N_31598,N_25327,N_28779);
nor U31599 (N_31599,N_29687,N_26486);
nor U31600 (N_31600,N_28894,N_28231);
nor U31601 (N_31601,N_29948,N_25091);
or U31602 (N_31602,N_29503,N_26764);
xnor U31603 (N_31603,N_29753,N_26190);
or U31604 (N_31604,N_25648,N_25983);
or U31605 (N_31605,N_25691,N_25701);
or U31606 (N_31606,N_25894,N_25464);
xnor U31607 (N_31607,N_26412,N_28834);
and U31608 (N_31608,N_26777,N_27949);
nand U31609 (N_31609,N_26063,N_25586);
and U31610 (N_31610,N_27305,N_29623);
or U31611 (N_31611,N_26104,N_28320);
nand U31612 (N_31612,N_27734,N_26117);
or U31613 (N_31613,N_29056,N_25732);
xor U31614 (N_31614,N_29165,N_26344);
nand U31615 (N_31615,N_28939,N_26142);
and U31616 (N_31616,N_29806,N_26744);
xnor U31617 (N_31617,N_27722,N_28630);
xnor U31618 (N_31618,N_26723,N_27496);
nor U31619 (N_31619,N_26436,N_29537);
nand U31620 (N_31620,N_26935,N_29602);
nor U31621 (N_31621,N_25061,N_26673);
nand U31622 (N_31622,N_27980,N_27604);
nand U31623 (N_31623,N_27829,N_28593);
or U31624 (N_31624,N_26728,N_25559);
or U31625 (N_31625,N_25230,N_28726);
nor U31626 (N_31626,N_25677,N_28827);
nand U31627 (N_31627,N_26375,N_29424);
nor U31628 (N_31628,N_29636,N_29283);
or U31629 (N_31629,N_28086,N_29473);
nand U31630 (N_31630,N_26087,N_27140);
and U31631 (N_31631,N_27191,N_26958);
xnor U31632 (N_31632,N_29783,N_26712);
and U31633 (N_31633,N_27035,N_29512);
nand U31634 (N_31634,N_26837,N_29260);
nand U31635 (N_31635,N_26322,N_28349);
nor U31636 (N_31636,N_29692,N_25039);
nor U31637 (N_31637,N_28198,N_27768);
and U31638 (N_31638,N_26897,N_29158);
nor U31639 (N_31639,N_26039,N_29820);
nor U31640 (N_31640,N_28239,N_25800);
nor U31641 (N_31641,N_27195,N_26829);
nand U31642 (N_31642,N_26088,N_29398);
nand U31643 (N_31643,N_28832,N_28147);
nor U31644 (N_31644,N_28439,N_25512);
and U31645 (N_31645,N_25319,N_25580);
or U31646 (N_31646,N_29543,N_25348);
nand U31647 (N_31647,N_25666,N_28277);
and U31648 (N_31648,N_26732,N_26441);
and U31649 (N_31649,N_27005,N_28197);
nand U31650 (N_31650,N_27794,N_25276);
xnor U31651 (N_31651,N_26939,N_29244);
nand U31652 (N_31652,N_28756,N_27873);
nand U31653 (N_31653,N_26511,N_28608);
nand U31654 (N_31654,N_28228,N_25073);
and U31655 (N_31655,N_28814,N_29603);
and U31656 (N_31656,N_29701,N_28119);
and U31657 (N_31657,N_28621,N_29462);
nand U31658 (N_31658,N_29230,N_28711);
nand U31659 (N_31659,N_25972,N_27231);
and U31660 (N_31660,N_26231,N_29258);
nor U31661 (N_31661,N_27711,N_27545);
and U31662 (N_31662,N_28739,N_26650);
nor U31663 (N_31663,N_25446,N_28488);
nor U31664 (N_31664,N_27977,N_25898);
nor U31665 (N_31665,N_27018,N_26578);
xnor U31666 (N_31666,N_29615,N_26618);
nand U31667 (N_31667,N_28980,N_27778);
and U31668 (N_31668,N_26266,N_29117);
and U31669 (N_31669,N_27559,N_26455);
or U31670 (N_31670,N_26991,N_28473);
and U31671 (N_31671,N_25385,N_26288);
and U31672 (N_31672,N_27319,N_28802);
and U31673 (N_31673,N_28419,N_28363);
nor U31674 (N_31674,N_25653,N_25974);
or U31675 (N_31675,N_26751,N_25275);
nor U31676 (N_31676,N_25790,N_26814);
nor U31677 (N_31677,N_29440,N_25763);
nand U31678 (N_31678,N_28022,N_28216);
nand U31679 (N_31679,N_28220,N_27495);
nor U31680 (N_31680,N_29831,N_29846);
nand U31681 (N_31681,N_28670,N_27912);
and U31682 (N_31682,N_27871,N_29550);
nor U31683 (N_31683,N_29466,N_26914);
nor U31684 (N_31684,N_26031,N_25619);
and U31685 (N_31685,N_26585,N_27089);
and U31686 (N_31686,N_27583,N_28911);
or U31687 (N_31687,N_28385,N_26980);
xnor U31688 (N_31688,N_29413,N_25846);
and U31689 (N_31689,N_26887,N_29364);
nor U31690 (N_31690,N_25871,N_29752);
or U31691 (N_31691,N_26115,N_28751);
xnor U31692 (N_31692,N_25386,N_26346);
nand U31693 (N_31693,N_26851,N_26319);
or U31694 (N_31694,N_26848,N_25833);
or U31695 (N_31695,N_28646,N_25964);
nor U31696 (N_31696,N_25583,N_28131);
xor U31697 (N_31697,N_25085,N_25657);
or U31698 (N_31698,N_28978,N_29607);
or U31699 (N_31699,N_29204,N_29917);
and U31700 (N_31700,N_27830,N_26359);
nor U31701 (N_31701,N_28292,N_28009);
nand U31702 (N_31702,N_25450,N_29800);
nor U31703 (N_31703,N_25594,N_29300);
xnor U31704 (N_31704,N_26586,N_29282);
nor U31705 (N_31705,N_26597,N_26858);
nor U31706 (N_31706,N_28556,N_26711);
xnor U31707 (N_31707,N_29275,N_28534);
nor U31708 (N_31708,N_27056,N_26497);
or U31709 (N_31709,N_25812,N_29361);
and U31710 (N_31710,N_26355,N_29169);
nor U31711 (N_31711,N_25786,N_28001);
nand U31712 (N_31712,N_29959,N_28514);
nand U31713 (N_31713,N_29303,N_26507);
or U31714 (N_31714,N_25504,N_29724);
or U31715 (N_31715,N_29770,N_28697);
nand U31716 (N_31716,N_29021,N_28984);
nor U31717 (N_31717,N_26509,N_28962);
and U31718 (N_31718,N_28517,N_27322);
nor U31719 (N_31719,N_26362,N_28041);
nand U31720 (N_31720,N_26999,N_27839);
xor U31721 (N_31721,N_29870,N_25617);
nor U31722 (N_31722,N_25239,N_27808);
nand U31723 (N_31723,N_26145,N_25168);
xor U31724 (N_31724,N_26278,N_27532);
nor U31725 (N_31725,N_25864,N_27484);
or U31726 (N_31726,N_29630,N_27235);
and U31727 (N_31727,N_29443,N_29605);
or U31728 (N_31728,N_29997,N_29217);
or U31729 (N_31729,N_25885,N_28276);
and U31730 (N_31730,N_26655,N_25948);
xnor U31731 (N_31731,N_27626,N_25185);
nand U31732 (N_31732,N_28958,N_28924);
nor U31733 (N_31733,N_29946,N_27371);
and U31734 (N_31734,N_26239,N_27515);
nand U31735 (N_31735,N_29357,N_26080);
nand U31736 (N_31736,N_25787,N_27024);
xor U31737 (N_31737,N_25998,N_29330);
nand U31738 (N_31738,N_26101,N_27031);
or U31739 (N_31739,N_25528,N_27510);
or U31740 (N_31740,N_25144,N_28254);
nand U31741 (N_31741,N_26609,N_25687);
and U31742 (N_31742,N_28123,N_28427);
nand U31743 (N_31743,N_29060,N_26408);
nor U31744 (N_31744,N_28042,N_28930);
xor U31745 (N_31745,N_27474,N_27771);
or U31746 (N_31746,N_28940,N_26049);
nor U31747 (N_31747,N_29765,N_28462);
nor U31748 (N_31748,N_26843,N_26445);
or U31749 (N_31749,N_26002,N_27390);
or U31750 (N_31750,N_28456,N_25125);
or U31751 (N_31751,N_25308,N_26888);
nand U31752 (N_31752,N_25907,N_29875);
or U31753 (N_31753,N_29246,N_28799);
and U31754 (N_31754,N_25863,N_25277);
or U31755 (N_31755,N_25163,N_26403);
nand U31756 (N_31756,N_29403,N_28242);
or U31757 (N_31757,N_26759,N_27757);
and U31758 (N_31758,N_29501,N_29441);
and U31759 (N_31759,N_26140,N_27321);
nand U31760 (N_31760,N_28769,N_26500);
nor U31761 (N_31761,N_25190,N_29444);
or U31762 (N_31762,N_27348,N_29393);
xnor U31763 (N_31763,N_25696,N_26567);
nand U31764 (N_31764,N_27579,N_27021);
or U31765 (N_31765,N_26765,N_29026);
and U31766 (N_31766,N_27358,N_25034);
xnor U31767 (N_31767,N_29711,N_25022);
nand U31768 (N_31768,N_27918,N_29662);
or U31769 (N_31769,N_28753,N_28700);
and U31770 (N_31770,N_26611,N_29480);
nor U31771 (N_31771,N_25480,N_28509);
xor U31772 (N_31772,N_25498,N_29668);
nor U31773 (N_31773,N_26185,N_27172);
nor U31774 (N_31774,N_28873,N_28935);
or U31775 (N_31775,N_25686,N_28661);
or U31776 (N_31776,N_27964,N_28187);
xnor U31777 (N_31777,N_26982,N_28720);
nand U31778 (N_31778,N_27196,N_26866);
and U31779 (N_31779,N_29825,N_26019);
and U31780 (N_31780,N_27334,N_29598);
xor U31781 (N_31781,N_27209,N_28070);
and U31782 (N_31782,N_27208,N_26388);
xnor U31783 (N_31783,N_26943,N_29788);
nor U31784 (N_31784,N_25908,N_28988);
xor U31785 (N_31785,N_28633,N_26217);
and U31786 (N_31786,N_29670,N_25773);
or U31787 (N_31787,N_25772,N_26672);
nor U31788 (N_31788,N_26581,N_28793);
and U31789 (N_31789,N_26390,N_25602);
nor U31790 (N_31790,N_29924,N_29601);
nor U31791 (N_31791,N_25548,N_29618);
nand U31792 (N_31792,N_28856,N_26989);
or U31793 (N_31793,N_27913,N_27824);
nand U31794 (N_31794,N_27239,N_26094);
nor U31795 (N_31795,N_29981,N_29896);
and U31796 (N_31796,N_25158,N_29053);
or U31797 (N_31797,N_26250,N_29496);
nand U31798 (N_31798,N_29679,N_26050);
nand U31799 (N_31799,N_26544,N_28732);
or U31800 (N_31800,N_28327,N_29037);
and U31801 (N_31801,N_27308,N_26584);
and U31802 (N_31802,N_29920,N_28874);
xnor U31803 (N_31803,N_27923,N_29681);
nand U31804 (N_31804,N_26472,N_28463);
or U31805 (N_31805,N_25768,N_26207);
and U31806 (N_31806,N_26492,N_25116);
nand U31807 (N_31807,N_25867,N_25367);
nand U31808 (N_31808,N_29384,N_29189);
nor U31809 (N_31809,N_29597,N_25662);
xnor U31810 (N_31810,N_26734,N_27646);
nand U31811 (N_31811,N_28200,N_25914);
and U31812 (N_31812,N_29780,N_26789);
and U31813 (N_31813,N_29349,N_29363);
or U31814 (N_31814,N_28928,N_26921);
and U31815 (N_31815,N_28431,N_29069);
and U31816 (N_31816,N_25995,N_28728);
and U31817 (N_31817,N_25644,N_27132);
or U31818 (N_31818,N_28632,N_26081);
xor U31819 (N_31819,N_29589,N_25735);
or U31820 (N_31820,N_25046,N_26008);
or U31821 (N_31821,N_28212,N_27407);
nor U31822 (N_31822,N_27622,N_25300);
nor U31823 (N_31823,N_29447,N_25749);
xnor U31824 (N_31824,N_28578,N_26725);
and U31825 (N_31825,N_29507,N_25702);
xnor U31826 (N_31826,N_27569,N_27998);
or U31827 (N_31827,N_25118,N_27364);
nand U31828 (N_31828,N_29655,N_29257);
and U31829 (N_31829,N_29259,N_27493);
xor U31830 (N_31830,N_29157,N_29738);
and U31831 (N_31831,N_28176,N_29652);
nand U31832 (N_31832,N_26696,N_28482);
nand U31833 (N_31833,N_28949,N_26841);
nand U31834 (N_31834,N_27575,N_25663);
and U31835 (N_31835,N_29055,N_27168);
xnor U31836 (N_31836,N_26681,N_29759);
nor U31837 (N_31837,N_29421,N_27872);
nor U31838 (N_31838,N_28794,N_28294);
or U31839 (N_31839,N_29025,N_26645);
and U31840 (N_31840,N_28909,N_29086);
or U31841 (N_31841,N_28511,N_29471);
nor U31842 (N_31842,N_27712,N_29900);
nand U31843 (N_31843,N_29878,N_27707);
xnor U31844 (N_31844,N_25161,N_27258);
nand U31845 (N_31845,N_27841,N_25301);
or U31846 (N_31846,N_26122,N_26541);
or U31847 (N_31847,N_26300,N_26983);
or U31848 (N_31848,N_26325,N_25257);
xnor U31849 (N_31849,N_25011,N_29067);
xnor U31850 (N_31850,N_28734,N_25142);
nand U31851 (N_31851,N_25099,N_25905);
and U31852 (N_31852,N_27660,N_28325);
and U31853 (N_31853,N_27064,N_29741);
nor U31854 (N_31854,N_25804,N_29813);
and U31855 (N_31855,N_29306,N_26026);
nor U31856 (N_31856,N_25302,N_26628);
nor U31857 (N_31857,N_29595,N_27782);
nand U31858 (N_31858,N_27260,N_27990);
and U31859 (N_31859,N_27184,N_27048);
or U31860 (N_31860,N_28409,N_29024);
nor U31861 (N_31861,N_28011,N_25077);
or U31862 (N_31862,N_25649,N_25297);
nor U31863 (N_31863,N_26857,N_29931);
nor U31864 (N_31864,N_27606,N_27290);
nor U31865 (N_31865,N_28652,N_25634);
xnor U31866 (N_31866,N_26004,N_28291);
nor U31867 (N_31867,N_26802,N_27279);
and U31868 (N_31868,N_25199,N_25282);
nand U31869 (N_31869,N_25103,N_27974);
and U31870 (N_31870,N_26490,N_26697);
or U31871 (N_31871,N_25656,N_28346);
nor U31872 (N_31872,N_26545,N_28882);
nand U31873 (N_31873,N_28623,N_29995);
or U31874 (N_31874,N_27386,N_27070);
or U31875 (N_31875,N_28343,N_25476);
nor U31876 (N_31876,N_29481,N_25334);
or U31877 (N_31877,N_29482,N_28487);
nand U31878 (N_31878,N_29438,N_27692);
xnor U31879 (N_31879,N_28737,N_26280);
xor U31880 (N_31880,N_28380,N_28440);
nand U31881 (N_31881,N_27561,N_26038);
or U31882 (N_31882,N_27811,N_26940);
nor U31883 (N_31883,N_27555,N_28379);
or U31884 (N_31884,N_27058,N_25798);
nor U31885 (N_31885,N_25181,N_28274);
xor U31886 (N_31886,N_27694,N_28965);
nor U31887 (N_31887,N_26714,N_25069);
and U31888 (N_31888,N_27731,N_27783);
and U31889 (N_31889,N_29122,N_25676);
nand U31890 (N_31890,N_25380,N_26589);
and U31891 (N_31891,N_28560,N_25936);
or U31892 (N_31892,N_29940,N_26761);
and U31893 (N_31893,N_28133,N_26330);
or U31894 (N_31894,N_29458,N_27795);
xnor U31895 (N_31895,N_29928,N_26822);
and U31896 (N_31896,N_28989,N_27130);
or U31897 (N_31897,N_25876,N_25286);
nor U31898 (N_31898,N_27814,N_26693);
nor U31899 (N_31899,N_28541,N_29977);
nand U31900 (N_31900,N_29090,N_28388);
or U31901 (N_31901,N_28367,N_29208);
xor U31902 (N_31902,N_28253,N_25516);
nor U31903 (N_31903,N_28059,N_27032);
or U31904 (N_31904,N_27991,N_27526);
xnor U31905 (N_31905,N_26414,N_26100);
and U31906 (N_31906,N_26109,N_26003);
or U31907 (N_31907,N_25946,N_27611);
nand U31908 (N_31908,N_26867,N_29745);
nor U31909 (N_31909,N_29214,N_26141);
and U31910 (N_31910,N_27907,N_25315);
or U31911 (N_31911,N_26488,N_27531);
and U31912 (N_31912,N_27223,N_25753);
or U31913 (N_31913,N_25950,N_25283);
or U31914 (N_31914,N_25620,N_26533);
nor U31915 (N_31915,N_27071,N_29845);
and U31916 (N_31916,N_28186,N_26400);
and U31917 (N_31917,N_25826,N_29898);
xor U31918 (N_31918,N_27925,N_29159);
or U31919 (N_31919,N_29490,N_26736);
or U31920 (N_31920,N_25985,N_29560);
nor U31921 (N_31921,N_27845,N_28111);
and U31922 (N_31922,N_28543,N_28663);
and U31923 (N_31923,N_29375,N_26978);
nor U31924 (N_31924,N_28806,N_28146);
nand U31925 (N_31925,N_26011,N_25596);
nand U31926 (N_31926,N_26493,N_26919);
xor U31927 (N_31927,N_28626,N_29880);
or U31928 (N_31928,N_28638,N_27458);
nand U31929 (N_31929,N_26304,N_25592);
or U31930 (N_31930,N_28004,N_29958);
nand U31931 (N_31931,N_26836,N_26798);
xnor U31932 (N_31932,N_28329,N_26413);
nor U31933 (N_31933,N_25058,N_29751);
and U31934 (N_31934,N_29218,N_27596);
or U31935 (N_31935,N_26502,N_28048);
or U31936 (N_31936,N_27435,N_25916);
nand U31937 (N_31937,N_29017,N_26463);
or U31938 (N_31938,N_27045,N_26106);
and U31939 (N_31939,N_26125,N_25294);
xor U31940 (N_31940,N_25440,N_26137);
nor U31941 (N_31941,N_26947,N_27374);
and U31942 (N_31942,N_28203,N_25265);
nand U31943 (N_31943,N_25870,N_28522);
or U31944 (N_31944,N_29559,N_26110);
nand U31945 (N_31945,N_29925,N_29359);
and U31946 (N_31946,N_25603,N_28580);
nand U31947 (N_31947,N_26477,N_27816);
or U31948 (N_31948,N_27131,N_27893);
nor U31949 (N_31949,N_26209,N_26677);
and U31950 (N_31950,N_26929,N_29386);
and U31951 (N_31951,N_26119,N_25502);
and U31952 (N_31952,N_29897,N_27155);
nand U31953 (N_31953,N_25038,N_27690);
or U31954 (N_31954,N_28333,N_29077);
and U31955 (N_31955,N_25233,N_25101);
or U31956 (N_31956,N_27107,N_25425);
or U31957 (N_31957,N_25311,N_25370);
and U31958 (N_31958,N_26889,N_27044);
nand U31959 (N_31959,N_25631,N_28332);
nand U31960 (N_31960,N_29683,N_28223);
or U31961 (N_31961,N_27217,N_27060);
nand U31962 (N_31962,N_25324,N_27950);
nand U31963 (N_31963,N_29028,N_25281);
nand U31964 (N_31964,N_25509,N_26526);
and U31965 (N_31965,N_29962,N_25187);
xor U31966 (N_31966,N_27887,N_29808);
xnor U31967 (N_31967,N_25741,N_28526);
xnor U31968 (N_31968,N_27929,N_28535);
and U31969 (N_31969,N_29201,N_29647);
and U31970 (N_31970,N_27932,N_29485);
and U31971 (N_31971,N_28342,N_28839);
nor U31972 (N_31972,N_27506,N_26971);
and U31973 (N_31973,N_27580,N_27188);
or U31974 (N_31974,N_25567,N_26382);
xnor U31975 (N_31975,N_28695,N_26287);
nor U31976 (N_31976,N_26904,N_27568);
and U31977 (N_31977,N_25153,N_29823);
nand U31978 (N_31978,N_29682,N_29558);
or U31979 (N_31979,N_29614,N_28283);
and U31980 (N_31980,N_29761,N_27788);
nor U31981 (N_31981,N_27224,N_25614);
or U31982 (N_31982,N_28612,N_29406);
or U31983 (N_31983,N_27880,N_29899);
or U31984 (N_31984,N_27121,N_29243);
nand U31985 (N_31985,N_28256,N_26350);
or U31986 (N_31986,N_25984,N_28820);
xor U31987 (N_31987,N_26323,N_28777);
and U31988 (N_31988,N_27082,N_25418);
and U31989 (N_31989,N_27851,N_29376);
or U31990 (N_31990,N_27666,N_26801);
and U31991 (N_31991,N_26035,N_26223);
nand U31992 (N_31992,N_26944,N_27434);
nor U31993 (N_31993,N_26791,N_27597);
nand U31994 (N_31994,N_27406,N_25462);
nand U31995 (N_31995,N_25899,N_28375);
nand U31996 (N_31996,N_29974,N_27197);
xor U31997 (N_31997,N_28703,N_29183);
or U31998 (N_31998,N_25481,N_29926);
nor U31999 (N_31999,N_25415,N_29127);
nor U32000 (N_32000,N_27136,N_26523);
and U32001 (N_32001,N_27901,N_25890);
nor U32002 (N_32002,N_29418,N_26668);
and U32003 (N_32003,N_27922,N_26112);
nand U32004 (N_32004,N_29130,N_29592);
or U32005 (N_32005,N_28950,N_25997);
nand U32006 (N_32006,N_27586,N_28548);
nor U32007 (N_32007,N_27123,N_25075);
xor U32008 (N_32008,N_29794,N_29700);
nand U32009 (N_32009,N_28725,N_26563);
nand U32010 (N_32010,N_27351,N_26787);
nor U32011 (N_32011,N_27668,N_29491);
and U32012 (N_32012,N_25169,N_29205);
nor U32013 (N_32013,N_25652,N_25441);
and U32014 (N_32014,N_27536,N_27519);
or U32015 (N_32015,N_28230,N_27699);
or U32016 (N_32016,N_27636,N_27192);
or U32017 (N_32017,N_27370,N_26752);
nor U32018 (N_32018,N_26716,N_25299);
or U32019 (N_32019,N_26525,N_27691);
nand U32020 (N_32020,N_28437,N_29186);
nand U32021 (N_32021,N_27275,N_29858);
xor U32022 (N_32022,N_25122,N_26178);
nand U32023 (N_32023,N_27769,N_29089);
nor U32024 (N_32024,N_27686,N_26920);
nor U32025 (N_32025,N_28020,N_27651);
or U32026 (N_32026,N_27436,N_27178);
nand U32027 (N_32027,N_29697,N_25782);
or U32028 (N_32028,N_29487,N_25363);
xor U32029 (N_32029,N_29514,N_29474);
nor U32030 (N_32030,N_25079,N_25979);
and U32031 (N_32031,N_26373,N_27079);
and U32032 (N_32032,N_25827,N_27921);
or U32033 (N_32033,N_28600,N_27868);
or U32034 (N_32034,N_25488,N_28758);
xor U32035 (N_32035,N_27629,N_29206);
and U32036 (N_32036,N_25123,N_27617);
nor U32037 (N_32037,N_28465,N_28692);
and U32038 (N_32038,N_26995,N_27463);
nor U32039 (N_32039,N_26894,N_28643);
and U32040 (N_32040,N_25435,N_25830);
and U32041 (N_32041,N_29182,N_25203);
nor U32042 (N_32042,N_25341,N_25309);
nand U32043 (N_32043,N_28731,N_26896);
and U32044 (N_32044,N_25994,N_27885);
or U32045 (N_32045,N_25693,N_25411);
and U32046 (N_32046,N_26262,N_26396);
nand U32047 (N_32047,N_29291,N_25305);
and U32048 (N_32048,N_26334,N_28891);
nand U32049 (N_32049,N_26055,N_27914);
nor U32050 (N_32050,N_25565,N_29734);
and U32051 (N_32051,N_26333,N_29468);
or U32052 (N_32052,N_28489,N_25379);
nor U32053 (N_32053,N_26421,N_29588);
nor U32054 (N_32054,N_26360,N_29587);
and U32055 (N_32055,N_29942,N_25076);
or U32056 (N_32056,N_29068,N_25934);
nand U32057 (N_32057,N_26748,N_28144);
nor U32058 (N_32058,N_26111,N_27449);
nand U32059 (N_32059,N_25845,N_29264);
and U32060 (N_32060,N_29139,N_25802);
or U32061 (N_32061,N_28122,N_29344);
nand U32062 (N_32062,N_28008,N_25514);
nor U32063 (N_32063,N_26877,N_28168);
xor U32064 (N_32064,N_26235,N_28425);
nand U32065 (N_32065,N_25566,N_27269);
xor U32066 (N_32066,N_26532,N_27466);
nand U32067 (N_32067,N_26556,N_27292);
and U32068 (N_32068,N_25520,N_27772);
nand U32069 (N_32069,N_27507,N_28520);
nand U32070 (N_32070,N_27502,N_27478);
nor U32071 (N_32071,N_28130,N_27509);
xnor U32072 (N_32072,N_26630,N_26827);
nor U32073 (N_32073,N_27010,N_26184);
nand U32074 (N_32074,N_26608,N_25562);
nand U32075 (N_32075,N_28736,N_25991);
or U32076 (N_32076,N_27678,N_25295);
or U32077 (N_32077,N_25909,N_27096);
xor U32078 (N_32078,N_27714,N_28597);
nand U32079 (N_32079,N_27341,N_25606);
nand U32080 (N_32080,N_28458,N_27530);
and U32081 (N_32081,N_26846,N_27119);
and U32082 (N_32082,N_25176,N_27790);
nor U32083 (N_32083,N_27013,N_29145);
xor U32084 (N_32084,N_25345,N_28901);
nand U32085 (N_32085,N_28100,N_25839);
xnor U32086 (N_32086,N_29379,N_28840);
nor U32087 (N_32087,N_27362,N_28819);
nor U32088 (N_32088,N_26909,N_29184);
xnor U32089 (N_32089,N_29706,N_27902);
nor U32090 (N_32090,N_27135,N_25328);
or U32091 (N_32091,N_25351,N_27713);
or U32092 (N_32092,N_26598,N_28946);
nor U32093 (N_32093,N_25202,N_25534);
nand U32094 (N_32094,N_27670,N_25003);
or U32095 (N_32095,N_26146,N_28860);
and U32096 (N_32096,N_27735,N_27919);
nand U32097 (N_32097,N_28330,N_25544);
nor U32098 (N_32098,N_27634,N_29742);
nand U32099 (N_32099,N_26746,N_29796);
nand U32100 (N_32100,N_27162,N_26709);
nor U32101 (N_32101,N_26780,N_28014);
nand U32102 (N_32102,N_25433,N_26582);
xnor U32103 (N_32103,N_25364,N_28326);
or U32104 (N_32104,N_25794,N_25066);
or U32105 (N_32105,N_29129,N_28812);
nor U32106 (N_32106,N_29704,N_25571);
nand U32107 (N_32107,N_28151,N_29331);
or U32108 (N_32108,N_26070,N_26121);
or U32109 (N_32109,N_27274,N_28195);
nand U32110 (N_32110,N_29152,N_26518);
or U32111 (N_32111,N_26933,N_26591);
nand U32112 (N_32112,N_27052,N_28261);
or U32113 (N_32113,N_29048,N_25369);
xnor U32114 (N_32114,N_27105,N_25331);
nand U32115 (N_32115,N_28286,N_25783);
or U32116 (N_32116,N_28246,N_27706);
nand U32117 (N_32117,N_28282,N_29016);
nor U32118 (N_32118,N_26644,N_25444);
nor U32119 (N_32119,N_26692,N_29029);
and U32120 (N_32120,N_29332,N_26058);
and U32121 (N_32121,N_26305,N_28145);
or U32122 (N_32122,N_25731,N_29574);
or U32123 (N_32123,N_29287,N_25106);
nand U32124 (N_32124,N_26968,N_29249);
xnor U32125 (N_32125,N_26254,N_26134);
or U32126 (N_32126,N_28281,N_29222);
nand U32127 (N_32127,N_26717,N_29125);
or U32128 (N_32128,N_29072,N_25259);
nand U32129 (N_32129,N_29632,N_29043);
and U32130 (N_32130,N_25670,N_25564);
xor U32131 (N_32131,N_28204,N_29110);
and U32132 (N_32132,N_29631,N_27075);
nor U32133 (N_32133,N_28871,N_26130);
nand U32134 (N_32134,N_28744,N_28539);
xor U32135 (N_32135,N_26954,N_26624);
nor U32136 (N_32136,N_26804,N_29834);
and U32137 (N_32137,N_25298,N_26391);
or U32138 (N_32138,N_28854,N_26702);
or U32139 (N_32139,N_25227,N_29309);
or U32140 (N_32140,N_26313,N_29840);
and U32141 (N_32141,N_25524,N_25321);
and U32142 (N_32142,N_27693,N_28913);
nor U32143 (N_32143,N_26747,N_27927);
xnor U32144 (N_32144,N_26970,N_29990);
nand U32145 (N_32145,N_27653,N_29420);
nand U32146 (N_32146,N_29014,N_27447);
nand U32147 (N_32147,N_27066,N_27160);
and U32148 (N_32148,N_27800,N_26386);
or U32149 (N_32149,N_26107,N_25332);
nand U32150 (N_32150,N_29710,N_26510);
nor U32151 (N_32151,N_28723,N_29949);
nor U32152 (N_32152,N_29953,N_28816);
nor U32153 (N_32153,N_25417,N_26384);
and U32154 (N_32154,N_28540,N_28992);
nand U32155 (N_32155,N_28969,N_25769);
nand U32156 (N_32156,N_26539,N_29101);
or U32157 (N_32157,N_29795,N_29427);
nand U32158 (N_32158,N_29951,N_29382);
or U32159 (N_32159,N_25483,N_27477);
or U32160 (N_32160,N_29255,N_25545);
nor U32161 (N_32161,N_27852,N_26797);
or U32162 (N_32162,N_27620,N_28781);
or U32163 (N_32163,N_27588,N_29155);
nor U32164 (N_32164,N_28389,N_25006);
nor U32165 (N_32165,N_28757,N_27972);
or U32166 (N_32166,N_28089,N_28285);
xnor U32167 (N_32167,N_26093,N_26023);
nand U32168 (N_32168,N_26135,N_25020);
or U32169 (N_32169,N_29578,N_28443);
nand U32170 (N_32170,N_27975,N_28925);
or U32171 (N_32171,N_29339,N_25127);
or U32172 (N_32172,N_28353,N_26064);
nor U32173 (N_32173,N_27423,N_27721);
nand U32174 (N_32174,N_25490,N_25814);
and U32175 (N_32175,N_29316,N_25805);
and U32176 (N_32176,N_29748,N_29521);
xnor U32177 (N_32177,N_29336,N_26865);
nor U32178 (N_32178,N_27015,N_27970);
xor U32179 (N_32179,N_27295,N_28273);
xor U32180 (N_32180,N_26279,N_26755);
or U32181 (N_32181,N_26228,N_28293);
nor U32182 (N_32182,N_28822,N_25650);
nor U32183 (N_32183,N_27971,N_28357);
or U32184 (N_32184,N_28618,N_26957);
nand U32185 (N_32185,N_26733,N_28995);
or U32186 (N_32186,N_25752,N_25680);
or U32187 (N_32187,N_25458,N_28313);
nor U32188 (N_32188,N_26392,N_29519);
or U32189 (N_32189,N_29012,N_26245);
xnor U32190 (N_32190,N_26770,N_25472);
or U32191 (N_32191,N_29437,N_26376);
and U32192 (N_32192,N_27581,N_28694);
or U32193 (N_32193,N_27992,N_28424);
xor U32194 (N_32194,N_25897,N_25258);
or U32195 (N_32195,N_25110,N_26264);
nand U32196 (N_32196,N_26559,N_27857);
or U32197 (N_32197,N_27294,N_25403);
and U32198 (N_32198,N_29889,N_28717);
xor U32199 (N_32199,N_27650,N_27087);
nand U32200 (N_32200,N_25556,N_27244);
nand U32201 (N_32201,N_28582,N_28446);
and U32202 (N_32202,N_26394,N_28317);
xor U32203 (N_32203,N_28420,N_27248);
or U32204 (N_32204,N_29882,N_26139);
nor U32205 (N_32205,N_29933,N_27095);
and U32206 (N_32206,N_26162,N_27310);
and U32207 (N_32207,N_29721,N_25669);
xor U32208 (N_32208,N_27398,N_25368);
or U32209 (N_32209,N_27892,N_25961);
nor U32210 (N_32210,N_29136,N_29992);
and U32211 (N_32211,N_29031,N_28944);
xnor U32212 (N_32212,N_25518,N_26934);
nand U32213 (N_32213,N_26086,N_26530);
nand U32214 (N_32214,N_25859,N_26029);
or U32215 (N_32215,N_26200,N_29439);
nor U32216 (N_32216,N_29033,N_28504);
and U32217 (N_32217,N_25951,N_25339);
and U32218 (N_32218,N_27612,N_25989);
nor U32219 (N_32219,N_27715,N_27257);
nand U32220 (N_32220,N_25613,N_27996);
nand U32221 (N_32221,N_25778,N_25949);
and U32222 (N_32222,N_29083,N_28622);
xor U32223 (N_32223,N_25322,N_29492);
and U32224 (N_32224,N_29431,N_25155);
nand U32225 (N_32225,N_27512,N_26739);
xnor U32226 (N_32226,N_28957,N_26385);
and U32227 (N_32227,N_28997,N_26328);
xor U32228 (N_32228,N_25848,N_27301);
and U32229 (N_32229,N_29534,N_25359);
or U32230 (N_32230,N_25437,N_27332);
or U32231 (N_32231,N_25817,N_28382);
or U32232 (N_32232,N_28124,N_26077);
nor U32233 (N_32233,N_26014,N_29351);
nor U32234 (N_32234,N_28416,N_29994);
xnor U32235 (N_32235,N_25292,N_29562);
or U32236 (N_32236,N_29591,N_25636);
xor U32237 (N_32237,N_26859,N_25718);
nor U32238 (N_32238,N_25711,N_26161);
nand U32239 (N_32239,N_25540,N_26269);
and U32240 (N_32240,N_26977,N_27683);
nor U32241 (N_32241,N_28687,N_27906);
nand U32242 (N_32242,N_27973,N_28886);
nor U32243 (N_32243,N_28955,N_28454);
and U32244 (N_32244,N_25784,N_26658);
nor U32245 (N_32245,N_25200,N_28975);
nand U32246 (N_32246,N_29610,N_25927);
nand U32247 (N_32247,N_26722,N_25618);
nor U32248 (N_32248,N_26123,N_25068);
nand U32249 (N_32249,N_26443,N_26898);
or U32250 (N_32250,N_27272,N_27416);
nor U32251 (N_32251,N_27667,N_29885);
and U32252 (N_32252,N_27669,N_25358);
nor U32253 (N_32253,N_29311,N_26636);
and U32254 (N_32254,N_27958,N_25470);
xor U32255 (N_32255,N_26295,N_25734);
and U32256 (N_32256,N_29310,N_28007);
nand U32257 (N_32257,N_26936,N_28654);
or U32258 (N_32258,N_26923,N_25382);
or U32259 (N_32259,N_25255,N_25508);
or U32260 (N_32260,N_28855,N_27249);
nor U32261 (N_32261,N_29178,N_25171);
nor U32262 (N_32262,N_28421,N_28538);
nor U32263 (N_32263,N_27798,N_29646);
or U32264 (N_32264,N_27562,N_29829);
or U32265 (N_32265,N_25408,N_28390);
nor U32266 (N_32266,N_25554,N_29173);
nor U32267 (N_32267,N_29886,N_27955);
or U32268 (N_32268,N_26964,N_27422);
nand U32269 (N_32269,N_29539,N_28497);
nor U32270 (N_32270,N_29176,N_28671);
and U32271 (N_32271,N_29895,N_27607);
nand U32272 (N_32272,N_25262,N_28305);
nand U32273 (N_32273,N_26434,N_28033);
or U32274 (N_32274,N_29561,N_28098);
or U32275 (N_32275,N_26248,N_28536);
nor U32276 (N_32276,N_28931,N_28183);
or U32277 (N_32277,N_27787,N_25396);
xnor U32278 (N_32278,N_25866,N_29986);
xor U32279 (N_32279,N_29304,N_28552);
nor U32280 (N_32280,N_28545,N_29781);
and U32281 (N_32281,N_27444,N_29525);
nor U32282 (N_32282,N_25453,N_28710);
xnor U32283 (N_32283,N_25459,N_29871);
and U32284 (N_32284,N_28472,N_28500);
xor U32285 (N_32285,N_28937,N_28404);
and U32286 (N_32286,N_26439,N_29188);
nor U32287 (N_32287,N_27491,N_27023);
and U32288 (N_32288,N_25938,N_26775);
and U32289 (N_32289,N_25645,N_28923);
and U32290 (N_32290,N_25134,N_26965);
and U32291 (N_32291,N_25913,N_27552);
and U32292 (N_32292,N_28708,N_25228);
nor U32293 (N_32293,N_28824,N_29837);
nor U32294 (N_32294,N_26479,N_28915);
and U32295 (N_32295,N_26926,N_29095);
xor U32296 (N_32296,N_28775,N_28474);
or U32297 (N_32297,N_29370,N_25655);
xor U32298 (N_32298,N_29677,N_27883);
xnor U32299 (N_32299,N_28056,N_28859);
or U32300 (N_32300,N_25853,N_28423);
nor U32301 (N_32301,N_27158,N_29672);
nand U32302 (N_32302,N_29366,N_27643);
xor U32303 (N_32303,N_28810,N_28184);
nand U32304 (N_32304,N_29383,N_29649);
or U32305 (N_32305,N_28315,N_29637);
and U32306 (N_32306,N_29340,N_27501);
or U32307 (N_32307,N_26160,N_26349);
nor U32308 (N_32308,N_25398,N_27941);
xnor U32309 (N_32309,N_27212,N_27126);
nand U32310 (N_32310,N_25577,N_26205);
or U32311 (N_32311,N_26873,N_28899);
and U32312 (N_32312,N_29527,N_27523);
nand U32313 (N_32313,N_27522,N_29254);
nand U32314 (N_32314,N_28976,N_27337);
nand U32315 (N_32315,N_29392,N_25496);
and U32316 (N_32316,N_27952,N_29766);
nor U32317 (N_32317,N_25552,N_25271);
nor U32318 (N_32318,N_25059,N_25090);
xnor U32319 (N_32319,N_26580,N_26501);
and U32320 (N_32320,N_25585,N_25261);
nor U32321 (N_32321,N_26704,N_29517);
or U32322 (N_32322,N_29528,N_26720);
and U32323 (N_32323,N_26524,N_26183);
nand U32324 (N_32324,N_26812,N_28767);
and U32325 (N_32325,N_26310,N_27273);
nor U32326 (N_32326,N_25426,N_27550);
nor U32327 (N_32327,N_26247,N_27065);
nand U32328 (N_32328,N_28973,N_27621);
and U32329 (N_32329,N_26536,N_25140);
nand U32330 (N_32330,N_29762,N_28457);
xor U32331 (N_32331,N_29844,N_25375);
and U32332 (N_32332,N_25576,N_25089);
and U32333 (N_32333,N_26495,N_29970);
or U32334 (N_32334,N_29355,N_26605);
nand U32335 (N_32335,N_26508,N_28811);
nor U32336 (N_32336,N_25033,N_25404);
xor U32337 (N_32337,N_28667,N_27413);
xor U32338 (N_32338,N_25536,N_26028);
nand U32339 (N_32339,N_28837,N_26188);
or U32340 (N_32340,N_29939,N_25032);
nor U32341 (N_32341,N_29133,N_27312);
nand U32342 (N_32342,N_27437,N_27793);
nand U32343 (N_32343,N_27896,N_25579);
nand U32344 (N_32344,N_28872,N_26984);
xnor U32345 (N_32345,N_27767,N_25917);
nor U32346 (N_32346,N_25466,N_29428);
nor U32347 (N_32347,N_29642,N_25511);
nand U32348 (N_32348,N_26922,N_28747);
and U32349 (N_32349,N_29929,N_25449);
and U32350 (N_32350,N_28863,N_29854);
and U32351 (N_32351,N_28252,N_29789);
and U32352 (N_32352,N_27372,N_27751);
and U32353 (N_32353,N_26422,N_28666);
nand U32354 (N_32354,N_27441,N_28365);
and U32355 (N_32355,N_28099,N_27558);
nand U32356 (N_32356,N_28845,N_26415);
or U32357 (N_32357,N_26849,N_25664);
and U32358 (N_32358,N_26057,N_25414);
nor U32359 (N_32359,N_29504,N_29278);
or U32360 (N_32360,N_26364,N_28650);
nand U32361 (N_32361,N_25269,N_26116);
nor U32362 (N_32362,N_25918,N_27218);
nor U32363 (N_32363,N_29045,N_29010);
nor U32364 (N_32364,N_25004,N_27609);
and U32365 (N_32365,N_29389,N_25546);
nand U32366 (N_32366,N_27271,N_29148);
or U32367 (N_32367,N_29975,N_29270);
nand U32368 (N_32368,N_28869,N_28095);
nand U32369 (N_32369,N_25975,N_29141);
xnor U32370 (N_32370,N_29020,N_27154);
or U32371 (N_32371,N_28217,N_28804);
nor U32372 (N_32372,N_26666,N_26749);
and U32373 (N_32373,N_28864,N_28677);
or U32374 (N_32374,N_29177,N_25886);
nand U32375 (N_32375,N_26275,N_28038);
and U32376 (N_32376,N_27585,N_29565);
and U32377 (N_32377,N_26061,N_27225);
nor U32378 (N_32378,N_27935,N_25889);
nand U32379 (N_32379,N_28025,N_27698);
nor U32380 (N_32380,N_27836,N_25744);
or U32381 (N_32381,N_27856,N_29841);
nand U32382 (N_32382,N_28101,N_25924);
nor U32383 (N_32383,N_26895,N_27242);
xnor U32384 (N_32384,N_26583,N_27720);
or U32385 (N_32385,N_27017,N_27655);
and U32386 (N_32386,N_29695,N_25429);
nor U32387 (N_32387,N_25139,N_25154);
and U32388 (N_32388,N_28449,N_26010);
or U32389 (N_32389,N_27748,N_29991);
and U32390 (N_32390,N_26006,N_26251);
or U32391 (N_32391,N_27345,N_28134);
nand U32392 (N_32392,N_25697,N_28918);
nand U32393 (N_32393,N_25723,N_25001);
nor U32394 (N_32394,N_27837,N_29976);
nor U32395 (N_32395,N_29323,N_28450);
or U32396 (N_32396,N_27202,N_29909);
nand U32397 (N_32397,N_29621,N_28907);
or U32398 (N_32398,N_26419,N_27897);
nor U32399 (N_32399,N_26819,N_25156);
xnor U32400 (N_32400,N_29625,N_28302);
or U32401 (N_32401,N_28106,N_26399);
nand U32402 (N_32402,N_26656,N_25157);
nor U32403 (N_32403,N_29096,N_29551);
xnor U32404 (N_32404,N_26564,N_29689);
xnor U32405 (N_32405,N_28087,N_29513);
nand U32406 (N_32406,N_26908,N_29735);
nand U32407 (N_32407,N_28105,N_26699);
and U32408 (N_32408,N_29567,N_27968);
nor U32409 (N_32409,N_27895,N_29293);
xnor U32410 (N_32410,N_28010,N_25615);
nor U32411 (N_32411,N_26715,N_25198);
nand U32412 (N_32412,N_25574,N_29372);
nand U32413 (N_32413,N_29126,N_25713);
and U32414 (N_32414,N_25117,N_29407);
or U32415 (N_32415,N_26193,N_26345);
nor U32416 (N_32416,N_29934,N_29147);
and U32417 (N_32417,N_25195,N_29744);
nand U32418 (N_32418,N_29600,N_26299);
or U32419 (N_32419,N_27826,N_25391);
nor U32420 (N_32420,N_28319,N_26573);
or U32421 (N_32421,N_27832,N_27630);
nor U32422 (N_32422,N_27228,N_29322);
and U32423 (N_32423,N_27193,N_26048);
nand U32424 (N_32424,N_26651,N_25138);
nand U32425 (N_32425,N_28244,N_29830);
nand U32426 (N_32426,N_27928,N_28519);
xnor U32427 (N_32427,N_28245,N_26517);
and U32428 (N_32428,N_25109,N_27641);
xnor U32429 (N_32429,N_27835,N_27143);
nor U32430 (N_32430,N_26976,N_29500);
or U32431 (N_32431,N_29399,N_29768);
nand U32432 (N_32432,N_25448,N_27904);
nor U32433 (N_32433,N_26265,N_25346);
or U32434 (N_32434,N_26148,N_28121);
nor U32435 (N_32435,N_26481,N_27676);
nor U32436 (N_32436,N_25388,N_29747);
and U32437 (N_32437,N_29947,N_25843);
nor U32438 (N_32438,N_27861,N_26788);
nor U32439 (N_32439,N_27252,N_29648);
or U32440 (N_32440,N_28620,N_25489);
nor U32441 (N_32441,N_29542,N_26643);
or U32442 (N_32442,N_27261,N_26127);
nor U32443 (N_32443,N_25881,N_29265);
nor U32444 (N_32444,N_29181,N_28604);
and U32445 (N_32445,N_29299,N_29192);
nor U32446 (N_32446,N_25044,N_25930);
and U32447 (N_32447,N_29725,N_28574);
and U32448 (N_32448,N_28304,N_26177);
or U32449 (N_32449,N_28324,N_26613);
or U32450 (N_32450,N_25823,N_25306);
nand U32451 (N_32451,N_26606,N_26649);
xor U32452 (N_32452,N_27898,N_29969);
xnor U32453 (N_32453,N_29790,N_27645);
or U32454 (N_32454,N_29179,N_26596);
nor U32455 (N_32455,N_25993,N_27059);
nand U32456 (N_32456,N_27339,N_25755);
nor U32457 (N_32457,N_25771,N_27812);
nor U32458 (N_32458,N_27363,N_29388);
nor U32459 (N_32459,N_28607,N_27739);
and U32460 (N_32460,N_25623,N_28698);
nor U32461 (N_32461,N_27590,N_26084);
or U32462 (N_32462,N_27026,N_28611);
or U32463 (N_32463,N_28154,N_29862);
and U32464 (N_32464,N_29459,N_26124);
xor U32465 (N_32465,N_27460,N_27702);
and U32466 (N_32466,N_25707,N_25241);
and U32467 (N_32467,N_28412,N_26956);
nand U32468 (N_32468,N_29242,N_26604);
nand U32469 (N_32469,N_25303,N_29639);
nand U32470 (N_32470,N_27097,N_25591);
and U32471 (N_32471,N_25688,N_29085);
and U32472 (N_32472,N_26120,N_27369);
and U32473 (N_32473,N_28707,N_25159);
nand U32474 (N_32474,N_28092,N_27979);
or U32475 (N_32475,N_29338,N_27916);
and U32476 (N_32476,N_26072,N_25009);
xor U32477 (N_32477,N_29062,N_29286);
nand U32478 (N_32478,N_27740,N_26860);
nor U32479 (N_32479,N_27847,N_26255);
nor U32480 (N_32480,N_26306,N_27953);
nor U32481 (N_32481,N_28537,N_28788);
nor U32482 (N_32482,N_29978,N_25024);
nor U32483 (N_32483,N_25970,N_29116);
nor U32484 (N_32484,N_27028,N_25925);
xnor U32485 (N_32485,N_28961,N_28977);
and U32486 (N_32486,N_28403,N_25189);
nand U32487 (N_32487,N_26037,N_26155);
nand U32488 (N_32488,N_28492,N_25177);
and U32489 (N_32489,N_25780,N_26963);
nor U32490 (N_32490,N_25807,N_29536);
and U32491 (N_32491,N_29454,N_28613);
nor U32492 (N_32492,N_26411,N_26409);
and U32493 (N_32493,N_29518,N_26365);
nor U32494 (N_32494,N_26191,N_25130);
xnor U32495 (N_32495,N_28112,N_28227);
nor U32496 (N_32496,N_25167,N_28815);
and U32497 (N_32497,N_27405,N_25986);
and U32498 (N_32498,N_28057,N_28826);
or U32499 (N_32499,N_29884,N_26113);
nand U32500 (N_32500,N_29497,N_29897);
nand U32501 (N_32501,N_27389,N_26674);
nor U32502 (N_32502,N_28531,N_25554);
and U32503 (N_32503,N_25739,N_29053);
or U32504 (N_32504,N_25222,N_26638);
and U32505 (N_32505,N_27979,N_25597);
xor U32506 (N_32506,N_28709,N_26332);
and U32507 (N_32507,N_29156,N_27603);
nand U32508 (N_32508,N_27534,N_29136);
nor U32509 (N_32509,N_27097,N_26863);
or U32510 (N_32510,N_29290,N_25345);
and U32511 (N_32511,N_29854,N_25224);
and U32512 (N_32512,N_28897,N_25912);
nor U32513 (N_32513,N_26775,N_27621);
nor U32514 (N_32514,N_29865,N_25388);
nand U32515 (N_32515,N_29349,N_27662);
nor U32516 (N_32516,N_25262,N_28588);
nor U32517 (N_32517,N_29491,N_25958);
or U32518 (N_32518,N_29772,N_28311);
and U32519 (N_32519,N_25328,N_26726);
nand U32520 (N_32520,N_26777,N_26936);
nand U32521 (N_32521,N_28428,N_25547);
or U32522 (N_32522,N_29485,N_28222);
nor U32523 (N_32523,N_25992,N_29415);
and U32524 (N_32524,N_27995,N_28194);
and U32525 (N_32525,N_29803,N_27676);
xor U32526 (N_32526,N_29742,N_27108);
nand U32527 (N_32527,N_29731,N_28146);
nor U32528 (N_32528,N_25453,N_28021);
and U32529 (N_32529,N_28272,N_28716);
or U32530 (N_32530,N_28819,N_25414);
nand U32531 (N_32531,N_28169,N_29738);
nor U32532 (N_32532,N_26897,N_25436);
nand U32533 (N_32533,N_26516,N_27100);
or U32534 (N_32534,N_29262,N_28093);
xor U32535 (N_32535,N_25678,N_28705);
nor U32536 (N_32536,N_27873,N_29493);
nor U32537 (N_32537,N_27485,N_29235);
nor U32538 (N_32538,N_28514,N_27449);
nor U32539 (N_32539,N_29140,N_25544);
and U32540 (N_32540,N_29219,N_28053);
nand U32541 (N_32541,N_27716,N_25864);
xor U32542 (N_32542,N_29441,N_25444);
nor U32543 (N_32543,N_28228,N_25982);
and U32544 (N_32544,N_29155,N_26176);
or U32545 (N_32545,N_29056,N_25709);
or U32546 (N_32546,N_27064,N_25336);
nand U32547 (N_32547,N_26245,N_28808);
and U32548 (N_32548,N_28031,N_27718);
nor U32549 (N_32549,N_27912,N_29981);
and U32550 (N_32550,N_25876,N_25239);
xor U32551 (N_32551,N_27443,N_26814);
nor U32552 (N_32552,N_28574,N_25653);
nand U32553 (N_32553,N_27350,N_29088);
or U32554 (N_32554,N_27472,N_29631);
nand U32555 (N_32555,N_29676,N_27121);
nor U32556 (N_32556,N_29092,N_27407);
or U32557 (N_32557,N_25432,N_27737);
nor U32558 (N_32558,N_29412,N_25227);
nor U32559 (N_32559,N_28357,N_28427);
nand U32560 (N_32560,N_25070,N_25056);
nand U32561 (N_32561,N_29526,N_26149);
and U32562 (N_32562,N_28003,N_27285);
xnor U32563 (N_32563,N_28474,N_26987);
and U32564 (N_32564,N_26842,N_26166);
nand U32565 (N_32565,N_29167,N_27968);
and U32566 (N_32566,N_25005,N_26953);
nand U32567 (N_32567,N_28565,N_28991);
or U32568 (N_32568,N_28737,N_25959);
or U32569 (N_32569,N_29925,N_27378);
nand U32570 (N_32570,N_26094,N_25766);
or U32571 (N_32571,N_25736,N_27995);
nand U32572 (N_32572,N_27804,N_29749);
nor U32573 (N_32573,N_29386,N_27301);
and U32574 (N_32574,N_28561,N_28186);
xnor U32575 (N_32575,N_28460,N_27551);
or U32576 (N_32576,N_29633,N_29122);
nor U32577 (N_32577,N_25402,N_26118);
nor U32578 (N_32578,N_27814,N_26944);
nand U32579 (N_32579,N_28458,N_26938);
or U32580 (N_32580,N_27591,N_26034);
and U32581 (N_32581,N_28587,N_25338);
nor U32582 (N_32582,N_27603,N_28700);
and U32583 (N_32583,N_27877,N_26568);
nor U32584 (N_32584,N_26707,N_28221);
and U32585 (N_32585,N_26673,N_27121);
and U32586 (N_32586,N_27528,N_25922);
or U32587 (N_32587,N_25599,N_26985);
or U32588 (N_32588,N_28811,N_26758);
or U32589 (N_32589,N_26392,N_29727);
and U32590 (N_32590,N_29642,N_26008);
or U32591 (N_32591,N_29143,N_25151);
nand U32592 (N_32592,N_26393,N_25315);
nand U32593 (N_32593,N_25491,N_29621);
and U32594 (N_32594,N_28495,N_26857);
xor U32595 (N_32595,N_28854,N_27509);
xnor U32596 (N_32596,N_29525,N_27498);
and U32597 (N_32597,N_25023,N_28986);
nand U32598 (N_32598,N_27728,N_25870);
nor U32599 (N_32599,N_27925,N_26010);
nand U32600 (N_32600,N_27295,N_28725);
nor U32601 (N_32601,N_25051,N_26144);
nand U32602 (N_32602,N_25403,N_25384);
and U32603 (N_32603,N_25949,N_27727);
or U32604 (N_32604,N_25372,N_26767);
nand U32605 (N_32605,N_26876,N_28267);
nor U32606 (N_32606,N_28724,N_27781);
and U32607 (N_32607,N_26803,N_28002);
and U32608 (N_32608,N_29450,N_25000);
or U32609 (N_32609,N_29413,N_25632);
nor U32610 (N_32610,N_25927,N_27106);
nor U32611 (N_32611,N_27860,N_25998);
nand U32612 (N_32612,N_27156,N_25540);
nand U32613 (N_32613,N_29481,N_26150);
and U32614 (N_32614,N_27095,N_27914);
nor U32615 (N_32615,N_28247,N_28585);
and U32616 (N_32616,N_29725,N_29032);
nand U32617 (N_32617,N_26258,N_27318);
and U32618 (N_32618,N_27930,N_26819);
nand U32619 (N_32619,N_28005,N_26579);
nor U32620 (N_32620,N_26772,N_26841);
nand U32621 (N_32621,N_28174,N_28207);
or U32622 (N_32622,N_27695,N_28803);
nand U32623 (N_32623,N_28298,N_28522);
and U32624 (N_32624,N_27360,N_26912);
nor U32625 (N_32625,N_27892,N_29211);
nand U32626 (N_32626,N_29533,N_26077);
and U32627 (N_32627,N_27107,N_25085);
nor U32628 (N_32628,N_27215,N_29984);
nor U32629 (N_32629,N_27564,N_25557);
nor U32630 (N_32630,N_28900,N_26091);
or U32631 (N_32631,N_26132,N_28854);
nand U32632 (N_32632,N_25716,N_27538);
nand U32633 (N_32633,N_27350,N_25538);
nand U32634 (N_32634,N_25352,N_27066);
nand U32635 (N_32635,N_25887,N_25118);
or U32636 (N_32636,N_25326,N_28340);
and U32637 (N_32637,N_28729,N_25014);
xnor U32638 (N_32638,N_27743,N_25245);
xor U32639 (N_32639,N_29138,N_29387);
xnor U32640 (N_32640,N_26539,N_29211);
nand U32641 (N_32641,N_27671,N_28239);
nor U32642 (N_32642,N_28189,N_28363);
and U32643 (N_32643,N_25875,N_26422);
xnor U32644 (N_32644,N_28105,N_26853);
or U32645 (N_32645,N_26760,N_29198);
nand U32646 (N_32646,N_29506,N_25867);
or U32647 (N_32647,N_26964,N_28593);
nor U32648 (N_32648,N_28615,N_27471);
nor U32649 (N_32649,N_27035,N_27014);
or U32650 (N_32650,N_28359,N_25939);
or U32651 (N_32651,N_29379,N_29652);
nor U32652 (N_32652,N_29043,N_29728);
nor U32653 (N_32653,N_25699,N_27884);
nor U32654 (N_32654,N_29410,N_29393);
nand U32655 (N_32655,N_25956,N_27511);
and U32656 (N_32656,N_29641,N_28488);
or U32657 (N_32657,N_29673,N_29410);
or U32658 (N_32658,N_29092,N_26967);
nand U32659 (N_32659,N_28562,N_28867);
or U32660 (N_32660,N_28718,N_25391);
nand U32661 (N_32661,N_29838,N_27677);
nor U32662 (N_32662,N_28279,N_29621);
nor U32663 (N_32663,N_28574,N_28255);
and U32664 (N_32664,N_26664,N_27191);
nor U32665 (N_32665,N_27714,N_26424);
or U32666 (N_32666,N_28218,N_29320);
or U32667 (N_32667,N_25742,N_29626);
and U32668 (N_32668,N_27162,N_25298);
nand U32669 (N_32669,N_27259,N_29459);
nor U32670 (N_32670,N_25455,N_28176);
or U32671 (N_32671,N_27189,N_26159);
nor U32672 (N_32672,N_26023,N_28367);
nor U32673 (N_32673,N_28286,N_29804);
nor U32674 (N_32674,N_26733,N_28724);
nand U32675 (N_32675,N_29163,N_28939);
or U32676 (N_32676,N_27417,N_29866);
nor U32677 (N_32677,N_25302,N_28248);
nor U32678 (N_32678,N_26088,N_25238);
and U32679 (N_32679,N_25375,N_28777);
or U32680 (N_32680,N_27767,N_28452);
nor U32681 (N_32681,N_25918,N_28365);
nand U32682 (N_32682,N_26848,N_26436);
and U32683 (N_32683,N_28871,N_27132);
nand U32684 (N_32684,N_28695,N_26806);
nor U32685 (N_32685,N_28263,N_26131);
nor U32686 (N_32686,N_28923,N_27858);
and U32687 (N_32687,N_29300,N_26139);
nor U32688 (N_32688,N_25871,N_25885);
nand U32689 (N_32689,N_26372,N_29871);
nor U32690 (N_32690,N_26764,N_28968);
or U32691 (N_32691,N_25614,N_26077);
nand U32692 (N_32692,N_25300,N_29382);
or U32693 (N_32693,N_25910,N_25598);
nand U32694 (N_32694,N_28069,N_28558);
and U32695 (N_32695,N_27257,N_28779);
or U32696 (N_32696,N_26855,N_27479);
nor U32697 (N_32697,N_26312,N_29661);
nor U32698 (N_32698,N_29697,N_28076);
and U32699 (N_32699,N_27765,N_28807);
nor U32700 (N_32700,N_29818,N_28266);
or U32701 (N_32701,N_29810,N_26290);
or U32702 (N_32702,N_28738,N_27743);
nand U32703 (N_32703,N_26794,N_25210);
or U32704 (N_32704,N_28078,N_25920);
nand U32705 (N_32705,N_25009,N_25501);
and U32706 (N_32706,N_29276,N_29110);
xor U32707 (N_32707,N_27693,N_25961);
nand U32708 (N_32708,N_28175,N_29663);
nor U32709 (N_32709,N_26480,N_27212);
or U32710 (N_32710,N_28952,N_27847);
xnor U32711 (N_32711,N_26548,N_25749);
nor U32712 (N_32712,N_25338,N_25703);
xor U32713 (N_32713,N_29992,N_29666);
xnor U32714 (N_32714,N_28654,N_25149);
xnor U32715 (N_32715,N_29778,N_26573);
nor U32716 (N_32716,N_27318,N_26034);
or U32717 (N_32717,N_25319,N_25221);
xor U32718 (N_32718,N_25108,N_26280);
nor U32719 (N_32719,N_29339,N_29658);
nand U32720 (N_32720,N_25453,N_28497);
or U32721 (N_32721,N_25659,N_28221);
nor U32722 (N_32722,N_26992,N_28073);
xor U32723 (N_32723,N_28097,N_26527);
and U32724 (N_32724,N_29460,N_27615);
xnor U32725 (N_32725,N_27786,N_28025);
nand U32726 (N_32726,N_27602,N_25241);
and U32727 (N_32727,N_25433,N_25079);
or U32728 (N_32728,N_25127,N_29275);
or U32729 (N_32729,N_27312,N_25648);
xnor U32730 (N_32730,N_28611,N_25488);
or U32731 (N_32731,N_29795,N_29024);
or U32732 (N_32732,N_29660,N_25611);
and U32733 (N_32733,N_27070,N_25191);
and U32734 (N_32734,N_27332,N_27808);
or U32735 (N_32735,N_25108,N_28155);
nand U32736 (N_32736,N_29209,N_25298);
and U32737 (N_32737,N_29446,N_26438);
and U32738 (N_32738,N_25234,N_29005);
and U32739 (N_32739,N_27244,N_29783);
nand U32740 (N_32740,N_25960,N_29239);
xnor U32741 (N_32741,N_26096,N_28181);
nand U32742 (N_32742,N_26997,N_29131);
nand U32743 (N_32743,N_26137,N_26984);
xnor U32744 (N_32744,N_28981,N_25956);
nor U32745 (N_32745,N_29197,N_25610);
and U32746 (N_32746,N_26660,N_25404);
or U32747 (N_32747,N_29749,N_29056);
or U32748 (N_32748,N_26082,N_28065);
nand U32749 (N_32749,N_29174,N_25972);
nand U32750 (N_32750,N_27465,N_29961);
nand U32751 (N_32751,N_28379,N_26939);
nor U32752 (N_32752,N_26955,N_25877);
nand U32753 (N_32753,N_25195,N_27896);
xnor U32754 (N_32754,N_28276,N_29549);
nand U32755 (N_32755,N_25427,N_29783);
and U32756 (N_32756,N_29233,N_26647);
xnor U32757 (N_32757,N_28770,N_29512);
nor U32758 (N_32758,N_25826,N_25063);
nand U32759 (N_32759,N_28337,N_26509);
and U32760 (N_32760,N_27430,N_25587);
or U32761 (N_32761,N_27795,N_27641);
nor U32762 (N_32762,N_29477,N_27791);
nand U32763 (N_32763,N_29001,N_29762);
nor U32764 (N_32764,N_26140,N_26852);
nor U32765 (N_32765,N_29652,N_25588);
nor U32766 (N_32766,N_29012,N_29051);
or U32767 (N_32767,N_26949,N_28462);
and U32768 (N_32768,N_26193,N_27616);
nor U32769 (N_32769,N_27167,N_29994);
or U32770 (N_32770,N_28607,N_25154);
nand U32771 (N_32771,N_27886,N_29239);
nand U32772 (N_32772,N_29425,N_27544);
and U32773 (N_32773,N_27965,N_25065);
nor U32774 (N_32774,N_26007,N_26578);
or U32775 (N_32775,N_25873,N_25013);
or U32776 (N_32776,N_28941,N_28594);
nand U32777 (N_32777,N_28543,N_28891);
and U32778 (N_32778,N_25418,N_25672);
and U32779 (N_32779,N_26440,N_26950);
and U32780 (N_32780,N_28588,N_25511);
nand U32781 (N_32781,N_28606,N_27274);
nand U32782 (N_32782,N_26308,N_29410);
and U32783 (N_32783,N_27975,N_29457);
nand U32784 (N_32784,N_28333,N_26693);
and U32785 (N_32785,N_28424,N_25472);
and U32786 (N_32786,N_29744,N_27467);
and U32787 (N_32787,N_26151,N_28081);
and U32788 (N_32788,N_25410,N_26314);
nand U32789 (N_32789,N_27715,N_27089);
or U32790 (N_32790,N_27826,N_28695);
nand U32791 (N_32791,N_29127,N_25142);
and U32792 (N_32792,N_26759,N_26827);
xnor U32793 (N_32793,N_27178,N_25693);
and U32794 (N_32794,N_29448,N_27009);
nand U32795 (N_32795,N_26167,N_27047);
xnor U32796 (N_32796,N_25015,N_25998);
and U32797 (N_32797,N_27984,N_29830);
or U32798 (N_32798,N_26944,N_26291);
and U32799 (N_32799,N_28268,N_29875);
xor U32800 (N_32800,N_25526,N_26565);
or U32801 (N_32801,N_25815,N_27599);
nand U32802 (N_32802,N_26672,N_27321);
nor U32803 (N_32803,N_25412,N_26224);
nand U32804 (N_32804,N_29984,N_29313);
and U32805 (N_32805,N_27642,N_25405);
nand U32806 (N_32806,N_28460,N_25152);
xor U32807 (N_32807,N_29594,N_28613);
or U32808 (N_32808,N_27470,N_29025);
and U32809 (N_32809,N_26847,N_26080);
nand U32810 (N_32810,N_29926,N_25406);
nor U32811 (N_32811,N_26503,N_25964);
xnor U32812 (N_32812,N_29786,N_26767);
or U32813 (N_32813,N_26877,N_28191);
and U32814 (N_32814,N_26092,N_29696);
or U32815 (N_32815,N_27423,N_29393);
nor U32816 (N_32816,N_29477,N_29011);
and U32817 (N_32817,N_25244,N_27385);
xor U32818 (N_32818,N_29491,N_29988);
nand U32819 (N_32819,N_27238,N_25907);
and U32820 (N_32820,N_26312,N_29477);
and U32821 (N_32821,N_25082,N_27943);
nand U32822 (N_32822,N_28881,N_28393);
nand U32823 (N_32823,N_29979,N_26666);
nor U32824 (N_32824,N_29658,N_26514);
nand U32825 (N_32825,N_29507,N_26657);
nand U32826 (N_32826,N_27320,N_29803);
xor U32827 (N_32827,N_28449,N_29504);
and U32828 (N_32828,N_29064,N_28891);
nand U32829 (N_32829,N_25701,N_28253);
and U32830 (N_32830,N_25775,N_29496);
nand U32831 (N_32831,N_27668,N_25999);
nand U32832 (N_32832,N_26709,N_27827);
nor U32833 (N_32833,N_29540,N_28035);
nor U32834 (N_32834,N_26786,N_26755);
nand U32835 (N_32835,N_27236,N_25045);
nor U32836 (N_32836,N_26960,N_28817);
and U32837 (N_32837,N_25629,N_27435);
nor U32838 (N_32838,N_28028,N_26970);
nor U32839 (N_32839,N_28457,N_28573);
nand U32840 (N_32840,N_29620,N_29022);
and U32841 (N_32841,N_26347,N_29178);
or U32842 (N_32842,N_26797,N_27956);
nand U32843 (N_32843,N_28405,N_26117);
xnor U32844 (N_32844,N_26184,N_26237);
and U32845 (N_32845,N_27078,N_25572);
or U32846 (N_32846,N_25749,N_25807);
nand U32847 (N_32847,N_29708,N_28811);
xor U32848 (N_32848,N_25134,N_26868);
nor U32849 (N_32849,N_26551,N_27361);
nor U32850 (N_32850,N_27916,N_27010);
nor U32851 (N_32851,N_25016,N_29826);
or U32852 (N_32852,N_27862,N_29725);
xnor U32853 (N_32853,N_29883,N_27385);
nor U32854 (N_32854,N_25319,N_27146);
nor U32855 (N_32855,N_25970,N_25220);
nand U32856 (N_32856,N_25909,N_26059);
and U32857 (N_32857,N_27317,N_29285);
nor U32858 (N_32858,N_26208,N_29051);
nor U32859 (N_32859,N_25934,N_25187);
and U32860 (N_32860,N_29194,N_28907);
nand U32861 (N_32861,N_26336,N_25276);
nor U32862 (N_32862,N_25890,N_29364);
nor U32863 (N_32863,N_25931,N_26164);
nor U32864 (N_32864,N_25851,N_27145);
xor U32865 (N_32865,N_26488,N_25933);
nor U32866 (N_32866,N_27341,N_26819);
xor U32867 (N_32867,N_29771,N_25256);
xnor U32868 (N_32868,N_28595,N_27527);
and U32869 (N_32869,N_29700,N_25095);
nor U32870 (N_32870,N_28978,N_29405);
and U32871 (N_32871,N_25220,N_29452);
or U32872 (N_32872,N_27013,N_26671);
and U32873 (N_32873,N_25793,N_25588);
and U32874 (N_32874,N_25491,N_25780);
nor U32875 (N_32875,N_28374,N_26416);
and U32876 (N_32876,N_28167,N_27702);
nand U32877 (N_32877,N_25601,N_25581);
nand U32878 (N_32878,N_29433,N_29488);
and U32879 (N_32879,N_27196,N_27882);
nand U32880 (N_32880,N_25804,N_25039);
or U32881 (N_32881,N_25818,N_29341);
or U32882 (N_32882,N_27927,N_26477);
xor U32883 (N_32883,N_25575,N_25435);
nand U32884 (N_32884,N_25429,N_26735);
and U32885 (N_32885,N_25640,N_26229);
nand U32886 (N_32886,N_28909,N_29862);
xnor U32887 (N_32887,N_29093,N_25466);
xnor U32888 (N_32888,N_25648,N_28021);
and U32889 (N_32889,N_28048,N_27513);
or U32890 (N_32890,N_29206,N_27388);
or U32891 (N_32891,N_29980,N_29628);
or U32892 (N_32892,N_25975,N_26622);
nand U32893 (N_32893,N_27019,N_28525);
nor U32894 (N_32894,N_28261,N_27385);
or U32895 (N_32895,N_25789,N_28352);
nand U32896 (N_32896,N_26506,N_26171);
nand U32897 (N_32897,N_29375,N_26521);
or U32898 (N_32898,N_27187,N_28983);
nand U32899 (N_32899,N_28944,N_29215);
nor U32900 (N_32900,N_27600,N_26193);
nand U32901 (N_32901,N_28786,N_26780);
xor U32902 (N_32902,N_26390,N_29716);
nand U32903 (N_32903,N_28949,N_25285);
or U32904 (N_32904,N_28823,N_26945);
nor U32905 (N_32905,N_28107,N_27793);
or U32906 (N_32906,N_26895,N_25731);
or U32907 (N_32907,N_28586,N_27389);
and U32908 (N_32908,N_27523,N_28759);
nand U32909 (N_32909,N_25700,N_28085);
nand U32910 (N_32910,N_25978,N_27583);
nor U32911 (N_32911,N_29896,N_27503);
or U32912 (N_32912,N_28513,N_27961);
and U32913 (N_32913,N_25400,N_28302);
nand U32914 (N_32914,N_25509,N_26878);
nor U32915 (N_32915,N_29186,N_25164);
or U32916 (N_32916,N_26683,N_28401);
nor U32917 (N_32917,N_25409,N_25264);
nor U32918 (N_32918,N_25008,N_29247);
nand U32919 (N_32919,N_25752,N_28262);
nand U32920 (N_32920,N_27190,N_28256);
nand U32921 (N_32921,N_25003,N_28842);
nand U32922 (N_32922,N_27793,N_28899);
and U32923 (N_32923,N_27317,N_27599);
and U32924 (N_32924,N_25712,N_26883);
and U32925 (N_32925,N_27587,N_26984);
or U32926 (N_32926,N_28197,N_28178);
nor U32927 (N_32927,N_28522,N_26163);
or U32928 (N_32928,N_26083,N_29839);
xnor U32929 (N_32929,N_28240,N_27882);
nor U32930 (N_32930,N_25149,N_28568);
and U32931 (N_32931,N_25882,N_25532);
or U32932 (N_32932,N_28560,N_29165);
nand U32933 (N_32933,N_29895,N_26009);
and U32934 (N_32934,N_27719,N_26447);
or U32935 (N_32935,N_25459,N_25196);
xor U32936 (N_32936,N_27759,N_25273);
nor U32937 (N_32937,N_29699,N_28404);
xnor U32938 (N_32938,N_26498,N_28861);
or U32939 (N_32939,N_25718,N_25147);
nand U32940 (N_32940,N_27636,N_29845);
or U32941 (N_32941,N_27305,N_26578);
nor U32942 (N_32942,N_27681,N_27606);
nor U32943 (N_32943,N_28930,N_28945);
nor U32944 (N_32944,N_25770,N_29069);
nand U32945 (N_32945,N_27800,N_25524);
nand U32946 (N_32946,N_27185,N_29477);
nand U32947 (N_32947,N_28007,N_29837);
nor U32948 (N_32948,N_26761,N_27242);
or U32949 (N_32949,N_28659,N_27431);
and U32950 (N_32950,N_27085,N_27747);
or U32951 (N_32951,N_26346,N_25276);
xnor U32952 (N_32952,N_25732,N_27147);
xnor U32953 (N_32953,N_26920,N_29455);
nor U32954 (N_32954,N_25211,N_25125);
nand U32955 (N_32955,N_25475,N_29726);
and U32956 (N_32956,N_29248,N_27443);
and U32957 (N_32957,N_28215,N_27714);
or U32958 (N_32958,N_27693,N_29845);
and U32959 (N_32959,N_29055,N_27326);
and U32960 (N_32960,N_25874,N_27701);
or U32961 (N_32961,N_25833,N_28360);
xnor U32962 (N_32962,N_25943,N_29248);
nand U32963 (N_32963,N_29635,N_26922);
or U32964 (N_32964,N_25874,N_29185);
or U32965 (N_32965,N_28866,N_27473);
and U32966 (N_32966,N_29271,N_29072);
nor U32967 (N_32967,N_28052,N_28191);
or U32968 (N_32968,N_27635,N_29537);
nor U32969 (N_32969,N_29359,N_29875);
nor U32970 (N_32970,N_28536,N_28411);
or U32971 (N_32971,N_27742,N_28106);
nand U32972 (N_32972,N_27158,N_25476);
nand U32973 (N_32973,N_27735,N_28511);
nand U32974 (N_32974,N_25842,N_27619);
xnor U32975 (N_32975,N_25730,N_29867);
or U32976 (N_32976,N_27776,N_28481);
and U32977 (N_32977,N_28564,N_28896);
and U32978 (N_32978,N_26434,N_27778);
nand U32979 (N_32979,N_28908,N_28292);
nor U32980 (N_32980,N_29767,N_27189);
nor U32981 (N_32981,N_29430,N_28894);
nand U32982 (N_32982,N_28294,N_29169);
or U32983 (N_32983,N_25943,N_26298);
and U32984 (N_32984,N_27612,N_26318);
or U32985 (N_32985,N_25069,N_29803);
nor U32986 (N_32986,N_29967,N_28031);
nand U32987 (N_32987,N_29261,N_27743);
or U32988 (N_32988,N_26303,N_25268);
xnor U32989 (N_32989,N_29148,N_29411);
nand U32990 (N_32990,N_26598,N_29582);
or U32991 (N_32991,N_28718,N_25681);
and U32992 (N_32992,N_26645,N_28816);
and U32993 (N_32993,N_25486,N_29857);
nand U32994 (N_32994,N_25403,N_26558);
nand U32995 (N_32995,N_26047,N_26458);
and U32996 (N_32996,N_27951,N_29386);
nor U32997 (N_32997,N_25252,N_26583);
nand U32998 (N_32998,N_26358,N_28516);
xnor U32999 (N_32999,N_28185,N_29946);
nor U33000 (N_33000,N_27342,N_27468);
xnor U33001 (N_33001,N_28461,N_29444);
and U33002 (N_33002,N_28271,N_26914);
xnor U33003 (N_33003,N_29979,N_29357);
nand U33004 (N_33004,N_28027,N_27544);
and U33005 (N_33005,N_27137,N_25095);
or U33006 (N_33006,N_25519,N_27935);
xnor U33007 (N_33007,N_25749,N_28706);
or U33008 (N_33008,N_26437,N_26688);
and U33009 (N_33009,N_26707,N_29821);
nor U33010 (N_33010,N_27248,N_26222);
nor U33011 (N_33011,N_27880,N_25240);
or U33012 (N_33012,N_29840,N_26548);
or U33013 (N_33013,N_26959,N_28785);
nand U33014 (N_33014,N_26110,N_29051);
nor U33015 (N_33015,N_26879,N_26157);
nor U33016 (N_33016,N_26621,N_27804);
nor U33017 (N_33017,N_28056,N_27785);
nor U33018 (N_33018,N_29715,N_27826);
and U33019 (N_33019,N_27167,N_27764);
and U33020 (N_33020,N_26306,N_28712);
nand U33021 (N_33021,N_29004,N_28785);
or U33022 (N_33022,N_28575,N_29535);
and U33023 (N_33023,N_29108,N_28266);
nand U33024 (N_33024,N_25479,N_27161);
and U33025 (N_33025,N_29049,N_27968);
nor U33026 (N_33026,N_29304,N_27830);
or U33027 (N_33027,N_28104,N_26940);
nand U33028 (N_33028,N_29908,N_25983);
and U33029 (N_33029,N_25731,N_28720);
and U33030 (N_33030,N_26123,N_26678);
or U33031 (N_33031,N_29397,N_29989);
or U33032 (N_33032,N_27905,N_29528);
nor U33033 (N_33033,N_26400,N_29316);
or U33034 (N_33034,N_29527,N_26652);
xnor U33035 (N_33035,N_28110,N_26716);
and U33036 (N_33036,N_25381,N_29372);
nand U33037 (N_33037,N_28103,N_26300);
or U33038 (N_33038,N_29830,N_25213);
nand U33039 (N_33039,N_28965,N_29413);
nor U33040 (N_33040,N_27544,N_27694);
and U33041 (N_33041,N_26989,N_25777);
nand U33042 (N_33042,N_29087,N_27468);
and U33043 (N_33043,N_25775,N_25528);
nand U33044 (N_33044,N_29718,N_25782);
and U33045 (N_33045,N_25384,N_28433);
and U33046 (N_33046,N_25506,N_26097);
xnor U33047 (N_33047,N_26570,N_28939);
nor U33048 (N_33048,N_27407,N_27991);
nor U33049 (N_33049,N_27704,N_27454);
nor U33050 (N_33050,N_25357,N_27307);
and U33051 (N_33051,N_28308,N_26718);
nor U33052 (N_33052,N_28517,N_29234);
or U33053 (N_33053,N_28354,N_29768);
and U33054 (N_33054,N_27982,N_27996);
nor U33055 (N_33055,N_27580,N_29672);
or U33056 (N_33056,N_28460,N_29827);
and U33057 (N_33057,N_29749,N_27001);
nand U33058 (N_33058,N_27616,N_29384);
nand U33059 (N_33059,N_26095,N_26696);
nor U33060 (N_33060,N_29021,N_26817);
nand U33061 (N_33061,N_27344,N_25916);
and U33062 (N_33062,N_25029,N_28013);
xnor U33063 (N_33063,N_27695,N_26806);
xnor U33064 (N_33064,N_26273,N_27358);
nand U33065 (N_33065,N_25184,N_28010);
and U33066 (N_33066,N_25463,N_27677);
and U33067 (N_33067,N_28563,N_26059);
nor U33068 (N_33068,N_28824,N_25514);
xnor U33069 (N_33069,N_26806,N_28469);
nor U33070 (N_33070,N_26045,N_26821);
nand U33071 (N_33071,N_25662,N_27050);
nand U33072 (N_33072,N_26267,N_25973);
nor U33073 (N_33073,N_29794,N_26958);
nor U33074 (N_33074,N_29205,N_28197);
and U33075 (N_33075,N_26404,N_28896);
nor U33076 (N_33076,N_29883,N_25755);
and U33077 (N_33077,N_29315,N_26634);
nor U33078 (N_33078,N_29121,N_29114);
nor U33079 (N_33079,N_29192,N_27805);
nor U33080 (N_33080,N_26064,N_27746);
nand U33081 (N_33081,N_27534,N_29140);
nor U33082 (N_33082,N_28767,N_26410);
nand U33083 (N_33083,N_29016,N_25051);
or U33084 (N_33084,N_25057,N_27021);
or U33085 (N_33085,N_28891,N_26704);
xor U33086 (N_33086,N_29363,N_29447);
nand U33087 (N_33087,N_25152,N_26199);
or U33088 (N_33088,N_25194,N_27066);
and U33089 (N_33089,N_29884,N_26521);
nand U33090 (N_33090,N_27563,N_27584);
nor U33091 (N_33091,N_26236,N_29408);
nand U33092 (N_33092,N_26278,N_28753);
xnor U33093 (N_33093,N_25496,N_26426);
nor U33094 (N_33094,N_25762,N_25889);
nand U33095 (N_33095,N_26192,N_27635);
nor U33096 (N_33096,N_29268,N_27450);
nand U33097 (N_33097,N_25858,N_29135);
and U33098 (N_33098,N_29825,N_28856);
nor U33099 (N_33099,N_29683,N_29909);
nor U33100 (N_33100,N_29063,N_26496);
nand U33101 (N_33101,N_29715,N_26968);
xnor U33102 (N_33102,N_27303,N_28555);
or U33103 (N_33103,N_28248,N_25621);
nor U33104 (N_33104,N_29637,N_27871);
xor U33105 (N_33105,N_28600,N_27233);
and U33106 (N_33106,N_26290,N_26544);
nand U33107 (N_33107,N_28832,N_28398);
and U33108 (N_33108,N_28050,N_27563);
nand U33109 (N_33109,N_27358,N_28068);
and U33110 (N_33110,N_26298,N_25619);
and U33111 (N_33111,N_29303,N_29980);
xor U33112 (N_33112,N_25797,N_26538);
and U33113 (N_33113,N_26087,N_25769);
and U33114 (N_33114,N_28685,N_28190);
xor U33115 (N_33115,N_28936,N_27936);
xnor U33116 (N_33116,N_28389,N_28150);
nand U33117 (N_33117,N_29305,N_25731);
nand U33118 (N_33118,N_29316,N_26359);
and U33119 (N_33119,N_25087,N_27673);
and U33120 (N_33120,N_25788,N_25072);
nor U33121 (N_33121,N_25118,N_27909);
and U33122 (N_33122,N_27196,N_26984);
or U33123 (N_33123,N_29054,N_28635);
and U33124 (N_33124,N_28090,N_25548);
and U33125 (N_33125,N_25459,N_28676);
or U33126 (N_33126,N_29642,N_25934);
nand U33127 (N_33127,N_28528,N_28493);
or U33128 (N_33128,N_28986,N_26450);
and U33129 (N_33129,N_26495,N_25532);
or U33130 (N_33130,N_28740,N_25921);
nor U33131 (N_33131,N_25680,N_29612);
xor U33132 (N_33132,N_29601,N_25381);
nand U33133 (N_33133,N_26154,N_29780);
xor U33134 (N_33134,N_25136,N_27790);
or U33135 (N_33135,N_26662,N_25482);
nand U33136 (N_33136,N_28789,N_26274);
nor U33137 (N_33137,N_29036,N_28230);
xnor U33138 (N_33138,N_26692,N_25158);
and U33139 (N_33139,N_28912,N_26713);
xnor U33140 (N_33140,N_28784,N_25915);
nor U33141 (N_33141,N_27709,N_29005);
nand U33142 (N_33142,N_26378,N_25952);
nor U33143 (N_33143,N_28880,N_28561);
or U33144 (N_33144,N_29851,N_25388);
and U33145 (N_33145,N_29515,N_25675);
or U33146 (N_33146,N_26819,N_28005);
nor U33147 (N_33147,N_26083,N_25700);
and U33148 (N_33148,N_26781,N_29989);
nor U33149 (N_33149,N_26664,N_25689);
xnor U33150 (N_33150,N_27894,N_26697);
or U33151 (N_33151,N_28450,N_27569);
nand U33152 (N_33152,N_25402,N_29029);
and U33153 (N_33153,N_28948,N_26738);
and U33154 (N_33154,N_28634,N_26887);
nand U33155 (N_33155,N_29188,N_25782);
nor U33156 (N_33156,N_28127,N_29715);
nand U33157 (N_33157,N_25715,N_29025);
nor U33158 (N_33158,N_27814,N_26480);
or U33159 (N_33159,N_28288,N_27348);
xor U33160 (N_33160,N_29074,N_28872);
or U33161 (N_33161,N_29750,N_26055);
nand U33162 (N_33162,N_28373,N_28622);
and U33163 (N_33163,N_26645,N_25093);
nand U33164 (N_33164,N_27371,N_25056);
or U33165 (N_33165,N_28245,N_25699);
nand U33166 (N_33166,N_25802,N_28873);
nand U33167 (N_33167,N_26551,N_27981);
nor U33168 (N_33168,N_28981,N_26421);
nor U33169 (N_33169,N_28536,N_27722);
and U33170 (N_33170,N_27930,N_28707);
xnor U33171 (N_33171,N_26507,N_25360);
nor U33172 (N_33172,N_28261,N_29505);
or U33173 (N_33173,N_26752,N_29416);
and U33174 (N_33174,N_29898,N_29822);
and U33175 (N_33175,N_25177,N_29144);
nand U33176 (N_33176,N_25977,N_26479);
and U33177 (N_33177,N_29638,N_27055);
nand U33178 (N_33178,N_26176,N_29325);
xor U33179 (N_33179,N_26295,N_28250);
or U33180 (N_33180,N_26449,N_29100);
or U33181 (N_33181,N_28726,N_25976);
nor U33182 (N_33182,N_29868,N_25890);
or U33183 (N_33183,N_27946,N_25792);
xnor U33184 (N_33184,N_29582,N_29261);
or U33185 (N_33185,N_25432,N_25563);
nor U33186 (N_33186,N_28322,N_29276);
xor U33187 (N_33187,N_26432,N_27936);
nand U33188 (N_33188,N_25663,N_28862);
xor U33189 (N_33189,N_29958,N_26205);
nand U33190 (N_33190,N_29642,N_29942);
or U33191 (N_33191,N_28311,N_25441);
nor U33192 (N_33192,N_27736,N_26884);
and U33193 (N_33193,N_28084,N_25895);
nand U33194 (N_33194,N_25459,N_27046);
or U33195 (N_33195,N_27370,N_25098);
nand U33196 (N_33196,N_25915,N_29851);
nor U33197 (N_33197,N_27092,N_29178);
and U33198 (N_33198,N_27845,N_26835);
nand U33199 (N_33199,N_26894,N_27147);
or U33200 (N_33200,N_25138,N_27200);
xnor U33201 (N_33201,N_28480,N_27234);
nor U33202 (N_33202,N_29182,N_29721);
or U33203 (N_33203,N_26589,N_29756);
and U33204 (N_33204,N_27701,N_25016);
and U33205 (N_33205,N_28776,N_25774);
and U33206 (N_33206,N_28470,N_26234);
and U33207 (N_33207,N_27175,N_28454);
and U33208 (N_33208,N_28639,N_26749);
nor U33209 (N_33209,N_29191,N_27105);
or U33210 (N_33210,N_25782,N_25570);
or U33211 (N_33211,N_26443,N_27681);
and U33212 (N_33212,N_27822,N_26123);
nand U33213 (N_33213,N_27617,N_27756);
or U33214 (N_33214,N_27421,N_29983);
or U33215 (N_33215,N_25467,N_28432);
nand U33216 (N_33216,N_25277,N_29116);
and U33217 (N_33217,N_27688,N_25207);
nor U33218 (N_33218,N_28074,N_29654);
nor U33219 (N_33219,N_27817,N_28108);
xor U33220 (N_33220,N_25811,N_28700);
and U33221 (N_33221,N_28420,N_29489);
nor U33222 (N_33222,N_28338,N_25675);
xnor U33223 (N_33223,N_27496,N_29172);
or U33224 (N_33224,N_25624,N_29862);
and U33225 (N_33225,N_26737,N_26539);
and U33226 (N_33226,N_27577,N_29592);
nand U33227 (N_33227,N_29218,N_29019);
or U33228 (N_33228,N_26092,N_27822);
or U33229 (N_33229,N_28769,N_29727);
nand U33230 (N_33230,N_26888,N_26600);
or U33231 (N_33231,N_25809,N_25467);
and U33232 (N_33232,N_29649,N_27934);
nand U33233 (N_33233,N_26945,N_29195);
nor U33234 (N_33234,N_29309,N_26044);
xnor U33235 (N_33235,N_27614,N_28491);
nand U33236 (N_33236,N_29462,N_28799);
nor U33237 (N_33237,N_29768,N_25738);
nor U33238 (N_33238,N_27095,N_26013);
xor U33239 (N_33239,N_25463,N_26545);
and U33240 (N_33240,N_27929,N_26978);
and U33241 (N_33241,N_26668,N_29618);
or U33242 (N_33242,N_27288,N_27148);
or U33243 (N_33243,N_26508,N_25132);
and U33244 (N_33244,N_26866,N_29809);
nand U33245 (N_33245,N_26958,N_27790);
nor U33246 (N_33246,N_25022,N_26063);
nand U33247 (N_33247,N_27137,N_26673);
or U33248 (N_33248,N_25809,N_28915);
nor U33249 (N_33249,N_29835,N_27377);
and U33250 (N_33250,N_26656,N_25897);
and U33251 (N_33251,N_29913,N_27293);
or U33252 (N_33252,N_25478,N_28967);
and U33253 (N_33253,N_28044,N_28663);
nand U33254 (N_33254,N_28597,N_26234);
or U33255 (N_33255,N_25191,N_29898);
or U33256 (N_33256,N_28866,N_26489);
nand U33257 (N_33257,N_28677,N_29952);
nand U33258 (N_33258,N_27522,N_28548);
and U33259 (N_33259,N_26712,N_29120);
and U33260 (N_33260,N_29150,N_27617);
nand U33261 (N_33261,N_29653,N_26251);
nand U33262 (N_33262,N_26524,N_27346);
and U33263 (N_33263,N_29963,N_26095);
and U33264 (N_33264,N_29282,N_25214);
nor U33265 (N_33265,N_29978,N_28158);
nand U33266 (N_33266,N_28011,N_27993);
or U33267 (N_33267,N_27938,N_26184);
nand U33268 (N_33268,N_27369,N_28968);
and U33269 (N_33269,N_26052,N_25875);
nor U33270 (N_33270,N_28383,N_27599);
nor U33271 (N_33271,N_25090,N_27508);
nand U33272 (N_33272,N_29576,N_26038);
or U33273 (N_33273,N_28428,N_29207);
nor U33274 (N_33274,N_29104,N_29623);
nor U33275 (N_33275,N_26625,N_25981);
nor U33276 (N_33276,N_27817,N_27623);
nor U33277 (N_33277,N_29411,N_25303);
and U33278 (N_33278,N_25248,N_28457);
nor U33279 (N_33279,N_29494,N_29175);
nor U33280 (N_33280,N_28070,N_25125);
and U33281 (N_33281,N_27847,N_28665);
and U33282 (N_33282,N_29589,N_29588);
or U33283 (N_33283,N_29324,N_28488);
xor U33284 (N_33284,N_27486,N_29558);
or U33285 (N_33285,N_29770,N_26212);
and U33286 (N_33286,N_29921,N_25567);
nand U33287 (N_33287,N_26729,N_25421);
nor U33288 (N_33288,N_29058,N_27370);
or U33289 (N_33289,N_28921,N_25573);
and U33290 (N_33290,N_27621,N_25340);
or U33291 (N_33291,N_27787,N_29739);
and U33292 (N_33292,N_27226,N_28901);
or U33293 (N_33293,N_27913,N_29774);
and U33294 (N_33294,N_26812,N_25953);
or U33295 (N_33295,N_27601,N_25043);
nand U33296 (N_33296,N_28138,N_28161);
nor U33297 (N_33297,N_28266,N_28770);
xnor U33298 (N_33298,N_28151,N_29214);
nand U33299 (N_33299,N_27035,N_28056);
nand U33300 (N_33300,N_29963,N_28777);
and U33301 (N_33301,N_28826,N_29105);
or U33302 (N_33302,N_29447,N_29056);
xor U33303 (N_33303,N_27044,N_26578);
and U33304 (N_33304,N_26637,N_27447);
nor U33305 (N_33305,N_25054,N_28804);
and U33306 (N_33306,N_26526,N_26951);
nand U33307 (N_33307,N_29062,N_28176);
or U33308 (N_33308,N_27525,N_26374);
nand U33309 (N_33309,N_25146,N_25632);
and U33310 (N_33310,N_28736,N_28019);
or U33311 (N_33311,N_29211,N_27191);
nor U33312 (N_33312,N_28054,N_28748);
xnor U33313 (N_33313,N_28931,N_26844);
and U33314 (N_33314,N_26375,N_25070);
xor U33315 (N_33315,N_25535,N_27547);
xnor U33316 (N_33316,N_25634,N_26642);
or U33317 (N_33317,N_25846,N_28239);
nand U33318 (N_33318,N_27769,N_27449);
or U33319 (N_33319,N_28827,N_27763);
xnor U33320 (N_33320,N_29674,N_28245);
nand U33321 (N_33321,N_25135,N_29651);
nand U33322 (N_33322,N_27260,N_29914);
nor U33323 (N_33323,N_26375,N_28985);
and U33324 (N_33324,N_28567,N_25914);
and U33325 (N_33325,N_28154,N_26708);
xor U33326 (N_33326,N_29241,N_26792);
nor U33327 (N_33327,N_26772,N_28910);
or U33328 (N_33328,N_25094,N_29644);
or U33329 (N_33329,N_26286,N_26018);
nor U33330 (N_33330,N_26945,N_27448);
nand U33331 (N_33331,N_25937,N_27321);
or U33332 (N_33332,N_27663,N_29914);
xor U33333 (N_33333,N_29224,N_25259);
nand U33334 (N_33334,N_25303,N_27048);
nor U33335 (N_33335,N_26811,N_27042);
nand U33336 (N_33336,N_28629,N_29209);
nand U33337 (N_33337,N_26089,N_27494);
and U33338 (N_33338,N_26798,N_29712);
or U33339 (N_33339,N_28139,N_29340);
and U33340 (N_33340,N_27911,N_25037);
nand U33341 (N_33341,N_29154,N_29117);
nand U33342 (N_33342,N_25038,N_26445);
nor U33343 (N_33343,N_28732,N_29191);
and U33344 (N_33344,N_27910,N_27859);
nand U33345 (N_33345,N_28590,N_27619);
nor U33346 (N_33346,N_29617,N_27453);
or U33347 (N_33347,N_28634,N_26346);
nor U33348 (N_33348,N_27313,N_26988);
and U33349 (N_33349,N_28287,N_27197);
xnor U33350 (N_33350,N_29756,N_27842);
nand U33351 (N_33351,N_29795,N_25958);
nor U33352 (N_33352,N_29248,N_28310);
or U33353 (N_33353,N_25361,N_25421);
or U33354 (N_33354,N_28457,N_27424);
nand U33355 (N_33355,N_28440,N_27725);
nor U33356 (N_33356,N_28382,N_29110);
nand U33357 (N_33357,N_29378,N_28334);
nand U33358 (N_33358,N_26110,N_27167);
nand U33359 (N_33359,N_26378,N_26465);
nand U33360 (N_33360,N_29708,N_26890);
nand U33361 (N_33361,N_26629,N_29613);
xor U33362 (N_33362,N_27299,N_28400);
nand U33363 (N_33363,N_25189,N_26844);
nand U33364 (N_33364,N_28413,N_26099);
or U33365 (N_33365,N_25419,N_27136);
nand U33366 (N_33366,N_29432,N_25077);
and U33367 (N_33367,N_25796,N_25893);
or U33368 (N_33368,N_28264,N_27971);
nand U33369 (N_33369,N_27964,N_29726);
nor U33370 (N_33370,N_28396,N_28361);
and U33371 (N_33371,N_27326,N_26456);
or U33372 (N_33372,N_26130,N_25584);
and U33373 (N_33373,N_28641,N_25471);
xor U33374 (N_33374,N_25346,N_28812);
nor U33375 (N_33375,N_27402,N_29845);
and U33376 (N_33376,N_29170,N_25207);
nand U33377 (N_33377,N_26382,N_26113);
or U33378 (N_33378,N_27806,N_29647);
and U33379 (N_33379,N_29994,N_27488);
or U33380 (N_33380,N_28221,N_28202);
or U33381 (N_33381,N_25864,N_29173);
nor U33382 (N_33382,N_26360,N_26250);
nand U33383 (N_33383,N_27790,N_26382);
nor U33384 (N_33384,N_25130,N_27471);
nand U33385 (N_33385,N_27255,N_28569);
nand U33386 (N_33386,N_29262,N_27409);
nand U33387 (N_33387,N_27716,N_29823);
nand U33388 (N_33388,N_25087,N_25225);
nand U33389 (N_33389,N_27630,N_26717);
or U33390 (N_33390,N_25687,N_26906);
xnor U33391 (N_33391,N_27695,N_26844);
and U33392 (N_33392,N_26687,N_25642);
or U33393 (N_33393,N_29500,N_28057);
and U33394 (N_33394,N_25505,N_28026);
xor U33395 (N_33395,N_25471,N_27132);
nor U33396 (N_33396,N_26831,N_26696);
or U33397 (N_33397,N_26567,N_26299);
nand U33398 (N_33398,N_28734,N_26539);
nor U33399 (N_33399,N_25804,N_25565);
and U33400 (N_33400,N_25079,N_28782);
xnor U33401 (N_33401,N_25825,N_26863);
or U33402 (N_33402,N_28221,N_25250);
or U33403 (N_33403,N_28219,N_28025);
and U33404 (N_33404,N_29331,N_27857);
and U33405 (N_33405,N_28304,N_27588);
nor U33406 (N_33406,N_28048,N_26560);
or U33407 (N_33407,N_26276,N_25976);
and U33408 (N_33408,N_27156,N_28605);
nand U33409 (N_33409,N_26065,N_28924);
xor U33410 (N_33410,N_29435,N_25407);
nand U33411 (N_33411,N_25889,N_25677);
and U33412 (N_33412,N_28944,N_29961);
nor U33413 (N_33413,N_29041,N_29760);
and U33414 (N_33414,N_27080,N_29149);
and U33415 (N_33415,N_25274,N_28925);
xor U33416 (N_33416,N_25774,N_29441);
nor U33417 (N_33417,N_29342,N_28931);
nor U33418 (N_33418,N_25397,N_28005);
xnor U33419 (N_33419,N_26868,N_27208);
and U33420 (N_33420,N_29266,N_26056);
and U33421 (N_33421,N_25630,N_25103);
xor U33422 (N_33422,N_27318,N_28915);
or U33423 (N_33423,N_25140,N_29945);
or U33424 (N_33424,N_25528,N_29078);
nor U33425 (N_33425,N_28966,N_27489);
nand U33426 (N_33426,N_28407,N_28941);
nand U33427 (N_33427,N_27799,N_27497);
nor U33428 (N_33428,N_29120,N_29509);
nor U33429 (N_33429,N_26199,N_25121);
or U33430 (N_33430,N_29033,N_27212);
nor U33431 (N_33431,N_25886,N_29217);
xor U33432 (N_33432,N_29696,N_29282);
nor U33433 (N_33433,N_27697,N_26860);
or U33434 (N_33434,N_25114,N_29859);
nor U33435 (N_33435,N_27581,N_28684);
and U33436 (N_33436,N_25912,N_29574);
nand U33437 (N_33437,N_27639,N_29787);
nand U33438 (N_33438,N_29459,N_25238);
or U33439 (N_33439,N_28857,N_29124);
or U33440 (N_33440,N_25054,N_29924);
or U33441 (N_33441,N_27433,N_26331);
nor U33442 (N_33442,N_27388,N_25864);
nand U33443 (N_33443,N_29649,N_25671);
or U33444 (N_33444,N_25628,N_29836);
or U33445 (N_33445,N_25430,N_29008);
or U33446 (N_33446,N_29230,N_29534);
nand U33447 (N_33447,N_27081,N_26896);
nand U33448 (N_33448,N_25536,N_27751);
nand U33449 (N_33449,N_28020,N_25295);
nor U33450 (N_33450,N_29510,N_25110);
xnor U33451 (N_33451,N_25565,N_26154);
nand U33452 (N_33452,N_25642,N_27570);
nand U33453 (N_33453,N_27130,N_28273);
nor U33454 (N_33454,N_28126,N_26162);
and U33455 (N_33455,N_28962,N_25551);
nand U33456 (N_33456,N_28058,N_25693);
nor U33457 (N_33457,N_28581,N_25391);
or U33458 (N_33458,N_28437,N_29397);
and U33459 (N_33459,N_29405,N_28903);
and U33460 (N_33460,N_27397,N_25638);
nor U33461 (N_33461,N_26180,N_27036);
or U33462 (N_33462,N_26438,N_26718);
or U33463 (N_33463,N_27767,N_27057);
nor U33464 (N_33464,N_28784,N_25522);
nand U33465 (N_33465,N_25195,N_28445);
nand U33466 (N_33466,N_29356,N_26634);
xor U33467 (N_33467,N_28386,N_28115);
nor U33468 (N_33468,N_27043,N_28576);
or U33469 (N_33469,N_25540,N_25764);
nand U33470 (N_33470,N_29626,N_25885);
and U33471 (N_33471,N_28315,N_26632);
or U33472 (N_33472,N_28618,N_27865);
nand U33473 (N_33473,N_29809,N_27824);
nor U33474 (N_33474,N_29981,N_29067);
and U33475 (N_33475,N_26129,N_26430);
nor U33476 (N_33476,N_26567,N_27454);
or U33477 (N_33477,N_26888,N_28136);
or U33478 (N_33478,N_25321,N_28977);
nor U33479 (N_33479,N_25730,N_26696);
or U33480 (N_33480,N_25276,N_28818);
or U33481 (N_33481,N_25991,N_26180);
and U33482 (N_33482,N_27959,N_29406);
nand U33483 (N_33483,N_25973,N_26583);
nand U33484 (N_33484,N_25314,N_25868);
and U33485 (N_33485,N_28044,N_27594);
and U33486 (N_33486,N_25058,N_28277);
or U33487 (N_33487,N_26352,N_29474);
xor U33488 (N_33488,N_27536,N_26190);
xnor U33489 (N_33489,N_26745,N_25786);
and U33490 (N_33490,N_29199,N_27585);
or U33491 (N_33491,N_25851,N_25065);
nor U33492 (N_33492,N_27864,N_26184);
or U33493 (N_33493,N_28467,N_25902);
or U33494 (N_33494,N_28177,N_26901);
or U33495 (N_33495,N_27865,N_29351);
nand U33496 (N_33496,N_27377,N_28449);
nor U33497 (N_33497,N_26660,N_28603);
nor U33498 (N_33498,N_27092,N_26945);
xnor U33499 (N_33499,N_28937,N_28158);
and U33500 (N_33500,N_27796,N_26165);
nor U33501 (N_33501,N_25212,N_26759);
nand U33502 (N_33502,N_28725,N_28857);
or U33503 (N_33503,N_25081,N_28937);
or U33504 (N_33504,N_27381,N_25474);
and U33505 (N_33505,N_28678,N_27066);
or U33506 (N_33506,N_28827,N_25319);
and U33507 (N_33507,N_28109,N_27856);
nor U33508 (N_33508,N_26866,N_29407);
and U33509 (N_33509,N_28966,N_28281);
xnor U33510 (N_33510,N_28120,N_26423);
or U33511 (N_33511,N_29488,N_25938);
xnor U33512 (N_33512,N_26525,N_25616);
nand U33513 (N_33513,N_29341,N_29919);
nand U33514 (N_33514,N_28720,N_28211);
or U33515 (N_33515,N_27670,N_26999);
xnor U33516 (N_33516,N_26562,N_29169);
nor U33517 (N_33517,N_27733,N_25154);
nor U33518 (N_33518,N_27781,N_27294);
or U33519 (N_33519,N_29358,N_25885);
nor U33520 (N_33520,N_29969,N_26861);
xor U33521 (N_33521,N_29552,N_25712);
and U33522 (N_33522,N_26341,N_26763);
nor U33523 (N_33523,N_29246,N_25344);
nor U33524 (N_33524,N_28416,N_27039);
xnor U33525 (N_33525,N_29905,N_25542);
nor U33526 (N_33526,N_27513,N_27048);
nand U33527 (N_33527,N_28722,N_27731);
nor U33528 (N_33528,N_27488,N_26603);
and U33529 (N_33529,N_28947,N_25732);
xnor U33530 (N_33530,N_26760,N_29939);
xnor U33531 (N_33531,N_25067,N_25467);
nand U33532 (N_33532,N_28115,N_28717);
xor U33533 (N_33533,N_27822,N_27661);
and U33534 (N_33534,N_25931,N_27685);
nand U33535 (N_33535,N_27324,N_27492);
or U33536 (N_33536,N_26571,N_29880);
or U33537 (N_33537,N_29548,N_25953);
nor U33538 (N_33538,N_27182,N_27315);
or U33539 (N_33539,N_27285,N_26073);
nand U33540 (N_33540,N_27656,N_27804);
and U33541 (N_33541,N_25773,N_27983);
and U33542 (N_33542,N_28600,N_25510);
or U33543 (N_33543,N_28621,N_29416);
nor U33544 (N_33544,N_28173,N_28526);
and U33545 (N_33545,N_25900,N_27090);
xor U33546 (N_33546,N_27372,N_29603);
nor U33547 (N_33547,N_28548,N_29790);
and U33548 (N_33548,N_28263,N_25232);
or U33549 (N_33549,N_28203,N_26475);
xnor U33550 (N_33550,N_27369,N_27928);
or U33551 (N_33551,N_26173,N_25365);
xnor U33552 (N_33552,N_27634,N_28797);
nand U33553 (N_33553,N_25609,N_29647);
and U33554 (N_33554,N_25247,N_25383);
xor U33555 (N_33555,N_28075,N_28699);
nand U33556 (N_33556,N_28496,N_27227);
nor U33557 (N_33557,N_28990,N_27222);
nor U33558 (N_33558,N_29544,N_25159);
nor U33559 (N_33559,N_26884,N_26406);
xor U33560 (N_33560,N_29515,N_26507);
nor U33561 (N_33561,N_25349,N_28727);
or U33562 (N_33562,N_27981,N_25029);
nor U33563 (N_33563,N_26430,N_29601);
and U33564 (N_33564,N_28007,N_28748);
nand U33565 (N_33565,N_25547,N_29999);
nand U33566 (N_33566,N_27978,N_26967);
or U33567 (N_33567,N_27005,N_25700);
nor U33568 (N_33568,N_29556,N_27606);
and U33569 (N_33569,N_27511,N_26793);
nor U33570 (N_33570,N_26822,N_27123);
and U33571 (N_33571,N_26672,N_28686);
and U33572 (N_33572,N_27435,N_26202);
nand U33573 (N_33573,N_28903,N_29039);
xor U33574 (N_33574,N_25545,N_25643);
nor U33575 (N_33575,N_29419,N_26531);
or U33576 (N_33576,N_25296,N_25172);
or U33577 (N_33577,N_29743,N_28949);
and U33578 (N_33578,N_26358,N_28551);
and U33579 (N_33579,N_28081,N_28700);
nor U33580 (N_33580,N_28333,N_29365);
and U33581 (N_33581,N_29074,N_29187);
and U33582 (N_33582,N_27248,N_25103);
nor U33583 (N_33583,N_26843,N_25785);
and U33584 (N_33584,N_29801,N_26541);
or U33585 (N_33585,N_25506,N_27497);
nor U33586 (N_33586,N_26055,N_27302);
or U33587 (N_33587,N_25562,N_28864);
and U33588 (N_33588,N_25790,N_28869);
or U33589 (N_33589,N_28942,N_26616);
or U33590 (N_33590,N_27077,N_28211);
xor U33591 (N_33591,N_25875,N_27201);
and U33592 (N_33592,N_26632,N_29635);
nor U33593 (N_33593,N_25871,N_28149);
nand U33594 (N_33594,N_26176,N_25359);
nor U33595 (N_33595,N_26195,N_27857);
and U33596 (N_33596,N_28822,N_27096);
nor U33597 (N_33597,N_25469,N_25698);
or U33598 (N_33598,N_28748,N_28037);
or U33599 (N_33599,N_28330,N_27794);
xor U33600 (N_33600,N_28957,N_28946);
nor U33601 (N_33601,N_28839,N_26851);
nor U33602 (N_33602,N_26473,N_29504);
nor U33603 (N_33603,N_29422,N_29651);
or U33604 (N_33604,N_26808,N_25602);
nor U33605 (N_33605,N_26302,N_25374);
nand U33606 (N_33606,N_28085,N_27342);
and U33607 (N_33607,N_28836,N_28278);
or U33608 (N_33608,N_26215,N_28558);
nand U33609 (N_33609,N_26128,N_25668);
and U33610 (N_33610,N_29929,N_26417);
or U33611 (N_33611,N_25753,N_29224);
nor U33612 (N_33612,N_28150,N_28305);
nor U33613 (N_33613,N_26602,N_28390);
nand U33614 (N_33614,N_26622,N_29382);
nor U33615 (N_33615,N_26939,N_28541);
and U33616 (N_33616,N_29132,N_26190);
or U33617 (N_33617,N_25858,N_29814);
nor U33618 (N_33618,N_26311,N_29020);
nand U33619 (N_33619,N_27914,N_28553);
and U33620 (N_33620,N_25145,N_25075);
and U33621 (N_33621,N_28454,N_28381);
nand U33622 (N_33622,N_25526,N_28584);
or U33623 (N_33623,N_28016,N_26342);
nor U33624 (N_33624,N_27601,N_26111);
or U33625 (N_33625,N_27531,N_26079);
or U33626 (N_33626,N_28967,N_27429);
or U33627 (N_33627,N_29374,N_26370);
and U33628 (N_33628,N_28349,N_26756);
xor U33629 (N_33629,N_29174,N_26329);
or U33630 (N_33630,N_25698,N_26052);
nor U33631 (N_33631,N_29982,N_28238);
nor U33632 (N_33632,N_29345,N_25045);
and U33633 (N_33633,N_29851,N_28863);
and U33634 (N_33634,N_25979,N_29547);
and U33635 (N_33635,N_29105,N_25468);
nand U33636 (N_33636,N_29392,N_29679);
or U33637 (N_33637,N_27658,N_27440);
and U33638 (N_33638,N_28736,N_26116);
or U33639 (N_33639,N_29548,N_25868);
and U33640 (N_33640,N_29061,N_27160);
nand U33641 (N_33641,N_28632,N_26784);
or U33642 (N_33642,N_28579,N_28630);
or U33643 (N_33643,N_28256,N_29987);
or U33644 (N_33644,N_27485,N_28478);
xnor U33645 (N_33645,N_25553,N_27845);
xnor U33646 (N_33646,N_29755,N_27007);
nand U33647 (N_33647,N_29291,N_27703);
nor U33648 (N_33648,N_27405,N_25362);
xnor U33649 (N_33649,N_28767,N_28335);
and U33650 (N_33650,N_29344,N_25906);
and U33651 (N_33651,N_28966,N_26429);
xor U33652 (N_33652,N_27959,N_27845);
nor U33653 (N_33653,N_25028,N_29673);
or U33654 (N_33654,N_29096,N_27374);
nor U33655 (N_33655,N_27856,N_28508);
nor U33656 (N_33656,N_27212,N_26297);
or U33657 (N_33657,N_25423,N_25641);
nor U33658 (N_33658,N_28055,N_25332);
nand U33659 (N_33659,N_26797,N_25773);
and U33660 (N_33660,N_27513,N_25407);
or U33661 (N_33661,N_28991,N_25895);
nor U33662 (N_33662,N_29627,N_25436);
or U33663 (N_33663,N_26048,N_29907);
nand U33664 (N_33664,N_27509,N_27516);
nor U33665 (N_33665,N_26191,N_27797);
and U33666 (N_33666,N_26429,N_25613);
and U33667 (N_33667,N_28770,N_28505);
nor U33668 (N_33668,N_26938,N_27565);
nand U33669 (N_33669,N_25989,N_28684);
and U33670 (N_33670,N_27858,N_25989);
xor U33671 (N_33671,N_25361,N_26049);
or U33672 (N_33672,N_25022,N_26597);
xor U33673 (N_33673,N_27952,N_28742);
and U33674 (N_33674,N_27755,N_25449);
nor U33675 (N_33675,N_29315,N_25958);
xor U33676 (N_33676,N_25430,N_28521);
and U33677 (N_33677,N_26315,N_25352);
or U33678 (N_33678,N_29163,N_25855);
and U33679 (N_33679,N_25092,N_29159);
nand U33680 (N_33680,N_25042,N_27207);
nand U33681 (N_33681,N_28257,N_29500);
nor U33682 (N_33682,N_27190,N_26727);
nor U33683 (N_33683,N_25635,N_29144);
and U33684 (N_33684,N_28351,N_27316);
and U33685 (N_33685,N_25750,N_27920);
nand U33686 (N_33686,N_26940,N_29788);
and U33687 (N_33687,N_26938,N_26266);
nor U33688 (N_33688,N_26664,N_27113);
and U33689 (N_33689,N_25974,N_27791);
or U33690 (N_33690,N_26456,N_26082);
nand U33691 (N_33691,N_28839,N_27407);
nor U33692 (N_33692,N_29010,N_27059);
and U33693 (N_33693,N_26714,N_26578);
xnor U33694 (N_33694,N_29154,N_27600);
nand U33695 (N_33695,N_29793,N_27609);
and U33696 (N_33696,N_28247,N_26932);
xnor U33697 (N_33697,N_25751,N_28339);
and U33698 (N_33698,N_28609,N_29843);
and U33699 (N_33699,N_26700,N_26501);
nor U33700 (N_33700,N_28380,N_27469);
nand U33701 (N_33701,N_29449,N_27877);
or U33702 (N_33702,N_27321,N_26178);
and U33703 (N_33703,N_27857,N_29921);
nor U33704 (N_33704,N_27179,N_27234);
nor U33705 (N_33705,N_25203,N_26962);
and U33706 (N_33706,N_28720,N_27809);
nor U33707 (N_33707,N_29530,N_29561);
or U33708 (N_33708,N_25868,N_25136);
or U33709 (N_33709,N_29846,N_29308);
and U33710 (N_33710,N_29542,N_25449);
and U33711 (N_33711,N_26892,N_26176);
nand U33712 (N_33712,N_28263,N_28503);
and U33713 (N_33713,N_28247,N_26668);
nand U33714 (N_33714,N_28480,N_27094);
or U33715 (N_33715,N_28679,N_25587);
or U33716 (N_33716,N_26320,N_25998);
or U33717 (N_33717,N_26824,N_25332);
nand U33718 (N_33718,N_26547,N_26140);
or U33719 (N_33719,N_29506,N_27924);
and U33720 (N_33720,N_29112,N_27205);
nor U33721 (N_33721,N_27431,N_25394);
xor U33722 (N_33722,N_26417,N_28260);
nor U33723 (N_33723,N_28058,N_28788);
nand U33724 (N_33724,N_26830,N_28571);
and U33725 (N_33725,N_27849,N_27868);
nand U33726 (N_33726,N_26262,N_27046);
and U33727 (N_33727,N_27613,N_29867);
nand U33728 (N_33728,N_29867,N_27990);
nand U33729 (N_33729,N_26675,N_25877);
xnor U33730 (N_33730,N_29738,N_28491);
xor U33731 (N_33731,N_27656,N_29134);
and U33732 (N_33732,N_25148,N_27945);
or U33733 (N_33733,N_26656,N_26449);
nand U33734 (N_33734,N_29797,N_28569);
nand U33735 (N_33735,N_25489,N_25224);
or U33736 (N_33736,N_28105,N_29414);
nor U33737 (N_33737,N_28841,N_28656);
nand U33738 (N_33738,N_27444,N_29645);
or U33739 (N_33739,N_26773,N_28470);
and U33740 (N_33740,N_25504,N_26912);
and U33741 (N_33741,N_28580,N_25745);
nand U33742 (N_33742,N_27650,N_26679);
or U33743 (N_33743,N_28054,N_27044);
nand U33744 (N_33744,N_27246,N_26285);
nor U33745 (N_33745,N_25213,N_28615);
and U33746 (N_33746,N_29087,N_29883);
nand U33747 (N_33747,N_25533,N_29398);
nor U33748 (N_33748,N_25639,N_27307);
or U33749 (N_33749,N_27877,N_29634);
nand U33750 (N_33750,N_27273,N_29937);
or U33751 (N_33751,N_28437,N_25697);
and U33752 (N_33752,N_27871,N_29281);
nor U33753 (N_33753,N_29741,N_25775);
nor U33754 (N_33754,N_27013,N_28728);
or U33755 (N_33755,N_29050,N_25341);
nor U33756 (N_33756,N_28135,N_26381);
and U33757 (N_33757,N_27008,N_27551);
or U33758 (N_33758,N_29237,N_28202);
or U33759 (N_33759,N_26389,N_25517);
nand U33760 (N_33760,N_28555,N_29734);
xor U33761 (N_33761,N_27974,N_28092);
and U33762 (N_33762,N_26644,N_28164);
and U33763 (N_33763,N_25292,N_29934);
xor U33764 (N_33764,N_28776,N_29370);
or U33765 (N_33765,N_26393,N_26795);
or U33766 (N_33766,N_27546,N_25382);
or U33767 (N_33767,N_26088,N_29340);
nor U33768 (N_33768,N_27841,N_27734);
nor U33769 (N_33769,N_26574,N_29454);
nor U33770 (N_33770,N_29856,N_29656);
nand U33771 (N_33771,N_28748,N_26323);
nor U33772 (N_33772,N_25371,N_27108);
or U33773 (N_33773,N_25224,N_27586);
nor U33774 (N_33774,N_29239,N_29945);
and U33775 (N_33775,N_29615,N_29873);
nand U33776 (N_33776,N_25171,N_27221);
xnor U33777 (N_33777,N_25895,N_25663);
nor U33778 (N_33778,N_28452,N_29051);
and U33779 (N_33779,N_28221,N_25907);
nand U33780 (N_33780,N_28378,N_26006);
nor U33781 (N_33781,N_27426,N_27827);
nand U33782 (N_33782,N_27169,N_27328);
xor U33783 (N_33783,N_29091,N_25907);
nor U33784 (N_33784,N_26373,N_29844);
nor U33785 (N_33785,N_29365,N_25758);
nand U33786 (N_33786,N_27827,N_28453);
nor U33787 (N_33787,N_29387,N_26721);
nand U33788 (N_33788,N_25131,N_29401);
or U33789 (N_33789,N_27097,N_27260);
nand U33790 (N_33790,N_26630,N_29424);
and U33791 (N_33791,N_27051,N_27414);
xor U33792 (N_33792,N_27110,N_26170);
nand U33793 (N_33793,N_27515,N_25174);
nor U33794 (N_33794,N_29904,N_25087);
nand U33795 (N_33795,N_27241,N_26031);
and U33796 (N_33796,N_25893,N_25245);
nor U33797 (N_33797,N_25770,N_28101);
and U33798 (N_33798,N_28261,N_25311);
nor U33799 (N_33799,N_27080,N_25636);
or U33800 (N_33800,N_28779,N_27252);
xnor U33801 (N_33801,N_28625,N_26317);
nand U33802 (N_33802,N_28078,N_25202);
xor U33803 (N_33803,N_28001,N_26023);
and U33804 (N_33804,N_28388,N_25413);
nor U33805 (N_33805,N_28722,N_29544);
nand U33806 (N_33806,N_28275,N_26217);
or U33807 (N_33807,N_27384,N_25776);
or U33808 (N_33808,N_28647,N_27037);
nand U33809 (N_33809,N_29716,N_29051);
nand U33810 (N_33810,N_26197,N_28127);
nor U33811 (N_33811,N_25231,N_28418);
or U33812 (N_33812,N_25573,N_27055);
and U33813 (N_33813,N_26275,N_25126);
nand U33814 (N_33814,N_29241,N_25542);
nor U33815 (N_33815,N_26673,N_29315);
and U33816 (N_33816,N_29653,N_27323);
nor U33817 (N_33817,N_26654,N_28785);
nand U33818 (N_33818,N_27123,N_25269);
nor U33819 (N_33819,N_29626,N_29995);
or U33820 (N_33820,N_29738,N_27279);
nand U33821 (N_33821,N_29453,N_28308);
or U33822 (N_33822,N_29538,N_27651);
or U33823 (N_33823,N_29610,N_26186);
nand U33824 (N_33824,N_29271,N_26537);
or U33825 (N_33825,N_28531,N_26677);
nand U33826 (N_33826,N_27323,N_27564);
or U33827 (N_33827,N_29482,N_28288);
or U33828 (N_33828,N_26466,N_29607);
and U33829 (N_33829,N_28409,N_25629);
xor U33830 (N_33830,N_25740,N_28643);
and U33831 (N_33831,N_28182,N_28047);
nor U33832 (N_33832,N_28139,N_28678);
nor U33833 (N_33833,N_29562,N_26081);
and U33834 (N_33834,N_25690,N_26586);
and U33835 (N_33835,N_28893,N_25712);
and U33836 (N_33836,N_27969,N_29073);
and U33837 (N_33837,N_26612,N_29727);
or U33838 (N_33838,N_27475,N_26574);
nor U33839 (N_33839,N_27364,N_27845);
and U33840 (N_33840,N_25806,N_27593);
and U33841 (N_33841,N_28851,N_29041);
and U33842 (N_33842,N_26765,N_29865);
or U33843 (N_33843,N_25076,N_28824);
or U33844 (N_33844,N_27580,N_27638);
or U33845 (N_33845,N_29695,N_29335);
or U33846 (N_33846,N_27746,N_28991);
and U33847 (N_33847,N_28200,N_25506);
nor U33848 (N_33848,N_26314,N_26869);
and U33849 (N_33849,N_28614,N_26765);
nand U33850 (N_33850,N_27648,N_27995);
or U33851 (N_33851,N_25900,N_29382);
and U33852 (N_33852,N_25939,N_27100);
or U33853 (N_33853,N_29027,N_27917);
xor U33854 (N_33854,N_27858,N_26995);
nand U33855 (N_33855,N_28743,N_29423);
and U33856 (N_33856,N_28550,N_28318);
and U33857 (N_33857,N_26154,N_28131);
and U33858 (N_33858,N_26286,N_28478);
and U33859 (N_33859,N_25923,N_27786);
nor U33860 (N_33860,N_28893,N_28554);
nor U33861 (N_33861,N_28411,N_25078);
nand U33862 (N_33862,N_26330,N_26450);
nor U33863 (N_33863,N_27006,N_28688);
or U33864 (N_33864,N_29876,N_26025);
or U33865 (N_33865,N_25868,N_25652);
nand U33866 (N_33866,N_25883,N_27935);
nand U33867 (N_33867,N_28998,N_26562);
nand U33868 (N_33868,N_27340,N_27589);
and U33869 (N_33869,N_25600,N_29361);
or U33870 (N_33870,N_26065,N_27994);
nor U33871 (N_33871,N_25772,N_28172);
nor U33872 (N_33872,N_25290,N_28937);
and U33873 (N_33873,N_26372,N_25532);
or U33874 (N_33874,N_27312,N_26730);
or U33875 (N_33875,N_25920,N_28261);
and U33876 (N_33876,N_27316,N_26198);
and U33877 (N_33877,N_28189,N_28185);
xor U33878 (N_33878,N_29018,N_26585);
nand U33879 (N_33879,N_28160,N_25754);
and U33880 (N_33880,N_27243,N_29181);
nand U33881 (N_33881,N_28746,N_26686);
nand U33882 (N_33882,N_27632,N_28237);
and U33883 (N_33883,N_26530,N_26804);
or U33884 (N_33884,N_27413,N_26361);
or U33885 (N_33885,N_25401,N_26556);
nor U33886 (N_33886,N_25746,N_28786);
nor U33887 (N_33887,N_25340,N_25850);
nand U33888 (N_33888,N_25700,N_29138);
or U33889 (N_33889,N_28042,N_27459);
or U33890 (N_33890,N_29683,N_29397);
or U33891 (N_33891,N_26762,N_28125);
and U33892 (N_33892,N_26355,N_27164);
nand U33893 (N_33893,N_29383,N_29736);
nand U33894 (N_33894,N_25429,N_29869);
xor U33895 (N_33895,N_27933,N_28505);
xor U33896 (N_33896,N_28168,N_25961);
and U33897 (N_33897,N_26335,N_27311);
and U33898 (N_33898,N_26869,N_25995);
nand U33899 (N_33899,N_25256,N_26204);
nor U33900 (N_33900,N_28815,N_28843);
and U33901 (N_33901,N_26017,N_27436);
or U33902 (N_33902,N_27532,N_27007);
nand U33903 (N_33903,N_27108,N_26502);
or U33904 (N_33904,N_25163,N_27985);
nor U33905 (N_33905,N_26300,N_28350);
and U33906 (N_33906,N_27135,N_27819);
xnor U33907 (N_33907,N_27455,N_26381);
and U33908 (N_33908,N_25684,N_28427);
and U33909 (N_33909,N_27771,N_29458);
nor U33910 (N_33910,N_25797,N_28852);
and U33911 (N_33911,N_26666,N_27193);
nand U33912 (N_33912,N_25964,N_26863);
xor U33913 (N_33913,N_27165,N_25835);
nor U33914 (N_33914,N_29134,N_26070);
nor U33915 (N_33915,N_28480,N_27042);
nor U33916 (N_33916,N_29208,N_28337);
or U33917 (N_33917,N_26803,N_28893);
or U33918 (N_33918,N_27894,N_26367);
and U33919 (N_33919,N_25699,N_26597);
nor U33920 (N_33920,N_28554,N_28637);
nand U33921 (N_33921,N_27889,N_25289);
nor U33922 (N_33922,N_26382,N_29929);
xnor U33923 (N_33923,N_26536,N_29139);
nor U33924 (N_33924,N_26258,N_25958);
and U33925 (N_33925,N_29533,N_28889);
and U33926 (N_33926,N_25701,N_26288);
nand U33927 (N_33927,N_28144,N_28074);
nand U33928 (N_33928,N_27445,N_27060);
nor U33929 (N_33929,N_26847,N_28545);
xnor U33930 (N_33930,N_27845,N_29883);
or U33931 (N_33931,N_29633,N_29446);
nor U33932 (N_33932,N_28935,N_25449);
nor U33933 (N_33933,N_28542,N_25040);
and U33934 (N_33934,N_26471,N_26918);
nand U33935 (N_33935,N_29869,N_29037);
or U33936 (N_33936,N_29900,N_25793);
nand U33937 (N_33937,N_25646,N_29831);
and U33938 (N_33938,N_29522,N_25904);
or U33939 (N_33939,N_29283,N_26887);
nand U33940 (N_33940,N_29884,N_25498);
nand U33941 (N_33941,N_25687,N_26553);
xnor U33942 (N_33942,N_29372,N_29100);
nand U33943 (N_33943,N_25053,N_29521);
nor U33944 (N_33944,N_26721,N_27580);
or U33945 (N_33945,N_29201,N_26204);
nor U33946 (N_33946,N_26814,N_26250);
nand U33947 (N_33947,N_29454,N_28670);
and U33948 (N_33948,N_29235,N_26483);
and U33949 (N_33949,N_25764,N_29298);
nand U33950 (N_33950,N_28889,N_28334);
and U33951 (N_33951,N_28278,N_27742);
nor U33952 (N_33952,N_29679,N_25823);
nor U33953 (N_33953,N_27353,N_26572);
and U33954 (N_33954,N_27636,N_27816);
nor U33955 (N_33955,N_25935,N_29847);
nand U33956 (N_33956,N_28563,N_25702);
nor U33957 (N_33957,N_29594,N_28717);
nor U33958 (N_33958,N_27133,N_25718);
or U33959 (N_33959,N_28212,N_26298);
nor U33960 (N_33960,N_29786,N_26455);
and U33961 (N_33961,N_27651,N_28464);
and U33962 (N_33962,N_29396,N_26054);
or U33963 (N_33963,N_28463,N_27221);
and U33964 (N_33964,N_25200,N_28254);
and U33965 (N_33965,N_28600,N_27397);
nand U33966 (N_33966,N_29345,N_26878);
and U33967 (N_33967,N_29290,N_27768);
or U33968 (N_33968,N_27131,N_29551);
and U33969 (N_33969,N_29876,N_26109);
nor U33970 (N_33970,N_26044,N_26745);
nand U33971 (N_33971,N_25698,N_28023);
nor U33972 (N_33972,N_26836,N_27459);
and U33973 (N_33973,N_26262,N_28973);
nand U33974 (N_33974,N_27024,N_27056);
nor U33975 (N_33975,N_26379,N_26626);
and U33976 (N_33976,N_28471,N_27724);
nor U33977 (N_33977,N_26929,N_25968);
nand U33978 (N_33978,N_26183,N_28375);
nor U33979 (N_33979,N_25328,N_29600);
nor U33980 (N_33980,N_27425,N_26961);
nor U33981 (N_33981,N_27151,N_28333);
and U33982 (N_33982,N_27310,N_29322);
or U33983 (N_33983,N_28963,N_25052);
or U33984 (N_33984,N_27059,N_26168);
xor U33985 (N_33985,N_28923,N_27262);
nand U33986 (N_33986,N_28767,N_25749);
or U33987 (N_33987,N_25171,N_26631);
and U33988 (N_33988,N_28117,N_27745);
and U33989 (N_33989,N_26214,N_28751);
nor U33990 (N_33990,N_26428,N_28023);
nand U33991 (N_33991,N_26669,N_26062);
and U33992 (N_33992,N_28473,N_28544);
nor U33993 (N_33993,N_29799,N_27319);
or U33994 (N_33994,N_26938,N_25458);
nor U33995 (N_33995,N_26435,N_28432);
and U33996 (N_33996,N_26868,N_28952);
xnor U33997 (N_33997,N_27982,N_28916);
or U33998 (N_33998,N_26687,N_29811);
nor U33999 (N_33999,N_28592,N_27480);
xnor U34000 (N_34000,N_26372,N_29911);
or U34001 (N_34001,N_28726,N_29631);
or U34002 (N_34002,N_26891,N_27976);
or U34003 (N_34003,N_27256,N_25433);
nand U34004 (N_34004,N_27446,N_29877);
or U34005 (N_34005,N_29792,N_26823);
or U34006 (N_34006,N_29862,N_25453);
nor U34007 (N_34007,N_28432,N_25920);
xnor U34008 (N_34008,N_25171,N_25748);
nor U34009 (N_34009,N_28159,N_25179);
and U34010 (N_34010,N_29916,N_26868);
nand U34011 (N_34011,N_29841,N_27681);
or U34012 (N_34012,N_28334,N_27500);
nor U34013 (N_34013,N_28343,N_27654);
and U34014 (N_34014,N_26465,N_28873);
or U34015 (N_34015,N_25941,N_29090);
or U34016 (N_34016,N_25276,N_25992);
and U34017 (N_34017,N_27785,N_26308);
nor U34018 (N_34018,N_27566,N_26340);
and U34019 (N_34019,N_25824,N_25097);
nand U34020 (N_34020,N_28845,N_27579);
or U34021 (N_34021,N_28997,N_27543);
nor U34022 (N_34022,N_29606,N_28774);
and U34023 (N_34023,N_25073,N_27528);
nor U34024 (N_34024,N_25090,N_25258);
and U34025 (N_34025,N_25367,N_28869);
and U34026 (N_34026,N_28419,N_27780);
nor U34027 (N_34027,N_28994,N_29598);
nand U34028 (N_34028,N_27071,N_29920);
and U34029 (N_34029,N_27596,N_29689);
nand U34030 (N_34030,N_28262,N_28197);
and U34031 (N_34031,N_25264,N_25969);
or U34032 (N_34032,N_26671,N_27719);
or U34033 (N_34033,N_25681,N_28856);
nand U34034 (N_34034,N_26246,N_28573);
nand U34035 (N_34035,N_27833,N_27939);
or U34036 (N_34036,N_29293,N_29057);
or U34037 (N_34037,N_29423,N_25078);
and U34038 (N_34038,N_26247,N_27662);
and U34039 (N_34039,N_27708,N_27311);
nor U34040 (N_34040,N_25926,N_26728);
or U34041 (N_34041,N_25960,N_27666);
nand U34042 (N_34042,N_26908,N_25330);
xnor U34043 (N_34043,N_26722,N_29459);
nor U34044 (N_34044,N_28113,N_26433);
or U34045 (N_34045,N_29764,N_28954);
nand U34046 (N_34046,N_28761,N_26810);
or U34047 (N_34047,N_29373,N_25814);
xnor U34048 (N_34048,N_28333,N_27520);
nand U34049 (N_34049,N_25474,N_28055);
or U34050 (N_34050,N_25327,N_26400);
nor U34051 (N_34051,N_27252,N_29508);
xor U34052 (N_34052,N_29545,N_27312);
or U34053 (N_34053,N_26865,N_27590);
or U34054 (N_34054,N_27638,N_25448);
xnor U34055 (N_34055,N_29190,N_27245);
and U34056 (N_34056,N_26686,N_28652);
and U34057 (N_34057,N_29353,N_27572);
nand U34058 (N_34058,N_27604,N_28472);
and U34059 (N_34059,N_25563,N_27224);
and U34060 (N_34060,N_26708,N_27313);
and U34061 (N_34061,N_26995,N_26078);
nand U34062 (N_34062,N_26735,N_29836);
nor U34063 (N_34063,N_28888,N_27955);
and U34064 (N_34064,N_26375,N_29638);
or U34065 (N_34065,N_27986,N_28099);
xnor U34066 (N_34066,N_27150,N_25007);
xor U34067 (N_34067,N_27685,N_28874);
nand U34068 (N_34068,N_26895,N_27517);
nand U34069 (N_34069,N_29387,N_29428);
or U34070 (N_34070,N_25076,N_27642);
nand U34071 (N_34071,N_26115,N_29479);
or U34072 (N_34072,N_25784,N_25909);
and U34073 (N_34073,N_27073,N_27358);
or U34074 (N_34074,N_25743,N_27363);
or U34075 (N_34075,N_25018,N_28096);
nand U34076 (N_34076,N_28352,N_26809);
nand U34077 (N_34077,N_26964,N_27042);
and U34078 (N_34078,N_28110,N_27907);
xor U34079 (N_34079,N_29489,N_28257);
nand U34080 (N_34080,N_29150,N_25059);
nand U34081 (N_34081,N_28103,N_27691);
nand U34082 (N_34082,N_27126,N_26265);
nand U34083 (N_34083,N_27021,N_28841);
and U34084 (N_34084,N_29595,N_29994);
nand U34085 (N_34085,N_27828,N_29081);
nand U34086 (N_34086,N_28786,N_26691);
xor U34087 (N_34087,N_29886,N_26296);
nand U34088 (N_34088,N_25436,N_28036);
nor U34089 (N_34089,N_26436,N_25206);
nor U34090 (N_34090,N_29465,N_26104);
and U34091 (N_34091,N_25614,N_29226);
nand U34092 (N_34092,N_29361,N_28169);
nor U34093 (N_34093,N_27751,N_27533);
xor U34094 (N_34094,N_25363,N_27742);
nand U34095 (N_34095,N_29307,N_28501);
and U34096 (N_34096,N_25533,N_29269);
and U34097 (N_34097,N_26811,N_27595);
xnor U34098 (N_34098,N_25448,N_25158);
and U34099 (N_34099,N_27894,N_27608);
nor U34100 (N_34100,N_27186,N_29419);
and U34101 (N_34101,N_29558,N_27581);
nand U34102 (N_34102,N_27096,N_29700);
or U34103 (N_34103,N_29906,N_27407);
nand U34104 (N_34104,N_26627,N_29410);
nand U34105 (N_34105,N_27578,N_26905);
and U34106 (N_34106,N_27082,N_28021);
and U34107 (N_34107,N_25724,N_25875);
xor U34108 (N_34108,N_28015,N_29899);
and U34109 (N_34109,N_26042,N_28252);
and U34110 (N_34110,N_28969,N_25469);
or U34111 (N_34111,N_26401,N_29959);
nor U34112 (N_34112,N_25567,N_25307);
nor U34113 (N_34113,N_25576,N_25908);
xor U34114 (N_34114,N_29097,N_28692);
nand U34115 (N_34115,N_28710,N_25965);
nor U34116 (N_34116,N_25828,N_26596);
and U34117 (N_34117,N_28954,N_25049);
nand U34118 (N_34118,N_25980,N_25834);
or U34119 (N_34119,N_27611,N_28444);
and U34120 (N_34120,N_26444,N_26501);
and U34121 (N_34121,N_29285,N_26545);
nor U34122 (N_34122,N_29482,N_26229);
or U34123 (N_34123,N_28224,N_27450);
or U34124 (N_34124,N_25827,N_26074);
and U34125 (N_34125,N_27826,N_27329);
or U34126 (N_34126,N_29335,N_25727);
or U34127 (N_34127,N_28095,N_29753);
nor U34128 (N_34128,N_25494,N_27267);
and U34129 (N_34129,N_25318,N_29950);
nand U34130 (N_34130,N_25595,N_29973);
or U34131 (N_34131,N_29373,N_26411);
xnor U34132 (N_34132,N_29937,N_25065);
or U34133 (N_34133,N_25883,N_25829);
nor U34134 (N_34134,N_28275,N_25088);
nor U34135 (N_34135,N_29022,N_28839);
xnor U34136 (N_34136,N_25947,N_28324);
or U34137 (N_34137,N_27110,N_28325);
nand U34138 (N_34138,N_28706,N_27650);
nor U34139 (N_34139,N_27639,N_29397);
and U34140 (N_34140,N_27223,N_28877);
and U34141 (N_34141,N_29713,N_28451);
or U34142 (N_34142,N_28000,N_25850);
nor U34143 (N_34143,N_28433,N_28266);
nand U34144 (N_34144,N_29695,N_29892);
and U34145 (N_34145,N_29771,N_28140);
and U34146 (N_34146,N_29036,N_26961);
nor U34147 (N_34147,N_27487,N_26208);
xor U34148 (N_34148,N_29930,N_25568);
nor U34149 (N_34149,N_27381,N_26224);
or U34150 (N_34150,N_25099,N_25054);
or U34151 (N_34151,N_27285,N_28873);
and U34152 (N_34152,N_26052,N_25448);
xor U34153 (N_34153,N_25968,N_26020);
nand U34154 (N_34154,N_27439,N_25936);
or U34155 (N_34155,N_28943,N_28699);
xnor U34156 (N_34156,N_26486,N_26758);
nand U34157 (N_34157,N_25562,N_26928);
and U34158 (N_34158,N_28364,N_28101);
xor U34159 (N_34159,N_28508,N_25235);
nand U34160 (N_34160,N_29503,N_25175);
nand U34161 (N_34161,N_28964,N_29968);
or U34162 (N_34162,N_29079,N_29938);
nor U34163 (N_34163,N_26254,N_27042);
or U34164 (N_34164,N_29999,N_29980);
or U34165 (N_34165,N_26812,N_26978);
or U34166 (N_34166,N_26314,N_26159);
nor U34167 (N_34167,N_27573,N_28641);
nor U34168 (N_34168,N_28713,N_27851);
or U34169 (N_34169,N_26911,N_29208);
nand U34170 (N_34170,N_28756,N_29775);
nor U34171 (N_34171,N_25377,N_26286);
nor U34172 (N_34172,N_26325,N_28389);
nor U34173 (N_34173,N_28329,N_26630);
nor U34174 (N_34174,N_27382,N_26367);
nand U34175 (N_34175,N_27905,N_26622);
nor U34176 (N_34176,N_25136,N_27740);
and U34177 (N_34177,N_28328,N_27490);
or U34178 (N_34178,N_26032,N_29413);
or U34179 (N_34179,N_29447,N_25845);
nand U34180 (N_34180,N_25972,N_28627);
xor U34181 (N_34181,N_27414,N_25153);
nand U34182 (N_34182,N_29008,N_29651);
nand U34183 (N_34183,N_25405,N_29279);
and U34184 (N_34184,N_26314,N_27724);
or U34185 (N_34185,N_29174,N_25008);
nor U34186 (N_34186,N_27281,N_29307);
and U34187 (N_34187,N_25249,N_29583);
and U34188 (N_34188,N_28873,N_28914);
or U34189 (N_34189,N_25740,N_27853);
nand U34190 (N_34190,N_27031,N_26645);
nor U34191 (N_34191,N_27636,N_25445);
nand U34192 (N_34192,N_28259,N_27795);
and U34193 (N_34193,N_26985,N_28894);
xnor U34194 (N_34194,N_29018,N_25954);
or U34195 (N_34195,N_29068,N_26325);
nor U34196 (N_34196,N_28704,N_29070);
or U34197 (N_34197,N_29764,N_28863);
or U34198 (N_34198,N_29884,N_27882);
or U34199 (N_34199,N_27237,N_28280);
nor U34200 (N_34200,N_26180,N_25660);
nor U34201 (N_34201,N_28611,N_28319);
and U34202 (N_34202,N_29115,N_29349);
xor U34203 (N_34203,N_28813,N_26801);
nor U34204 (N_34204,N_29153,N_29646);
nor U34205 (N_34205,N_25163,N_28963);
and U34206 (N_34206,N_29034,N_26455);
or U34207 (N_34207,N_27949,N_28077);
nand U34208 (N_34208,N_26685,N_26484);
nand U34209 (N_34209,N_28721,N_28977);
and U34210 (N_34210,N_25266,N_29092);
xnor U34211 (N_34211,N_25210,N_26354);
nand U34212 (N_34212,N_28544,N_29522);
or U34213 (N_34213,N_26083,N_28492);
nor U34214 (N_34214,N_26531,N_28195);
nand U34215 (N_34215,N_29005,N_28666);
and U34216 (N_34216,N_29328,N_28387);
nand U34217 (N_34217,N_25499,N_29986);
nor U34218 (N_34218,N_27220,N_27608);
nor U34219 (N_34219,N_26434,N_26275);
and U34220 (N_34220,N_29078,N_25411);
nor U34221 (N_34221,N_26175,N_27505);
xnor U34222 (N_34222,N_29207,N_27274);
or U34223 (N_34223,N_29053,N_29281);
nand U34224 (N_34224,N_28880,N_29523);
nor U34225 (N_34225,N_26738,N_27926);
nor U34226 (N_34226,N_27305,N_27292);
nand U34227 (N_34227,N_28496,N_29085);
and U34228 (N_34228,N_25037,N_26595);
xnor U34229 (N_34229,N_27534,N_26071);
nor U34230 (N_34230,N_26952,N_27366);
and U34231 (N_34231,N_27723,N_29627);
or U34232 (N_34232,N_26616,N_29833);
or U34233 (N_34233,N_26204,N_26140);
nand U34234 (N_34234,N_27223,N_25968);
or U34235 (N_34235,N_29722,N_29402);
or U34236 (N_34236,N_27083,N_28639);
nand U34237 (N_34237,N_25265,N_27363);
or U34238 (N_34238,N_26848,N_29664);
or U34239 (N_34239,N_27800,N_26930);
or U34240 (N_34240,N_29635,N_28034);
and U34241 (N_34241,N_29632,N_25408);
or U34242 (N_34242,N_25877,N_26907);
nand U34243 (N_34243,N_28207,N_28486);
and U34244 (N_34244,N_25011,N_28872);
nand U34245 (N_34245,N_26715,N_26658);
and U34246 (N_34246,N_27723,N_28667);
nor U34247 (N_34247,N_28484,N_28995);
or U34248 (N_34248,N_26931,N_26716);
or U34249 (N_34249,N_26121,N_25965);
nor U34250 (N_34250,N_27810,N_28645);
nor U34251 (N_34251,N_25030,N_26396);
nand U34252 (N_34252,N_25151,N_28592);
or U34253 (N_34253,N_26489,N_29334);
and U34254 (N_34254,N_26515,N_25186);
or U34255 (N_34255,N_29352,N_28566);
and U34256 (N_34256,N_29413,N_26116);
or U34257 (N_34257,N_26643,N_28779);
nor U34258 (N_34258,N_26389,N_26999);
nand U34259 (N_34259,N_27478,N_29547);
xor U34260 (N_34260,N_27099,N_28849);
nor U34261 (N_34261,N_27093,N_26627);
or U34262 (N_34262,N_29470,N_27000);
or U34263 (N_34263,N_26512,N_26993);
nor U34264 (N_34264,N_26446,N_27513);
nor U34265 (N_34265,N_26954,N_26055);
and U34266 (N_34266,N_27191,N_27337);
xnor U34267 (N_34267,N_26476,N_27716);
xor U34268 (N_34268,N_27707,N_29686);
nor U34269 (N_34269,N_29600,N_26136);
nand U34270 (N_34270,N_27587,N_25260);
nand U34271 (N_34271,N_27365,N_27537);
nand U34272 (N_34272,N_26856,N_27450);
or U34273 (N_34273,N_25302,N_27448);
nor U34274 (N_34274,N_29076,N_28606);
and U34275 (N_34275,N_25832,N_26372);
nor U34276 (N_34276,N_26932,N_29119);
or U34277 (N_34277,N_26001,N_27241);
xor U34278 (N_34278,N_25243,N_29238);
nor U34279 (N_34279,N_26050,N_25433);
nand U34280 (N_34280,N_27558,N_28257);
or U34281 (N_34281,N_29558,N_27159);
or U34282 (N_34282,N_29159,N_25147);
nor U34283 (N_34283,N_27099,N_29619);
nor U34284 (N_34284,N_25460,N_26056);
nand U34285 (N_34285,N_28190,N_29135);
and U34286 (N_34286,N_26530,N_25599);
nor U34287 (N_34287,N_26641,N_25829);
nor U34288 (N_34288,N_26239,N_26413);
nor U34289 (N_34289,N_29328,N_27000);
or U34290 (N_34290,N_28416,N_25274);
or U34291 (N_34291,N_25604,N_26787);
and U34292 (N_34292,N_27307,N_29214);
xor U34293 (N_34293,N_26122,N_29062);
xnor U34294 (N_34294,N_25492,N_25270);
or U34295 (N_34295,N_25079,N_26785);
nand U34296 (N_34296,N_27348,N_26650);
or U34297 (N_34297,N_29944,N_26234);
or U34298 (N_34298,N_25896,N_25195);
nand U34299 (N_34299,N_26199,N_25312);
xor U34300 (N_34300,N_28436,N_28197);
nand U34301 (N_34301,N_29646,N_27869);
nand U34302 (N_34302,N_27722,N_25412);
and U34303 (N_34303,N_25887,N_26684);
nor U34304 (N_34304,N_27666,N_28931);
or U34305 (N_34305,N_29863,N_28334);
nand U34306 (N_34306,N_28054,N_27874);
nand U34307 (N_34307,N_26911,N_28007);
nand U34308 (N_34308,N_29781,N_25687);
or U34309 (N_34309,N_27286,N_29864);
nor U34310 (N_34310,N_29273,N_29605);
and U34311 (N_34311,N_26557,N_25073);
and U34312 (N_34312,N_25972,N_26474);
nor U34313 (N_34313,N_29904,N_25013);
or U34314 (N_34314,N_29962,N_26153);
xnor U34315 (N_34315,N_28521,N_26297);
and U34316 (N_34316,N_26618,N_29323);
nand U34317 (N_34317,N_28130,N_25843);
xnor U34318 (N_34318,N_27790,N_27725);
or U34319 (N_34319,N_28629,N_26576);
nor U34320 (N_34320,N_26491,N_26854);
xnor U34321 (N_34321,N_29173,N_25577);
xor U34322 (N_34322,N_27678,N_28114);
nor U34323 (N_34323,N_28187,N_27864);
xor U34324 (N_34324,N_29822,N_26373);
nor U34325 (N_34325,N_28446,N_27981);
nand U34326 (N_34326,N_28346,N_29946);
or U34327 (N_34327,N_26310,N_28716);
nor U34328 (N_34328,N_27666,N_28586);
nand U34329 (N_34329,N_28348,N_28016);
xor U34330 (N_34330,N_25456,N_25390);
xnor U34331 (N_34331,N_26702,N_28849);
xnor U34332 (N_34332,N_29917,N_27059);
nor U34333 (N_34333,N_25630,N_28705);
and U34334 (N_34334,N_28574,N_29493);
or U34335 (N_34335,N_27799,N_28183);
nor U34336 (N_34336,N_28544,N_27707);
or U34337 (N_34337,N_27979,N_27649);
nand U34338 (N_34338,N_29704,N_28647);
nor U34339 (N_34339,N_29333,N_26964);
or U34340 (N_34340,N_28939,N_29122);
or U34341 (N_34341,N_26519,N_29401);
and U34342 (N_34342,N_28362,N_29494);
or U34343 (N_34343,N_27367,N_27531);
nand U34344 (N_34344,N_28448,N_28184);
or U34345 (N_34345,N_26955,N_27243);
nand U34346 (N_34346,N_28337,N_27646);
or U34347 (N_34347,N_28285,N_26467);
nor U34348 (N_34348,N_28495,N_26748);
nand U34349 (N_34349,N_29305,N_28075);
nor U34350 (N_34350,N_26474,N_29688);
xor U34351 (N_34351,N_27728,N_26817);
nand U34352 (N_34352,N_25993,N_26601);
or U34353 (N_34353,N_27594,N_27661);
or U34354 (N_34354,N_29852,N_27811);
nand U34355 (N_34355,N_29496,N_28372);
nand U34356 (N_34356,N_29930,N_28511);
xor U34357 (N_34357,N_27152,N_27442);
xnor U34358 (N_34358,N_27704,N_29088);
nand U34359 (N_34359,N_29136,N_27112);
nor U34360 (N_34360,N_26804,N_26575);
xor U34361 (N_34361,N_26404,N_28103);
and U34362 (N_34362,N_29577,N_25936);
nand U34363 (N_34363,N_27998,N_26570);
xor U34364 (N_34364,N_28915,N_27574);
or U34365 (N_34365,N_29753,N_27176);
or U34366 (N_34366,N_25678,N_28445);
and U34367 (N_34367,N_27507,N_26914);
nand U34368 (N_34368,N_28729,N_25012);
and U34369 (N_34369,N_29290,N_27258);
xnor U34370 (N_34370,N_25938,N_27153);
nor U34371 (N_34371,N_25918,N_28132);
nor U34372 (N_34372,N_26446,N_27426);
and U34373 (N_34373,N_27537,N_25405);
nor U34374 (N_34374,N_28661,N_28937);
nand U34375 (N_34375,N_26000,N_27831);
and U34376 (N_34376,N_26185,N_25042);
nand U34377 (N_34377,N_26121,N_26650);
or U34378 (N_34378,N_29343,N_25623);
and U34379 (N_34379,N_28668,N_29480);
nor U34380 (N_34380,N_28240,N_27764);
nor U34381 (N_34381,N_27551,N_28786);
nand U34382 (N_34382,N_26425,N_29638);
xor U34383 (N_34383,N_26009,N_28653);
nor U34384 (N_34384,N_28517,N_25117);
or U34385 (N_34385,N_26644,N_27290);
xor U34386 (N_34386,N_27513,N_25416);
xnor U34387 (N_34387,N_27477,N_25396);
and U34388 (N_34388,N_28594,N_27626);
nand U34389 (N_34389,N_25690,N_26913);
or U34390 (N_34390,N_29105,N_28909);
and U34391 (N_34391,N_29046,N_28634);
nand U34392 (N_34392,N_28214,N_27193);
or U34393 (N_34393,N_28697,N_25214);
nor U34394 (N_34394,N_28114,N_26461);
and U34395 (N_34395,N_25759,N_29316);
or U34396 (N_34396,N_25306,N_29983);
nand U34397 (N_34397,N_29964,N_25823);
nor U34398 (N_34398,N_25125,N_28356);
or U34399 (N_34399,N_27604,N_27721);
or U34400 (N_34400,N_28567,N_27872);
nor U34401 (N_34401,N_26634,N_25673);
and U34402 (N_34402,N_25432,N_25132);
nor U34403 (N_34403,N_26886,N_26593);
or U34404 (N_34404,N_29015,N_26365);
nand U34405 (N_34405,N_29081,N_25553);
nand U34406 (N_34406,N_25147,N_26137);
and U34407 (N_34407,N_26214,N_28565);
and U34408 (N_34408,N_29766,N_29941);
and U34409 (N_34409,N_26908,N_28760);
nand U34410 (N_34410,N_27949,N_27924);
nand U34411 (N_34411,N_28892,N_25812);
nand U34412 (N_34412,N_25154,N_27936);
nand U34413 (N_34413,N_27076,N_28005);
or U34414 (N_34414,N_28655,N_29274);
nor U34415 (N_34415,N_28686,N_29518);
or U34416 (N_34416,N_26159,N_26712);
and U34417 (N_34417,N_28180,N_29424);
nand U34418 (N_34418,N_26024,N_26334);
nor U34419 (N_34419,N_28056,N_27376);
nand U34420 (N_34420,N_27901,N_28349);
nand U34421 (N_34421,N_27860,N_29643);
nand U34422 (N_34422,N_29650,N_28613);
or U34423 (N_34423,N_27667,N_26536);
and U34424 (N_34424,N_27038,N_28045);
or U34425 (N_34425,N_25233,N_29118);
and U34426 (N_34426,N_26013,N_27006);
or U34427 (N_34427,N_27188,N_29032);
nor U34428 (N_34428,N_28922,N_25356);
nor U34429 (N_34429,N_26522,N_27441);
and U34430 (N_34430,N_27841,N_27687);
or U34431 (N_34431,N_29100,N_25026);
and U34432 (N_34432,N_25496,N_27709);
or U34433 (N_34433,N_26553,N_29074);
and U34434 (N_34434,N_25364,N_27945);
nor U34435 (N_34435,N_28179,N_28767);
nor U34436 (N_34436,N_25537,N_26906);
and U34437 (N_34437,N_29101,N_28034);
and U34438 (N_34438,N_29120,N_27790);
or U34439 (N_34439,N_29177,N_27629);
xnor U34440 (N_34440,N_25043,N_26602);
and U34441 (N_34441,N_28896,N_29925);
nor U34442 (N_34442,N_25719,N_25937);
nor U34443 (N_34443,N_28390,N_25368);
nand U34444 (N_34444,N_26621,N_28585);
xor U34445 (N_34445,N_27993,N_26446);
nor U34446 (N_34446,N_29780,N_29082);
or U34447 (N_34447,N_29029,N_25047);
nor U34448 (N_34448,N_27787,N_25414);
nand U34449 (N_34449,N_27936,N_26844);
nor U34450 (N_34450,N_25107,N_26907);
nand U34451 (N_34451,N_26381,N_26742);
and U34452 (N_34452,N_25867,N_26534);
nand U34453 (N_34453,N_27993,N_25508);
nor U34454 (N_34454,N_29294,N_26927);
nor U34455 (N_34455,N_26095,N_29042);
and U34456 (N_34456,N_29358,N_25855);
xnor U34457 (N_34457,N_28567,N_25722);
xor U34458 (N_34458,N_29886,N_26713);
xor U34459 (N_34459,N_28686,N_27013);
or U34460 (N_34460,N_27633,N_27085);
nor U34461 (N_34461,N_25444,N_28863);
nand U34462 (N_34462,N_29074,N_25203);
and U34463 (N_34463,N_25553,N_26996);
nand U34464 (N_34464,N_28416,N_26032);
and U34465 (N_34465,N_25321,N_25921);
nand U34466 (N_34466,N_25767,N_29771);
and U34467 (N_34467,N_26340,N_28290);
nand U34468 (N_34468,N_25300,N_27429);
and U34469 (N_34469,N_29307,N_25328);
nand U34470 (N_34470,N_28354,N_27080);
or U34471 (N_34471,N_26433,N_27066);
or U34472 (N_34472,N_26564,N_28983);
nand U34473 (N_34473,N_27125,N_27652);
nand U34474 (N_34474,N_25717,N_28784);
nor U34475 (N_34475,N_27803,N_29190);
and U34476 (N_34476,N_29632,N_29863);
nand U34477 (N_34477,N_27267,N_26338);
nor U34478 (N_34478,N_28074,N_29645);
xnor U34479 (N_34479,N_27935,N_29748);
nor U34480 (N_34480,N_29598,N_29733);
or U34481 (N_34481,N_29611,N_27644);
nand U34482 (N_34482,N_26216,N_28088);
or U34483 (N_34483,N_26468,N_26240);
nor U34484 (N_34484,N_28948,N_25356);
and U34485 (N_34485,N_26100,N_29531);
nor U34486 (N_34486,N_26298,N_27670);
nor U34487 (N_34487,N_27135,N_26193);
nor U34488 (N_34488,N_26849,N_27056);
and U34489 (N_34489,N_26120,N_25700);
or U34490 (N_34490,N_25601,N_27643);
or U34491 (N_34491,N_26679,N_26442);
or U34492 (N_34492,N_29914,N_27531);
nand U34493 (N_34493,N_29526,N_28215);
xor U34494 (N_34494,N_29052,N_28768);
xnor U34495 (N_34495,N_28364,N_26762);
nand U34496 (N_34496,N_25629,N_29775);
nor U34497 (N_34497,N_27868,N_27125);
nand U34498 (N_34498,N_25312,N_25978);
xnor U34499 (N_34499,N_25904,N_26608);
nand U34500 (N_34500,N_25454,N_27862);
or U34501 (N_34501,N_28619,N_27231);
or U34502 (N_34502,N_25412,N_28416);
and U34503 (N_34503,N_25016,N_28064);
or U34504 (N_34504,N_26346,N_28208);
and U34505 (N_34505,N_28994,N_28481);
and U34506 (N_34506,N_28144,N_25314);
and U34507 (N_34507,N_26795,N_26775);
or U34508 (N_34508,N_26530,N_28885);
nand U34509 (N_34509,N_28228,N_28483);
xnor U34510 (N_34510,N_29931,N_27247);
xnor U34511 (N_34511,N_27007,N_26282);
nor U34512 (N_34512,N_25906,N_25444);
nor U34513 (N_34513,N_27810,N_27174);
and U34514 (N_34514,N_26826,N_26809);
or U34515 (N_34515,N_29762,N_26123);
nor U34516 (N_34516,N_25193,N_28968);
nand U34517 (N_34517,N_29073,N_25383);
nor U34518 (N_34518,N_29020,N_25477);
or U34519 (N_34519,N_25602,N_26193);
nand U34520 (N_34520,N_29807,N_26574);
nand U34521 (N_34521,N_26538,N_25253);
and U34522 (N_34522,N_25954,N_25045);
or U34523 (N_34523,N_28770,N_29676);
or U34524 (N_34524,N_27775,N_27218);
and U34525 (N_34525,N_25133,N_27061);
nor U34526 (N_34526,N_27014,N_28445);
nor U34527 (N_34527,N_25785,N_25948);
xor U34528 (N_34528,N_27823,N_29985);
nor U34529 (N_34529,N_29276,N_27496);
and U34530 (N_34530,N_26640,N_26295);
and U34531 (N_34531,N_26351,N_25928);
or U34532 (N_34532,N_27796,N_26851);
or U34533 (N_34533,N_29922,N_29775);
nor U34534 (N_34534,N_26706,N_27576);
or U34535 (N_34535,N_29356,N_27065);
and U34536 (N_34536,N_29592,N_28392);
nand U34537 (N_34537,N_25194,N_27915);
nor U34538 (N_34538,N_27469,N_27535);
xor U34539 (N_34539,N_28015,N_27819);
nor U34540 (N_34540,N_26499,N_28175);
nor U34541 (N_34541,N_28033,N_28481);
or U34542 (N_34542,N_28600,N_26489);
xnor U34543 (N_34543,N_28146,N_27656);
and U34544 (N_34544,N_29810,N_27627);
and U34545 (N_34545,N_29443,N_29924);
and U34546 (N_34546,N_25594,N_29494);
nand U34547 (N_34547,N_27081,N_28279);
nand U34548 (N_34548,N_27113,N_26039);
and U34549 (N_34549,N_29610,N_25404);
or U34550 (N_34550,N_27574,N_28267);
or U34551 (N_34551,N_27144,N_28131);
nand U34552 (N_34552,N_29429,N_26796);
nand U34553 (N_34553,N_27552,N_28310);
nand U34554 (N_34554,N_27812,N_25579);
and U34555 (N_34555,N_27367,N_27959);
nand U34556 (N_34556,N_27340,N_28661);
nor U34557 (N_34557,N_27074,N_26523);
nand U34558 (N_34558,N_25173,N_29829);
xnor U34559 (N_34559,N_28570,N_27564);
nand U34560 (N_34560,N_29283,N_26869);
nand U34561 (N_34561,N_26584,N_27525);
nor U34562 (N_34562,N_25734,N_28054);
and U34563 (N_34563,N_28534,N_27382);
nand U34564 (N_34564,N_25447,N_27279);
and U34565 (N_34565,N_27369,N_25991);
or U34566 (N_34566,N_29738,N_25372);
xor U34567 (N_34567,N_25488,N_29463);
and U34568 (N_34568,N_26161,N_28143);
nor U34569 (N_34569,N_27729,N_28831);
and U34570 (N_34570,N_29017,N_25448);
nand U34571 (N_34571,N_26622,N_25864);
nor U34572 (N_34572,N_26591,N_26840);
and U34573 (N_34573,N_29049,N_28058);
and U34574 (N_34574,N_29933,N_26884);
nand U34575 (N_34575,N_29728,N_26804);
or U34576 (N_34576,N_27447,N_27255);
and U34577 (N_34577,N_29630,N_27122);
xnor U34578 (N_34578,N_28614,N_29942);
and U34579 (N_34579,N_27377,N_25925);
or U34580 (N_34580,N_26586,N_27604);
and U34581 (N_34581,N_26914,N_27714);
xnor U34582 (N_34582,N_27342,N_29980);
nor U34583 (N_34583,N_25342,N_25116);
nor U34584 (N_34584,N_29950,N_27412);
or U34585 (N_34585,N_27354,N_26884);
nor U34586 (N_34586,N_25486,N_28981);
or U34587 (N_34587,N_29121,N_25867);
nand U34588 (N_34588,N_29472,N_29181);
or U34589 (N_34589,N_29887,N_29091);
nor U34590 (N_34590,N_25098,N_27166);
and U34591 (N_34591,N_27318,N_29570);
nand U34592 (N_34592,N_29603,N_29283);
nor U34593 (N_34593,N_27921,N_25451);
nor U34594 (N_34594,N_29236,N_25186);
or U34595 (N_34595,N_29073,N_25672);
xor U34596 (N_34596,N_25882,N_26373);
and U34597 (N_34597,N_27469,N_28868);
or U34598 (N_34598,N_25860,N_29437);
and U34599 (N_34599,N_25195,N_29463);
or U34600 (N_34600,N_25176,N_25196);
nor U34601 (N_34601,N_26692,N_27060);
and U34602 (N_34602,N_28961,N_29669);
and U34603 (N_34603,N_27464,N_28448);
or U34604 (N_34604,N_27315,N_29023);
or U34605 (N_34605,N_27822,N_25128);
and U34606 (N_34606,N_26609,N_25722);
or U34607 (N_34607,N_27901,N_27722);
xor U34608 (N_34608,N_29031,N_25071);
or U34609 (N_34609,N_28165,N_25655);
or U34610 (N_34610,N_25504,N_28759);
and U34611 (N_34611,N_28702,N_27763);
nor U34612 (N_34612,N_29907,N_27503);
and U34613 (N_34613,N_29838,N_28571);
and U34614 (N_34614,N_25154,N_26438);
nand U34615 (N_34615,N_29466,N_27486);
and U34616 (N_34616,N_25228,N_29132);
nor U34617 (N_34617,N_28572,N_25106);
nand U34618 (N_34618,N_25724,N_25846);
or U34619 (N_34619,N_28050,N_26475);
nand U34620 (N_34620,N_26392,N_27796);
and U34621 (N_34621,N_26807,N_27510);
or U34622 (N_34622,N_25494,N_28438);
xor U34623 (N_34623,N_29104,N_26069);
nand U34624 (N_34624,N_27886,N_28457);
and U34625 (N_34625,N_25008,N_27325);
or U34626 (N_34626,N_29443,N_28120);
nor U34627 (N_34627,N_26697,N_25740);
nor U34628 (N_34628,N_26391,N_27656);
or U34629 (N_34629,N_26466,N_25169);
or U34630 (N_34630,N_28290,N_25757);
nor U34631 (N_34631,N_27382,N_28213);
and U34632 (N_34632,N_26430,N_25307);
and U34633 (N_34633,N_26281,N_29076);
nand U34634 (N_34634,N_29881,N_28980);
nor U34635 (N_34635,N_26906,N_29149);
nor U34636 (N_34636,N_26231,N_25406);
nand U34637 (N_34637,N_28454,N_25159);
xnor U34638 (N_34638,N_26538,N_26095);
nor U34639 (N_34639,N_25218,N_27260);
or U34640 (N_34640,N_29236,N_25114);
or U34641 (N_34641,N_28515,N_25987);
nor U34642 (N_34642,N_28580,N_29772);
nor U34643 (N_34643,N_25078,N_28502);
and U34644 (N_34644,N_27137,N_27676);
or U34645 (N_34645,N_27671,N_29735);
nor U34646 (N_34646,N_25327,N_26980);
nand U34647 (N_34647,N_29041,N_28384);
and U34648 (N_34648,N_28363,N_29698);
nand U34649 (N_34649,N_26428,N_29191);
or U34650 (N_34650,N_26874,N_27457);
nor U34651 (N_34651,N_27067,N_25093);
or U34652 (N_34652,N_27063,N_25246);
xor U34653 (N_34653,N_25647,N_25846);
nor U34654 (N_34654,N_28362,N_25219);
or U34655 (N_34655,N_27274,N_28423);
and U34656 (N_34656,N_25435,N_28266);
or U34657 (N_34657,N_26807,N_29002);
xor U34658 (N_34658,N_29967,N_29984);
nand U34659 (N_34659,N_29107,N_27429);
and U34660 (N_34660,N_25244,N_28408);
or U34661 (N_34661,N_25195,N_27511);
and U34662 (N_34662,N_25628,N_29074);
nor U34663 (N_34663,N_25753,N_27924);
nor U34664 (N_34664,N_28132,N_29460);
nand U34665 (N_34665,N_25240,N_26706);
and U34666 (N_34666,N_27119,N_26383);
xor U34667 (N_34667,N_25127,N_27956);
nor U34668 (N_34668,N_27569,N_29177);
or U34669 (N_34669,N_28865,N_27860);
or U34670 (N_34670,N_29093,N_28528);
nor U34671 (N_34671,N_28679,N_28799);
or U34672 (N_34672,N_28149,N_29678);
nor U34673 (N_34673,N_25420,N_25314);
or U34674 (N_34674,N_25648,N_27721);
xor U34675 (N_34675,N_26915,N_29595);
nand U34676 (N_34676,N_27797,N_27166);
nand U34677 (N_34677,N_29931,N_29901);
nand U34678 (N_34678,N_26404,N_28111);
and U34679 (N_34679,N_25019,N_26941);
nand U34680 (N_34680,N_25940,N_26737);
xnor U34681 (N_34681,N_26305,N_25224);
or U34682 (N_34682,N_25878,N_28228);
nand U34683 (N_34683,N_27477,N_26732);
or U34684 (N_34684,N_29457,N_25945);
and U34685 (N_34685,N_25016,N_25924);
nor U34686 (N_34686,N_26791,N_25946);
nand U34687 (N_34687,N_28536,N_27994);
nand U34688 (N_34688,N_26481,N_29009);
nand U34689 (N_34689,N_28439,N_28275);
nand U34690 (N_34690,N_27992,N_27851);
nand U34691 (N_34691,N_29427,N_25538);
nand U34692 (N_34692,N_26340,N_27639);
xnor U34693 (N_34693,N_27649,N_27487);
or U34694 (N_34694,N_28560,N_26502);
nor U34695 (N_34695,N_27889,N_26815);
xnor U34696 (N_34696,N_27487,N_28757);
and U34697 (N_34697,N_27509,N_29851);
xnor U34698 (N_34698,N_25847,N_27115);
nor U34699 (N_34699,N_25658,N_29121);
and U34700 (N_34700,N_25461,N_28205);
and U34701 (N_34701,N_28254,N_25269);
and U34702 (N_34702,N_25142,N_27754);
nand U34703 (N_34703,N_28805,N_26654);
nor U34704 (N_34704,N_29224,N_27230);
nor U34705 (N_34705,N_29493,N_28801);
or U34706 (N_34706,N_26546,N_28083);
or U34707 (N_34707,N_28951,N_25543);
nor U34708 (N_34708,N_28442,N_27856);
nand U34709 (N_34709,N_25429,N_27849);
nor U34710 (N_34710,N_27206,N_25011);
or U34711 (N_34711,N_25696,N_27162);
xor U34712 (N_34712,N_26084,N_28072);
and U34713 (N_34713,N_26334,N_25627);
nand U34714 (N_34714,N_29159,N_27004);
nor U34715 (N_34715,N_25938,N_28904);
or U34716 (N_34716,N_28759,N_28180);
nand U34717 (N_34717,N_28679,N_26348);
nand U34718 (N_34718,N_29859,N_26257);
nand U34719 (N_34719,N_25178,N_26656);
nand U34720 (N_34720,N_26722,N_27878);
nor U34721 (N_34721,N_26422,N_26133);
nand U34722 (N_34722,N_26772,N_29448);
nand U34723 (N_34723,N_27106,N_29156);
or U34724 (N_34724,N_26133,N_26114);
xnor U34725 (N_34725,N_28614,N_27982);
nor U34726 (N_34726,N_27328,N_26050);
xor U34727 (N_34727,N_27594,N_27557);
nand U34728 (N_34728,N_29495,N_25779);
nand U34729 (N_34729,N_25258,N_29151);
and U34730 (N_34730,N_29492,N_27649);
or U34731 (N_34731,N_27170,N_27344);
and U34732 (N_34732,N_27803,N_29759);
nor U34733 (N_34733,N_28860,N_25759);
and U34734 (N_34734,N_26161,N_25470);
and U34735 (N_34735,N_29832,N_28814);
nand U34736 (N_34736,N_29072,N_29593);
nor U34737 (N_34737,N_29429,N_28930);
and U34738 (N_34738,N_26020,N_27895);
or U34739 (N_34739,N_29065,N_29581);
xnor U34740 (N_34740,N_26983,N_27928);
or U34741 (N_34741,N_28622,N_26196);
nand U34742 (N_34742,N_27311,N_26445);
and U34743 (N_34743,N_29958,N_29342);
nand U34744 (N_34744,N_25069,N_26402);
nor U34745 (N_34745,N_29028,N_26969);
or U34746 (N_34746,N_29202,N_27646);
nand U34747 (N_34747,N_26452,N_29837);
or U34748 (N_34748,N_28457,N_25806);
nor U34749 (N_34749,N_27737,N_25958);
or U34750 (N_34750,N_28504,N_26485);
xor U34751 (N_34751,N_27053,N_26101);
nand U34752 (N_34752,N_28314,N_27913);
xnor U34753 (N_34753,N_26968,N_26916);
nor U34754 (N_34754,N_26691,N_27291);
and U34755 (N_34755,N_27722,N_27227);
nor U34756 (N_34756,N_29971,N_27710);
or U34757 (N_34757,N_25321,N_26151);
nor U34758 (N_34758,N_25166,N_25155);
xor U34759 (N_34759,N_29357,N_27220);
nor U34760 (N_34760,N_28790,N_26417);
and U34761 (N_34761,N_29953,N_25977);
or U34762 (N_34762,N_25838,N_25411);
and U34763 (N_34763,N_27651,N_29042);
xnor U34764 (N_34764,N_28991,N_28937);
nand U34765 (N_34765,N_25196,N_28300);
and U34766 (N_34766,N_29328,N_28285);
nor U34767 (N_34767,N_25801,N_28477);
nand U34768 (N_34768,N_28723,N_29589);
and U34769 (N_34769,N_29801,N_28229);
nand U34770 (N_34770,N_28273,N_28846);
or U34771 (N_34771,N_29933,N_28223);
xor U34772 (N_34772,N_27399,N_25957);
nor U34773 (N_34773,N_26591,N_27613);
and U34774 (N_34774,N_29478,N_29855);
and U34775 (N_34775,N_27975,N_27727);
and U34776 (N_34776,N_27268,N_28436);
or U34777 (N_34777,N_27369,N_28521);
or U34778 (N_34778,N_29573,N_25808);
or U34779 (N_34779,N_28475,N_29696);
nand U34780 (N_34780,N_28635,N_29368);
or U34781 (N_34781,N_29215,N_29743);
nor U34782 (N_34782,N_29122,N_27052);
or U34783 (N_34783,N_29433,N_27778);
xor U34784 (N_34784,N_29465,N_26634);
or U34785 (N_34785,N_28956,N_28217);
nor U34786 (N_34786,N_26302,N_27631);
nor U34787 (N_34787,N_26845,N_29211);
nor U34788 (N_34788,N_28305,N_26532);
and U34789 (N_34789,N_26853,N_29292);
and U34790 (N_34790,N_29568,N_25719);
and U34791 (N_34791,N_29081,N_26916);
or U34792 (N_34792,N_28632,N_29669);
xnor U34793 (N_34793,N_25978,N_28447);
nand U34794 (N_34794,N_25089,N_25756);
nand U34795 (N_34795,N_28701,N_29763);
and U34796 (N_34796,N_25192,N_27291);
nand U34797 (N_34797,N_28408,N_28404);
nand U34798 (N_34798,N_27381,N_27412);
and U34799 (N_34799,N_26852,N_29448);
and U34800 (N_34800,N_27323,N_29094);
xnor U34801 (N_34801,N_28381,N_29768);
nand U34802 (N_34802,N_27228,N_28908);
nand U34803 (N_34803,N_27259,N_25104);
nor U34804 (N_34804,N_29196,N_28054);
nand U34805 (N_34805,N_29311,N_27432);
and U34806 (N_34806,N_29216,N_28775);
xnor U34807 (N_34807,N_25758,N_29295);
nand U34808 (N_34808,N_25752,N_26411);
or U34809 (N_34809,N_29648,N_27115);
or U34810 (N_34810,N_28891,N_28892);
nor U34811 (N_34811,N_26346,N_25331);
nand U34812 (N_34812,N_29831,N_29492);
nor U34813 (N_34813,N_27799,N_28874);
and U34814 (N_34814,N_27487,N_29301);
or U34815 (N_34815,N_28398,N_25940);
or U34816 (N_34816,N_25358,N_29416);
and U34817 (N_34817,N_27015,N_29680);
and U34818 (N_34818,N_25240,N_28869);
nor U34819 (N_34819,N_26151,N_27803);
nor U34820 (N_34820,N_27776,N_28580);
and U34821 (N_34821,N_27161,N_27920);
or U34822 (N_34822,N_27700,N_25446);
or U34823 (N_34823,N_29128,N_29809);
nor U34824 (N_34824,N_26318,N_28961);
and U34825 (N_34825,N_26111,N_25934);
nand U34826 (N_34826,N_27145,N_26608);
or U34827 (N_34827,N_29621,N_28310);
or U34828 (N_34828,N_26097,N_28396);
nand U34829 (N_34829,N_26187,N_28504);
and U34830 (N_34830,N_29420,N_28724);
nand U34831 (N_34831,N_25647,N_28909);
and U34832 (N_34832,N_25150,N_27745);
nor U34833 (N_34833,N_27962,N_28297);
xnor U34834 (N_34834,N_28104,N_26423);
or U34835 (N_34835,N_29135,N_27555);
nand U34836 (N_34836,N_27532,N_25429);
nand U34837 (N_34837,N_26085,N_27554);
or U34838 (N_34838,N_25262,N_29093);
or U34839 (N_34839,N_27514,N_29442);
nor U34840 (N_34840,N_26031,N_27815);
nor U34841 (N_34841,N_26138,N_29414);
and U34842 (N_34842,N_27258,N_28080);
or U34843 (N_34843,N_27813,N_26463);
and U34844 (N_34844,N_28167,N_28156);
nand U34845 (N_34845,N_27894,N_25838);
xnor U34846 (N_34846,N_28735,N_29985);
nor U34847 (N_34847,N_26509,N_27401);
nand U34848 (N_34848,N_28761,N_28049);
nor U34849 (N_34849,N_25463,N_25585);
or U34850 (N_34850,N_27051,N_26239);
nand U34851 (N_34851,N_27426,N_28346);
nor U34852 (N_34852,N_28805,N_25399);
nor U34853 (N_34853,N_27614,N_28616);
nor U34854 (N_34854,N_28428,N_27716);
nand U34855 (N_34855,N_25392,N_26433);
or U34856 (N_34856,N_29464,N_28511);
nand U34857 (N_34857,N_27314,N_27732);
or U34858 (N_34858,N_28617,N_29093);
nand U34859 (N_34859,N_25897,N_25329);
nor U34860 (N_34860,N_28532,N_28361);
nor U34861 (N_34861,N_29815,N_28472);
and U34862 (N_34862,N_25270,N_29177);
xnor U34863 (N_34863,N_29128,N_29501);
nand U34864 (N_34864,N_26779,N_26496);
nand U34865 (N_34865,N_28302,N_29063);
nor U34866 (N_34866,N_29870,N_26292);
and U34867 (N_34867,N_26006,N_27740);
xnor U34868 (N_34868,N_28855,N_29647);
and U34869 (N_34869,N_29872,N_29901);
nand U34870 (N_34870,N_29945,N_27991);
and U34871 (N_34871,N_25441,N_27504);
nand U34872 (N_34872,N_27386,N_27950);
and U34873 (N_34873,N_25807,N_26125);
and U34874 (N_34874,N_26495,N_26467);
nor U34875 (N_34875,N_28748,N_26290);
xor U34876 (N_34876,N_25019,N_27766);
nand U34877 (N_34877,N_29407,N_27636);
or U34878 (N_34878,N_25202,N_27223);
nand U34879 (N_34879,N_28830,N_29563);
nand U34880 (N_34880,N_28607,N_27573);
nand U34881 (N_34881,N_27319,N_29169);
nand U34882 (N_34882,N_28312,N_29176);
and U34883 (N_34883,N_28729,N_28942);
nor U34884 (N_34884,N_28903,N_26701);
nand U34885 (N_34885,N_29514,N_28790);
nor U34886 (N_34886,N_26051,N_26254);
and U34887 (N_34887,N_28384,N_27843);
or U34888 (N_34888,N_26599,N_28067);
and U34889 (N_34889,N_29968,N_27038);
or U34890 (N_34890,N_28768,N_26256);
and U34891 (N_34891,N_27383,N_27783);
nor U34892 (N_34892,N_27262,N_27806);
xnor U34893 (N_34893,N_27106,N_26196);
and U34894 (N_34894,N_26166,N_27355);
nor U34895 (N_34895,N_28665,N_26887);
and U34896 (N_34896,N_27203,N_27052);
and U34897 (N_34897,N_25372,N_28892);
nor U34898 (N_34898,N_26089,N_26694);
or U34899 (N_34899,N_27611,N_26507);
nor U34900 (N_34900,N_27933,N_29773);
xor U34901 (N_34901,N_27367,N_25501);
nor U34902 (N_34902,N_28696,N_26613);
or U34903 (N_34903,N_28377,N_27579);
nand U34904 (N_34904,N_26748,N_29213);
nand U34905 (N_34905,N_29088,N_26941);
nor U34906 (N_34906,N_25997,N_27040);
or U34907 (N_34907,N_27178,N_26267);
nand U34908 (N_34908,N_27545,N_28166);
xnor U34909 (N_34909,N_28355,N_29964);
or U34910 (N_34910,N_25818,N_28430);
xor U34911 (N_34911,N_26560,N_27031);
xnor U34912 (N_34912,N_25028,N_26570);
or U34913 (N_34913,N_25291,N_27711);
nand U34914 (N_34914,N_29921,N_25289);
and U34915 (N_34915,N_25654,N_29934);
or U34916 (N_34916,N_26172,N_28445);
or U34917 (N_34917,N_28294,N_27459);
nor U34918 (N_34918,N_29875,N_26714);
nand U34919 (N_34919,N_25125,N_28976);
and U34920 (N_34920,N_26525,N_25314);
or U34921 (N_34921,N_25649,N_26695);
nor U34922 (N_34922,N_27387,N_25361);
and U34923 (N_34923,N_28428,N_28023);
nand U34924 (N_34924,N_25848,N_27904);
nor U34925 (N_34925,N_29718,N_27179);
nor U34926 (N_34926,N_28976,N_28713);
or U34927 (N_34927,N_28250,N_27993);
or U34928 (N_34928,N_29977,N_27601);
nor U34929 (N_34929,N_27521,N_29472);
nor U34930 (N_34930,N_28931,N_26868);
xor U34931 (N_34931,N_25840,N_26464);
or U34932 (N_34932,N_25271,N_27792);
nor U34933 (N_34933,N_29623,N_28399);
and U34934 (N_34934,N_25551,N_27881);
nor U34935 (N_34935,N_26295,N_29926);
or U34936 (N_34936,N_28200,N_29670);
and U34937 (N_34937,N_26762,N_27411);
or U34938 (N_34938,N_29618,N_26140);
or U34939 (N_34939,N_28642,N_26072);
nor U34940 (N_34940,N_29779,N_27386);
and U34941 (N_34941,N_26048,N_25118);
nand U34942 (N_34942,N_27040,N_26850);
nor U34943 (N_34943,N_29446,N_28938);
or U34944 (N_34944,N_27767,N_28608);
xor U34945 (N_34945,N_26192,N_27472);
and U34946 (N_34946,N_25527,N_27742);
and U34947 (N_34947,N_28566,N_25375);
nor U34948 (N_34948,N_25811,N_27166);
and U34949 (N_34949,N_29347,N_26617);
nor U34950 (N_34950,N_29251,N_27559);
nor U34951 (N_34951,N_26156,N_29124);
nor U34952 (N_34952,N_26695,N_28902);
xor U34953 (N_34953,N_27854,N_27262);
nand U34954 (N_34954,N_25923,N_28750);
or U34955 (N_34955,N_25580,N_28809);
and U34956 (N_34956,N_26611,N_29965);
or U34957 (N_34957,N_29296,N_27246);
nor U34958 (N_34958,N_26820,N_29438);
nand U34959 (N_34959,N_27703,N_28660);
and U34960 (N_34960,N_29324,N_28745);
and U34961 (N_34961,N_27080,N_25275);
nor U34962 (N_34962,N_29699,N_25974);
nor U34963 (N_34963,N_25098,N_28009);
nor U34964 (N_34964,N_25772,N_25481);
and U34965 (N_34965,N_27160,N_29042);
nand U34966 (N_34966,N_28877,N_27891);
nor U34967 (N_34967,N_26929,N_26540);
or U34968 (N_34968,N_26830,N_26791);
and U34969 (N_34969,N_26585,N_28187);
nor U34970 (N_34970,N_26538,N_25827);
nor U34971 (N_34971,N_28884,N_29793);
and U34972 (N_34972,N_26775,N_25797);
or U34973 (N_34973,N_28139,N_29818);
nand U34974 (N_34974,N_29387,N_29781);
nand U34975 (N_34975,N_28129,N_27685);
or U34976 (N_34976,N_28949,N_25242);
nor U34977 (N_34977,N_28323,N_28919);
and U34978 (N_34978,N_29844,N_27256);
nand U34979 (N_34979,N_27301,N_28279);
and U34980 (N_34980,N_25246,N_26532);
or U34981 (N_34981,N_25697,N_27233);
or U34982 (N_34982,N_29931,N_28498);
nor U34983 (N_34983,N_29195,N_29737);
nor U34984 (N_34984,N_25604,N_26124);
and U34985 (N_34985,N_27643,N_25771);
nor U34986 (N_34986,N_27615,N_25583);
or U34987 (N_34987,N_28661,N_27125);
nand U34988 (N_34988,N_28907,N_25557);
nand U34989 (N_34989,N_27789,N_29314);
or U34990 (N_34990,N_25037,N_25092);
or U34991 (N_34991,N_29543,N_29711);
or U34992 (N_34992,N_27875,N_25664);
nor U34993 (N_34993,N_26929,N_25030);
nand U34994 (N_34994,N_25968,N_26228);
nor U34995 (N_34995,N_29232,N_27263);
or U34996 (N_34996,N_26286,N_27775);
and U34997 (N_34997,N_29543,N_26959);
and U34998 (N_34998,N_28353,N_27429);
nor U34999 (N_34999,N_27848,N_29451);
xor U35000 (N_35000,N_33267,N_31904);
nand U35001 (N_35001,N_30792,N_33025);
or U35002 (N_35002,N_32031,N_30323);
nand U35003 (N_35003,N_34037,N_31032);
and U35004 (N_35004,N_34072,N_34721);
or U35005 (N_35005,N_30953,N_34320);
and U35006 (N_35006,N_31274,N_31792);
and U35007 (N_35007,N_30506,N_32619);
nand U35008 (N_35008,N_33389,N_34515);
xnor U35009 (N_35009,N_30771,N_33910);
and U35010 (N_35010,N_33824,N_30108);
nand U35011 (N_35011,N_34796,N_30615);
nand U35012 (N_35012,N_30082,N_32608);
nand U35013 (N_35013,N_34305,N_34651);
or U35014 (N_35014,N_34707,N_32664);
or U35015 (N_35015,N_32679,N_30408);
nor U35016 (N_35016,N_34917,N_32676);
nand U35017 (N_35017,N_31950,N_30701);
nor U35018 (N_35018,N_33643,N_34311);
xor U35019 (N_35019,N_33754,N_33807);
nor U35020 (N_35020,N_34230,N_31307);
nor U35021 (N_35021,N_33164,N_31087);
or U35022 (N_35022,N_34246,N_33054);
nand U35023 (N_35023,N_32897,N_33001);
and U35024 (N_35024,N_34384,N_32372);
nor U35025 (N_35025,N_33798,N_30420);
and U35026 (N_35026,N_31101,N_34885);
nor U35027 (N_35027,N_32161,N_31786);
and U35028 (N_35028,N_33848,N_33293);
or U35029 (N_35029,N_32121,N_33426);
and U35030 (N_35030,N_33612,N_33773);
xor U35031 (N_35031,N_32934,N_30929);
nand U35032 (N_35032,N_32385,N_30919);
nor U35033 (N_35033,N_32929,N_31612);
nor U35034 (N_35034,N_33526,N_33353);
or U35035 (N_35035,N_34097,N_34465);
or U35036 (N_35036,N_33682,N_31934);
and U35037 (N_35037,N_30072,N_31668);
and U35038 (N_35038,N_33912,N_32413);
nor U35039 (N_35039,N_31316,N_31319);
nand U35040 (N_35040,N_30634,N_31893);
or U35041 (N_35041,N_33181,N_32744);
or U35042 (N_35042,N_30227,N_30350);
or U35043 (N_35043,N_31938,N_30503);
or U35044 (N_35044,N_31590,N_32133);
and U35045 (N_35045,N_32292,N_34418);
or U35046 (N_35046,N_34929,N_31839);
xor U35047 (N_35047,N_31824,N_33958);
nand U35048 (N_35048,N_31991,N_33387);
nor U35049 (N_35049,N_31091,N_31565);
nor U35050 (N_35050,N_31752,N_30572);
or U35051 (N_35051,N_30830,N_30294);
and U35052 (N_35052,N_33925,N_32347);
and U35053 (N_35053,N_34074,N_30641);
nand U35054 (N_35054,N_33457,N_34837);
or U35055 (N_35055,N_30902,N_34294);
nand U35056 (N_35056,N_34836,N_34626);
nor U35057 (N_35057,N_30221,N_33927);
nor U35058 (N_35058,N_32730,N_34889);
and U35059 (N_35059,N_31369,N_34611);
nand U35060 (N_35060,N_34233,N_34965);
nor U35061 (N_35061,N_30692,N_32505);
and U35062 (N_35062,N_31981,N_30988);
nand U35063 (N_35063,N_34582,N_32850);
nand U35064 (N_35064,N_32531,N_31331);
and U35065 (N_35065,N_33407,N_33760);
xor U35066 (N_35066,N_31190,N_33627);
nor U35067 (N_35067,N_31017,N_31096);
and U35068 (N_35068,N_32311,N_30728);
or U35069 (N_35069,N_32200,N_33514);
xnor U35070 (N_35070,N_30275,N_33364);
nand U35071 (N_35071,N_30022,N_31621);
or U35072 (N_35072,N_30473,N_33215);
and U35073 (N_35073,N_31700,N_30693);
and U35074 (N_35074,N_31855,N_31488);
nand U35075 (N_35075,N_31348,N_30242);
nand U35076 (N_35076,N_30786,N_33665);
xor U35077 (N_35077,N_30265,N_31215);
nand U35078 (N_35078,N_33883,N_30211);
or U35079 (N_35079,N_33314,N_32651);
and U35080 (N_35080,N_32454,N_33484);
nand U35081 (N_35081,N_33712,N_33330);
and U35082 (N_35082,N_33495,N_32891);
and U35083 (N_35083,N_34143,N_30984);
nor U35084 (N_35084,N_33413,N_32403);
or U35085 (N_35085,N_31601,N_33605);
nand U35086 (N_35086,N_33108,N_31733);
xor U35087 (N_35087,N_33995,N_31437);
xnor U35088 (N_35088,N_31715,N_34194);
nor U35089 (N_35089,N_34962,N_32696);
and U35090 (N_35090,N_30854,N_32177);
and U35091 (N_35091,N_32665,N_32969);
nor U35092 (N_35092,N_34124,N_30811);
nor U35093 (N_35093,N_32108,N_34270);
nand U35094 (N_35094,N_33060,N_30458);
nand U35095 (N_35095,N_32958,N_34617);
nor U35096 (N_35096,N_33897,N_31294);
or U35097 (N_35097,N_33736,N_32309);
nand U35098 (N_35098,N_34785,N_30038);
xor U35099 (N_35099,N_31254,N_33171);
and U35100 (N_35100,N_31907,N_34927);
nand U35101 (N_35101,N_33519,N_32760);
nor U35102 (N_35102,N_31647,N_32642);
or U35103 (N_35103,N_33951,N_33621);
and U35104 (N_35104,N_34653,N_33151);
and U35105 (N_35105,N_31238,N_30455);
nor U35106 (N_35106,N_31526,N_33147);
or U35107 (N_35107,N_30307,N_33074);
and U35108 (N_35108,N_33355,N_33078);
xnor U35109 (N_35109,N_30036,N_31471);
and U35110 (N_35110,N_34736,N_32545);
and U35111 (N_35111,N_34869,N_31035);
nor U35112 (N_35112,N_34844,N_33812);
and U35113 (N_35113,N_30710,N_33220);
and U35114 (N_35114,N_32089,N_31843);
or U35115 (N_35115,N_34379,N_32908);
and U35116 (N_35116,N_31756,N_33296);
xnor U35117 (N_35117,N_34047,N_31131);
and U35118 (N_35118,N_34782,N_31969);
nand U35119 (N_35119,N_31246,N_30126);
xor U35120 (N_35120,N_32553,N_34870);
nor U35121 (N_35121,N_31566,N_34952);
nand U35122 (N_35122,N_33663,N_30181);
or U35123 (N_35123,N_31518,N_32128);
nand U35124 (N_35124,N_34671,N_34549);
or U35125 (N_35125,N_31684,N_30763);
and U35126 (N_35126,N_33004,N_33163);
xor U35127 (N_35127,N_31745,N_30869);
xor U35128 (N_35128,N_33709,N_33844);
nor U35129 (N_35129,N_32020,N_31941);
or U35130 (N_35130,N_34352,N_34073);
and U35131 (N_35131,N_32497,N_31311);
xor U35132 (N_35132,N_31944,N_30065);
or U35133 (N_35133,N_32291,N_32228);
and U35134 (N_35134,N_34968,N_30399);
nor U35135 (N_35135,N_32455,N_33072);
nand U35136 (N_35136,N_30421,N_32968);
nor U35137 (N_35137,N_30633,N_31758);
and U35138 (N_35138,N_33962,N_31722);
nor U35139 (N_35139,N_32517,N_32254);
nor U35140 (N_35140,N_34601,N_30248);
nand U35141 (N_35141,N_31396,N_33036);
or U35142 (N_35142,N_34413,N_32075);
or U35143 (N_35143,N_33153,N_32667);
nor U35144 (N_35144,N_31270,N_34499);
or U35145 (N_35145,N_32150,N_30303);
nand U35146 (N_35146,N_33752,N_32209);
nor U35147 (N_35147,N_31485,N_31736);
and U35148 (N_35148,N_32337,N_30779);
and U35149 (N_35149,N_30379,N_33565);
or U35150 (N_35150,N_32600,N_30289);
or U35151 (N_35151,N_33056,N_32474);
nor U35152 (N_35152,N_32388,N_32876);
nand U35153 (N_35153,N_30435,N_33188);
or U35154 (N_35154,N_33370,N_30066);
or U35155 (N_35155,N_31321,N_34300);
nor U35156 (N_35156,N_34242,N_32016);
and U35157 (N_35157,N_32123,N_34309);
and U35158 (N_35158,N_34620,N_34477);
or U35159 (N_35159,N_33698,N_34361);
or U35160 (N_35160,N_31070,N_31025);
nand U35161 (N_35161,N_34659,N_30921);
and U35162 (N_35162,N_31961,N_34062);
nand U35163 (N_35163,N_30247,N_33801);
or U35164 (N_35164,N_34520,N_34524);
and U35165 (N_35165,N_32858,N_30497);
xor U35166 (N_35166,N_34825,N_33743);
or U35167 (N_35167,N_30551,N_32794);
xnor U35168 (N_35168,N_32831,N_32686);
or U35169 (N_35169,N_31018,N_31469);
nor U35170 (N_35170,N_31408,N_32728);
nor U35171 (N_35171,N_34119,N_31995);
and U35172 (N_35172,N_31155,N_34888);
and U35173 (N_35173,N_34328,N_33491);
or U35174 (N_35174,N_31492,N_31891);
and U35175 (N_35175,N_34541,N_31126);
nor U35176 (N_35176,N_31506,N_31209);
and U35177 (N_35177,N_34843,N_33249);
or U35178 (N_35178,N_33438,N_32045);
nor U35179 (N_35179,N_30286,N_31329);
nor U35180 (N_35180,N_30282,N_34264);
nor U35181 (N_35181,N_32591,N_34356);
nand U35182 (N_35182,N_34061,N_34387);
nand U35183 (N_35183,N_30164,N_33795);
or U35184 (N_35184,N_34807,N_32606);
nor U35185 (N_35185,N_34219,N_33977);
nor U35186 (N_35186,N_33536,N_32350);
or U35187 (N_35187,N_32453,N_32787);
nor U35188 (N_35188,N_30196,N_33862);
and U35189 (N_35189,N_30872,N_30552);
nand U35190 (N_35190,N_31418,N_33778);
and U35191 (N_35191,N_32614,N_33434);
or U35192 (N_35192,N_34934,N_33369);
or U35193 (N_35193,N_30907,N_34731);
nor U35194 (N_35194,N_30646,N_30269);
and U35195 (N_35195,N_32539,N_30782);
xnor U35196 (N_35196,N_34853,N_33646);
or U35197 (N_35197,N_30881,N_31704);
xnor U35198 (N_35198,N_31744,N_33750);
nor U35199 (N_35199,N_33919,N_30474);
or U35200 (N_35200,N_30115,N_30146);
and U35201 (N_35201,N_34067,N_34148);
nor U35202 (N_35202,N_32776,N_34471);
nor U35203 (N_35203,N_32759,N_30610);
or U35204 (N_35204,N_30833,N_34110);
xor U35205 (N_35205,N_32640,N_33562);
nor U35206 (N_35206,N_32697,N_34406);
xor U35207 (N_35207,N_31439,N_30536);
nand U35208 (N_35208,N_31218,N_31364);
or U35209 (N_35209,N_31800,N_31508);
nor U35210 (N_35210,N_32765,N_32285);
and U35211 (N_35211,N_30026,N_33437);
and U35212 (N_35212,N_31498,N_32513);
nand U35213 (N_35213,N_34021,N_33974);
and U35214 (N_35214,N_33990,N_32083);
and U35215 (N_35215,N_33606,N_34318);
and U35216 (N_35216,N_33602,N_30824);
nor U35217 (N_35217,N_34377,N_33041);
or U35218 (N_35218,N_32426,N_32241);
and U35219 (N_35219,N_34269,N_33430);
and U35220 (N_35220,N_31873,N_32305);
or U35221 (N_35221,N_31521,N_33936);
and U35222 (N_35222,N_32992,N_34569);
nor U35223 (N_35223,N_30570,N_31985);
or U35224 (N_35224,N_30481,N_32826);
or U35225 (N_35225,N_34289,N_30186);
nor U35226 (N_35226,N_30228,N_32297);
nor U35227 (N_35227,N_31347,N_31415);
nand U35228 (N_35228,N_33961,N_30918);
nand U35229 (N_35229,N_30237,N_31936);
nand U35230 (N_35230,N_30512,N_32470);
and U35231 (N_35231,N_31504,N_33303);
nor U35232 (N_35232,N_34660,N_30301);
and U35233 (N_35233,N_33989,N_34223);
nor U35234 (N_35234,N_34057,N_31421);
and U35235 (N_35235,N_33329,N_33265);
nand U35236 (N_35236,N_30487,N_30057);
and U35237 (N_35237,N_30808,N_30518);
and U35238 (N_35238,N_30417,N_34459);
nand U35239 (N_35239,N_33386,N_31996);
and U35240 (N_35240,N_30983,N_34804);
and U35241 (N_35241,N_31987,N_30719);
nor U35242 (N_35242,N_30324,N_30097);
nor U35243 (N_35243,N_32152,N_32562);
or U35244 (N_35244,N_32515,N_30740);
nand U35245 (N_35245,N_30171,N_33288);
nor U35246 (N_35246,N_32536,N_32047);
or U35247 (N_35247,N_32360,N_31925);
nor U35248 (N_35248,N_31856,N_31646);
and U35249 (N_35249,N_30908,N_34226);
nand U35250 (N_35250,N_31636,N_30510);
and U35251 (N_35251,N_33779,N_31496);
or U35252 (N_35252,N_34537,N_30114);
and U35253 (N_35253,N_30790,N_31284);
xnor U35254 (N_35254,N_31906,N_34069);
or U35255 (N_35255,N_30606,N_33931);
nor U35256 (N_35256,N_33318,N_33367);
or U35257 (N_35257,N_31681,N_31105);
or U35258 (N_35258,N_34429,N_34939);
nand U35259 (N_35259,N_33639,N_33493);
and U35260 (N_35260,N_33737,N_30046);
or U35261 (N_35261,N_34603,N_33679);
or U35262 (N_35262,N_34724,N_32986);
nor U35263 (N_35263,N_32756,N_34393);
nand U35264 (N_35264,N_30488,N_34370);
nand U35265 (N_35265,N_33228,N_31483);
and U35266 (N_35266,N_33906,N_30004);
and U35267 (N_35267,N_30280,N_32815);
nand U35268 (N_35268,N_31477,N_30681);
nand U35269 (N_35269,N_32954,N_31540);
nor U35270 (N_35270,N_30684,N_34200);
nand U35271 (N_35271,N_30622,N_33282);
nor U35272 (N_35272,N_30911,N_33687);
nand U35273 (N_35273,N_34894,N_32140);
or U35274 (N_35274,N_32709,N_30575);
or U35275 (N_35275,N_34241,N_32037);
nand U35276 (N_35276,N_34507,N_31200);
and U35277 (N_35277,N_32137,N_33494);
nand U35278 (N_35278,N_34977,N_32871);
or U35279 (N_35279,N_31472,N_33622);
and U35280 (N_35280,N_30637,N_32859);
and U35281 (N_35281,N_31179,N_34616);
nand U35282 (N_35282,N_32516,N_30620);
or U35283 (N_35283,N_33062,N_30434);
and U35284 (N_35284,N_33258,N_30699);
nor U35285 (N_35285,N_30479,N_34262);
nor U35286 (N_35286,N_32499,N_30729);
nand U35287 (N_35287,N_30224,N_30652);
nor U35288 (N_35288,N_31291,N_32861);
and U35289 (N_35289,N_32567,N_34704);
nor U35290 (N_35290,N_30745,N_31788);
or U35291 (N_35291,N_34739,N_33653);
xor U35292 (N_35292,N_33816,N_33098);
nor U35293 (N_35293,N_31805,N_31862);
nand U35294 (N_35294,N_31427,N_33713);
or U35295 (N_35295,N_31253,N_31196);
nand U35296 (N_35296,N_31442,N_34763);
nor U35297 (N_35297,N_34364,N_33261);
or U35298 (N_35298,N_30849,N_32912);
nor U35299 (N_35299,N_31440,N_33205);
and U35300 (N_35300,N_33269,N_32713);
xnor U35301 (N_35301,N_31860,N_34841);
nor U35302 (N_35302,N_30631,N_33866);
nand U35303 (N_35303,N_31631,N_30314);
or U35304 (N_35304,N_34938,N_34316);
nor U35305 (N_35305,N_30347,N_33811);
or U35306 (N_35306,N_34277,N_33231);
xor U35307 (N_35307,N_30217,N_31964);
or U35308 (N_35308,N_31114,N_32789);
and U35309 (N_35309,N_33143,N_33738);
and U35310 (N_35310,N_30612,N_33049);
or U35311 (N_35311,N_32232,N_32535);
and U35312 (N_35312,N_34622,N_31702);
or U35313 (N_35313,N_32638,N_32077);
nand U35314 (N_35314,N_30850,N_30353);
and U35315 (N_35315,N_33826,N_34455);
and U35316 (N_35316,N_32288,N_31771);
nor U35317 (N_35317,N_31512,N_31072);
and U35318 (N_35318,N_31108,N_33131);
or U35319 (N_35319,N_33260,N_34470);
nand U35320 (N_35320,N_32508,N_32219);
nand U35321 (N_35321,N_31455,N_32593);
and U35322 (N_35322,N_30851,N_33822);
nand U35323 (N_35323,N_32503,N_33206);
nor U35324 (N_35324,N_30152,N_33864);
or U35325 (N_35325,N_34913,N_31341);
nand U35326 (N_35326,N_33214,N_33075);
or U35327 (N_35327,N_32715,N_32702);
and U35328 (N_35328,N_30187,N_34845);
nor U35329 (N_35329,N_34243,N_32964);
or U35330 (N_35330,N_30590,N_30376);
and U35331 (N_35331,N_34967,N_33462);
xor U35332 (N_35332,N_33630,N_34166);
xnor U35333 (N_35333,N_32468,N_34907);
and U35334 (N_35334,N_34991,N_32883);
and U35335 (N_35335,N_32893,N_32681);
nor U35336 (N_35336,N_33672,N_33292);
nor U35337 (N_35337,N_32376,N_34754);
nor U35338 (N_35338,N_34390,N_32084);
nor U35339 (N_35339,N_33574,N_32420);
nand U35340 (N_35340,N_32576,N_31664);
nand U35341 (N_35341,N_34041,N_31393);
nand U35342 (N_35342,N_34705,N_31001);
nor U35343 (N_35343,N_31153,N_32641);
nand U35344 (N_35344,N_31659,N_34564);
nand U35345 (N_35345,N_34697,N_30039);
nor U35346 (N_35346,N_30493,N_32362);
nor U35347 (N_35347,N_33478,N_31333);
and U35348 (N_35348,N_30844,N_33327);
nand U35349 (N_35349,N_34102,N_32646);
nor U35350 (N_35350,N_34481,N_30125);
and U35351 (N_35351,N_33944,N_33764);
and U35352 (N_35352,N_34127,N_32845);
xor U35353 (N_35353,N_32913,N_33673);
or U35354 (N_35354,N_30313,N_30653);
and U35355 (N_35355,N_34497,N_31557);
and U35356 (N_35356,N_33928,N_34798);
nor U35357 (N_35357,N_33831,N_31342);
nand U35358 (N_35358,N_34975,N_33103);
nor U35359 (N_35359,N_30985,N_34900);
nor U35360 (N_35360,N_30885,N_33090);
or U35361 (N_35361,N_30132,N_34107);
or U35362 (N_35362,N_30522,N_32189);
and U35363 (N_35363,N_30501,N_33800);
or U35364 (N_35364,N_30962,N_33290);
or U35365 (N_35365,N_33027,N_30414);
nand U35366 (N_35366,N_32999,N_30588);
nand U35367 (N_35367,N_31021,N_32684);
xnor U35368 (N_35368,N_30975,N_33092);
and U35369 (N_35369,N_33112,N_31394);
and U35370 (N_35370,N_32587,N_32119);
and U35371 (N_35371,N_34872,N_31561);
or U35372 (N_35372,N_31592,N_32415);
nor U35373 (N_35373,N_32381,N_33350);
and U35374 (N_35374,N_30776,N_32449);
nor U35375 (N_35375,N_32772,N_32923);
nand U35376 (N_35376,N_33842,N_33654);
nor U35377 (N_35377,N_30725,N_31619);
nand U35378 (N_35378,N_30624,N_32570);
nand U35379 (N_35379,N_32579,N_30793);
or U35380 (N_35380,N_30024,N_30268);
and U35381 (N_35381,N_32452,N_33408);
nand U35382 (N_35382,N_33308,N_32537);
nor U35383 (N_35383,N_30932,N_34452);
or U35384 (N_35384,N_32844,N_33200);
or U35385 (N_35385,N_34522,N_33182);
nor U35386 (N_35386,N_34024,N_33028);
or U35387 (N_35387,N_31336,N_32936);
xor U35388 (N_35388,N_32563,N_34442);
and U35389 (N_35389,N_32661,N_33130);
nor U35390 (N_35390,N_32314,N_33052);
and U35391 (N_35391,N_30753,N_34932);
or U35392 (N_35392,N_33344,N_32690);
nand U35393 (N_35393,N_33575,N_32252);
nand U35394 (N_35394,N_31059,N_33813);
nand U35395 (N_35395,N_34883,N_32012);
nand U35396 (N_35396,N_33730,N_33359);
xnor U35397 (N_35397,N_30581,N_31167);
or U35398 (N_35398,N_33005,N_34279);
nor U35399 (N_35399,N_31337,N_31379);
or U35400 (N_35400,N_34528,N_30466);
and U35401 (N_35401,N_34086,N_34420);
nor U35402 (N_35402,N_33357,N_31470);
nand U35403 (N_35403,N_33063,N_30917);
and U35404 (N_35404,N_31199,N_30069);
and U35405 (N_35405,N_32321,N_31711);
xor U35406 (N_35406,N_31147,N_30866);
nand U35407 (N_35407,N_34084,N_32157);
xor U35408 (N_35408,N_30156,N_31320);
nor U35409 (N_35409,N_34447,N_30337);
nand U35410 (N_35410,N_34985,N_34192);
nor U35411 (N_35411,N_32941,N_33416);
xor U35412 (N_35412,N_31334,N_30320);
nor U35413 (N_35413,N_32990,N_31881);
nor U35414 (N_35414,N_31391,N_30863);
xnor U35415 (N_35415,N_32026,N_32338);
nand U35416 (N_35416,N_31064,N_31271);
or U35417 (N_35417,N_30386,N_32771);
xor U35418 (N_35418,N_31958,N_34218);
nor U35419 (N_35419,N_31529,N_34039);
or U35420 (N_35420,N_31296,N_32530);
nand U35421 (N_35421,N_32906,N_34635);
nand U35422 (N_35422,N_33058,N_34983);
and U35423 (N_35423,N_30101,N_30560);
nor U35424 (N_35424,N_31276,N_30475);
xnor U35425 (N_35425,N_31494,N_34656);
nor U35426 (N_35426,N_33414,N_32983);
nand U35427 (N_35427,N_32168,N_30516);
nand U35428 (N_35428,N_31088,N_30179);
or U35429 (N_35429,N_32721,N_32129);
or U35430 (N_35430,N_31830,N_31380);
nor U35431 (N_35431,N_32754,N_31520);
nand U35432 (N_35432,N_31546,N_31292);
nor U35433 (N_35433,N_32096,N_32618);
nor U35434 (N_35434,N_31463,N_33032);
and U35435 (N_35435,N_33235,N_33262);
nor U35436 (N_35436,N_31008,N_32616);
or U35437 (N_35437,N_33583,N_34164);
and U35438 (N_35438,N_32926,N_33875);
nor U35439 (N_35439,N_34467,N_34299);
nand U35440 (N_35440,N_31986,N_33920);
and U35441 (N_35441,N_34347,N_30713);
or U35442 (N_35442,N_33594,N_31825);
or U35443 (N_35443,N_33867,N_30822);
nand U35444 (N_35444,N_33655,N_30812);
nor U35445 (N_35445,N_32821,N_31970);
nand U35446 (N_35446,N_33502,N_34901);
and U35447 (N_35447,N_34899,N_32743);
and U35448 (N_35448,N_32708,N_31759);
nor U35449 (N_35449,N_33008,N_32741);
and U35450 (N_35450,N_32577,N_34823);
nand U35451 (N_35451,N_31029,N_34634);
nand U35452 (N_35452,N_30766,N_30075);
or U35453 (N_35453,N_30029,N_33211);
nor U35454 (N_35454,N_33899,N_34065);
nor U35455 (N_35455,N_31648,N_34648);
nand U35456 (N_35456,N_32827,N_31544);
and U35457 (N_35457,N_32528,N_32175);
xnor U35458 (N_35458,N_30138,N_34698);
or U35459 (N_35459,N_32431,N_33134);
nor U35460 (N_35460,N_31791,N_33194);
and U35461 (N_35461,N_34990,N_30912);
and U35462 (N_35462,N_32610,N_34291);
or U35463 (N_35463,N_30051,N_30131);
and U35464 (N_35464,N_32746,N_33320);
nand U35465 (N_35465,N_30044,N_33497);
or U35466 (N_35466,N_31318,N_30019);
or U35467 (N_35467,N_32590,N_33395);
nand U35468 (N_35468,N_30914,N_32205);
nand U35469 (N_35469,N_30695,N_30768);
nand U35470 (N_35470,N_34593,N_32120);
and U35471 (N_35471,N_33588,N_30220);
nand U35472 (N_35472,N_31921,N_32764);
or U35473 (N_35473,N_33522,N_30616);
nor U35474 (N_35474,N_31890,N_30368);
nand U35475 (N_35475,N_31812,N_31446);
or U35476 (N_35476,N_32199,N_31589);
nor U35477 (N_35477,N_30299,N_32341);
or U35478 (N_35478,N_34592,N_33294);
nor U35479 (N_35479,N_34994,N_34020);
xor U35480 (N_35480,N_33446,N_31650);
nand U35481 (N_35481,N_34474,N_34822);
nand U35482 (N_35482,N_31766,N_31849);
and U35483 (N_35483,N_31845,N_34397);
or U35484 (N_35484,N_30548,N_33037);
nand U35485 (N_35485,N_34163,N_33139);
and U35486 (N_35486,N_33718,N_32597);
and U35487 (N_35487,N_32324,N_32330);
and U35488 (N_35488,N_31283,N_30859);
nand U35489 (N_35489,N_32411,N_32304);
nand U35490 (N_35490,N_31382,N_33374);
and U35491 (N_35491,N_32255,N_30883);
xnor U35492 (N_35492,N_30091,N_31116);
and U35493 (N_35493,N_34700,N_30149);
xor U35494 (N_35494,N_34147,N_32757);
xor U35495 (N_35495,N_34898,N_31997);
xnor U35496 (N_35496,N_33635,N_33666);
nor U35497 (N_35497,N_34896,N_33585);
or U35498 (N_35498,N_32186,N_33753);
and U35499 (N_35499,N_33162,N_32498);
and U35500 (N_35500,N_31273,N_33530);
xnor U35501 (N_35501,N_34684,N_32215);
nand U35502 (N_35502,N_31407,N_34123);
nand U35503 (N_35503,N_31086,N_31490);
nand U35504 (N_35504,N_31607,N_32048);
and U35505 (N_35505,N_34551,N_31878);
and U35506 (N_35506,N_32176,N_34773);
and U35507 (N_35507,N_30317,N_30950);
nor U35508 (N_35508,N_31136,N_33084);
xor U35509 (N_35509,N_34966,N_30216);
or U35510 (N_35510,N_31339,N_34574);
nand U35511 (N_35511,N_30553,N_34909);
nand U35512 (N_35512,N_32406,N_32910);
xnor U35513 (N_35513,N_30671,N_33420);
nand U35514 (N_35514,N_34742,N_32072);
nand U35515 (N_35515,N_33378,N_31499);
and U35516 (N_35516,N_34842,N_34175);
or U35517 (N_35517,N_34193,N_33399);
nor U35518 (N_35518,N_30165,N_33289);
or U35519 (N_35519,N_31553,N_34605);
and U35520 (N_35520,N_32359,N_33007);
or U35521 (N_35521,N_32617,N_31489);
nand U35522 (N_35522,N_30327,N_32272);
nor U35523 (N_35523,N_31265,N_33264);
and U35524 (N_35524,N_30549,N_34645);
or U35525 (N_35525,N_30331,N_34469);
nand U35526 (N_35526,N_31068,N_30702);
nand U35527 (N_35527,N_31482,N_33109);
or U35528 (N_35528,N_30439,N_33472);
nand U35529 (N_35529,N_31295,N_33129);
nand U35530 (N_35530,N_34920,N_33154);
xnor U35531 (N_35531,N_34411,N_31783);
xor U35532 (N_35532,N_30965,N_31627);
nand U35533 (N_35533,N_31836,N_33298);
xnor U35534 (N_35534,N_31450,N_30129);
xor U35535 (N_35535,N_33706,N_32933);
or U35536 (N_35536,N_32685,N_32817);
nor U35537 (N_35537,N_32416,N_32706);
nand U35538 (N_35538,N_30948,N_31010);
and U35539 (N_35539,N_31299,N_32339);
nor U35540 (N_35540,N_31063,N_32396);
or U35541 (N_35541,N_31887,N_30613);
or U35542 (N_35542,N_33617,N_34797);
nor U35543 (N_35543,N_33216,N_32391);
xnor U35544 (N_35544,N_30712,N_31898);
nand U35545 (N_35545,N_31831,N_30055);
nand U35546 (N_35546,N_31288,N_34871);
nor U35547 (N_35547,N_31678,N_32125);
or U35548 (N_35548,N_33785,N_34506);
or U35549 (N_35549,N_33696,N_32509);
nor U35550 (N_35550,N_32393,N_32962);
and U35551 (N_35551,N_34235,N_31360);
or U35552 (N_35552,N_34744,N_31661);
xor U35553 (N_35553,N_32250,N_32568);
xnor U35554 (N_35554,N_34012,N_30400);
nand U35555 (N_35555,N_30178,N_33968);
nand U35556 (N_35556,N_33365,N_31539);
and U35557 (N_35557,N_34500,N_34591);
and U35558 (N_35558,N_30843,N_31857);
nor U35559 (N_35559,N_32107,N_30901);
or U35560 (N_35560,N_30664,N_34771);
xnor U35561 (N_35561,N_33034,N_32966);
nor U35562 (N_35562,N_33721,N_30159);
nor U35563 (N_35563,N_33015,N_31356);
or U35564 (N_35564,N_30489,N_31819);
nand U35565 (N_35565,N_34234,N_30047);
and U35566 (N_35566,N_32780,N_32633);
or U35567 (N_35567,N_33383,N_32830);
nand U35568 (N_35568,N_34115,N_31901);
nand U35569 (N_35569,N_32162,N_31312);
or U35570 (N_35570,N_34979,N_34006);
and U35571 (N_35571,N_33933,N_32081);
and U35572 (N_35572,N_30173,N_33723);
and U35573 (N_35573,N_33513,N_30764);
nor U35574 (N_35574,N_30384,N_30166);
and U35575 (N_35575,N_34863,N_30875);
nand U35576 (N_35576,N_32087,N_30504);
or U35577 (N_35577,N_31864,N_34876);
nor U35578 (N_35578,N_31868,N_33343);
nand U35579 (N_35579,N_30690,N_31576);
or U35580 (N_35580,N_30926,N_33789);
and U35581 (N_35581,N_34516,N_33337);
or U35582 (N_35582,N_33805,N_33498);
nand U35583 (N_35583,N_31110,N_33879);
nand U35584 (N_35584,N_32445,N_33548);
xor U35585 (N_35585,N_32857,N_33878);
or U35586 (N_35586,N_31642,N_31412);
nor U35587 (N_35587,N_34441,N_34079);
nor U35588 (N_35588,N_32058,N_34414);
and U35589 (N_35589,N_31840,N_30405);
nand U35590 (N_35590,N_32972,N_33043);
nand U35591 (N_35591,N_33031,N_33448);
or U35592 (N_35592,N_32496,N_32011);
or U35593 (N_35593,N_32507,N_32626);
or U35594 (N_35594,N_31821,N_30060);
nand U35595 (N_35595,N_30201,N_31575);
or U35596 (N_35596,N_33984,N_30632);
and U35597 (N_35597,N_31537,N_32578);
and U35598 (N_35598,N_32332,N_31534);
nand U35599 (N_35599,N_31327,N_33393);
nand U35600 (N_35600,N_33882,N_33379);
nand U35601 (N_35601,N_30325,N_30717);
xnor U35602 (N_35602,N_34421,N_30463);
or U35603 (N_35603,N_30083,N_34172);
or U35604 (N_35604,N_31798,N_31066);
and U35605 (N_35605,N_34519,N_30896);
or U35606 (N_35606,N_31889,N_31028);
nor U35607 (N_35607,N_34566,N_34632);
nor U35608 (N_35608,N_34596,N_34273);
nor U35609 (N_35609,N_31712,N_34112);
or U35610 (N_35610,N_30663,N_31676);
and U35611 (N_35611,N_31143,N_34360);
nand U35612 (N_35612,N_34867,N_33244);
and U35613 (N_35613,N_31027,N_34747);
nor U35614 (N_35614,N_34369,N_33368);
or U35615 (N_35615,N_32996,N_32274);
or U35616 (N_35616,N_30449,N_33700);
or U35617 (N_35617,N_30566,N_31198);
xor U35618 (N_35618,N_33888,N_30003);
and U35619 (N_35619,N_30571,N_33949);
and U35620 (N_35620,N_31757,N_34717);
nand U35621 (N_35621,N_31127,N_31653);
or U35622 (N_35622,N_31183,N_34891);
or U35623 (N_35623,N_34525,N_34854);
or U35624 (N_35624,N_32064,N_33546);
and U35625 (N_35625,N_34495,N_32034);
and U35626 (N_35626,N_34729,N_33595);
or U35627 (N_35627,N_30234,N_30261);
or U35628 (N_35628,N_32653,N_30255);
or U35629 (N_35629,N_34159,N_34090);
nand U35630 (N_35630,N_32703,N_34770);
and U35631 (N_35631,N_34325,N_32798);
nand U35632 (N_35632,N_30599,N_32985);
nor U35633 (N_35633,N_30876,N_31024);
nand U35634 (N_35634,N_31614,N_33468);
nor U35635 (N_35635,N_34054,N_34160);
and U35636 (N_35636,N_31789,N_32588);
and U35637 (N_35637,N_34788,N_31883);
and U35638 (N_35638,N_33719,N_31809);
xor U35639 (N_35639,N_30730,N_31509);
nand U35640 (N_35640,N_32649,N_30938);
nor U35641 (N_35641,N_34426,N_30727);
and U35642 (N_35642,N_31924,N_34004);
nor U35643 (N_35643,N_32183,N_30021);
or U35644 (N_35644,N_30651,N_33473);
nand U35645 (N_35645,N_31967,N_30805);
and U35646 (N_35646,N_31252,N_33576);
and U35647 (N_35647,N_33509,N_32289);
and U35648 (N_35648,N_30398,N_32778);
nor U35649 (N_35649,N_33083,N_30388);
and U35650 (N_35650,N_33450,N_31236);
nand U35651 (N_35651,N_32342,N_30429);
or U35652 (N_35652,N_32313,N_33953);
nor U35653 (N_35653,N_33891,N_32417);
nor U35654 (N_35654,N_34093,N_30202);
xnor U35655 (N_35655,N_31381,N_31402);
or U35656 (N_35656,N_31569,N_34131);
or U35657 (N_35657,N_33219,N_34443);
nand U35658 (N_35658,N_34475,N_30836);
or U35659 (N_35659,N_34278,N_33642);
nor U35660 (N_35660,N_34096,N_31572);
nand U35661 (N_35661,N_32694,N_31806);
nor U35662 (N_35662,N_32447,N_30470);
nand U35663 (N_35663,N_33207,N_32148);
and U35664 (N_35664,N_30576,N_34662);
nor U35665 (N_35665,N_34586,N_32253);
or U35666 (N_35666,N_32434,N_32278);
nand U35667 (N_35667,N_33222,N_33894);
xor U35668 (N_35668,N_32796,N_31502);
nor U35669 (N_35669,N_33212,N_33384);
and U35670 (N_35670,N_33312,N_32574);
nor U35671 (N_35671,N_32755,N_31014);
nor U35672 (N_35672,N_32572,N_30333);
nand U35673 (N_35673,N_33628,N_31876);
nor U35674 (N_35674,N_30419,N_30991);
or U35675 (N_35675,N_34126,N_31187);
and U35676 (N_35676,N_32622,N_30751);
and U35677 (N_35677,N_34085,N_32580);
or U35678 (N_35678,N_31383,N_34231);
nand U35679 (N_35679,N_33417,N_31326);
and U35680 (N_35680,N_33676,N_33396);
nand U35681 (N_35681,N_34002,N_34022);
and U35682 (N_35682,N_31674,N_33144);
and U35683 (N_35683,N_31213,N_31909);
nand U35684 (N_35684,N_33578,N_33853);
nor U35685 (N_35685,N_31444,N_33118);
nand U35686 (N_35686,N_30415,N_34196);
nor U35687 (N_35687,N_33451,N_31903);
xor U35688 (N_35688,N_32837,N_32479);
and U35689 (N_35689,N_33846,N_32950);
nand U35690 (N_35690,N_33507,N_31740);
nand U35691 (N_35691,N_30349,N_30521);
nor U35692 (N_35692,N_30193,N_31303);
xor U35693 (N_35693,N_32957,N_32904);
or U35694 (N_35694,N_32557,N_31117);
or U35695 (N_35695,N_31036,N_32290);
and U35696 (N_35696,N_34982,N_32334);
and U35697 (N_35697,N_34879,N_33184);
and U35698 (N_35698,N_34327,N_34448);
or U35699 (N_35699,N_34178,N_33896);
and U35700 (N_35700,N_30832,N_32004);
or U35701 (N_35701,N_32522,N_33952);
xor U35702 (N_35702,N_30140,N_30053);
or U35703 (N_35703,N_33053,N_31655);
xnor U35704 (N_35704,N_31181,N_31940);
and U35705 (N_35705,N_30568,N_31401);
or U35706 (N_35706,N_33756,N_33599);
nand U35707 (N_35707,N_32367,N_34388);
nand U35708 (N_35708,N_34639,N_34557);
nand U35709 (N_35709,N_33667,N_32000);
nor U35710 (N_35710,N_32639,N_30428);
nor U35711 (N_35711,N_30078,N_30177);
nand U35712 (N_35712,N_30931,N_33030);
or U35713 (N_35713,N_31808,N_31031);
or U35714 (N_35714,N_32870,N_34669);
or U35715 (N_35715,N_33814,N_32541);
nand U35716 (N_35716,N_33113,N_33339);
nor U35717 (N_35717,N_33326,N_33740);
nor U35718 (N_35718,N_31658,N_33088);
nor U35719 (N_35719,N_34733,N_32989);
nand U35720 (N_35720,N_30994,N_31106);
nand U35721 (N_35721,N_32864,N_31097);
and U35722 (N_35722,N_33690,N_34827);
nor U35723 (N_35723,N_33918,N_31080);
or U35724 (N_35724,N_30977,N_30054);
and U35725 (N_35725,N_32261,N_32548);
and U35726 (N_35726,N_31582,N_30297);
or U35727 (N_35727,N_30370,N_30540);
and U35728 (N_35728,N_34070,N_31829);
nor U35729 (N_35729,N_30121,N_32840);
or U35730 (N_35730,N_34741,N_31794);
and U35731 (N_35731,N_31611,N_34458);
and U35732 (N_35732,N_30093,N_30290);
nor U35733 (N_35733,N_34158,N_32774);
nor U35734 (N_35734,N_31892,N_33189);
nand U35735 (N_35735,N_34017,N_31870);
nor U35736 (N_35736,N_33999,N_30531);
or U35737 (N_35737,N_34001,N_32273);
or U35738 (N_35738,N_30444,N_32566);
nand U35739 (N_35739,N_33726,N_31052);
or U35740 (N_35740,N_34964,N_32738);
and U35741 (N_35741,N_31375,N_33568);
or U35742 (N_35742,N_32753,N_33237);
xnor U35743 (N_35743,N_33523,N_31905);
nand U35744 (N_35744,N_32280,N_34274);
and U35745 (N_35745,N_31416,N_33914);
nor U35746 (N_35746,N_34280,N_32412);
or U35747 (N_35747,N_31042,N_34378);
nor U35748 (N_35748,N_31047,N_31998);
nand U35749 (N_35749,N_34439,N_31573);
nand U35750 (N_35750,N_31932,N_31847);
nor U35751 (N_35751,N_34402,N_30711);
or U35752 (N_35752,N_33688,N_33481);
nor U35753 (N_35753,N_30395,N_30076);
nand U35754 (N_35754,N_33983,N_31053);
or U35755 (N_35755,N_30033,N_32491);
nor U35756 (N_35756,N_34025,N_32216);
and U35757 (N_35757,N_33540,N_31208);
and U35758 (N_35758,N_34758,N_31773);
or U35759 (N_35759,N_31204,N_34599);
or U35760 (N_35760,N_31739,N_34535);
or U35761 (N_35761,N_32807,N_33381);
or U35762 (N_35762,N_30781,N_31784);
nand U35763 (N_35763,N_32101,N_33475);
nand U35764 (N_35764,N_34944,N_33987);
and U35765 (N_35765,N_33537,N_31130);
and U35766 (N_35766,N_31464,N_30554);
nand U35767 (N_35767,N_31268,N_31507);
or U35768 (N_35768,N_32097,N_33124);
and U35769 (N_35769,N_33463,N_34567);
and U35770 (N_35770,N_31092,N_34946);
nand U35771 (N_35771,N_31962,N_31657);
nor U35772 (N_35772,N_30180,N_34137);
or U35773 (N_35773,N_30241,N_32243);
and U35774 (N_35774,N_33645,N_31388);
or U35775 (N_35775,N_30025,N_33942);
and U35776 (N_35776,N_30007,N_34957);
or U35777 (N_35777,N_30966,N_30192);
nor U35778 (N_35778,N_33963,N_31956);
or U35779 (N_35779,N_30453,N_30445);
and U35780 (N_35780,N_33636,N_33998);
nor U35781 (N_35781,N_31206,N_31656);
nand U35782 (N_35782,N_34980,N_30604);
nor U35783 (N_35783,N_34116,N_32422);
nand U35784 (N_35784,N_30956,N_32663);
xnor U35785 (N_35785,N_31933,N_31803);
or U35786 (N_35786,N_31229,N_33877);
or U35787 (N_35787,N_33981,N_34348);
nand U35788 (N_35788,N_33133,N_32955);
and U35789 (N_35789,N_30813,N_32630);
or U35790 (N_35790,N_32856,N_33305);
nor U35791 (N_35791,N_32841,N_32322);
nand U35792 (N_35792,N_33767,N_31785);
nand U35793 (N_35793,N_33404,N_30794);
nand U35794 (N_35794,N_31527,N_32407);
nand U35795 (N_35795,N_31767,N_30035);
or U35796 (N_35796,N_31168,N_32432);
or U35797 (N_35797,N_30527,N_33142);
nor U35798 (N_35798,N_33657,N_30204);
nor U35799 (N_35799,N_32224,N_34009);
nor U35800 (N_35800,N_33234,N_34308);
xor U35801 (N_35801,N_33804,N_30422);
nand U35802 (N_35802,N_34383,N_31165);
nor U35803 (N_35803,N_30592,N_30535);
nor U35804 (N_35804,N_34170,N_30697);
and U35805 (N_35805,N_34799,N_31201);
nand U35806 (N_35806,N_31974,N_33994);
xor U35807 (N_35807,N_34678,N_32799);
and U35808 (N_35808,N_31353,N_31620);
or U35809 (N_35809,N_34333,N_30184);
and U35810 (N_35810,N_31652,N_33851);
nor U35811 (N_35811,N_33900,N_30706);
and U35812 (N_35812,N_32111,N_32940);
and U35813 (N_35813,N_32596,N_31811);
or U35814 (N_35814,N_30170,N_33930);
xnor U35815 (N_35815,N_33500,N_32204);
nor U35816 (N_35816,N_32269,N_31282);
or U35817 (N_35817,N_31603,N_33973);
nor U35818 (N_35818,N_34408,N_34996);
or U35819 (N_35819,N_30015,N_31564);
nand U35820 (N_35820,N_33570,N_31026);
and U35821 (N_35821,N_31691,N_30245);
and U35822 (N_35822,N_34859,N_32458);
or U35823 (N_35823,N_32398,N_30432);
nand U35824 (N_35824,N_30890,N_34546);
and U35825 (N_35825,N_30904,N_33669);
nand U35826 (N_35826,N_32803,N_33202);
nor U35827 (N_35827,N_34314,N_34734);
nand U35828 (N_35828,N_34831,N_31929);
and U35829 (N_35829,N_32784,N_32029);
and U35830 (N_35830,N_30979,N_32364);
or U35831 (N_35831,N_33796,N_32854);
and U35832 (N_35832,N_34708,N_31872);
nand U35833 (N_35833,N_30582,N_34410);
nand U35834 (N_35834,N_30351,N_34556);
nand U35835 (N_35835,N_33427,N_30773);
xor U35836 (N_35836,N_31751,N_31467);
nand U35837 (N_35837,N_33317,N_31366);
nand U35838 (N_35838,N_31119,N_32900);
or U35839 (N_35839,N_34892,N_32259);
and U35840 (N_35840,N_31447,N_34304);
and U35841 (N_35841,N_34517,N_33016);
or U35842 (N_35842,N_30666,N_34565);
nor U35843 (N_35843,N_30529,N_33823);
nand U35844 (N_35844,N_32249,N_32720);
xnor U35845 (N_35845,N_33436,N_32325);
nand U35846 (N_35846,N_30837,N_33122);
nor U35847 (N_35847,N_34628,N_32700);
nand U35848 (N_35848,N_32716,N_33782);
and U35849 (N_35849,N_34083,N_31445);
nor U35850 (N_35850,N_32404,N_33309);
xor U35851 (N_35851,N_31184,N_34679);
and U35852 (N_35852,N_32266,N_30998);
nand U35853 (N_35853,N_34214,N_30650);
or U35854 (N_35854,N_32010,N_33071);
nor U35855 (N_35855,N_32783,N_31625);
and U35856 (N_35856,N_34464,N_31006);
or U35857 (N_35857,N_32980,N_34908);
and U35858 (N_35858,N_31135,N_33658);
or U35859 (N_35859,N_34607,N_34190);
and U35860 (N_35860,N_31721,N_31977);
nor U35861 (N_35861,N_33566,N_30311);
or U35862 (N_35862,N_34285,N_34512);
or U35863 (N_35863,N_31071,N_30110);
nand U35864 (N_35864,N_32418,N_30785);
nand U35865 (N_35865,N_33735,N_30084);
nor U35866 (N_35866,N_34375,N_33978);
or U35867 (N_35867,N_32085,N_30657);
xnor U35868 (N_35868,N_32549,N_30716);
and U35869 (N_35869,N_31043,N_34761);
or U35870 (N_35870,N_34059,N_31133);
and U35871 (N_35871,N_30480,N_30981);
nand U35872 (N_35872,N_30380,N_34256);
nor U35873 (N_35873,N_31920,N_30274);
nor U35874 (N_35874,N_30922,N_31604);
and U35875 (N_35875,N_30064,N_31263);
and U35876 (N_35876,N_31765,N_34727);
nor U35877 (N_35877,N_31615,N_33018);
nand U35878 (N_35878,N_31129,N_31816);
and U35879 (N_35879,N_34915,N_32217);
and U35880 (N_35880,N_31525,N_34578);
nor U35881 (N_35881,N_33429,N_33114);
nor U35882 (N_35882,N_30667,N_34051);
or U35883 (N_35883,N_34014,N_33059);
and U35884 (N_35884,N_32003,N_30243);
or U35885 (N_35885,N_33203,N_33401);
and U35886 (N_35886,N_33300,N_34094);
xor U35887 (N_35887,N_34210,N_30880);
or U35888 (N_35888,N_33020,N_31062);
or U35889 (N_35889,N_34904,N_31041);
or U35890 (N_35890,N_31144,N_34202);
nand U35891 (N_35891,N_31384,N_33757);
nor U35892 (N_35892,N_33400,N_32511);
xor U35893 (N_35893,N_33940,N_32206);
or U35894 (N_35894,N_33023,N_31164);
nand U35895 (N_35895,N_31984,N_31448);
and U35896 (N_35896,N_30279,N_32922);
and U35897 (N_35897,N_32005,N_33405);
and U35898 (N_35898,N_31731,N_33937);
or U35899 (N_35899,N_30155,N_32191);
nand U35900 (N_35900,N_33567,N_33745);
or U35901 (N_35901,N_33677,N_32512);
or U35902 (N_35902,N_34857,N_32182);
and U35903 (N_35903,N_34737,N_31244);
and U35904 (N_35904,N_33104,N_30968);
nor U35905 (N_35905,N_33397,N_30256);
nand U35906 (N_35906,N_30997,N_33233);
nand U35907 (N_35907,N_32308,N_33901);
and U35908 (N_35908,N_33648,N_30617);
or U35909 (N_35909,N_30250,N_32239);
or U35910 (N_35910,N_34502,N_33835);
or U35911 (N_35911,N_32355,N_32220);
or U35912 (N_35912,N_33115,N_30120);
and U35913 (N_35913,N_31769,N_32915);
and U35914 (N_35914,N_33550,N_32258);
xnor U35915 (N_35915,N_31665,N_34716);
nand U35916 (N_35916,N_32053,N_32550);
or U35917 (N_35917,N_32810,N_32546);
nor U35918 (N_35918,N_34437,N_31972);
or U35919 (N_35919,N_30189,N_30360);
and U35920 (N_35920,N_32820,N_33571);
xnor U35921 (N_35921,N_32762,N_34066);
nand U35922 (N_35922,N_30049,N_30796);
and U35923 (N_35923,N_33554,N_30731);
nand U35924 (N_35924,N_30485,N_30462);
nand U35925 (N_35925,N_33670,N_32523);
and U35926 (N_35926,N_31491,N_34394);
nor U35927 (N_35927,N_32993,N_32899);
or U35928 (N_35928,N_30490,N_31355);
or U35929 (N_35929,N_30591,N_31854);
or U35930 (N_35930,N_32874,N_33534);
nor U35931 (N_35931,N_33176,N_34181);
or U35932 (N_35932,N_32295,N_30119);
nor U35933 (N_35933,N_34179,N_34434);
and U35934 (N_35934,N_34817,N_31719);
and U35935 (N_35935,N_31523,N_34819);
or U35936 (N_35936,N_32331,N_32648);
xnor U35937 (N_35937,N_31581,N_31373);
or U35938 (N_35938,N_33165,N_31528);
and U35939 (N_35939,N_34189,N_34366);
or U35940 (N_35940,N_31703,N_31515);
nand U35941 (N_35941,N_30879,N_31699);
nand U35942 (N_35942,N_33347,N_30647);
and U35943 (N_35943,N_30969,N_33573);
and U35944 (N_35944,N_30361,N_31927);
nand U35945 (N_35945,N_34527,N_33342);
or U35946 (N_35946,N_31227,N_31205);
nand U35947 (N_35947,N_33232,N_31597);
nand U35948 (N_35948,N_31828,N_33774);
nor U35949 (N_35949,N_33418,N_34776);
and U35950 (N_35950,N_34453,N_30541);
nor U35951 (N_35951,N_31154,N_30532);
nand U35952 (N_35952,N_32154,N_34775);
or U35953 (N_35953,N_31695,N_30112);
nand U35954 (N_35954,N_33455,N_34229);
and U35955 (N_35955,N_33302,N_30680);
xnor U35956 (N_35956,N_34132,N_31701);
or U35957 (N_35957,N_31677,N_31170);
nor U35958 (N_35958,N_33861,N_33615);
nor U35959 (N_35959,N_30446,N_30980);
and U35960 (N_35960,N_32822,N_31988);
nand U35961 (N_35961,N_31365,N_33067);
and U35962 (N_35962,N_32863,N_31641);
nor U35963 (N_35963,N_33452,N_31708);
xnor U35964 (N_35964,N_33556,N_31145);
and U35965 (N_35965,N_34583,N_34532);
and U35966 (N_35966,N_31007,N_34133);
and U35967 (N_35967,N_31166,N_32423);
and U35968 (N_35968,N_34625,N_33932);
and U35969 (N_35969,N_34306,N_32440);
nand U35970 (N_35970,N_32282,N_30841);
xor U35971 (N_35971,N_33935,N_30157);
and U35972 (N_35972,N_32547,N_32818);
nor U35973 (N_35973,N_31637,N_33652);
xor U35974 (N_35974,N_31411,N_31842);
and U35975 (N_35975,N_30744,N_33517);
nand U35976 (N_35976,N_30334,N_33093);
or U35977 (N_35977,N_32173,N_33501);
nor U35978 (N_35978,N_31367,N_30277);
nor U35979 (N_35979,N_34213,N_34293);
or U35980 (N_35980,N_34005,N_32677);
xor U35981 (N_35981,N_33884,N_32998);
and U35982 (N_35982,N_34676,N_31937);
and U35983 (N_35983,N_31214,N_33227);
nand U35984 (N_35984,N_32124,N_34034);
nor U35985 (N_35985,N_33777,N_31189);
nor U35986 (N_35986,N_30798,N_33499);
or U35987 (N_35987,N_31245,N_32581);
nor U35988 (N_35988,N_33166,N_34992);
or U35989 (N_35989,N_33872,N_33744);
and U35990 (N_35990,N_34511,N_31774);
nand U35991 (N_35991,N_33997,N_33678);
and U35992 (N_35992,N_33209,N_33225);
or U35993 (N_35993,N_34030,N_31137);
nand U35994 (N_35994,N_32802,N_32067);
and U35995 (N_35995,N_32098,N_30579);
nor U35996 (N_35996,N_32055,N_31858);
and U35997 (N_35997,N_32654,N_31458);
nand U35998 (N_35998,N_32271,N_34600);
nor U35999 (N_35999,N_31192,N_30509);
and U36000 (N_36000,N_34743,N_33443);
nand U36001 (N_36001,N_32773,N_34813);
nand U36002 (N_36002,N_34301,N_31049);
nor U36003 (N_36003,N_34960,N_34263);
nor U36004 (N_36004,N_31345,N_34560);
or U36005 (N_36005,N_34696,N_33366);
or U36006 (N_36006,N_34088,N_30203);
and U36007 (N_36007,N_34673,N_32866);
and U36008 (N_36008,N_33727,N_32211);
xor U36009 (N_36009,N_31980,N_33287);
and U36010 (N_36010,N_31406,N_34445);
nor U36011 (N_36011,N_34345,N_34203);
nand U36012 (N_36012,N_34454,N_30212);
xor U36013 (N_36013,N_30649,N_34663);
nor U36014 (N_36014,N_34312,N_32666);
and U36015 (N_36015,N_33348,N_33082);
nand U36016 (N_36016,N_31662,N_34064);
nand U36017 (N_36017,N_33693,N_34355);
and U36018 (N_36018,N_33471,N_30803);
nand U36019 (N_36019,N_31436,N_34482);
nor U36020 (N_36020,N_31242,N_32327);
and U36021 (N_36021,N_30477,N_33254);
nand U36022 (N_36022,N_30134,N_32264);
and U36023 (N_36023,N_34198,N_30341);
nand U36024 (N_36024,N_33694,N_30668);
and U36025 (N_36025,N_32749,N_31241);
xnor U36026 (N_36026,N_30978,N_33749);
or U36027 (N_36027,N_30639,N_31738);
and U36028 (N_36028,N_30209,N_34503);
nor U36029 (N_36029,N_33352,N_32878);
or U36030 (N_36030,N_31362,N_32939);
or U36031 (N_36031,N_33240,N_31960);
nor U36032 (N_36032,N_31219,N_31543);
or U36033 (N_36033,N_34440,N_34473);
nand U36034 (N_36034,N_32298,N_33715);
nand U36035 (N_36035,N_34665,N_30263);
and U36036 (N_36036,N_34045,N_32573);
nor U36037 (N_36037,N_32143,N_32905);
and U36038 (N_36038,N_31571,N_34856);
or U36039 (N_36039,N_31022,N_33871);
and U36040 (N_36040,N_30726,N_32660);
or U36041 (N_36041,N_32707,N_32178);
xor U36042 (N_36042,N_32268,N_34284);
nor U36043 (N_36043,N_34321,N_30011);
nor U36044 (N_36044,N_34138,N_34550);
nand U36045 (N_36045,N_33415,N_34809);
and U36046 (N_36046,N_33541,N_31484);
and U36047 (N_36047,N_31742,N_32044);
or U36048 (N_36048,N_34694,N_33532);
and U36049 (N_36049,N_34689,N_33604);
or U36050 (N_36050,N_32435,N_33250);
xor U36051 (N_36051,N_30139,N_30464);
nor U36052 (N_36052,N_32126,N_32758);
nand U36053 (N_36053,N_30642,N_31250);
and U36054 (N_36054,N_32689,N_32932);
or U36055 (N_36055,N_33126,N_33299);
or U36056 (N_36056,N_30063,N_33029);
nor U36057 (N_36057,N_33771,N_30748);
nand U36058 (N_36058,N_32808,N_33533);
nand U36059 (N_36059,N_34861,N_30696);
nand U36060 (N_36060,N_33986,N_30061);
nand U36061 (N_36061,N_34236,N_31182);
or U36062 (N_36062,N_31317,N_31827);
and U36063 (N_36063,N_34476,N_34650);
nor U36064 (N_36064,N_31138,N_30989);
and U36065 (N_36065,N_32604,N_33068);
nor U36066 (N_36066,N_31163,N_34998);
nand U36067 (N_36067,N_33903,N_34319);
nor U36068 (N_36068,N_32971,N_32049);
xnor U36069 (N_36069,N_31034,N_34906);
nor U36070 (N_36070,N_32819,N_34399);
xnor U36071 (N_36071,N_31413,N_34307);
or U36072 (N_36072,N_33385,N_33346);
and U36073 (N_36073,N_32166,N_31709);
nor U36074 (N_36074,N_33284,N_32534);
and U36075 (N_36075,N_30611,N_32698);
nand U36076 (N_36076,N_30372,N_33923);
nor U36077 (N_36077,N_33629,N_31804);
or U36078 (N_36078,N_32387,N_34646);
or U36079 (N_36079,N_33821,N_34780);
and U36080 (N_36080,N_34412,N_33283);
xnor U36081 (N_36081,N_31005,N_31954);
or U36082 (N_36082,N_32227,N_32144);
nand U36083 (N_36083,N_33638,N_31949);
and U36084 (N_36084,N_31610,N_33685);
nand U36085 (N_36085,N_31844,N_32556);
or U36086 (N_36086,N_32172,N_32234);
nor U36087 (N_36087,N_31567,N_31928);
nand U36088 (N_36088,N_34658,N_33453);
nor U36089 (N_36089,N_34485,N_34884);
nand U36090 (N_36090,N_34334,N_34423);
and U36091 (N_36091,N_34349,N_32742);
xor U36092 (N_36092,N_30974,N_34351);
nand U36093 (N_36093,N_33137,N_31726);
and U36094 (N_36094,N_33857,N_31149);
xor U36095 (N_36095,N_31570,N_32343);
nand U36096 (N_36096,N_31966,N_30257);
and U36097 (N_36097,N_32804,N_32062);
and U36098 (N_36098,N_32456,N_32256);
or U36099 (N_36099,N_30957,N_30842);
or U36100 (N_36100,N_33263,N_32382);
nand U36101 (N_36101,N_34409,N_34222);
or U36102 (N_36102,N_32611,N_33160);
nand U36103 (N_36103,N_33858,N_32267);
and U36104 (N_36104,N_31037,N_34156);
xor U36105 (N_36105,N_34128,N_30636);
nor U36106 (N_36106,N_34933,N_33692);
nor U36107 (N_36107,N_32340,N_30402);
xnor U36108 (N_36108,N_31780,N_32222);
nor U36109 (N_36109,N_30831,N_30448);
and U36110 (N_36110,N_31826,N_33335);
xor U36111 (N_36111,N_31171,N_33065);
or U36112 (N_36112,N_32717,N_31501);
nand U36113 (N_36113,N_30098,N_30893);
xnor U36114 (N_36114,N_30659,N_34768);
nor U36115 (N_36115,N_34250,N_31896);
nor U36116 (N_36116,N_33549,N_33279);
nand U36117 (N_36117,N_33634,N_32726);
nor U36118 (N_36118,N_34487,N_32683);
nand U36119 (N_36119,N_34790,N_34810);
nand U36120 (N_36120,N_33921,N_32747);
nor U36121 (N_36121,N_31778,N_32039);
and U36122 (N_36122,N_30742,N_30465);
nor U36123 (N_36123,N_32208,N_31083);
or U36124 (N_36124,N_30229,N_32401);
and U36125 (N_36125,N_32761,N_30963);
or U36126 (N_36126,N_31343,N_32357);
and U36127 (N_36127,N_32492,N_31125);
nor U36128 (N_36128,N_33208,N_32093);
nor U36129 (N_36129,N_33409,N_32210);
nor U36130 (N_36130,N_34637,N_33145);
nand U36131 (N_36131,N_31056,N_33524);
nand U36132 (N_36132,N_34139,N_31989);
or U36133 (N_36133,N_32984,N_32947);
and U36134 (N_36134,N_32843,N_34713);
nand U36135 (N_36135,N_30447,N_31272);
and U36136 (N_36136,N_30747,N_33431);
or U36137 (N_36137,N_31435,N_31667);
nand U36138 (N_36138,N_31481,N_31095);
nand U36139 (N_36139,N_34752,N_32131);
nand U36140 (N_36140,N_31161,N_33569);
nand U36141 (N_36141,N_31983,N_32655);
and U36142 (N_36142,N_31207,N_33490);
nand U36143 (N_36143,N_30378,N_30769);
or U36144 (N_36144,N_30635,N_33332);
nor U36145 (N_36145,N_30427,N_32345);
xor U36146 (N_36146,N_31583,N_30927);
nor U36147 (N_36147,N_32270,N_34466);
and U36148 (N_36148,N_33506,N_33177);
nand U36149 (N_36149,N_32066,N_30625);
or U36150 (N_36150,N_31796,N_33376);
nor U36151 (N_36151,N_34923,N_31814);
nor U36152 (N_36152,N_33581,N_31790);
and U36153 (N_36153,N_34935,N_31817);
xnor U36154 (N_36154,N_33057,N_30825);
nor U36155 (N_36155,N_31728,N_33600);
nand U36156 (N_36156,N_32564,N_30218);
nor U36157 (N_36157,N_30213,N_34217);
and U36158 (N_36158,N_30705,N_31454);
xnor U36159 (N_36159,N_31511,N_31850);
nor U36160 (N_36160,N_30045,N_33040);
or U36161 (N_36161,N_32192,N_34740);
or U36162 (N_36162,N_30043,N_34880);
nand U36163 (N_36163,N_32935,N_32620);
nand U36164 (N_36164,N_30393,N_33913);
nor U36165 (N_36165,N_32475,N_34205);
and U36166 (N_36166,N_30559,N_34275);
nand U36167 (N_36167,N_34288,N_30087);
and U36168 (N_36168,N_30339,N_31643);
nand U36169 (N_36169,N_30525,N_31424);
or U36170 (N_36170,N_32995,N_30732);
and U36171 (N_36171,N_32410,N_33580);
and U36172 (N_36172,N_34873,N_31420);
or U36173 (N_36173,N_33223,N_33086);
nand U36174 (N_36174,N_34864,N_30877);
nor U36175 (N_36175,N_33046,N_32699);
xnor U36176 (N_36176,N_32790,N_33909);
and U36177 (N_36177,N_32732,N_31749);
or U36178 (N_36178,N_33808,N_31867);
and U36179 (N_36179,N_31239,N_32961);
nand U36180 (N_36180,N_32246,N_34922);
nand U36181 (N_36181,N_33766,N_32095);
and U36182 (N_36182,N_32867,N_34259);
or U36183 (N_36183,N_34168,N_30235);
nor U36184 (N_36184,N_30442,N_31012);
or U36185 (N_36185,N_34011,N_30430);
and U36186 (N_36186,N_32953,N_32248);
and U36187 (N_36187,N_34833,N_33887);
xor U36188 (N_36188,N_30829,N_30498);
nor U36189 (N_36189,N_32136,N_33422);
or U36190 (N_36190,N_31449,N_34816);
and U36191 (N_36191,N_34834,N_34690);
or U36192 (N_36192,N_31076,N_31073);
nand U36193 (N_36193,N_34918,N_32520);
or U36194 (N_36194,N_30806,N_32911);
or U36195 (N_36195,N_34342,N_33492);
or U36196 (N_36196,N_34220,N_30924);
nor U36197 (N_36197,N_34675,N_33535);
nand U36198 (N_36198,N_34403,N_32718);
nand U36199 (N_36199,N_31743,N_31630);
and U36200 (N_36200,N_33746,N_31223);
nor U36201 (N_36201,N_31524,N_30809);
xor U36202 (N_36202,N_32017,N_31452);
or U36203 (N_36203,N_33589,N_30276);
nand U36204 (N_36204,N_31081,N_30909);
nand U36205 (N_36205,N_33880,N_34498);
xnor U36206 (N_36206,N_33881,N_34405);
nand U36207 (N_36207,N_30107,N_32378);
nand U36208 (N_36208,N_31915,N_31562);
and U36209 (N_36209,N_31926,N_30080);
nor U36210 (N_36210,N_33256,N_30865);
nor U36211 (N_36211,N_34038,N_30578);
nand U36212 (N_36212,N_32533,N_31574);
and U36213 (N_36213,N_34563,N_30500);
or U36214 (N_36214,N_32920,N_31859);
and U36215 (N_36215,N_33793,N_31880);
nand U36216 (N_36216,N_33286,N_32307);
or U36217 (N_36217,N_34255,N_32811);
and U36218 (N_36218,N_30147,N_32544);
or U36219 (N_36219,N_34109,N_34396);
or U36220 (N_36220,N_31750,N_34091);
nor U36221 (N_36221,N_30362,N_34769);
nor U36222 (N_36222,N_33097,N_31871);
or U36223 (N_36223,N_34281,N_33839);
and U36224 (N_36224,N_30534,N_33827);
and U36225 (N_36225,N_34433,N_30772);
xnor U36226 (N_36226,N_31633,N_34882);
or U36227 (N_36227,N_30971,N_34677);
nand U36228 (N_36228,N_30721,N_31663);
xnor U36229 (N_36229,N_34941,N_30357);
or U36230 (N_36230,N_31203,N_34446);
nand U36231 (N_36231,N_34478,N_30654);
xnor U36232 (N_36232,N_34121,N_32901);
or U36233 (N_36233,N_31776,N_33840);
or U36234 (N_36234,N_34183,N_33560);
xor U36235 (N_36235,N_31599,N_31579);
or U36236 (N_36236,N_30467,N_31912);
and U36237 (N_36237,N_32519,N_31060);
and U36238 (N_36238,N_33849,N_31863);
nor U36239 (N_36239,N_30452,N_32476);
xnor U36240 (N_36240,N_31755,N_31993);
and U36241 (N_36241,N_30864,N_33647);
nor U36242 (N_36242,N_31698,N_32028);
nor U36243 (N_36243,N_32443,N_30797);
nand U36244 (N_36244,N_34211,N_34513);
and U36245 (N_36245,N_30150,N_30715);
nor U36246 (N_36246,N_33614,N_30648);
nor U36247 (N_36247,N_30205,N_32791);
nor U36248 (N_36248,N_34559,N_30834);
and U36249 (N_36249,N_34971,N_30226);
nand U36250 (N_36250,N_33229,N_30113);
or U36251 (N_36251,N_32959,N_32484);
and U36252 (N_36252,N_34529,N_30780);
nand U36253 (N_36253,N_32433,N_32895);
or U36254 (N_36254,N_30888,N_33832);
nor U36255 (N_36255,N_30102,N_34693);
nand U36256 (N_36256,N_31232,N_34268);
or U36257 (N_36257,N_32240,N_33341);
or U36258 (N_36258,N_33869,N_32518);
nor U36259 (N_36259,N_30310,N_32631);
nand U36260 (N_36260,N_34614,N_34674);
nor U36261 (N_36261,N_34297,N_34173);
nor U36262 (N_36262,N_31902,N_34523);
xnor U36263 (N_36263,N_30374,N_30088);
nand U36264 (N_36264,N_31015,N_32319);
or U36265 (N_36265,N_30686,N_33127);
or U36266 (N_36266,N_33683,N_32361);
nand U36267 (N_36267,N_30640,N_30660);
xor U36268 (N_36268,N_31587,N_31802);
nand U36269 (N_36269,N_32158,N_34749);
and U36270 (N_36270,N_32659,N_33725);
nand U36271 (N_36271,N_32214,N_30367);
or U36272 (N_36272,N_31350,N_31478);
and U36273 (N_36273,N_33971,N_33631);
nor U36274 (N_36274,N_30530,N_34260);
nor U36275 (N_36275,N_30638,N_32383);
nor U36276 (N_36276,N_31957,N_33070);
nand U36277 (N_36277,N_30206,N_32705);
and U36278 (N_36278,N_30949,N_30267);
xnor U36279 (N_36279,N_33948,N_34672);
nand U36280 (N_36280,N_31228,N_34575);
and U36281 (N_36281,N_32457,N_32488);
nand U36282 (N_36282,N_33239,N_31221);
xor U36283 (N_36283,N_31266,N_31293);
or U36284 (N_36284,N_34926,N_31335);
or U36285 (N_36285,N_31799,N_32938);
and U36286 (N_36286,N_30321,N_33338);
nand U36287 (N_36287,N_32834,N_31720);
nand U36288 (N_36288,N_32160,N_30006);
nand U36289 (N_36289,N_31474,N_33487);
nor U36290 (N_36290,N_30214,N_32428);
nor U36291 (N_36291,N_34814,N_30135);
nand U36292 (N_36292,N_34850,N_32287);
nor U36293 (N_36293,N_34815,N_33543);
xnor U36294 (N_36294,N_32300,N_30390);
and U36295 (N_36295,N_32559,N_33295);
or U36296 (N_36296,N_33183,N_31351);
or U36297 (N_36297,N_30172,N_30600);
and U36298 (N_36298,N_30459,N_30223);
nor U36299 (N_36299,N_34023,N_34577);
nand U36300 (N_36300,N_33221,N_32982);
and U36301 (N_36301,N_33128,N_34292);
or U36302 (N_36302,N_31249,N_31818);
nor U36303 (N_36303,N_34188,N_33132);
or U36304 (N_36304,N_34585,N_31098);
and U36305 (N_36305,N_33802,N_32977);
xnor U36306 (N_36306,N_34382,N_32397);
nor U36307 (N_36307,N_31300,N_33095);
nor U36308 (N_36308,N_33035,N_31233);
nand U36309 (N_36309,N_30739,N_33758);
and U36310 (N_36310,N_34629,N_30345);
and U36311 (N_36311,N_32729,N_34692);
nor U36312 (N_36312,N_34953,N_31810);
or U36313 (N_36313,N_30117,N_32242);
or U36314 (N_36314,N_30787,N_30593);
xor U36315 (N_36315,N_30312,N_32632);
or U36316 (N_36316,N_30677,N_33742);
nor U36317 (N_36317,N_30665,N_30925);
or U36318 (N_36318,N_30608,N_33868);
and U36319 (N_36319,N_30507,N_30898);
nor U36320 (N_36320,N_34792,N_33003);
nor U36321 (N_36321,N_30905,N_34961);
or U36322 (N_36322,N_33388,N_30058);
and U36323 (N_36323,N_34018,N_34555);
and U36324 (N_36324,N_33625,N_31465);
nand U36325 (N_36325,N_33195,N_34636);
xor U36326 (N_36326,N_31359,N_30743);
nor U36327 (N_36327,N_31724,N_33424);
nand U36328 (N_36328,N_33019,N_31279);
nand U36329 (N_36329,N_31823,N_31772);
or U36330 (N_36330,N_30937,N_30930);
or U36331 (N_36331,N_30068,N_31099);
or U36332 (N_36332,N_32179,N_34258);
nor U36333 (N_36333,N_32769,N_33557);
nand U36334 (N_36334,N_30012,N_31462);
nand U36335 (N_36335,N_30698,N_33825);
and U36336 (N_36336,N_32658,N_32021);
and U36337 (N_36337,N_34618,N_33281);
and U36338 (N_36338,N_30392,N_32465);
and U36339 (N_36339,N_31886,N_32988);
or U36340 (N_36340,N_33380,N_33632);
nand U36341 (N_36341,N_34240,N_31476);
nand U36342 (N_36342,N_30673,N_32390);
or U36343 (N_36343,N_31103,N_30239);
xor U36344 (N_36344,N_32276,N_31522);
nor U36345 (N_36345,N_33623,N_30010);
nor U36346 (N_36346,N_30778,N_32296);
and U36347 (N_36347,N_30894,N_32825);
nor U36348 (N_36348,N_30258,N_32634);
nand U36349 (N_36349,N_33765,N_31990);
xnor U36350 (N_36350,N_32197,N_30109);
xnor U36351 (N_36351,N_34951,N_34584);
and U36352 (N_36352,N_34766,N_33817);
or U36353 (N_36353,N_34794,N_33970);
and U36354 (N_36354,N_32970,N_30607);
nand U36355 (N_36355,N_31340,N_34490);
nor U36356 (N_36356,N_34104,N_31169);
and U36357 (N_36357,N_33140,N_31315);
or U36358 (N_36358,N_34652,N_33373);
and U36359 (N_36359,N_32855,N_33845);
nand U36360 (N_36360,N_30283,N_30515);
nand U36361 (N_36361,N_34245,N_31685);
nand U36362 (N_36362,N_33255,N_33272);
nor U36363 (N_36363,N_33559,N_31085);
and U36364 (N_36364,N_30982,N_34514);
xnor U36365 (N_36365,N_33428,N_32680);
xnor U36366 (N_36366,N_34595,N_30158);
nand U36367 (N_36367,N_34374,N_30086);
nand U36368 (N_36368,N_32719,N_33939);
and U36369 (N_36369,N_32481,N_34509);
or U36370 (N_36370,N_32842,N_33959);
or U36371 (N_36371,N_30557,N_32656);
nor U36372 (N_36372,N_34779,N_34483);
or U36373 (N_36373,N_32812,N_32896);
or U36374 (N_36374,N_32069,N_31580);
xnor U36375 (N_36375,N_32650,N_34886);
nand U36376 (N_36376,N_34791,N_30694);
or U36377 (N_36377,N_34594,N_34313);
and U36378 (N_36378,N_33852,N_31951);
nand U36379 (N_36379,N_30707,N_30584);
and U36380 (N_36380,N_34043,N_32190);
nor U36381 (N_36381,N_33747,N_34337);
nand U36382 (N_36382,N_34921,N_34385);
nor U36383 (N_36383,N_30198,N_32647);
and U36384 (N_36384,N_33781,N_31175);
xor U36385 (N_36385,N_33390,N_34602);
nor U36386 (N_36386,N_31919,N_31235);
and U36387 (N_36387,N_30708,N_30236);
nor U36388 (N_36388,N_34542,N_33377);
nor U36389 (N_36389,N_34140,N_32196);
and U36390 (N_36390,N_31513,N_31275);
nor U36391 (N_36391,N_32038,N_33945);
or U36392 (N_36392,N_34201,N_33336);
or U36393 (N_36393,N_33439,N_31234);
or U36394 (N_36394,N_31922,N_33893);
xor U36395 (N_36395,N_32147,N_34157);
nand U36396 (N_36396,N_33503,N_30626);
and U36397 (N_36397,N_32586,N_30176);
and U36398 (N_36398,N_32092,N_30861);
or U36399 (N_36399,N_32019,N_33584);
nand U36400 (N_36400,N_34504,N_31503);
and U36401 (N_36401,N_34078,N_30704);
and U36402 (N_36402,N_33345,N_32960);
nor U36403 (N_36403,N_31180,N_32007);
nand U36404 (N_36404,N_30222,N_34435);
or U36405 (N_36405,N_33094,N_30961);
and U36406 (N_36406,N_31185,N_32921);
or U36407 (N_36407,N_33590,N_30502);
and U36408 (N_36408,N_31044,N_31459);
nor U36409 (N_36409,N_33855,N_31309);
nand U36410 (N_36410,N_33425,N_33762);
or U36411 (N_36411,N_33204,N_33433);
and U36412 (N_36412,N_34613,N_31077);
or U36413 (N_36413,N_34046,N_30853);
or U36414 (N_36414,N_34155,N_31779);
nor U36415 (N_36415,N_32846,N_32056);
nand U36416 (N_36416,N_32030,N_31162);
nand U36417 (N_36417,N_30724,N_34101);
and U36418 (N_36418,N_33358,N_30305);
and U36419 (N_36419,N_32472,N_30308);
xnor U36420 (N_36420,N_34936,N_34451);
and U36421 (N_36421,N_30118,N_33792);
nand U36422 (N_36422,N_30528,N_34135);
nor U36423 (N_36423,N_33192,N_32310);
or U36424 (N_36424,N_33440,N_34630);
nor U36425 (N_36425,N_34571,N_33156);
and U36426 (N_36426,N_31838,N_34253);
and U36427 (N_36427,N_32805,N_32245);
and U36428 (N_36428,N_31016,N_32363);
xor U36429 (N_36429,N_31952,N_33199);
xnor U36430 (N_36430,N_33874,N_31510);
xnor U36431 (N_36431,N_31629,N_32061);
nor U36432 (N_36432,N_34533,N_30903);
or U36433 (N_36433,N_32770,N_31332);
and U36434 (N_36434,N_32226,N_30761);
or U36435 (N_36435,N_31594,N_33252);
or U36436 (N_36436,N_31550,N_34099);
nor U36437 (N_36437,N_31945,N_33477);
nand U36438 (N_36438,N_33876,N_33664);
nand U36439 (N_36439,N_30580,N_34199);
nand U36440 (N_36440,N_34714,N_30100);
nor U36441 (N_36441,N_32370,N_30952);
or U36442 (N_36442,N_32462,N_33729);
nor U36443 (N_36443,N_32425,N_30685);
xnor U36444 (N_36444,N_33674,N_31914);
or U36445 (N_36445,N_34916,N_31555);
or U36446 (N_36446,N_31908,N_31371);
nor U36447 (N_36447,N_33432,N_30852);
or U36448 (N_36448,N_33064,N_30389);
nor U36449 (N_36449,N_30056,N_34680);
or U36450 (N_36450,N_31953,N_30383);
nand U36451 (N_36451,N_31694,N_34832);
xnor U36452 (N_36452,N_32975,N_33141);
nor U36453 (N_36453,N_34130,N_30799);
nor U36454 (N_36454,N_31417,N_34531);
nor U36455 (N_36455,N_34619,N_34683);
nand U36456 (N_36456,N_30478,N_33701);
nor U36457 (N_36457,N_30827,N_31730);
nand U36458 (N_36458,N_34553,N_30095);
and U36459 (N_36459,N_30441,N_32106);
xnor U36460 (N_36460,N_30363,N_31298);
nor U36461 (N_36461,N_32695,N_34425);
nand U36462 (N_36462,N_33120,N_30630);
and U36463 (N_36463,N_31453,N_32032);
nor U36464 (N_36464,N_31979,N_31618);
nand U36465 (N_36465,N_30783,N_30154);
or U36466 (N_36466,N_30067,N_30471);
and U36467 (N_36467,N_31461,N_34783);
xnor U36468 (N_36468,N_34978,N_31023);
xnor U36469 (N_36469,N_30545,N_31626);
nor U36470 (N_36470,N_33905,N_33485);
and U36471 (N_36471,N_34161,N_31094);
nand U36472 (N_36472,N_32952,N_33854);
nor U36473 (N_36473,N_34145,N_32991);
nor U36474 (N_36474,N_30511,N_30800);
nor U36475 (N_36475,N_31222,N_34897);
nand U36476 (N_36476,N_32260,N_33105);
xor U36477 (N_36477,N_34986,N_32916);
nor U36478 (N_36478,N_33297,N_33268);
nand U36479 (N_36479,N_33946,N_32115);
nand U36480 (N_36480,N_33929,N_34969);
nor U36481 (N_36481,N_32601,N_30319);
or U36482 (N_36482,N_31054,N_33924);
or U36483 (N_36483,N_32014,N_30153);
or U36484 (N_36484,N_33601,N_31820);
nand U36485 (N_36485,N_30491,N_33587);
nor U36486 (N_36486,N_31428,N_31306);
nand U36487 (N_36487,N_31122,N_31240);
nor U36488 (N_36488,N_30352,N_30913);
or U36489 (N_36489,N_34685,N_34272);
and U36490 (N_36490,N_31913,N_32329);
and U36491 (N_36491,N_33553,N_32116);
nand U36492 (N_36492,N_32203,N_32080);
and U36493 (N_36493,N_32483,N_33895);
or U36494 (N_36494,N_32185,N_32070);
and U36495 (N_36495,N_34186,N_30148);
nor U36496 (N_36496,N_31994,N_33226);
and U36497 (N_36497,N_31632,N_33819);
nand U36498 (N_36498,N_31256,N_34510);
and U36499 (N_36499,N_33763,N_30348);
nand U36500 (N_36500,N_32607,N_30770);
or U36501 (N_36501,N_32286,N_34460);
nor U36502 (N_36502,N_31982,N_33818);
nor U36503 (N_36503,N_32076,N_33843);
or U36504 (N_36504,N_34786,N_33847);
xor U36505 (N_36505,N_34075,N_33734);
nand U36506 (N_36506,N_32781,N_34463);
nand U36507 (N_36507,N_31815,N_34860);
or U36508 (N_36508,N_32375,N_33175);
and U36509 (N_36509,N_32543,N_31217);
or U36510 (N_36510,N_31911,N_34249);
or U36511 (N_36511,N_32502,N_31533);
or U36512 (N_36512,N_30411,N_32023);
and U36513 (N_36513,N_32354,N_33941);
nor U36514 (N_36514,N_30795,N_33489);
nand U36515 (N_36515,N_32436,N_34803);
or U36516 (N_36516,N_34644,N_33656);
nand U36517 (N_36517,N_34027,N_32015);
nor U36518 (N_36518,N_30619,N_33323);
or U36519 (N_36519,N_30200,N_32949);
and U36520 (N_36520,N_34174,N_30300);
and U36521 (N_36521,N_31549,N_33979);
nand U36522 (N_36522,N_32937,N_33266);
nor U36523 (N_36523,N_32373,N_31361);
nand U36524 (N_36524,N_30871,N_30366);
and U36525 (N_36525,N_34805,N_31150);
nor U36526 (N_36526,N_32643,N_32221);
nand U36527 (N_36527,N_30440,N_30886);
xor U36528 (N_36528,N_32117,N_30718);
or U36529 (N_36529,N_34238,N_34060);
or U36530 (N_36530,N_31568,N_34195);
and U36531 (N_36531,N_34344,N_31639);
nor U36532 (N_36532,N_33423,N_33447);
or U36533 (N_36533,N_33456,N_31475);
nor U36534 (N_36534,N_31392,N_32657);
or U36535 (N_36535,N_30942,N_30451);
or U36536 (N_36536,N_30484,N_31939);
nor U36537 (N_36537,N_34928,N_30030);
or U36538 (N_36538,N_31714,N_32480);
and U36539 (N_36539,N_34422,N_32344);
nand U36540 (N_36540,N_33026,N_33392);
or U36541 (N_36541,N_32139,N_33196);
nor U36542 (N_36542,N_31609,N_34610);
or U36543 (N_36543,N_30499,N_30508);
and U36544 (N_36544,N_32079,N_33442);
and U36545 (N_36545,N_33607,N_30754);
or U36546 (N_36546,N_32202,N_32025);
or U36547 (N_36547,N_32853,N_32281);
xor U36548 (N_36548,N_34225,N_32482);
xnor U36549 (N_36549,N_31211,N_33975);
nand U36550 (N_36550,N_32869,N_31142);
nor U36551 (N_36551,N_31848,N_31923);
nor U36552 (N_36552,N_33467,N_34457);
nor U36553 (N_36553,N_32275,N_34609);
and U36554 (N_36554,N_33486,N_30967);
and U36555 (N_36555,N_34449,N_34354);
nor U36556 (N_36556,N_32112,N_32928);
and U36557 (N_36557,N_33836,N_31735);
and U36558 (N_36558,N_30005,N_34106);
xnor U36559 (N_36559,N_31090,N_33334);
nand U36560 (N_36560,N_30329,N_32265);
nor U36561 (N_36561,N_30460,N_32623);
and U36562 (N_36562,N_34955,N_30185);
nor U36563 (N_36563,N_33926,N_32529);
nand U36564 (N_36564,N_34398,N_32979);
and U36565 (N_36565,N_34003,N_34604);
and U36566 (N_36566,N_30840,N_30814);
and U36567 (N_36567,N_32052,N_31781);
xnor U36568 (N_36568,N_33100,N_32925);
nor U36569 (N_36569,N_33412,N_30784);
or U36570 (N_36570,N_30096,N_32441);
xnor U36571 (N_36571,N_34795,N_30343);
nor U36572 (N_36572,N_30394,N_30688);
or U36573 (N_36573,N_34216,N_31176);
and U36574 (N_36574,N_34835,N_33148);
xnor U36575 (N_36575,N_30401,N_31545);
nand U36576 (N_36576,N_31451,N_34558);
and U36577 (N_36577,N_31531,N_33659);
or U36578 (N_36578,N_32645,N_32946);
and U36579 (N_36579,N_30207,N_30359);
nand U36580 (N_36580,N_30028,N_33479);
nor U36581 (N_36581,N_31763,N_34608);
xor U36582 (N_36582,N_34606,N_34924);
nand U36583 (N_36583,N_33174,N_31959);
and U36584 (N_36584,N_31675,N_30573);
nor U36585 (N_36585,N_33797,N_31634);
xor U36586 (N_36586,N_32489,N_31640);
and U36587 (N_36587,N_31931,N_32813);
or U36588 (N_36588,N_31660,N_30315);
and U36589 (N_36589,N_30759,N_34134);
nor U36590 (N_36590,N_31947,N_32068);
nor U36591 (N_36591,N_30296,N_34777);
nor U36592 (N_36592,N_33538,N_33582);
and U36593 (N_36593,N_31822,N_34122);
nor U36594 (N_36594,N_31853,N_32594);
nand U36595 (N_36595,N_33917,N_33885);
nor U36596 (N_36596,N_32598,N_33248);
or U36597 (N_36597,N_31669,N_32380);
and U36598 (N_36598,N_32997,N_30547);
nand U36599 (N_36599,N_32132,N_31267);
nor U36600 (N_36600,N_30208,N_31586);
nand U36601 (N_36601,N_33591,N_30944);
nand U36602 (N_36602,N_30801,N_30137);
or U36603 (N_36603,N_32366,N_34641);
xnor U36604 (N_36604,N_31596,N_34389);
or U36605 (N_36605,N_30679,N_30168);
and U36606 (N_36606,N_31322,N_32109);
and U36607 (N_36607,N_34948,N_34208);
nand U36608 (N_36608,N_34049,N_31807);
xnor U36609 (N_36609,N_32752,N_31753);
and U36610 (N_36610,N_33322,N_31386);
or U36611 (N_36611,N_34670,N_30476);
nand U36612 (N_36612,N_31264,N_33982);
or U36613 (N_36613,N_31177,N_34709);
nand U36614 (N_36614,N_32612,N_32427);
and U36615 (N_36615,N_31100,N_30496);
xnor U36616 (N_36616,N_31120,N_31231);
nor U36617 (N_36617,N_31139,N_31875);
nand U36618 (N_36618,N_31865,N_33547);
and U36619 (N_36619,N_32671,N_30767);
or U36620 (N_36620,N_31330,N_30910);
or U36621 (N_36621,N_33613,N_34521);
nand U36622 (N_36622,N_32504,N_30855);
nand U36623 (N_36623,N_33794,N_34942);
nor U36624 (N_36624,N_30412,N_31157);
or U36625 (N_36625,N_34930,N_31174);
nor U36626 (N_36626,N_30847,N_31216);
and U36627 (N_36627,N_34974,N_32525);
and U36628 (N_36628,N_32486,N_32102);
nand U36629 (N_36629,N_32629,N_31297);
nor U36630 (N_36630,N_34237,N_31955);
and U36631 (N_36631,N_34191,N_33610);
or U36632 (N_36632,N_32727,N_33915);
nor U36633 (N_36633,N_32711,N_33096);
nor U36634 (N_36634,N_30958,N_34579);
xnor U36635 (N_36635,N_34910,N_33671);
and U36636 (N_36636,N_30335,N_30523);
nand U36637 (N_36637,N_33755,N_30031);
nand U36638 (N_36638,N_33382,N_30433);
xor U36639 (N_36639,N_31040,N_31186);
xnor U36640 (N_36640,N_30397,N_33544);
nand U36641 (N_36641,N_32824,N_34013);
nand U36642 (N_36642,N_34753,N_30899);
nor U36643 (N_36643,N_32035,N_33640);
xnor U36644 (N_36644,N_30344,N_30627);
or U36645 (N_36645,N_30835,N_32613);
xnor U36646 (N_36646,N_34824,N_30870);
and U36647 (N_36647,N_30437,N_34949);
or U36648 (N_36648,N_34912,N_31713);
nor U36649 (N_36649,N_30326,N_30438);
and U36650 (N_36650,N_31074,N_32187);
nor U36651 (N_36651,N_30586,N_32477);
nand U36652 (N_36652,N_32231,N_32615);
xor U36653 (N_36653,N_30387,N_33178);
nor U36654 (N_36654,N_31410,N_33616);
nor U36655 (N_36655,N_32006,N_30062);
or U36656 (N_36656,N_32552,N_32165);
and U36657 (N_36657,N_32605,N_34987);
and U36658 (N_36658,N_30703,N_34764);
nand U36659 (N_36659,N_30346,N_30273);
and U36660 (N_36660,N_33714,N_33247);
or U36661 (N_36661,N_32444,N_33044);
and U36662 (N_36662,N_34432,N_30935);
nor U36663 (N_36663,N_33916,N_32723);
nor U36664 (N_36664,N_30494,N_34212);
or U36665 (N_36665,N_30486,N_30190);
or U36666 (N_36666,N_31777,N_30828);
or U36667 (N_36667,N_33277,N_31039);
nand U36668 (N_36668,N_33988,N_30519);
xor U36669 (N_36669,N_31030,N_33354);
and U36670 (N_36670,N_34667,N_33902);
xnor U36671 (N_36671,N_33315,N_30676);
nor U36672 (N_36672,N_30816,N_30556);
or U36673 (N_36673,N_33790,N_31884);
nor U36674 (N_36674,N_30542,N_32751);
and U36675 (N_36675,N_32130,N_34568);
nor U36676 (N_36676,N_34276,N_30757);
nand U36677 (N_36677,N_32223,N_34787);
xor U36678 (N_36678,N_31616,N_31707);
nor U36679 (N_36679,N_33806,N_31050);
or U36680 (N_36680,N_30089,N_32071);
nor U36681 (N_36681,N_34180,N_31628);
and U36682 (N_36682,N_34806,N_31251);
nor U36683 (N_36683,N_32057,N_32027);
nor U36684 (N_36684,N_31585,N_31357);
or U36685 (N_36685,N_34839,N_34152);
nor U36686 (N_36686,N_34840,N_31899);
nor U36687 (N_36687,N_34381,N_30071);
or U36688 (N_36688,N_32585,N_31258);
or U36689 (N_36689,N_34295,N_34919);
nand U36690 (N_36690,N_31055,N_33224);
xnor U36691 (N_36691,N_31747,N_30774);
nand U36692 (N_36692,N_34643,N_30550);
nor U36693 (N_36693,N_32201,N_33011);
and U36694 (N_36694,N_31795,N_33363);
xnor U36695 (N_36695,N_33280,N_30947);
nand U36696 (N_36696,N_31917,N_31045);
xnor U36697 (N_36697,N_32315,N_31692);
nand U36698 (N_36698,N_34875,N_34956);
and U36699 (N_36699,N_30999,N_33830);
and U36700 (N_36700,N_31212,N_34703);
nand U36701 (N_36701,N_30199,N_34668);
and U36702 (N_36702,N_32712,N_31885);
and U36703 (N_36703,N_34244,N_33708);
nand U36704 (N_36704,N_31441,N_30167);
and U36705 (N_36705,N_33892,N_30403);
or U36706 (N_36706,N_34627,N_34491);
nor U36707 (N_36707,N_32786,N_34711);
and U36708 (N_36708,N_31600,N_34855);
nor U36709 (N_36709,N_30240,N_32914);
nor U36710 (N_36710,N_32438,N_32890);
and U36711 (N_36711,N_33045,N_34373);
or U36712 (N_36712,N_33991,N_32907);
and U36713 (N_36713,N_33960,N_31399);
nor U36714 (N_36714,N_31787,N_31305);
or U36715 (N_36715,N_34881,N_34655);
nor U36716 (N_36716,N_31197,N_32888);
and U36717 (N_36717,N_34376,N_31727);
nand U36718 (N_36718,N_30672,N_30020);
and U36719 (N_36719,N_30354,N_30373);
or U36720 (N_36720,N_33889,N_34114);
and U36721 (N_36721,N_34182,N_34247);
and U36722 (N_36722,N_31584,N_31079);
nor U36723 (N_36723,N_30587,N_32386);
and U36724 (N_36724,N_31259,N_34778);
xnor U36725 (N_36725,N_32943,N_30658);
nand U36726 (N_36726,N_33684,N_32527);
nor U36727 (N_36727,N_32151,N_33066);
or U36728 (N_36728,N_30032,N_33611);
nand U36729 (N_36729,N_34098,N_34581);
and U36730 (N_36730,N_31519,N_31768);
nand U36731 (N_36731,N_33783,N_33316);
and U36732 (N_36732,N_31278,N_30669);
or U36733 (N_36733,N_31468,N_32141);
nor U36734 (N_36734,N_30259,N_30406);
nor U36735 (N_36735,N_32668,N_30569);
or U36736 (N_36736,N_33454,N_33731);
nand U36737 (N_36737,N_34937,N_33886);
nor U36738 (N_36738,N_33608,N_31195);
xnor U36739 (N_36739,N_33555,N_34322);
nor U36740 (N_36740,N_31389,N_31457);
or U36741 (N_36741,N_33080,N_32365);
and U36742 (N_36742,N_30598,N_33505);
nor U36743 (N_36743,N_31304,N_33351);
or U36744 (N_36744,N_30472,N_30804);
nor U36745 (N_36745,N_33421,N_30336);
nor U36746 (N_36746,N_30996,N_33964);
nand U36747 (N_36747,N_31113,N_32510);
nand U36748 (N_36748,N_32886,N_31710);
or U36749 (N_36749,N_34117,N_30561);
or U36750 (N_36750,N_32473,N_32963);
xnor U36751 (N_36751,N_33480,N_33010);
xor U36752 (N_36752,N_32540,N_32828);
nand U36753 (N_36753,N_33856,N_31837);
and U36754 (N_36754,N_34838,N_30085);
and U36755 (N_36755,N_34589,N_34419);
nor U36756 (N_36756,N_32782,N_30330);
or U36757 (N_36757,N_31376,N_32212);
nand U36758 (N_36758,N_34765,N_31430);
nand U36759 (N_36759,N_30018,N_30306);
nor U36760 (N_36760,N_32652,N_33592);
or U36761 (N_36761,N_31942,N_33704);
xnor U36762 (N_36762,N_33586,N_34151);
nor U36763 (N_36763,N_32009,N_33972);
nand U36764 (N_36764,N_31999,N_31115);
nor U36765 (N_36765,N_32377,N_32584);
nor U36766 (N_36766,N_31514,N_34686);
and U36767 (N_36767,N_32163,N_30309);
nor U36768 (N_36768,N_30810,N_32013);
nor U36769 (N_36769,N_33251,N_32024);
nand U36770 (N_36770,N_32688,N_33661);
nor U36771 (N_36771,N_30169,N_31943);
nor U36772 (N_36772,N_31372,N_30163);
nand U36773 (N_36773,N_30741,N_33504);
and U36774 (N_36774,N_30577,N_30629);
xnor U36775 (N_36775,N_34598,N_32094);
nand U36776 (N_36776,N_33079,N_32424);
nand U36777 (N_36777,N_31194,N_33596);
or U36778 (N_36778,N_32156,N_32134);
or U36779 (N_36779,N_32207,N_31754);
or U36780 (N_36780,N_31225,N_30094);
nor U36781 (N_36781,N_32251,N_34735);
or U36782 (N_36782,N_30141,N_32589);
nor U36783 (N_36783,N_33651,N_32213);
and U36784 (N_36784,N_30298,N_30285);
nor U36785 (N_36785,N_34638,N_34315);
nand U36786 (N_36786,N_30818,N_34080);
xnor U36787 (N_36787,N_32785,N_30070);
nor U36788 (N_36788,N_34878,N_33470);
and U36789 (N_36789,N_33048,N_34732);
or U36790 (N_36790,N_32930,N_34082);
nand U36791 (N_36791,N_34468,N_32320);
nand U36792 (N_36792,N_30073,N_32554);
nor U36793 (N_36793,N_34063,N_33372);
nand U36794 (N_36794,N_31541,N_33784);
and U36795 (N_36795,N_30251,N_30891);
or U36796 (N_36796,N_30823,N_33271);
nor U36797 (N_36797,N_31084,N_32450);
and U36798 (N_36798,N_30954,N_33791);
nand U36799 (N_36799,N_33403,N_34095);
xnor U36800 (N_36800,N_32521,N_30385);
and U36801 (N_36801,N_30425,N_33938);
and U36802 (N_36802,N_34751,N_34353);
nor U36803 (N_36803,N_31132,N_31682);
xnor U36804 (N_36804,N_34954,N_34544);
nor U36805 (N_36805,N_32389,N_34868);
nor U36806 (N_36806,N_30099,N_30188);
xor U36807 (N_36807,N_30720,N_34150);
nor U36808 (N_36808,N_32501,N_34461);
and U36809 (N_36809,N_30355,N_32022);
xor U36810 (N_36810,N_30789,N_30175);
and U36811 (N_36811,N_32218,N_30736);
or U36812 (N_36812,N_32575,N_31123);
xor U36813 (N_36813,N_32236,N_32777);
nor U36814 (N_36814,N_31148,N_30762);
and U36815 (N_36815,N_30884,N_31973);
xor U36816 (N_36816,N_34427,N_31971);
nand U36817 (N_36817,N_30288,N_33270);
and U36818 (N_36818,N_32490,N_34489);
nor U36819 (N_36819,N_34111,N_30483);
or U36820 (N_36820,N_31349,N_33246);
and U36821 (N_36821,N_33201,N_32942);
nor U36822 (N_36822,N_31737,N_34615);
nor U36823 (N_36823,N_32149,N_34100);
xnor U36824 (N_36824,N_33720,N_30304);
nor U36825 (N_36825,N_30558,N_31429);
and U36826 (N_36826,N_31644,N_30270);
nand U36827 (N_36827,N_30868,N_32725);
nand U36828 (N_36828,N_34993,N_30143);
and U36829 (N_36829,N_34793,N_30645);
nand U36830 (N_36830,N_32724,N_30450);
nand U36831 (N_36831,N_32104,N_31617);
and U36832 (N_36832,N_31328,N_33545);
nand U36833 (N_36833,N_30819,N_33012);
or U36834 (N_36834,N_34989,N_34501);
nor U36835 (N_36835,N_32860,N_32602);
nor U36836 (N_36836,N_32538,N_33087);
and U36837 (N_36837,N_33278,N_34136);
nand U36838 (N_36838,N_30381,N_34326);
and U36839 (N_36839,N_32847,N_34570);
or U36840 (N_36840,N_33768,N_30737);
xnor U36841 (N_36841,N_32277,N_30272);
or U36842 (N_36842,N_31895,N_32181);
or U36843 (N_36843,N_30596,N_32155);
nor U36844 (N_36844,N_31456,N_30262);
or U36845 (N_36845,N_32670,N_30603);
nand U36846 (N_36846,N_34404,N_32919);
and U36847 (N_36847,N_30424,N_32621);
or U36848 (N_36848,N_33458,N_34950);
or U36849 (N_36849,N_31390,N_31443);
nor U36850 (N_36850,N_33911,N_31237);
nand U36851 (N_36851,N_32312,N_30594);
or U36852 (N_36852,N_33890,N_34858);
nor U36853 (N_36853,N_33922,N_32687);
and U36854 (N_36854,N_30013,N_30675);
and U36855 (N_36855,N_30563,N_30643);
nor U36856 (N_36856,N_30601,N_33077);
nor U36857 (N_36857,N_30008,N_34028);
or U36858 (N_36858,N_30623,N_31672);
nor U36859 (N_36859,N_31078,N_33274);
xor U36860 (N_36860,N_32195,N_32110);
or U36861 (N_36861,N_32238,N_31622);
xor U36862 (N_36862,N_30017,N_30041);
nand U36863 (N_36863,N_30081,N_30123);
nand U36864 (N_36864,N_32346,N_31874);
or U36865 (N_36865,N_32795,N_33699);
nor U36866 (N_36866,N_33850,N_30889);
or U36867 (N_36867,N_34943,N_30431);
or U36868 (N_36868,N_33013,N_34340);
or U36869 (N_36869,N_33014,N_33967);
nor U36870 (N_36870,N_33273,N_30090);
and U36871 (N_36871,N_33803,N_32180);
or U36872 (N_36872,N_32225,N_30897);
nor U36873 (N_36873,N_31262,N_33515);
xnor U36874 (N_36874,N_32739,N_33061);
or U36875 (N_36875,N_32257,N_31801);
and U36876 (N_36876,N_30457,N_32247);
nand U36877 (N_36877,N_33943,N_33441);
nand U36878 (N_36878,N_33110,N_30752);
xor U36879 (N_36879,N_33076,N_32873);
and U36880 (N_36880,N_33739,N_31344);
nor U36881 (N_36881,N_32918,N_30691);
nand U36882 (N_36882,N_34358,N_31281);
nand U36883 (N_36883,N_31352,N_30941);
nor U36884 (N_36884,N_32351,N_34821);
nor U36885 (N_36885,N_30106,N_31946);
nor U36886 (N_36886,N_32001,N_30407);
or U36887 (N_36887,N_33950,N_33787);
and U36888 (N_36888,N_32682,N_30264);
or U36889 (N_36889,N_30520,N_30788);
xor U36890 (N_36890,N_34547,N_34959);
or U36891 (N_36891,N_31869,N_30733);
nand U36892 (N_36892,N_33898,N_32797);
nand U36893 (N_36893,N_31935,N_30856);
or U36894 (N_36894,N_31374,N_32674);
and U36895 (N_36895,N_33150,N_32429);
or U36896 (N_36896,N_33179,N_34902);
nand U36897 (N_36897,N_30318,N_32463);
or U36898 (N_36898,N_33449,N_32526);
nand U36899 (N_36899,N_33091,N_34647);
and U36900 (N_36900,N_33445,N_32973);
and U36901 (N_36901,N_34722,N_32293);
and U36902 (N_36902,N_33117,N_34661);
xnor U36903 (N_36903,N_32399,N_32892);
nand U36904 (N_36904,N_34552,N_30271);
and U36905 (N_36905,N_33474,N_32194);
nand U36906 (N_36906,N_30016,N_34772);
or U36907 (N_36907,N_34981,N_32965);
or U36908 (N_36908,N_31287,N_32446);
nand U36909 (N_36909,N_32333,N_30371);
or U36910 (N_36910,N_34032,N_32100);
nor U36911 (N_36911,N_31852,N_30765);
nor U36912 (N_36912,N_34362,N_34296);
nor U36913 (N_36913,N_33050,N_33980);
or U36914 (N_36914,N_33660,N_31422);
nand U36915 (N_36915,N_33733,N_31202);
nor U36916 (N_36916,N_32135,N_30364);
nand U36917 (N_36917,N_34176,N_30970);
nand U36918 (N_36918,N_34759,N_34699);
nor U36919 (N_36919,N_34719,N_30846);
nand U36920 (N_36920,N_31992,N_32091);
nand U36921 (N_36921,N_33402,N_32627);
and U36922 (N_36922,N_31536,N_32951);
nand U36923 (N_36923,N_33106,N_33024);
or U36924 (N_36924,N_30230,N_33976);
nand U36925 (N_36925,N_34745,N_34682);
nor U36926 (N_36926,N_30750,N_31065);
and U36927 (N_36927,N_34129,N_31671);
and U36928 (N_36928,N_31577,N_30295);
and U36929 (N_36929,N_31687,N_32599);
nor U36930 (N_36930,N_30160,N_34789);
nand U36931 (N_36931,N_31431,N_32188);
or U36932 (N_36932,N_34391,N_34530);
nand U36933 (N_36933,N_33241,N_34811);
and U36934 (N_36934,N_32532,N_31409);
or U36935 (N_36935,N_33675,N_34456);
nor U36936 (N_36936,N_32722,N_34371);
nand U36937 (N_36937,N_32731,N_31748);
nand U36938 (N_36938,N_33907,N_33525);
nand U36939 (N_36939,N_31965,N_34750);
nor U36940 (N_36940,N_31613,N_33724);
nand U36941 (N_36941,N_30543,N_31554);
or U36942 (N_36942,N_31224,N_34252);
or U36943 (N_36943,N_33934,N_32036);
nand U36944 (N_36944,N_33697,N_32122);
nor U36945 (N_36945,N_32849,N_31118);
nor U36946 (N_36946,N_31061,N_34621);
and U36947 (N_36947,N_32198,N_30238);
or U36948 (N_36948,N_34496,N_31505);
nand U36949 (N_36949,N_31595,N_30103);
or U36950 (N_36950,N_34573,N_31793);
nand U36951 (N_36951,N_30858,N_31011);
and U36952 (N_36952,N_33728,N_30838);
xor U36953 (N_36953,N_33510,N_31354);
or U36954 (N_36954,N_33152,N_34925);
and U36955 (N_36955,N_32046,N_30735);
or U36956 (N_36956,N_34077,N_31020);
and U36957 (N_36957,N_34505,N_32583);
nand U36958 (N_36958,N_34756,N_33180);
nand U36959 (N_36959,N_31038,N_33301);
and U36960 (N_36960,N_30807,N_31813);
and U36961 (N_36961,N_34357,N_32851);
or U36962 (N_36962,N_32931,N_32829);
nand U36963 (N_36963,N_33620,N_30943);
or U36964 (N_36964,N_32848,N_31159);
and U36965 (N_36965,N_34290,N_32644);
or U36966 (N_36966,N_33820,N_34995);
nor U36967 (N_36967,N_34561,N_32442);
and U36968 (N_36968,N_32262,N_30195);
xnor U36969 (N_36969,N_31226,N_32898);
and U36970 (N_36970,N_32073,N_34781);
nand U36971 (N_36971,N_32823,N_34808);
or U36972 (N_36972,N_34087,N_30145);
and U36973 (N_36973,N_30959,N_31002);
nand U36974 (N_36974,N_31683,N_30413);
and U36975 (N_36975,N_34548,N_33644);
nand U36976 (N_36976,N_30723,N_31623);
and U36977 (N_36977,N_33238,N_30404);
and U36978 (N_36978,N_30589,N_30050);
nor U36979 (N_36979,N_34331,N_34849);
or U36980 (N_36980,N_34338,N_31775);
xor U36981 (N_36981,N_33218,N_34691);
nor U36982 (N_36982,N_31762,N_31729);
or U36983 (N_36983,N_30934,N_32635);
nor U36984 (N_36984,N_33081,N_32495);
nor U36985 (N_36985,N_30328,N_33681);
and U36986 (N_36986,N_33870,N_33170);
and U36987 (N_36987,N_31841,N_33349);
nor U36988 (N_36988,N_34488,N_34113);
nand U36989 (N_36989,N_30225,N_34317);
nand U36990 (N_36990,N_30042,N_33276);
nand U36991 (N_36991,N_34287,N_31879);
and U36992 (N_36992,N_32592,N_33815);
and U36993 (N_36993,N_31560,N_34911);
or U36994 (N_36994,N_31378,N_31230);
nor U36995 (N_36995,N_34612,N_30946);
or U36996 (N_36996,N_34812,N_33444);
and U36997 (N_36997,N_30104,N_34187);
nand U36998 (N_36998,N_30987,N_31542);
nor U36999 (N_36999,N_32303,N_34372);
nand U37000 (N_37000,N_32033,N_32145);
or U37001 (N_37001,N_30105,N_30416);
or U37002 (N_37002,N_34169,N_30900);
and U37003 (N_37003,N_32565,N_32040);
or U37004 (N_37004,N_33572,N_34283);
nand U37005 (N_37005,N_34826,N_31466);
nor U37006 (N_37006,N_33285,N_32839);
and U37007 (N_37007,N_31051,N_31882);
or U37008 (N_37008,N_32171,N_30133);
nor U37009 (N_37009,N_32099,N_34232);
nor U37010 (N_37010,N_33102,N_34945);
nor U37011 (N_37011,N_30505,N_30955);
and U37012 (N_37012,N_31426,N_31432);
xnor U37013 (N_37013,N_34681,N_32909);
and U37014 (N_37014,N_30358,N_34239);
nand U37015 (N_37015,N_32294,N_34339);
or U37016 (N_37016,N_31134,N_32041);
nand U37017 (N_37017,N_30027,N_34407);
and U37018 (N_37018,N_34695,N_34118);
nand U37019 (N_37019,N_33776,N_32672);
and U37020 (N_37020,N_34738,N_34486);
and U37021 (N_37021,N_30986,N_32560);
and U37022 (N_37022,N_32692,N_33123);
and U37023 (N_37023,N_32678,N_32349);
nand U37024 (N_37024,N_34893,N_34450);
nand U37025 (N_37025,N_33099,N_31651);
nor U37026 (N_37026,N_30533,N_31552);
and U37027 (N_37027,N_32184,N_30034);
or U37028 (N_37028,N_32944,N_30746);
nand U37029 (N_37029,N_31308,N_31588);
nor U37030 (N_37030,N_33306,N_32317);
nor U37031 (N_37031,N_30839,N_31846);
and U37032 (N_37032,N_30873,N_30574);
or U37033 (N_37033,N_33253,N_34261);
and U37034 (N_37034,N_30023,N_31210);
or U37035 (N_37035,N_31067,N_32336);
or U37036 (N_37036,N_34141,N_30162);
or U37037 (N_37037,N_34623,N_34518);
and U37038 (N_37038,N_34332,N_30678);
or U37039 (N_37039,N_31338,N_32691);
xnor U37040 (N_37040,N_31082,N_34746);
nor U37041 (N_37041,N_30683,N_31591);
nand U37042 (N_37042,N_32409,N_30332);
and U37043 (N_37043,N_33482,N_34044);
nor U37044 (N_37044,N_30052,N_31188);
or U37045 (N_37045,N_31602,N_31152);
or U37046 (N_37046,N_32832,N_34350);
and U37047 (N_37047,N_31140,N_31680);
and U37048 (N_37048,N_30565,N_33111);
xor U37049 (N_37049,N_32114,N_32323);
or U37050 (N_37050,N_34702,N_31473);
nand U37051 (N_37051,N_31000,N_34251);
nand U37052 (N_37052,N_30130,N_30161);
and U37053 (N_37053,N_32306,N_33552);
or U37054 (N_37054,N_31500,N_32500);
nand U37055 (N_37055,N_33021,N_31009);
and U37056 (N_37056,N_33837,N_33325);
and U37057 (N_37057,N_32775,N_33561);
xnor U37058 (N_37058,N_31666,N_31363);
nand U37059 (N_37059,N_32882,N_30356);
nor U37060 (N_37060,N_33135,N_32704);
or U37061 (N_37061,N_32042,N_33197);
or U37062 (N_37062,N_32414,N_31004);
or U37063 (N_37063,N_33786,N_34438);
nand U37064 (N_37064,N_33732,N_30048);
or U37065 (N_37065,N_32459,N_30538);
xor U37066 (N_37066,N_33158,N_33985);
and U37067 (N_37067,N_30618,N_33770);
and U37068 (N_37068,N_33780,N_30936);
or U37069 (N_37069,N_34649,N_34055);
nand U37070 (N_37070,N_31593,N_34266);
nor U37071 (N_37071,N_34016,N_31075);
nand U37072 (N_37072,N_33307,N_32924);
and U37073 (N_37073,N_34221,N_31257);
and U37074 (N_37074,N_30233,N_32750);
or U37075 (N_37075,N_34493,N_33313);
nor U37076 (N_37076,N_30895,N_33529);
and U37077 (N_37077,N_34359,N_34462);
nand U37078 (N_37078,N_30409,N_30609);
nor U37079 (N_37079,N_33577,N_31834);
xnor U37080 (N_37080,N_32059,N_34830);
or U37081 (N_37081,N_31608,N_33419);
nor U37082 (N_37082,N_32127,N_31910);
and U37083 (N_37083,N_30597,N_31260);
or U37084 (N_37084,N_31033,N_30628);
nor U37085 (N_37085,N_32976,N_33435);
xnor U37086 (N_37086,N_34162,N_34865);
xnor U37087 (N_37087,N_34963,N_30396);
xnor U37088 (N_37088,N_32430,N_30562);
nor U37089 (N_37089,N_30194,N_34363);
nor U37090 (N_37090,N_33173,N_33038);
and U37091 (N_37091,N_33516,N_34480);
and U37092 (N_37092,N_32371,N_30661);
nor U37093 (N_37093,N_31495,N_30738);
nand U37094 (N_37094,N_32074,N_31548);
nand U37095 (N_37095,N_30674,N_34597);
xor U37096 (N_37096,N_33116,N_34036);
nor U37097 (N_37097,N_32551,N_34428);
nand U37098 (N_37098,N_30197,N_32793);
and U37099 (N_37099,N_32485,N_34976);
nor U37100 (N_37100,N_30848,N_30253);
and U37101 (N_37101,N_33761,N_31425);
or U37102 (N_37102,N_32872,N_32043);
and U37103 (N_37103,N_33865,N_32174);
nand U37104 (N_37104,N_33751,N_33810);
nor U37105 (N_37105,N_33155,N_31404);
or U37106 (N_37106,N_31414,N_32809);
nand U37107 (N_37107,N_30231,N_33101);
nor U37108 (N_37108,N_32301,N_30621);
xor U37109 (N_37109,N_31797,N_31377);
nor U37110 (N_37110,N_30482,N_31530);
nor U37111 (N_37111,N_31706,N_34624);
xnor U37112 (N_37112,N_33362,N_33508);
or U37113 (N_37113,N_31243,N_33371);
nor U37114 (N_37114,N_34042,N_31930);
nor U37115 (N_37115,N_32740,N_32318);
or U37116 (N_37116,N_32478,N_32881);
nand U37117 (N_37117,N_32701,N_31487);
and U37118 (N_37118,N_32662,N_31247);
or U37119 (N_37119,N_32302,N_30662);
xor U37120 (N_37120,N_32903,N_31178);
nand U37121 (N_37121,N_30111,N_32887);
xnor U37122 (N_37122,N_30689,N_34197);
and U37123 (N_37123,N_30342,N_33668);
xor U37124 (N_37124,N_31734,N_32571);
nor U37125 (N_37125,N_34801,N_30232);
or U37126 (N_37126,N_33275,N_34657);
nand U37127 (N_37127,N_33466,N_34310);
or U37128 (N_37128,N_34712,N_34947);
or U37129 (N_37129,N_30287,N_33460);
nor U37130 (N_37130,N_30939,N_33033);
or U37131 (N_37131,N_34050,N_33242);
nor U37132 (N_37132,N_32400,N_34015);
nand U37133 (N_37133,N_30734,N_33741);
nand U37134 (N_37134,N_33361,N_34590);
nor U37135 (N_37135,N_33695,N_33039);
nand U37136 (N_37136,N_32816,N_33398);
nand U37137 (N_37137,N_34847,N_33521);
or U37138 (N_37138,N_32086,N_34395);
or U37139 (N_37139,N_30369,N_34092);
nand U37140 (N_37140,N_34545,N_31111);
nand U37141 (N_37141,N_34484,N_32814);
or U37142 (N_37142,N_34730,N_30375);
or U37143 (N_37143,N_33597,N_31556);
or U37144 (N_37144,N_31370,N_33860);
and U37145 (N_37145,N_30760,N_34818);
nor U37146 (N_37146,N_32316,N_31419);
and U37147 (N_37147,N_32469,N_32353);
and U37148 (N_37148,N_31438,N_30878);
and U37149 (N_37149,N_32555,N_31089);
and U37150 (N_37150,N_34755,N_32792);
nand U37151 (N_37151,N_30923,N_31057);
nor U37152 (N_37152,N_34149,N_33069);
or U37153 (N_37153,N_34184,N_34424);
nor U37154 (N_37154,N_34784,N_31058);
and U37155 (N_37155,N_31395,N_34171);
nor U37156 (N_37156,N_30964,N_33711);
nor U37157 (N_37157,N_31963,N_30539);
nand U37158 (N_37158,N_32461,N_33579);
or U37159 (N_37159,N_34341,N_30916);
xnor U37160 (N_37160,N_32063,N_34688);
nand U37161 (N_37161,N_32230,N_33965);
nor U37162 (N_37162,N_34177,N_34008);
nand U37163 (N_37163,N_34204,N_32235);
or U37164 (N_37164,N_30316,N_33410);
xnor U37165 (N_37165,N_30817,N_33119);
nor U37166 (N_37166,N_31624,N_32779);
xor U37167 (N_37167,N_31547,N_33996);
and U37168 (N_37168,N_30585,N_33828);
or U37169 (N_37169,N_32279,N_33531);
nand U37170 (N_37170,N_32244,N_34903);
and U37171 (N_37171,N_32956,N_30291);
and U37172 (N_37172,N_31638,N_32806);
nor U37173 (N_37173,N_33469,N_34701);
nand U37174 (N_37174,N_33213,N_34076);
nand U37175 (N_37175,N_33411,N_31423);
nor U37176 (N_37176,N_32421,N_32733);
nor U37177 (N_37177,N_34931,N_34820);
and U37178 (N_37178,N_31761,N_30077);
and U37179 (N_37179,N_31723,N_32146);
or U37180 (N_37180,N_30544,N_34416);
and U37181 (N_37181,N_31696,N_30495);
xor U37182 (N_37182,N_34227,N_32852);
nor U37183 (N_37183,N_30302,N_32439);
nor U37184 (N_37184,N_30174,N_34538);
or U37185 (N_37185,N_32636,N_34444);
nor U37186 (N_37186,N_34706,N_31289);
nor U37187 (N_37187,N_32002,N_32263);
and U37188 (N_37188,N_32763,N_32609);
and U37189 (N_37189,N_33187,N_33637);
nor U37190 (N_37190,N_34081,N_31220);
and U37191 (N_37191,N_33356,N_32894);
and U37192 (N_37192,N_33488,N_32369);
and U37193 (N_37193,N_30882,N_34029);
and U37194 (N_37194,N_32090,N_31093);
nor U37195 (N_37195,N_33841,N_31689);
and U37196 (N_37196,N_32736,N_31285);
and U37197 (N_37197,N_31497,N_34654);
or U37198 (N_37198,N_33310,N_31948);
or U37199 (N_37199,N_30142,N_30040);
nand U37200 (N_37200,N_34999,N_32514);
nor U37201 (N_37201,N_33710,N_31673);
nand U37202 (N_37202,N_32494,N_34209);
nand U37203 (N_37203,N_33257,N_33799);
xnor U37204 (N_37204,N_34723,N_31109);
nor U37205 (N_37205,N_33649,N_32460);
or U37206 (N_37206,N_34329,N_34386);
nand U37207 (N_37207,N_32467,N_31325);
nor U37208 (N_37208,N_32875,N_33051);
and U37209 (N_37209,N_33321,N_31385);
nand U37210 (N_37210,N_33689,N_31368);
and U37211 (N_37211,N_32927,N_34282);
xnor U37212 (N_37212,N_32884,N_31532);
or U37213 (N_37213,N_32877,N_30555);
or U37214 (N_37214,N_33190,N_32159);
nor U37215 (N_37215,N_30454,N_31741);
and U37216 (N_37216,N_34687,N_30815);
and U37217 (N_37217,N_30915,N_34760);
or U37218 (N_37218,N_32506,N_34007);
nor U37219 (N_37219,N_34973,N_31121);
and U37220 (N_37220,N_33603,N_31832);
nor U37221 (N_37221,N_31277,N_30526);
nor U37222 (N_37222,N_31649,N_31538);
nor U37223 (N_37223,N_34215,N_34554);
nor U37224 (N_37224,N_34890,N_32879);
and U37225 (N_37225,N_34848,N_33459);
and U37226 (N_37226,N_32328,N_30791);
nor U37227 (N_37227,N_34802,N_33149);
or U37228 (N_37228,N_33527,N_34048);
xor U37229 (N_37229,N_30749,N_30410);
nand U37230 (N_37230,N_33465,N_30906);
nand U37231 (N_37231,N_30074,N_32193);
nand U37232 (N_37232,N_34368,N_34762);
or U37233 (N_37233,N_34543,N_33703);
nor U37234 (N_37234,N_30059,N_30254);
nor U37235 (N_37235,N_33245,N_33551);
and U37236 (N_37236,N_30246,N_31261);
or U37237 (N_37237,N_30418,N_34035);
xor U37238 (N_37238,N_32524,N_33833);
or U37239 (N_37239,N_33161,N_30514);
or U37240 (N_37240,N_32788,N_30820);
nand U37241 (N_37241,N_31558,N_32748);
or U37242 (N_37242,N_30990,N_30513);
and U37243 (N_37243,N_34336,N_30260);
nor U37244 (N_37244,N_30845,N_32767);
nand U37245 (N_37245,N_32766,N_34997);
nor U37246 (N_37246,N_34829,N_32603);
xnor U37247 (N_37247,N_34380,N_34972);
nor U37248 (N_37248,N_34877,N_31897);
nor U37249 (N_37249,N_31104,N_32060);
and U37250 (N_37250,N_34958,N_34895);
nor U37251 (N_37251,N_33662,N_31645);
nand U37252 (N_37252,N_33375,N_34154);
or U37253 (N_37253,N_33406,N_32737);
xnor U37254 (N_37254,N_32451,N_31286);
or U37255 (N_37255,N_33333,N_33476);
nand U37256 (N_37256,N_33243,N_30777);
nor U37257 (N_37257,N_31479,N_32335);
nand U37258 (N_37258,N_31697,N_33809);
and U37259 (N_37259,N_31894,N_32167);
nor U37260 (N_37260,N_31635,N_33705);
xnor U37261 (N_37261,N_33558,N_30338);
and U37262 (N_37262,N_34108,N_33542);
nand U37263 (N_37263,N_33461,N_30960);
nor U37264 (N_37264,N_30976,N_33304);
or U37265 (N_37265,N_33748,N_33956);
nor U37266 (N_37266,N_34105,N_34153);
or U37267 (N_37267,N_32103,N_30215);
nor U37268 (N_37268,N_34089,N_32408);
nor U37269 (N_37269,N_30000,N_30517);
or U37270 (N_37270,N_33157,N_34970);
and U37271 (N_37271,N_30644,N_30365);
or U37272 (N_37272,N_33564,N_32402);
or U37273 (N_37273,N_33957,N_32987);
nor U37274 (N_37274,N_34286,N_33259);
and U37275 (N_37275,N_34536,N_32967);
and U37276 (N_37276,N_34052,N_34640);
nor U37277 (N_37277,N_31480,N_31433);
or U37278 (N_37278,N_34323,N_30758);
nand U37279 (N_37279,N_32113,N_32018);
or U37280 (N_37280,N_34874,N_34539);
nor U37281 (N_37281,N_30920,N_32714);
or U37282 (N_37282,N_30537,N_31717);
nor U37283 (N_37283,N_33311,N_30144);
or U37284 (N_37284,N_33512,N_34572);
or U37285 (N_37285,N_33626,N_33125);
nor U37286 (N_37286,N_33121,N_33716);
nand U37287 (N_37287,N_30322,N_31877);
nand U37288 (N_37288,N_32582,N_31918);
nand U37289 (N_37289,N_30583,N_33511);
or U37290 (N_37290,N_31716,N_34851);
or U37291 (N_37291,N_31013,N_31146);
nor U37292 (N_37292,N_32673,N_34103);
nand U37293 (N_37293,N_34303,N_32801);
or U37294 (N_37294,N_34026,N_34914);
xor U37295 (N_37295,N_32569,N_32051);
or U37296 (N_37296,N_32628,N_32865);
and U37297 (N_37297,N_33772,N_30001);
and U37298 (N_37298,N_32561,N_30775);
nor U37299 (N_37299,N_32142,N_30564);
nor U37300 (N_37300,N_30456,N_31670);
and U37301 (N_37301,N_32237,N_32595);
or U37302 (N_37302,N_31517,N_32710);
and U37303 (N_37303,N_30014,N_33759);
and U37304 (N_37304,N_31400,N_30614);
or U37305 (N_37305,N_31158,N_33691);
nand U37306 (N_37306,N_32978,N_30862);
and U37307 (N_37307,N_33167,N_34862);
nor U37308 (N_37308,N_31160,N_33609);
nor U37309 (N_37309,N_32487,N_32624);
nand U37310 (N_37310,N_32153,N_33686);
nand U37311 (N_37311,N_30933,N_34298);
nand U37312 (N_37312,N_32283,N_33483);
nor U37313 (N_37313,N_31976,N_30992);
or U37314 (N_37314,N_31069,N_33722);
and U37315 (N_37315,N_34887,N_30210);
xor U37316 (N_37316,N_34492,N_31833);
or U37317 (N_37317,N_32138,N_31310);
nor U37318 (N_37318,N_34852,N_31705);
or U37319 (N_37319,N_31686,N_32437);
nor U37320 (N_37320,N_34058,N_32448);
nand U37321 (N_37321,N_34415,N_33138);
nand U37322 (N_37322,N_33236,N_31156);
nand U37323 (N_37323,N_30461,N_34576);
or U37324 (N_37324,N_34185,N_30682);
and U37325 (N_37325,N_32358,N_30826);
xnor U37326 (N_37326,N_34056,N_32917);
nor U37327 (N_37327,N_30284,N_31968);
or U37328 (N_37328,N_31046,N_33159);
and U37329 (N_37329,N_33520,N_32734);
and U37330 (N_37330,N_31690,N_34666);
or U37331 (N_37331,N_34165,N_33047);
nor U37332 (N_37332,N_30892,N_33528);
nor U37333 (N_37333,N_30278,N_30127);
or U37334 (N_37334,N_31688,N_30709);
and U37335 (N_37335,N_30656,N_30546);
nor U37336 (N_37336,N_32164,N_33496);
xor U37337 (N_37337,N_33539,N_34071);
and U37338 (N_37338,N_32885,N_34265);
nand U37339 (N_37339,N_30151,N_30469);
nor U37340 (N_37340,N_30281,N_32800);
nor U37341 (N_37341,N_32994,N_30687);
xnor U37342 (N_37342,N_32379,N_33633);
nor U37343 (N_37343,N_33834,N_30874);
nand U37344 (N_37344,N_33191,N_34846);
nand U37345 (N_37345,N_32880,N_32105);
nor U37346 (N_37346,N_31280,N_31598);
nor U37347 (N_37347,N_31314,N_30655);
nor U37348 (N_37348,N_31434,N_30183);
nor U37349 (N_37349,N_30116,N_30567);
and U37350 (N_37350,N_34343,N_34866);
xnor U37351 (N_37351,N_34346,N_31563);
or U37352 (N_37352,N_34633,N_30292);
and U37353 (N_37353,N_30945,N_31048);
nor U37354 (N_37354,N_31397,N_32395);
or U37355 (N_37355,N_32669,N_30266);
and U37356 (N_37356,N_32229,N_31124);
nand U37357 (N_37357,N_34146,N_32082);
and U37358 (N_37358,N_31107,N_32299);
and U37359 (N_37359,N_33006,N_31112);
or U37360 (N_37360,N_34040,N_33017);
and U37361 (N_37361,N_34144,N_30252);
nor U37362 (N_37362,N_34228,N_30973);
or U37363 (N_37363,N_31764,N_33198);
or U37364 (N_37364,N_30124,N_34728);
or U37365 (N_37365,N_33136,N_33022);
nand U37366 (N_37366,N_31387,N_32945);
nand U37367 (N_37367,N_30972,N_31782);
and U37368 (N_37368,N_34031,N_30887);
nor U37369 (N_37369,N_32889,N_30249);
nand U37370 (N_37370,N_34142,N_33331);
and U37371 (N_37371,N_33873,N_34748);
nand U37372 (N_37372,N_34417,N_34392);
nor U37373 (N_37373,N_34508,N_34715);
nand U37374 (N_37374,N_34302,N_31313);
or U37375 (N_37375,N_32374,N_33955);
nor U37376 (N_37376,N_34033,N_30340);
or U37377 (N_37377,N_31978,N_31606);
xor U37378 (N_37378,N_33000,N_31003);
nand U37379 (N_37379,N_31141,N_30009);
nand U37380 (N_37380,N_30443,N_31861);
and U37381 (N_37381,N_31191,N_31102);
xor U37382 (N_37382,N_33641,N_34587);
nand U37383 (N_37383,N_30595,N_31173);
and U37384 (N_37384,N_34365,N_32170);
xor U37385 (N_37385,N_32088,N_30492);
and U37386 (N_37386,N_33089,N_34767);
or U37387 (N_37387,N_34726,N_34367);
nand U37388 (N_37388,N_33291,N_31301);
nand U37389 (N_37389,N_33168,N_34984);
and U37390 (N_37390,N_31172,N_33464);
or U37391 (N_37391,N_32833,N_33769);
nand U37392 (N_37392,N_34710,N_32348);
or U37393 (N_37393,N_32352,N_32394);
or U37394 (N_37394,N_32405,N_30293);
or U37395 (N_37395,N_34828,N_32768);
xnor U37396 (N_37396,N_32675,N_32065);
and U37397 (N_37397,N_33328,N_31888);
nor U37398 (N_37398,N_33230,N_32838);
nor U37399 (N_37399,N_30468,N_34330);
nand U37400 (N_37400,N_32471,N_31324);
nor U37401 (N_37401,N_34534,N_31302);
or U37402 (N_37402,N_33829,N_34248);
nor U37403 (N_37403,N_31654,N_31151);
xnor U37404 (N_37404,N_30860,N_32868);
nor U37405 (N_37405,N_34494,N_33085);
nor U37406 (N_37406,N_33319,N_34271);
or U37407 (N_37407,N_33993,N_30714);
nor U37408 (N_37408,N_33908,N_32558);
and U37409 (N_37409,N_33707,N_30857);
nand U37410 (N_37410,N_31866,N_32326);
or U37411 (N_37411,N_33394,N_31398);
nand U37412 (N_37412,N_34580,N_32836);
nor U37413 (N_37413,N_31551,N_31269);
and U37414 (N_37414,N_30244,N_33360);
and U37415 (N_37415,N_31193,N_33992);
or U37416 (N_37416,N_34000,N_33185);
nand U37417 (N_37417,N_33969,N_30722);
and U37418 (N_37418,N_32392,N_34053);
and U37419 (N_37419,N_32384,N_33210);
xor U37420 (N_37420,N_32368,N_30191);
nand U37421 (N_37421,N_33598,N_31493);
or U37422 (N_37422,N_33619,N_31732);
nor U37423 (N_37423,N_34019,N_34720);
and U37424 (N_37424,N_30122,N_31346);
xnor U37425 (N_37425,N_33966,N_34588);
xnor U37426 (N_37426,N_33107,N_33391);
nand U37427 (N_37427,N_30602,N_34257);
and U37428 (N_37428,N_31358,N_30940);
nor U37429 (N_37429,N_32835,N_33055);
and U37430 (N_37430,N_34335,N_32625);
nand U37431 (N_37431,N_32981,N_34940);
or U37432 (N_37432,N_33904,N_32050);
nor U37433 (N_37433,N_31578,N_33042);
xor U37434 (N_37434,N_34167,N_31403);
nor U37435 (N_37435,N_31128,N_33518);
nand U37436 (N_37436,N_32902,N_33324);
xor U37437 (N_37437,N_31460,N_34267);
nand U37438 (N_37438,N_34800,N_32542);
or U37439 (N_37439,N_31725,N_30219);
nor U37440 (N_37440,N_30436,N_30426);
nand U37441 (N_37441,N_33775,N_30377);
xnor U37442 (N_37442,N_33838,N_34472);
nand U37443 (N_37443,N_31718,N_34401);
and U37444 (N_37444,N_34757,N_32466);
xnor U37445 (N_37445,N_34010,N_32464);
nor U37446 (N_37446,N_30867,N_30423);
nand U37447 (N_37447,N_34905,N_32948);
and U37448 (N_37448,N_32169,N_30092);
nand U37449 (N_37449,N_32419,N_30756);
nor U37450 (N_37450,N_33788,N_31405);
nor U37451 (N_37451,N_34125,N_34431);
nand U37452 (N_37452,N_34988,N_34068);
nor U37453 (N_37453,N_34207,N_34718);
xor U37454 (N_37454,N_34436,N_33169);
or U37455 (N_37455,N_32735,N_33172);
nand U37456 (N_37456,N_31248,N_34224);
and U37457 (N_37457,N_31770,N_30382);
and U37458 (N_37458,N_30700,N_33618);
nor U37459 (N_37459,N_32693,N_32493);
nor U37460 (N_37460,N_33717,N_32078);
and U37461 (N_37461,N_33186,N_32284);
nor U37462 (N_37462,N_31760,N_34526);
nor U37463 (N_37463,N_33217,N_32637);
and U37464 (N_37464,N_34254,N_31559);
xnor U37465 (N_37465,N_34479,N_30182);
or U37466 (N_37466,N_30951,N_34206);
nor U37467 (N_37467,N_33680,N_34120);
or U37468 (N_37468,N_31835,N_30524);
nand U37469 (N_37469,N_33009,N_34400);
and U37470 (N_37470,N_30605,N_31535);
and U37471 (N_37471,N_30821,N_30755);
nor U37472 (N_37472,N_34642,N_30928);
and U37473 (N_37473,N_31975,N_32054);
and U37474 (N_37474,N_34631,N_32862);
and U37475 (N_37475,N_32745,N_33193);
nand U37476 (N_37476,N_30136,N_33146);
nand U37477 (N_37477,N_30993,N_32974);
and U37478 (N_37478,N_34664,N_31516);
or U37479 (N_37479,N_34430,N_34774);
nor U37480 (N_37480,N_33563,N_32233);
nor U37481 (N_37481,N_31916,N_31679);
nand U37482 (N_37482,N_34324,N_30391);
nand U37483 (N_37483,N_32356,N_30802);
nor U37484 (N_37484,N_32118,N_33593);
nor U37485 (N_37485,N_31290,N_31693);
nand U37486 (N_37486,N_31851,N_31255);
nor U37487 (N_37487,N_30128,N_33702);
nand U37488 (N_37488,N_31323,N_31605);
or U37489 (N_37489,N_31486,N_34562);
xnor U37490 (N_37490,N_33624,N_33947);
and U37491 (N_37491,N_33002,N_33859);
and U37492 (N_37492,N_33340,N_31900);
or U37493 (N_37493,N_31746,N_34540);
nand U37494 (N_37494,N_30670,N_30079);
xor U37495 (N_37495,N_33863,N_30995);
or U37496 (N_37496,N_33650,N_34725);
or U37497 (N_37497,N_32008,N_31019);
xor U37498 (N_37498,N_30037,N_33073);
nand U37499 (N_37499,N_33954,N_30002);
and U37500 (N_37500,N_33875,N_34936);
xor U37501 (N_37501,N_34075,N_30662);
and U37502 (N_37502,N_32491,N_34773);
nand U37503 (N_37503,N_34775,N_30295);
and U37504 (N_37504,N_34692,N_34886);
nor U37505 (N_37505,N_31921,N_34205);
nor U37506 (N_37506,N_34646,N_33237);
or U37507 (N_37507,N_30534,N_31607);
or U37508 (N_37508,N_32841,N_32386);
nor U37509 (N_37509,N_30587,N_34321);
or U37510 (N_37510,N_30034,N_31452);
or U37511 (N_37511,N_34878,N_33500);
nand U37512 (N_37512,N_31440,N_33452);
nand U37513 (N_37513,N_30974,N_34729);
nor U37514 (N_37514,N_33594,N_31412);
nor U37515 (N_37515,N_30936,N_32630);
and U37516 (N_37516,N_33316,N_33231);
or U37517 (N_37517,N_32517,N_32101);
and U37518 (N_37518,N_34234,N_31950);
xor U37519 (N_37519,N_31050,N_34361);
and U37520 (N_37520,N_33533,N_30161);
and U37521 (N_37521,N_32495,N_33039);
nand U37522 (N_37522,N_33484,N_32820);
nor U37523 (N_37523,N_31074,N_34602);
nand U37524 (N_37524,N_31827,N_31097);
nand U37525 (N_37525,N_33127,N_30229);
xnor U37526 (N_37526,N_34599,N_31012);
nand U37527 (N_37527,N_31421,N_33235);
nor U37528 (N_37528,N_31716,N_32172);
nor U37529 (N_37529,N_31658,N_31744);
nand U37530 (N_37530,N_31422,N_30098);
and U37531 (N_37531,N_34238,N_32498);
nand U37532 (N_37532,N_30416,N_30007);
and U37533 (N_37533,N_34432,N_32908);
nand U37534 (N_37534,N_33109,N_31481);
nand U37535 (N_37535,N_33016,N_31852);
or U37536 (N_37536,N_30128,N_30326);
nand U37537 (N_37537,N_33512,N_34649);
nor U37538 (N_37538,N_32030,N_30455);
nand U37539 (N_37539,N_30468,N_33307);
nor U37540 (N_37540,N_30519,N_34027);
or U37541 (N_37541,N_32987,N_31016);
and U37542 (N_37542,N_33431,N_32224);
and U37543 (N_37543,N_30501,N_31074);
nor U37544 (N_37544,N_32850,N_30943);
nand U37545 (N_37545,N_34934,N_30018);
and U37546 (N_37546,N_33894,N_31613);
nor U37547 (N_37547,N_32966,N_33038);
or U37548 (N_37548,N_34300,N_33118);
or U37549 (N_37549,N_31283,N_32014);
or U37550 (N_37550,N_34609,N_30522);
nor U37551 (N_37551,N_32472,N_32903);
or U37552 (N_37552,N_30623,N_34830);
xor U37553 (N_37553,N_34671,N_30592);
or U37554 (N_37554,N_34092,N_32153);
nand U37555 (N_37555,N_31483,N_31552);
nor U37556 (N_37556,N_31724,N_30025);
and U37557 (N_37557,N_30388,N_34940);
nand U37558 (N_37558,N_31601,N_33138);
nor U37559 (N_37559,N_32123,N_33206);
or U37560 (N_37560,N_31109,N_34984);
and U37561 (N_37561,N_33782,N_31885);
or U37562 (N_37562,N_32766,N_33211);
or U37563 (N_37563,N_31768,N_30064);
and U37564 (N_37564,N_34238,N_34572);
nand U37565 (N_37565,N_33400,N_33208);
and U37566 (N_37566,N_34225,N_33590);
xor U37567 (N_37567,N_34903,N_30594);
nor U37568 (N_37568,N_33110,N_33441);
nor U37569 (N_37569,N_34889,N_31224);
or U37570 (N_37570,N_32318,N_34206);
nand U37571 (N_37571,N_30558,N_33762);
nor U37572 (N_37572,N_30229,N_34741);
nor U37573 (N_37573,N_32205,N_30721);
nand U37574 (N_37574,N_34665,N_32626);
and U37575 (N_37575,N_31121,N_34827);
and U37576 (N_37576,N_30229,N_31350);
or U37577 (N_37577,N_30832,N_30104);
nor U37578 (N_37578,N_33483,N_34361);
nand U37579 (N_37579,N_33375,N_34519);
nand U37580 (N_37580,N_33820,N_31198);
nand U37581 (N_37581,N_32663,N_32513);
and U37582 (N_37582,N_31290,N_33587);
or U37583 (N_37583,N_32033,N_33400);
and U37584 (N_37584,N_34744,N_33123);
nor U37585 (N_37585,N_30642,N_34382);
and U37586 (N_37586,N_30461,N_32985);
or U37587 (N_37587,N_33233,N_33100);
nand U37588 (N_37588,N_30124,N_34315);
and U37589 (N_37589,N_34105,N_33944);
or U37590 (N_37590,N_32288,N_33178);
or U37591 (N_37591,N_31344,N_33027);
nand U37592 (N_37592,N_30817,N_30513);
nand U37593 (N_37593,N_31671,N_33535);
nor U37594 (N_37594,N_34536,N_32002);
nor U37595 (N_37595,N_32490,N_31553);
and U37596 (N_37596,N_34146,N_30797);
nand U37597 (N_37597,N_34196,N_33871);
nand U37598 (N_37598,N_30762,N_31789);
nand U37599 (N_37599,N_33469,N_34985);
and U37600 (N_37600,N_33465,N_33372);
nor U37601 (N_37601,N_34839,N_34803);
or U37602 (N_37602,N_32360,N_32869);
or U37603 (N_37603,N_32366,N_33475);
nand U37604 (N_37604,N_31689,N_31678);
nor U37605 (N_37605,N_32604,N_32584);
and U37606 (N_37606,N_33524,N_32787);
or U37607 (N_37607,N_33299,N_32396);
nand U37608 (N_37608,N_33830,N_33821);
and U37609 (N_37609,N_33005,N_32209);
and U37610 (N_37610,N_31155,N_33823);
nand U37611 (N_37611,N_33666,N_30158);
xor U37612 (N_37612,N_34096,N_31269);
nor U37613 (N_37613,N_30365,N_30185);
nand U37614 (N_37614,N_30728,N_33587);
and U37615 (N_37615,N_31292,N_30324);
or U37616 (N_37616,N_34180,N_34377);
nand U37617 (N_37617,N_34085,N_31200);
nor U37618 (N_37618,N_32831,N_34668);
or U37619 (N_37619,N_33883,N_30542);
nor U37620 (N_37620,N_30974,N_31201);
nor U37621 (N_37621,N_33038,N_34921);
or U37622 (N_37622,N_34260,N_33990);
and U37623 (N_37623,N_32140,N_30504);
xor U37624 (N_37624,N_33754,N_34763);
nor U37625 (N_37625,N_32563,N_32490);
or U37626 (N_37626,N_31808,N_30122);
nor U37627 (N_37627,N_30667,N_33692);
or U37628 (N_37628,N_30104,N_34645);
or U37629 (N_37629,N_33976,N_32602);
nand U37630 (N_37630,N_30928,N_31880);
and U37631 (N_37631,N_31470,N_32038);
or U37632 (N_37632,N_32336,N_31563);
nor U37633 (N_37633,N_33704,N_33393);
nor U37634 (N_37634,N_31760,N_34303);
nor U37635 (N_37635,N_30832,N_30582);
nand U37636 (N_37636,N_33067,N_33400);
nand U37637 (N_37637,N_31439,N_34483);
nor U37638 (N_37638,N_31278,N_30554);
or U37639 (N_37639,N_33783,N_31011);
nor U37640 (N_37640,N_30220,N_33014);
or U37641 (N_37641,N_34956,N_32622);
nor U37642 (N_37642,N_31297,N_33324);
nand U37643 (N_37643,N_30709,N_32011);
or U37644 (N_37644,N_30048,N_33752);
or U37645 (N_37645,N_30908,N_30524);
or U37646 (N_37646,N_31589,N_32546);
and U37647 (N_37647,N_33624,N_30291);
nand U37648 (N_37648,N_33118,N_34110);
or U37649 (N_37649,N_31766,N_31862);
nand U37650 (N_37650,N_34176,N_31485);
and U37651 (N_37651,N_34107,N_30314);
nor U37652 (N_37652,N_34228,N_33959);
xor U37653 (N_37653,N_33733,N_33997);
or U37654 (N_37654,N_31184,N_30771);
and U37655 (N_37655,N_31761,N_30147);
nand U37656 (N_37656,N_34475,N_33688);
or U37657 (N_37657,N_34704,N_31190);
or U37658 (N_37658,N_30975,N_33211);
and U37659 (N_37659,N_34888,N_30827);
nor U37660 (N_37660,N_32010,N_34819);
xnor U37661 (N_37661,N_30773,N_33108);
nand U37662 (N_37662,N_30204,N_30381);
nor U37663 (N_37663,N_31263,N_32815);
nor U37664 (N_37664,N_30215,N_31525);
xnor U37665 (N_37665,N_30231,N_30279);
or U37666 (N_37666,N_31478,N_33649);
nor U37667 (N_37667,N_30267,N_32217);
nor U37668 (N_37668,N_33506,N_31906);
or U37669 (N_37669,N_32740,N_33534);
and U37670 (N_37670,N_31869,N_31085);
or U37671 (N_37671,N_30264,N_32402);
nand U37672 (N_37672,N_34533,N_34466);
nand U37673 (N_37673,N_32911,N_34116);
and U37674 (N_37674,N_33401,N_31932);
nor U37675 (N_37675,N_32409,N_34286);
and U37676 (N_37676,N_32683,N_34481);
or U37677 (N_37677,N_32373,N_32301);
nor U37678 (N_37678,N_34847,N_34606);
and U37679 (N_37679,N_33062,N_33371);
or U37680 (N_37680,N_30341,N_33450);
nor U37681 (N_37681,N_30785,N_33828);
nor U37682 (N_37682,N_33541,N_30898);
nor U37683 (N_37683,N_30500,N_34846);
nand U37684 (N_37684,N_33243,N_32774);
or U37685 (N_37685,N_30405,N_32948);
or U37686 (N_37686,N_33935,N_32127);
and U37687 (N_37687,N_30530,N_30527);
nand U37688 (N_37688,N_33504,N_30965);
nor U37689 (N_37689,N_31958,N_30226);
or U37690 (N_37690,N_34778,N_34623);
nand U37691 (N_37691,N_31175,N_33141);
nor U37692 (N_37692,N_31647,N_31357);
xor U37693 (N_37693,N_34188,N_34759);
xnor U37694 (N_37694,N_33397,N_33790);
nor U37695 (N_37695,N_34965,N_33477);
or U37696 (N_37696,N_31725,N_34015);
nand U37697 (N_37697,N_31724,N_34673);
and U37698 (N_37698,N_34512,N_31250);
or U37699 (N_37699,N_30557,N_30822);
or U37700 (N_37700,N_30145,N_34659);
nand U37701 (N_37701,N_30209,N_30792);
or U37702 (N_37702,N_30151,N_31751);
nand U37703 (N_37703,N_33794,N_34016);
nand U37704 (N_37704,N_31130,N_33706);
nor U37705 (N_37705,N_31758,N_33763);
nor U37706 (N_37706,N_32419,N_31763);
nand U37707 (N_37707,N_33860,N_32044);
or U37708 (N_37708,N_33547,N_31590);
xor U37709 (N_37709,N_32758,N_33799);
nor U37710 (N_37710,N_31373,N_34698);
xor U37711 (N_37711,N_30779,N_33316);
xor U37712 (N_37712,N_33981,N_31374);
nor U37713 (N_37713,N_32682,N_34029);
xnor U37714 (N_37714,N_30189,N_30366);
nor U37715 (N_37715,N_31144,N_30991);
xnor U37716 (N_37716,N_32939,N_31948);
nand U37717 (N_37717,N_34622,N_32819);
and U37718 (N_37718,N_33364,N_34925);
nand U37719 (N_37719,N_30786,N_31930);
nand U37720 (N_37720,N_30399,N_34548);
nand U37721 (N_37721,N_31246,N_32628);
or U37722 (N_37722,N_33525,N_31389);
or U37723 (N_37723,N_34560,N_30474);
nand U37724 (N_37724,N_33316,N_32383);
nand U37725 (N_37725,N_30234,N_32799);
and U37726 (N_37726,N_30076,N_32176);
or U37727 (N_37727,N_30841,N_33673);
nor U37728 (N_37728,N_30121,N_31644);
and U37729 (N_37729,N_30236,N_31885);
nand U37730 (N_37730,N_33580,N_30918);
and U37731 (N_37731,N_31618,N_33807);
or U37732 (N_37732,N_33449,N_34481);
and U37733 (N_37733,N_30557,N_31579);
nand U37734 (N_37734,N_30595,N_34089);
and U37735 (N_37735,N_32445,N_34785);
nand U37736 (N_37736,N_31767,N_31204);
xnor U37737 (N_37737,N_32745,N_32285);
and U37738 (N_37738,N_30670,N_32120);
nor U37739 (N_37739,N_34712,N_31359);
xor U37740 (N_37740,N_33593,N_32246);
nor U37741 (N_37741,N_34398,N_32975);
or U37742 (N_37742,N_31766,N_30991);
and U37743 (N_37743,N_32413,N_31316);
nand U37744 (N_37744,N_34826,N_33832);
or U37745 (N_37745,N_31715,N_30766);
nor U37746 (N_37746,N_30057,N_30879);
xor U37747 (N_37747,N_33881,N_32654);
or U37748 (N_37748,N_30553,N_32361);
and U37749 (N_37749,N_31174,N_30017);
nor U37750 (N_37750,N_30628,N_31201);
nand U37751 (N_37751,N_30535,N_32663);
and U37752 (N_37752,N_31905,N_33422);
nand U37753 (N_37753,N_34748,N_34485);
and U37754 (N_37754,N_30023,N_33082);
nand U37755 (N_37755,N_34385,N_32606);
nor U37756 (N_37756,N_32548,N_30423);
and U37757 (N_37757,N_30550,N_32002);
nor U37758 (N_37758,N_32938,N_30917);
nand U37759 (N_37759,N_34209,N_30386);
and U37760 (N_37760,N_30371,N_30109);
and U37761 (N_37761,N_34362,N_32750);
nand U37762 (N_37762,N_32999,N_34414);
nand U37763 (N_37763,N_33306,N_34522);
and U37764 (N_37764,N_31864,N_31408);
and U37765 (N_37765,N_32413,N_31391);
and U37766 (N_37766,N_31883,N_33799);
and U37767 (N_37767,N_31645,N_30980);
and U37768 (N_37768,N_33233,N_30981);
or U37769 (N_37769,N_34876,N_34237);
and U37770 (N_37770,N_34350,N_31761);
and U37771 (N_37771,N_31985,N_31399);
and U37772 (N_37772,N_30543,N_30054);
and U37773 (N_37773,N_31488,N_33206);
and U37774 (N_37774,N_34215,N_30940);
xor U37775 (N_37775,N_31474,N_34839);
or U37776 (N_37776,N_30412,N_34089);
or U37777 (N_37777,N_33533,N_33140);
nand U37778 (N_37778,N_33969,N_32359);
and U37779 (N_37779,N_34698,N_34826);
nor U37780 (N_37780,N_33949,N_31445);
and U37781 (N_37781,N_31134,N_30850);
nand U37782 (N_37782,N_30273,N_32471);
xnor U37783 (N_37783,N_34354,N_34375);
nor U37784 (N_37784,N_31480,N_32975);
or U37785 (N_37785,N_30334,N_32456);
nand U37786 (N_37786,N_30178,N_33275);
or U37787 (N_37787,N_34928,N_32484);
and U37788 (N_37788,N_34562,N_34195);
or U37789 (N_37789,N_33472,N_34995);
or U37790 (N_37790,N_33803,N_30591);
nor U37791 (N_37791,N_34552,N_34566);
and U37792 (N_37792,N_32857,N_34285);
nand U37793 (N_37793,N_30781,N_32979);
and U37794 (N_37794,N_31120,N_31026);
xor U37795 (N_37795,N_34625,N_33284);
nand U37796 (N_37796,N_34444,N_32190);
or U37797 (N_37797,N_31581,N_33498);
or U37798 (N_37798,N_31512,N_34869);
nand U37799 (N_37799,N_33299,N_33320);
nor U37800 (N_37800,N_30624,N_31135);
xor U37801 (N_37801,N_30135,N_32253);
nor U37802 (N_37802,N_30069,N_33485);
or U37803 (N_37803,N_31701,N_32099);
or U37804 (N_37804,N_33312,N_31278);
nor U37805 (N_37805,N_32253,N_30618);
or U37806 (N_37806,N_32345,N_32647);
nand U37807 (N_37807,N_34316,N_32180);
nand U37808 (N_37808,N_31519,N_31230);
and U37809 (N_37809,N_34128,N_30397);
and U37810 (N_37810,N_34698,N_32234);
nor U37811 (N_37811,N_30183,N_34109);
or U37812 (N_37812,N_32087,N_34627);
and U37813 (N_37813,N_33458,N_30074);
xnor U37814 (N_37814,N_31367,N_30228);
and U37815 (N_37815,N_34367,N_31342);
and U37816 (N_37816,N_34188,N_32781);
xor U37817 (N_37817,N_34322,N_34263);
nand U37818 (N_37818,N_30893,N_34890);
and U37819 (N_37819,N_31575,N_31129);
or U37820 (N_37820,N_31181,N_32474);
nor U37821 (N_37821,N_34057,N_31574);
and U37822 (N_37822,N_33021,N_31760);
or U37823 (N_37823,N_31371,N_34628);
nor U37824 (N_37824,N_31123,N_32285);
nand U37825 (N_37825,N_30847,N_34776);
nor U37826 (N_37826,N_30085,N_31615);
or U37827 (N_37827,N_33042,N_30831);
and U37828 (N_37828,N_34706,N_33673);
and U37829 (N_37829,N_30530,N_32263);
or U37830 (N_37830,N_34430,N_34608);
nor U37831 (N_37831,N_34580,N_32970);
nor U37832 (N_37832,N_34764,N_32283);
or U37833 (N_37833,N_31976,N_31847);
nand U37834 (N_37834,N_30319,N_30949);
and U37835 (N_37835,N_33130,N_30966);
nor U37836 (N_37836,N_30428,N_32878);
nand U37837 (N_37837,N_30980,N_30315);
nor U37838 (N_37838,N_32411,N_31819);
nor U37839 (N_37839,N_33284,N_33402);
nand U37840 (N_37840,N_32434,N_31075);
nor U37841 (N_37841,N_32763,N_33192);
nor U37842 (N_37842,N_34188,N_31825);
nand U37843 (N_37843,N_30036,N_31440);
nor U37844 (N_37844,N_32833,N_34212);
nand U37845 (N_37845,N_31008,N_34108);
xor U37846 (N_37846,N_30820,N_34274);
and U37847 (N_37847,N_34694,N_30006);
and U37848 (N_37848,N_31212,N_30259);
nand U37849 (N_37849,N_32291,N_33497);
or U37850 (N_37850,N_30300,N_32927);
or U37851 (N_37851,N_32090,N_30904);
or U37852 (N_37852,N_34111,N_33049);
xnor U37853 (N_37853,N_32392,N_32680);
and U37854 (N_37854,N_33050,N_33226);
nor U37855 (N_37855,N_31333,N_31401);
and U37856 (N_37856,N_32161,N_30079);
or U37857 (N_37857,N_34394,N_31382);
nor U37858 (N_37858,N_30633,N_34546);
and U37859 (N_37859,N_33534,N_31824);
nor U37860 (N_37860,N_30591,N_32428);
nand U37861 (N_37861,N_32853,N_34614);
nand U37862 (N_37862,N_31741,N_31245);
xor U37863 (N_37863,N_34603,N_30903);
or U37864 (N_37864,N_31825,N_32087);
and U37865 (N_37865,N_30452,N_33892);
nand U37866 (N_37866,N_33275,N_31128);
and U37867 (N_37867,N_31185,N_33376);
xor U37868 (N_37868,N_31896,N_30499);
and U37869 (N_37869,N_33332,N_34467);
xor U37870 (N_37870,N_32242,N_32689);
xor U37871 (N_37871,N_33792,N_33401);
and U37872 (N_37872,N_34508,N_32152);
and U37873 (N_37873,N_33188,N_30885);
nand U37874 (N_37874,N_30366,N_32684);
nor U37875 (N_37875,N_33344,N_30457);
or U37876 (N_37876,N_33251,N_31138);
nor U37877 (N_37877,N_31876,N_31960);
nand U37878 (N_37878,N_33299,N_30489);
nand U37879 (N_37879,N_34536,N_33176);
nand U37880 (N_37880,N_33197,N_30826);
xnor U37881 (N_37881,N_33465,N_32940);
and U37882 (N_37882,N_34878,N_33142);
or U37883 (N_37883,N_33336,N_33217);
and U37884 (N_37884,N_33540,N_31416);
and U37885 (N_37885,N_33016,N_34806);
nand U37886 (N_37886,N_31035,N_34515);
and U37887 (N_37887,N_34723,N_32511);
or U37888 (N_37888,N_30959,N_33619);
and U37889 (N_37889,N_33135,N_34911);
nand U37890 (N_37890,N_30349,N_33812);
and U37891 (N_37891,N_32442,N_32057);
and U37892 (N_37892,N_31091,N_33382);
xor U37893 (N_37893,N_33110,N_32529);
nor U37894 (N_37894,N_32871,N_34652);
and U37895 (N_37895,N_34311,N_31711);
and U37896 (N_37896,N_32321,N_30506);
or U37897 (N_37897,N_32451,N_32372);
or U37898 (N_37898,N_32182,N_32575);
nor U37899 (N_37899,N_32003,N_32612);
and U37900 (N_37900,N_30893,N_34465);
or U37901 (N_37901,N_34994,N_32316);
or U37902 (N_37902,N_32387,N_30828);
xor U37903 (N_37903,N_30998,N_33124);
nand U37904 (N_37904,N_30601,N_32200);
xor U37905 (N_37905,N_34185,N_34275);
or U37906 (N_37906,N_33693,N_34826);
nor U37907 (N_37907,N_32001,N_30946);
and U37908 (N_37908,N_31761,N_30196);
and U37909 (N_37909,N_30135,N_33022);
and U37910 (N_37910,N_31932,N_34715);
nand U37911 (N_37911,N_34342,N_32897);
and U37912 (N_37912,N_33242,N_32737);
nand U37913 (N_37913,N_32466,N_30906);
nor U37914 (N_37914,N_32206,N_32048);
xnor U37915 (N_37915,N_32597,N_32940);
and U37916 (N_37916,N_31606,N_30554);
nand U37917 (N_37917,N_32085,N_30099);
or U37918 (N_37918,N_32272,N_32877);
and U37919 (N_37919,N_31690,N_31862);
nand U37920 (N_37920,N_30499,N_31800);
nor U37921 (N_37921,N_30514,N_33968);
xnor U37922 (N_37922,N_34806,N_34366);
or U37923 (N_37923,N_31467,N_34564);
nand U37924 (N_37924,N_32820,N_33933);
and U37925 (N_37925,N_31665,N_30720);
or U37926 (N_37926,N_31697,N_30680);
nand U37927 (N_37927,N_32055,N_32597);
nand U37928 (N_37928,N_31914,N_34897);
and U37929 (N_37929,N_31943,N_32613);
and U37930 (N_37930,N_33622,N_34898);
and U37931 (N_37931,N_30663,N_34617);
and U37932 (N_37932,N_32714,N_32266);
xnor U37933 (N_37933,N_34816,N_33068);
nor U37934 (N_37934,N_30369,N_31645);
nor U37935 (N_37935,N_34238,N_33029);
nand U37936 (N_37936,N_33404,N_33003);
and U37937 (N_37937,N_34464,N_32664);
and U37938 (N_37938,N_32491,N_32639);
xnor U37939 (N_37939,N_31728,N_31903);
nor U37940 (N_37940,N_33410,N_31133);
nor U37941 (N_37941,N_31703,N_30582);
xor U37942 (N_37942,N_32378,N_34709);
nor U37943 (N_37943,N_30203,N_34497);
or U37944 (N_37944,N_33041,N_30917);
or U37945 (N_37945,N_30148,N_32626);
or U37946 (N_37946,N_30830,N_33309);
or U37947 (N_37947,N_30585,N_34900);
or U37948 (N_37948,N_32937,N_34827);
and U37949 (N_37949,N_34288,N_33208);
nor U37950 (N_37950,N_31173,N_34880);
and U37951 (N_37951,N_33077,N_30141);
nand U37952 (N_37952,N_30784,N_34499);
and U37953 (N_37953,N_34698,N_31976);
nand U37954 (N_37954,N_32211,N_33716);
xor U37955 (N_37955,N_30866,N_33413);
nor U37956 (N_37956,N_32423,N_33329);
nand U37957 (N_37957,N_33929,N_34689);
xnor U37958 (N_37958,N_32682,N_31848);
nand U37959 (N_37959,N_32795,N_31083);
nor U37960 (N_37960,N_32497,N_34747);
nor U37961 (N_37961,N_30174,N_31379);
or U37962 (N_37962,N_33110,N_31187);
and U37963 (N_37963,N_30928,N_32904);
nor U37964 (N_37964,N_33208,N_33272);
or U37965 (N_37965,N_34593,N_32858);
and U37966 (N_37966,N_33189,N_31680);
xnor U37967 (N_37967,N_33230,N_34087);
or U37968 (N_37968,N_30721,N_30976);
or U37969 (N_37969,N_31964,N_32389);
and U37970 (N_37970,N_32571,N_32574);
nor U37971 (N_37971,N_31647,N_34084);
or U37972 (N_37972,N_32148,N_30521);
nand U37973 (N_37973,N_30275,N_30609);
and U37974 (N_37974,N_33440,N_34558);
and U37975 (N_37975,N_33422,N_34532);
or U37976 (N_37976,N_32447,N_31771);
xnor U37977 (N_37977,N_32486,N_31028);
nor U37978 (N_37978,N_33828,N_31173);
and U37979 (N_37979,N_32134,N_34606);
or U37980 (N_37980,N_34847,N_30727);
nand U37981 (N_37981,N_34783,N_34142);
nor U37982 (N_37982,N_30549,N_33407);
xnor U37983 (N_37983,N_31120,N_31209);
nand U37984 (N_37984,N_33179,N_34316);
or U37985 (N_37985,N_34575,N_31272);
and U37986 (N_37986,N_30612,N_31941);
and U37987 (N_37987,N_30332,N_32205);
xor U37988 (N_37988,N_30787,N_32107);
nand U37989 (N_37989,N_33627,N_32274);
and U37990 (N_37990,N_30558,N_33091);
or U37991 (N_37991,N_33144,N_30426);
nor U37992 (N_37992,N_30283,N_34922);
nand U37993 (N_37993,N_34285,N_30554);
nor U37994 (N_37994,N_30557,N_31751);
or U37995 (N_37995,N_30733,N_32546);
nand U37996 (N_37996,N_34553,N_32215);
nor U37997 (N_37997,N_33386,N_33744);
nor U37998 (N_37998,N_31764,N_34443);
or U37999 (N_37999,N_34055,N_30372);
nand U38000 (N_38000,N_30097,N_34703);
nand U38001 (N_38001,N_30392,N_32235);
nand U38002 (N_38002,N_32462,N_33863);
or U38003 (N_38003,N_33083,N_33443);
or U38004 (N_38004,N_32973,N_34226);
nand U38005 (N_38005,N_33552,N_30995);
and U38006 (N_38006,N_33771,N_33095);
xor U38007 (N_38007,N_34292,N_33429);
or U38008 (N_38008,N_32594,N_32283);
nand U38009 (N_38009,N_30783,N_31894);
nand U38010 (N_38010,N_34392,N_34708);
nor U38011 (N_38011,N_34869,N_32818);
nor U38012 (N_38012,N_34587,N_34432);
nand U38013 (N_38013,N_34639,N_30644);
or U38014 (N_38014,N_32879,N_34388);
nor U38015 (N_38015,N_31491,N_31177);
nor U38016 (N_38016,N_31217,N_31240);
nor U38017 (N_38017,N_31977,N_30164);
nor U38018 (N_38018,N_31272,N_34692);
and U38019 (N_38019,N_31052,N_31160);
or U38020 (N_38020,N_34994,N_32027);
xor U38021 (N_38021,N_32013,N_33892);
nor U38022 (N_38022,N_31922,N_34375);
nor U38023 (N_38023,N_30401,N_30327);
nor U38024 (N_38024,N_34301,N_34560);
nor U38025 (N_38025,N_32802,N_31214);
and U38026 (N_38026,N_31231,N_31500);
nand U38027 (N_38027,N_31806,N_34073);
or U38028 (N_38028,N_33971,N_32710);
and U38029 (N_38029,N_31302,N_30926);
nor U38030 (N_38030,N_33843,N_32985);
nor U38031 (N_38031,N_30408,N_30108);
nor U38032 (N_38032,N_33873,N_33466);
xor U38033 (N_38033,N_31287,N_32725);
and U38034 (N_38034,N_34818,N_32933);
nand U38035 (N_38035,N_34142,N_33484);
or U38036 (N_38036,N_31998,N_32993);
nor U38037 (N_38037,N_34960,N_33121);
or U38038 (N_38038,N_33368,N_30753);
or U38039 (N_38039,N_34386,N_34152);
nor U38040 (N_38040,N_34514,N_31222);
xnor U38041 (N_38041,N_33718,N_32100);
xnor U38042 (N_38042,N_33958,N_30565);
or U38043 (N_38043,N_33280,N_30682);
nor U38044 (N_38044,N_30447,N_31507);
xor U38045 (N_38045,N_31199,N_34653);
nand U38046 (N_38046,N_34318,N_32122);
nor U38047 (N_38047,N_34594,N_30907);
nor U38048 (N_38048,N_30376,N_30479);
xnor U38049 (N_38049,N_30484,N_33119);
nor U38050 (N_38050,N_32133,N_30162);
nor U38051 (N_38051,N_33832,N_30169);
nand U38052 (N_38052,N_34723,N_34067);
xor U38053 (N_38053,N_34908,N_34318);
nor U38054 (N_38054,N_31750,N_31280);
nand U38055 (N_38055,N_32398,N_34862);
or U38056 (N_38056,N_30699,N_34237);
nand U38057 (N_38057,N_32941,N_32677);
nand U38058 (N_38058,N_30734,N_32028);
nand U38059 (N_38059,N_33398,N_34759);
nor U38060 (N_38060,N_31922,N_33810);
or U38061 (N_38061,N_34988,N_34646);
or U38062 (N_38062,N_32628,N_33916);
nand U38063 (N_38063,N_33387,N_32628);
and U38064 (N_38064,N_31862,N_32658);
or U38065 (N_38065,N_31153,N_34134);
and U38066 (N_38066,N_33680,N_32803);
or U38067 (N_38067,N_32395,N_31460);
nand U38068 (N_38068,N_32471,N_30952);
and U38069 (N_38069,N_33412,N_33980);
nand U38070 (N_38070,N_32247,N_32262);
nand U38071 (N_38071,N_34420,N_33044);
nand U38072 (N_38072,N_33880,N_30310);
nand U38073 (N_38073,N_32946,N_34570);
or U38074 (N_38074,N_33646,N_32766);
nor U38075 (N_38075,N_32968,N_30623);
xor U38076 (N_38076,N_34629,N_31882);
xor U38077 (N_38077,N_33187,N_34624);
or U38078 (N_38078,N_33661,N_33294);
or U38079 (N_38079,N_34227,N_30527);
and U38080 (N_38080,N_31496,N_30377);
xor U38081 (N_38081,N_34220,N_34739);
or U38082 (N_38082,N_30284,N_30682);
or U38083 (N_38083,N_31828,N_32220);
nand U38084 (N_38084,N_34094,N_33776);
or U38085 (N_38085,N_32560,N_31479);
and U38086 (N_38086,N_32879,N_31472);
and U38087 (N_38087,N_30403,N_30274);
and U38088 (N_38088,N_32524,N_32108);
or U38089 (N_38089,N_33213,N_30550);
nor U38090 (N_38090,N_30845,N_33248);
nor U38091 (N_38091,N_30525,N_32791);
nor U38092 (N_38092,N_34788,N_30526);
or U38093 (N_38093,N_31086,N_33614);
xnor U38094 (N_38094,N_32967,N_34564);
and U38095 (N_38095,N_33808,N_33999);
nor U38096 (N_38096,N_30267,N_30031);
xnor U38097 (N_38097,N_30573,N_33875);
nand U38098 (N_38098,N_32898,N_34885);
or U38099 (N_38099,N_32094,N_30349);
nand U38100 (N_38100,N_32933,N_31827);
nand U38101 (N_38101,N_33430,N_32889);
nand U38102 (N_38102,N_33146,N_34744);
nand U38103 (N_38103,N_30670,N_31232);
and U38104 (N_38104,N_33873,N_30919);
nor U38105 (N_38105,N_33375,N_30627);
xor U38106 (N_38106,N_34173,N_31579);
and U38107 (N_38107,N_34656,N_32342);
nand U38108 (N_38108,N_31133,N_30970);
nor U38109 (N_38109,N_30566,N_34530);
or U38110 (N_38110,N_30399,N_33555);
nor U38111 (N_38111,N_31257,N_31149);
nand U38112 (N_38112,N_32982,N_30300);
nor U38113 (N_38113,N_31978,N_31118);
nor U38114 (N_38114,N_31802,N_34949);
and U38115 (N_38115,N_33319,N_33989);
or U38116 (N_38116,N_30832,N_33550);
or U38117 (N_38117,N_33789,N_34371);
and U38118 (N_38118,N_33658,N_34358);
nand U38119 (N_38119,N_32772,N_33325);
xor U38120 (N_38120,N_33648,N_31504);
and U38121 (N_38121,N_31301,N_31895);
or U38122 (N_38122,N_34132,N_34769);
nand U38123 (N_38123,N_30334,N_32124);
or U38124 (N_38124,N_34567,N_32002);
or U38125 (N_38125,N_34045,N_31246);
or U38126 (N_38126,N_33355,N_34903);
xor U38127 (N_38127,N_32384,N_31488);
or U38128 (N_38128,N_31621,N_32520);
nand U38129 (N_38129,N_31888,N_32604);
xor U38130 (N_38130,N_31127,N_34300);
xnor U38131 (N_38131,N_31336,N_30095);
and U38132 (N_38132,N_31647,N_33334);
nor U38133 (N_38133,N_31920,N_32646);
nand U38134 (N_38134,N_30914,N_33202);
or U38135 (N_38135,N_30743,N_32799);
and U38136 (N_38136,N_30419,N_33621);
and U38137 (N_38137,N_31721,N_33024);
nor U38138 (N_38138,N_32113,N_30099);
or U38139 (N_38139,N_32545,N_31832);
and U38140 (N_38140,N_30295,N_34981);
or U38141 (N_38141,N_31854,N_33731);
xnor U38142 (N_38142,N_32077,N_33810);
nand U38143 (N_38143,N_33698,N_31925);
nand U38144 (N_38144,N_32163,N_32326);
nor U38145 (N_38145,N_31029,N_32177);
nand U38146 (N_38146,N_32251,N_32258);
or U38147 (N_38147,N_34795,N_30935);
nand U38148 (N_38148,N_31066,N_32099);
nor U38149 (N_38149,N_30899,N_33287);
or U38150 (N_38150,N_33264,N_32645);
nand U38151 (N_38151,N_34195,N_34799);
and U38152 (N_38152,N_33990,N_32476);
nand U38153 (N_38153,N_32343,N_32724);
or U38154 (N_38154,N_30182,N_32776);
and U38155 (N_38155,N_32419,N_31792);
nor U38156 (N_38156,N_32244,N_33298);
nand U38157 (N_38157,N_32104,N_31732);
and U38158 (N_38158,N_33199,N_31285);
or U38159 (N_38159,N_34582,N_34341);
nand U38160 (N_38160,N_31321,N_32728);
and U38161 (N_38161,N_34113,N_34802);
nor U38162 (N_38162,N_31708,N_34468);
xor U38163 (N_38163,N_30392,N_32510);
or U38164 (N_38164,N_32079,N_32635);
xnor U38165 (N_38165,N_32212,N_32215);
or U38166 (N_38166,N_32414,N_33495);
nand U38167 (N_38167,N_33799,N_31581);
nand U38168 (N_38168,N_33262,N_30887);
nor U38169 (N_38169,N_33160,N_30120);
nand U38170 (N_38170,N_34328,N_31960);
and U38171 (N_38171,N_34065,N_32466);
nand U38172 (N_38172,N_34579,N_33246);
nor U38173 (N_38173,N_32228,N_33696);
or U38174 (N_38174,N_33700,N_30088);
nand U38175 (N_38175,N_32408,N_33835);
or U38176 (N_38176,N_33112,N_31902);
nand U38177 (N_38177,N_31400,N_33008);
or U38178 (N_38178,N_32965,N_32411);
nand U38179 (N_38179,N_31170,N_34265);
nand U38180 (N_38180,N_31288,N_32797);
xor U38181 (N_38181,N_32243,N_31643);
nor U38182 (N_38182,N_34686,N_30572);
and U38183 (N_38183,N_31679,N_32593);
or U38184 (N_38184,N_33223,N_30782);
nand U38185 (N_38185,N_32885,N_32832);
or U38186 (N_38186,N_30794,N_32704);
and U38187 (N_38187,N_34174,N_34410);
nand U38188 (N_38188,N_31132,N_30475);
or U38189 (N_38189,N_32923,N_32167);
nor U38190 (N_38190,N_32365,N_33579);
nand U38191 (N_38191,N_30415,N_33672);
xor U38192 (N_38192,N_30262,N_34189);
and U38193 (N_38193,N_31958,N_32835);
nor U38194 (N_38194,N_33535,N_32698);
or U38195 (N_38195,N_34656,N_31261);
and U38196 (N_38196,N_32083,N_32155);
and U38197 (N_38197,N_31317,N_34318);
xnor U38198 (N_38198,N_33533,N_32384);
xnor U38199 (N_38199,N_34214,N_34024);
nand U38200 (N_38200,N_34676,N_33967);
and U38201 (N_38201,N_32294,N_30466);
xor U38202 (N_38202,N_34173,N_33805);
or U38203 (N_38203,N_30535,N_31262);
or U38204 (N_38204,N_33358,N_33093);
nand U38205 (N_38205,N_31590,N_31013);
nand U38206 (N_38206,N_34026,N_30516);
nor U38207 (N_38207,N_32552,N_30754);
nor U38208 (N_38208,N_31048,N_34848);
nor U38209 (N_38209,N_34552,N_30843);
nor U38210 (N_38210,N_34362,N_34248);
nand U38211 (N_38211,N_34279,N_31650);
or U38212 (N_38212,N_30978,N_34266);
nor U38213 (N_38213,N_31440,N_32773);
nor U38214 (N_38214,N_32450,N_31306);
nor U38215 (N_38215,N_32316,N_31955);
nor U38216 (N_38216,N_32245,N_30990);
nor U38217 (N_38217,N_32064,N_30100);
nor U38218 (N_38218,N_33568,N_31178);
or U38219 (N_38219,N_31014,N_34421);
nor U38220 (N_38220,N_32332,N_30581);
nor U38221 (N_38221,N_30165,N_32377);
nand U38222 (N_38222,N_31194,N_33557);
nor U38223 (N_38223,N_32241,N_34730);
and U38224 (N_38224,N_32057,N_30776);
nand U38225 (N_38225,N_33306,N_34821);
or U38226 (N_38226,N_31108,N_31355);
or U38227 (N_38227,N_32040,N_32097);
xor U38228 (N_38228,N_32587,N_34321);
xor U38229 (N_38229,N_30150,N_32852);
nand U38230 (N_38230,N_31542,N_34958);
nor U38231 (N_38231,N_32100,N_34427);
or U38232 (N_38232,N_32957,N_30123);
nand U38233 (N_38233,N_34285,N_34770);
nor U38234 (N_38234,N_31729,N_32545);
and U38235 (N_38235,N_30626,N_32833);
or U38236 (N_38236,N_33800,N_34642);
nor U38237 (N_38237,N_32379,N_30080);
nand U38238 (N_38238,N_34295,N_33512);
or U38239 (N_38239,N_31621,N_30372);
nor U38240 (N_38240,N_31986,N_31966);
nor U38241 (N_38241,N_31415,N_32034);
xnor U38242 (N_38242,N_34342,N_32295);
and U38243 (N_38243,N_30073,N_30049);
or U38244 (N_38244,N_31530,N_31764);
nand U38245 (N_38245,N_32724,N_30486);
nand U38246 (N_38246,N_31693,N_32601);
or U38247 (N_38247,N_34095,N_32217);
nor U38248 (N_38248,N_30637,N_34746);
and U38249 (N_38249,N_33696,N_32726);
xnor U38250 (N_38250,N_30789,N_30179);
nor U38251 (N_38251,N_33330,N_31111);
and U38252 (N_38252,N_34419,N_31433);
or U38253 (N_38253,N_34535,N_33703);
nand U38254 (N_38254,N_33958,N_33892);
nand U38255 (N_38255,N_32731,N_33080);
or U38256 (N_38256,N_33693,N_33824);
nor U38257 (N_38257,N_32635,N_30966);
and U38258 (N_38258,N_31609,N_31868);
nand U38259 (N_38259,N_30487,N_34281);
or U38260 (N_38260,N_34116,N_30883);
or U38261 (N_38261,N_32143,N_32932);
and U38262 (N_38262,N_30739,N_34488);
or U38263 (N_38263,N_34663,N_30662);
and U38264 (N_38264,N_34375,N_30088);
and U38265 (N_38265,N_34144,N_33224);
or U38266 (N_38266,N_33642,N_34785);
and U38267 (N_38267,N_33412,N_30961);
and U38268 (N_38268,N_30713,N_31211);
xor U38269 (N_38269,N_31071,N_32697);
nand U38270 (N_38270,N_34085,N_34895);
nand U38271 (N_38271,N_32913,N_30924);
or U38272 (N_38272,N_33583,N_34627);
and U38273 (N_38273,N_33859,N_33528);
nor U38274 (N_38274,N_32255,N_30740);
or U38275 (N_38275,N_30282,N_32040);
and U38276 (N_38276,N_31359,N_32750);
nor U38277 (N_38277,N_34059,N_32543);
or U38278 (N_38278,N_32012,N_33735);
nor U38279 (N_38279,N_32218,N_34753);
xnor U38280 (N_38280,N_32969,N_34617);
xnor U38281 (N_38281,N_31154,N_33237);
xor U38282 (N_38282,N_31724,N_34653);
nor U38283 (N_38283,N_31714,N_34765);
xor U38284 (N_38284,N_31340,N_30694);
nand U38285 (N_38285,N_30980,N_30402);
nor U38286 (N_38286,N_32794,N_31084);
or U38287 (N_38287,N_30349,N_31826);
nand U38288 (N_38288,N_33238,N_32543);
nor U38289 (N_38289,N_34467,N_31921);
nor U38290 (N_38290,N_33665,N_31105);
or U38291 (N_38291,N_32401,N_31028);
or U38292 (N_38292,N_31831,N_30755);
xor U38293 (N_38293,N_34863,N_32409);
nor U38294 (N_38294,N_33692,N_30574);
xnor U38295 (N_38295,N_31913,N_31401);
nand U38296 (N_38296,N_30717,N_34641);
nor U38297 (N_38297,N_33511,N_33002);
nand U38298 (N_38298,N_33247,N_32904);
nand U38299 (N_38299,N_32871,N_30691);
nor U38300 (N_38300,N_33871,N_32094);
and U38301 (N_38301,N_32864,N_33128);
or U38302 (N_38302,N_32295,N_32735);
nand U38303 (N_38303,N_32569,N_31922);
nand U38304 (N_38304,N_31158,N_30873);
nor U38305 (N_38305,N_34665,N_31471);
and U38306 (N_38306,N_33628,N_33578);
xor U38307 (N_38307,N_34463,N_34486);
nor U38308 (N_38308,N_30201,N_33238);
nor U38309 (N_38309,N_31270,N_30035);
or U38310 (N_38310,N_33153,N_31548);
nand U38311 (N_38311,N_32239,N_34552);
or U38312 (N_38312,N_34848,N_30139);
nand U38313 (N_38313,N_34702,N_31482);
nand U38314 (N_38314,N_30037,N_32501);
nand U38315 (N_38315,N_31709,N_33991);
nor U38316 (N_38316,N_32921,N_33770);
nand U38317 (N_38317,N_34816,N_32728);
nand U38318 (N_38318,N_32690,N_31757);
or U38319 (N_38319,N_33212,N_33108);
xor U38320 (N_38320,N_33402,N_33868);
nand U38321 (N_38321,N_32448,N_34365);
nor U38322 (N_38322,N_31464,N_31158);
or U38323 (N_38323,N_34124,N_34683);
xor U38324 (N_38324,N_31706,N_30734);
and U38325 (N_38325,N_32795,N_33182);
or U38326 (N_38326,N_33030,N_30156);
and U38327 (N_38327,N_34085,N_31115);
and U38328 (N_38328,N_33342,N_31542);
nand U38329 (N_38329,N_30215,N_34144);
or U38330 (N_38330,N_32746,N_33042);
nor U38331 (N_38331,N_30717,N_33840);
and U38332 (N_38332,N_34998,N_34352);
nand U38333 (N_38333,N_30362,N_30511);
or U38334 (N_38334,N_32761,N_30710);
nand U38335 (N_38335,N_30091,N_30208);
or U38336 (N_38336,N_31459,N_32670);
nand U38337 (N_38337,N_32257,N_33081);
nor U38338 (N_38338,N_33114,N_34285);
xnor U38339 (N_38339,N_31261,N_32660);
and U38340 (N_38340,N_30676,N_31811);
nor U38341 (N_38341,N_33595,N_31722);
and U38342 (N_38342,N_32154,N_34004);
and U38343 (N_38343,N_33624,N_31006);
or U38344 (N_38344,N_32199,N_34886);
xor U38345 (N_38345,N_30313,N_34174);
xnor U38346 (N_38346,N_33053,N_33459);
nor U38347 (N_38347,N_30384,N_32147);
nor U38348 (N_38348,N_30004,N_32011);
nand U38349 (N_38349,N_32173,N_32067);
xnor U38350 (N_38350,N_33458,N_31012);
nand U38351 (N_38351,N_30313,N_30390);
nand U38352 (N_38352,N_34648,N_34940);
or U38353 (N_38353,N_32551,N_33191);
nand U38354 (N_38354,N_33985,N_31274);
nor U38355 (N_38355,N_31156,N_32751);
or U38356 (N_38356,N_30010,N_30943);
nand U38357 (N_38357,N_34954,N_33059);
or U38358 (N_38358,N_30729,N_30177);
or U38359 (N_38359,N_32142,N_32964);
nor U38360 (N_38360,N_34649,N_33749);
and U38361 (N_38361,N_32433,N_30844);
nand U38362 (N_38362,N_30106,N_34986);
nand U38363 (N_38363,N_32507,N_34559);
and U38364 (N_38364,N_32896,N_30975);
nor U38365 (N_38365,N_33659,N_32760);
nand U38366 (N_38366,N_32134,N_31686);
and U38367 (N_38367,N_30380,N_31308);
xor U38368 (N_38368,N_30647,N_34669);
nand U38369 (N_38369,N_33695,N_31351);
and U38370 (N_38370,N_33116,N_33574);
nor U38371 (N_38371,N_31436,N_32943);
nor U38372 (N_38372,N_31526,N_34219);
or U38373 (N_38373,N_33098,N_30053);
or U38374 (N_38374,N_32542,N_33697);
nand U38375 (N_38375,N_32910,N_34908);
xnor U38376 (N_38376,N_34239,N_30221);
or U38377 (N_38377,N_34982,N_34922);
nand U38378 (N_38378,N_34749,N_32454);
nand U38379 (N_38379,N_33798,N_30484);
xnor U38380 (N_38380,N_31008,N_31463);
and U38381 (N_38381,N_32893,N_30001);
or U38382 (N_38382,N_31043,N_31007);
nand U38383 (N_38383,N_34578,N_33528);
or U38384 (N_38384,N_31152,N_31730);
and U38385 (N_38385,N_34789,N_32348);
nor U38386 (N_38386,N_30853,N_31588);
nand U38387 (N_38387,N_33048,N_32123);
nand U38388 (N_38388,N_31426,N_34368);
nor U38389 (N_38389,N_33923,N_33642);
and U38390 (N_38390,N_30091,N_33865);
nand U38391 (N_38391,N_30530,N_31653);
nand U38392 (N_38392,N_33832,N_33503);
nor U38393 (N_38393,N_33164,N_30545);
or U38394 (N_38394,N_34795,N_30212);
and U38395 (N_38395,N_30267,N_30458);
xnor U38396 (N_38396,N_30727,N_30657);
nor U38397 (N_38397,N_34298,N_30785);
nor U38398 (N_38398,N_34106,N_34223);
nor U38399 (N_38399,N_32602,N_34342);
nand U38400 (N_38400,N_34361,N_33795);
nor U38401 (N_38401,N_32246,N_32480);
or U38402 (N_38402,N_31336,N_30558);
or U38403 (N_38403,N_31892,N_33383);
nand U38404 (N_38404,N_32959,N_34333);
or U38405 (N_38405,N_34457,N_32242);
and U38406 (N_38406,N_32923,N_32960);
nand U38407 (N_38407,N_33631,N_32821);
nand U38408 (N_38408,N_33254,N_32948);
and U38409 (N_38409,N_31925,N_31989);
nor U38410 (N_38410,N_32230,N_30636);
nor U38411 (N_38411,N_31149,N_30082);
and U38412 (N_38412,N_34878,N_34433);
and U38413 (N_38413,N_31524,N_32558);
or U38414 (N_38414,N_30163,N_30333);
nand U38415 (N_38415,N_31093,N_34458);
or U38416 (N_38416,N_32159,N_31951);
or U38417 (N_38417,N_31938,N_34391);
nor U38418 (N_38418,N_30795,N_30088);
and U38419 (N_38419,N_31937,N_30098);
nand U38420 (N_38420,N_30061,N_30811);
or U38421 (N_38421,N_32847,N_31912);
xnor U38422 (N_38422,N_31656,N_33619);
nor U38423 (N_38423,N_34090,N_30697);
nand U38424 (N_38424,N_30011,N_30465);
nand U38425 (N_38425,N_32950,N_34890);
and U38426 (N_38426,N_34445,N_31803);
and U38427 (N_38427,N_34565,N_34872);
and U38428 (N_38428,N_32382,N_31346);
nand U38429 (N_38429,N_30311,N_30510);
and U38430 (N_38430,N_33892,N_34932);
nor U38431 (N_38431,N_30357,N_32818);
or U38432 (N_38432,N_31631,N_33670);
xor U38433 (N_38433,N_33974,N_33789);
or U38434 (N_38434,N_32747,N_34951);
and U38435 (N_38435,N_33095,N_30547);
and U38436 (N_38436,N_31001,N_30665);
or U38437 (N_38437,N_34002,N_30157);
or U38438 (N_38438,N_32015,N_33790);
xor U38439 (N_38439,N_33505,N_32640);
nand U38440 (N_38440,N_33396,N_33131);
and U38441 (N_38441,N_31470,N_33492);
and U38442 (N_38442,N_31277,N_32073);
or U38443 (N_38443,N_33110,N_30810);
or U38444 (N_38444,N_30494,N_32603);
and U38445 (N_38445,N_30767,N_30329);
nand U38446 (N_38446,N_30215,N_32424);
xor U38447 (N_38447,N_34769,N_34062);
or U38448 (N_38448,N_34442,N_34797);
and U38449 (N_38449,N_30341,N_33221);
and U38450 (N_38450,N_30346,N_32950);
nor U38451 (N_38451,N_34735,N_34497);
and U38452 (N_38452,N_34456,N_32764);
and U38453 (N_38453,N_33220,N_33251);
nand U38454 (N_38454,N_34980,N_30661);
nand U38455 (N_38455,N_31650,N_34749);
or U38456 (N_38456,N_32432,N_30001);
and U38457 (N_38457,N_34476,N_30277);
or U38458 (N_38458,N_33418,N_30467);
xor U38459 (N_38459,N_32888,N_34045);
xor U38460 (N_38460,N_30354,N_33963);
or U38461 (N_38461,N_34248,N_34401);
nor U38462 (N_38462,N_33145,N_30605);
or U38463 (N_38463,N_31223,N_33560);
xnor U38464 (N_38464,N_31823,N_32028);
and U38465 (N_38465,N_34758,N_33004);
and U38466 (N_38466,N_31544,N_30154);
or U38467 (N_38467,N_33147,N_30158);
and U38468 (N_38468,N_34468,N_32873);
nand U38469 (N_38469,N_33066,N_34706);
nor U38470 (N_38470,N_33456,N_31463);
and U38471 (N_38471,N_32001,N_31827);
or U38472 (N_38472,N_34045,N_32736);
nand U38473 (N_38473,N_33712,N_33970);
nor U38474 (N_38474,N_30649,N_31995);
nand U38475 (N_38475,N_32353,N_32459);
nor U38476 (N_38476,N_32956,N_31944);
nor U38477 (N_38477,N_30908,N_33661);
or U38478 (N_38478,N_30518,N_30714);
nand U38479 (N_38479,N_34417,N_32721);
nand U38480 (N_38480,N_33976,N_30834);
and U38481 (N_38481,N_30439,N_33434);
nand U38482 (N_38482,N_33325,N_30567);
or U38483 (N_38483,N_30175,N_33132);
xor U38484 (N_38484,N_30298,N_31020);
or U38485 (N_38485,N_32726,N_31831);
nand U38486 (N_38486,N_30683,N_30501);
and U38487 (N_38487,N_33995,N_32830);
nor U38488 (N_38488,N_32033,N_34475);
and U38489 (N_38489,N_34520,N_33489);
or U38490 (N_38490,N_33427,N_33738);
or U38491 (N_38491,N_32904,N_32502);
nand U38492 (N_38492,N_34391,N_30319);
nand U38493 (N_38493,N_30382,N_34923);
xnor U38494 (N_38494,N_30599,N_33156);
nand U38495 (N_38495,N_32294,N_32836);
or U38496 (N_38496,N_33082,N_34877);
and U38497 (N_38497,N_32244,N_34475);
and U38498 (N_38498,N_31278,N_31905);
nand U38499 (N_38499,N_34408,N_33628);
nor U38500 (N_38500,N_33556,N_30885);
nand U38501 (N_38501,N_31957,N_31782);
nor U38502 (N_38502,N_32314,N_31005);
xnor U38503 (N_38503,N_33803,N_31163);
or U38504 (N_38504,N_33582,N_30558);
nor U38505 (N_38505,N_33327,N_33549);
nor U38506 (N_38506,N_30460,N_32916);
or U38507 (N_38507,N_33981,N_33115);
nand U38508 (N_38508,N_31738,N_31858);
or U38509 (N_38509,N_34210,N_34632);
nand U38510 (N_38510,N_31991,N_31379);
and U38511 (N_38511,N_31563,N_34089);
and U38512 (N_38512,N_32843,N_33508);
nand U38513 (N_38513,N_32384,N_34457);
xnor U38514 (N_38514,N_30463,N_32855);
nor U38515 (N_38515,N_34786,N_30693);
xor U38516 (N_38516,N_33128,N_31575);
and U38517 (N_38517,N_33427,N_34235);
and U38518 (N_38518,N_31041,N_33542);
and U38519 (N_38519,N_32649,N_34353);
nand U38520 (N_38520,N_30747,N_30139);
and U38521 (N_38521,N_30134,N_31114);
nor U38522 (N_38522,N_31221,N_32117);
nand U38523 (N_38523,N_33392,N_30379);
nand U38524 (N_38524,N_33830,N_32365);
nand U38525 (N_38525,N_30303,N_31309);
nand U38526 (N_38526,N_33446,N_32075);
nor U38527 (N_38527,N_32664,N_30912);
xnor U38528 (N_38528,N_31031,N_33019);
nor U38529 (N_38529,N_32234,N_30298);
nand U38530 (N_38530,N_31800,N_31284);
nand U38531 (N_38531,N_32515,N_34932);
nand U38532 (N_38532,N_32557,N_30603);
and U38533 (N_38533,N_31236,N_34162);
or U38534 (N_38534,N_32485,N_32508);
nand U38535 (N_38535,N_30460,N_32120);
or U38536 (N_38536,N_31978,N_34024);
xor U38537 (N_38537,N_34519,N_34308);
nand U38538 (N_38538,N_34602,N_32885);
nor U38539 (N_38539,N_30295,N_30658);
nor U38540 (N_38540,N_30912,N_33888);
xor U38541 (N_38541,N_32038,N_33390);
and U38542 (N_38542,N_33231,N_30658);
or U38543 (N_38543,N_34035,N_33312);
nand U38544 (N_38544,N_32882,N_32821);
or U38545 (N_38545,N_31718,N_33386);
nand U38546 (N_38546,N_31705,N_33977);
nor U38547 (N_38547,N_31154,N_33305);
nor U38548 (N_38548,N_33804,N_32439);
nor U38549 (N_38549,N_31303,N_31905);
nand U38550 (N_38550,N_31186,N_31778);
and U38551 (N_38551,N_30218,N_30892);
nor U38552 (N_38552,N_34798,N_30040);
or U38553 (N_38553,N_34693,N_31768);
and U38554 (N_38554,N_34216,N_34738);
nor U38555 (N_38555,N_34459,N_31880);
nor U38556 (N_38556,N_31118,N_32798);
nor U38557 (N_38557,N_32084,N_31966);
xor U38558 (N_38558,N_34028,N_34015);
xnor U38559 (N_38559,N_32599,N_33833);
and U38560 (N_38560,N_34089,N_32059);
and U38561 (N_38561,N_33717,N_33348);
or U38562 (N_38562,N_32556,N_31559);
nand U38563 (N_38563,N_30596,N_31179);
nor U38564 (N_38564,N_32685,N_34046);
and U38565 (N_38565,N_32541,N_30766);
and U38566 (N_38566,N_34244,N_31573);
or U38567 (N_38567,N_31828,N_33591);
nand U38568 (N_38568,N_34932,N_32648);
and U38569 (N_38569,N_31036,N_31692);
and U38570 (N_38570,N_32962,N_32813);
nand U38571 (N_38571,N_33181,N_33500);
and U38572 (N_38572,N_32020,N_30354);
or U38573 (N_38573,N_30973,N_32085);
or U38574 (N_38574,N_30031,N_34322);
nor U38575 (N_38575,N_33731,N_32434);
and U38576 (N_38576,N_33702,N_32909);
and U38577 (N_38577,N_30115,N_32986);
nor U38578 (N_38578,N_31252,N_31094);
or U38579 (N_38579,N_31386,N_32078);
and U38580 (N_38580,N_30852,N_34675);
nand U38581 (N_38581,N_32246,N_32603);
or U38582 (N_38582,N_33274,N_31740);
nand U38583 (N_38583,N_30497,N_30839);
xnor U38584 (N_38584,N_31059,N_30365);
nor U38585 (N_38585,N_34505,N_32203);
nand U38586 (N_38586,N_30784,N_31276);
nor U38587 (N_38587,N_33126,N_30453);
nand U38588 (N_38588,N_34072,N_34511);
nor U38589 (N_38589,N_31632,N_32109);
nand U38590 (N_38590,N_30400,N_30999);
or U38591 (N_38591,N_30474,N_34226);
nand U38592 (N_38592,N_30464,N_32742);
or U38593 (N_38593,N_34563,N_30083);
and U38594 (N_38594,N_32446,N_30093);
nor U38595 (N_38595,N_34509,N_32439);
nand U38596 (N_38596,N_34083,N_32829);
or U38597 (N_38597,N_34764,N_31416);
or U38598 (N_38598,N_33062,N_34709);
nor U38599 (N_38599,N_32910,N_31394);
or U38600 (N_38600,N_32428,N_34258);
nor U38601 (N_38601,N_32235,N_31686);
nand U38602 (N_38602,N_34241,N_30602);
or U38603 (N_38603,N_34908,N_33630);
nand U38604 (N_38604,N_34725,N_32059);
nor U38605 (N_38605,N_32850,N_34046);
and U38606 (N_38606,N_34376,N_31263);
and U38607 (N_38607,N_34780,N_32049);
nand U38608 (N_38608,N_34054,N_30497);
or U38609 (N_38609,N_33165,N_34536);
and U38610 (N_38610,N_32159,N_30971);
and U38611 (N_38611,N_33088,N_31464);
nor U38612 (N_38612,N_31875,N_31289);
nor U38613 (N_38613,N_32686,N_30216);
nand U38614 (N_38614,N_34948,N_33906);
and U38615 (N_38615,N_31937,N_34759);
nor U38616 (N_38616,N_31307,N_31567);
nor U38617 (N_38617,N_32429,N_33544);
nor U38618 (N_38618,N_34442,N_30601);
nor U38619 (N_38619,N_34689,N_32073);
nand U38620 (N_38620,N_30979,N_32359);
xor U38621 (N_38621,N_33778,N_34665);
or U38622 (N_38622,N_30761,N_32915);
nor U38623 (N_38623,N_30427,N_32813);
nand U38624 (N_38624,N_31025,N_32501);
nor U38625 (N_38625,N_32215,N_33783);
and U38626 (N_38626,N_33267,N_33390);
nor U38627 (N_38627,N_32688,N_34595);
or U38628 (N_38628,N_31374,N_32103);
nand U38629 (N_38629,N_34091,N_30179);
nand U38630 (N_38630,N_34101,N_33803);
nand U38631 (N_38631,N_33675,N_32457);
nor U38632 (N_38632,N_32471,N_30586);
or U38633 (N_38633,N_34971,N_32070);
nor U38634 (N_38634,N_32349,N_31844);
or U38635 (N_38635,N_33607,N_32068);
xnor U38636 (N_38636,N_32325,N_31687);
nand U38637 (N_38637,N_32066,N_30330);
xnor U38638 (N_38638,N_30794,N_32281);
or U38639 (N_38639,N_34172,N_33986);
nor U38640 (N_38640,N_34329,N_33473);
or U38641 (N_38641,N_34579,N_34679);
or U38642 (N_38642,N_30204,N_30082);
and U38643 (N_38643,N_30756,N_32368);
nor U38644 (N_38644,N_33174,N_33691);
nand U38645 (N_38645,N_31071,N_30107);
nand U38646 (N_38646,N_34330,N_30246);
and U38647 (N_38647,N_30525,N_31036);
or U38648 (N_38648,N_31884,N_32337);
or U38649 (N_38649,N_34739,N_30748);
nand U38650 (N_38650,N_34843,N_30318);
and U38651 (N_38651,N_33053,N_34247);
xnor U38652 (N_38652,N_33371,N_32080);
nand U38653 (N_38653,N_34522,N_34735);
and U38654 (N_38654,N_30673,N_32756);
and U38655 (N_38655,N_32276,N_31572);
and U38656 (N_38656,N_31734,N_32238);
or U38657 (N_38657,N_32320,N_33761);
nand U38658 (N_38658,N_32905,N_34060);
and U38659 (N_38659,N_32163,N_30476);
or U38660 (N_38660,N_31326,N_34459);
or U38661 (N_38661,N_30107,N_32788);
nor U38662 (N_38662,N_34439,N_31048);
nand U38663 (N_38663,N_30312,N_33115);
and U38664 (N_38664,N_34101,N_32758);
nor U38665 (N_38665,N_30992,N_33608);
and U38666 (N_38666,N_31671,N_33893);
xor U38667 (N_38667,N_30712,N_31559);
nor U38668 (N_38668,N_34254,N_34342);
nor U38669 (N_38669,N_30464,N_33048);
nand U38670 (N_38670,N_33788,N_32446);
and U38671 (N_38671,N_31757,N_33586);
nor U38672 (N_38672,N_34870,N_30738);
and U38673 (N_38673,N_30111,N_30514);
nor U38674 (N_38674,N_34297,N_31955);
nor U38675 (N_38675,N_33965,N_31634);
nand U38676 (N_38676,N_30581,N_34506);
or U38677 (N_38677,N_34575,N_30388);
and U38678 (N_38678,N_30248,N_32000);
and U38679 (N_38679,N_31847,N_33526);
or U38680 (N_38680,N_30516,N_30592);
nand U38681 (N_38681,N_34949,N_34024);
or U38682 (N_38682,N_34797,N_31214);
and U38683 (N_38683,N_32430,N_33118);
xnor U38684 (N_38684,N_32003,N_34960);
nor U38685 (N_38685,N_33735,N_34469);
or U38686 (N_38686,N_33265,N_32616);
or U38687 (N_38687,N_31823,N_32655);
and U38688 (N_38688,N_30435,N_32139);
or U38689 (N_38689,N_30147,N_32407);
nand U38690 (N_38690,N_31699,N_31168);
and U38691 (N_38691,N_32948,N_34597);
nand U38692 (N_38692,N_32075,N_31751);
and U38693 (N_38693,N_32916,N_31595);
xnor U38694 (N_38694,N_34364,N_31071);
xnor U38695 (N_38695,N_31075,N_33038);
or U38696 (N_38696,N_30981,N_34043);
xor U38697 (N_38697,N_32011,N_33816);
or U38698 (N_38698,N_31824,N_33610);
xor U38699 (N_38699,N_30483,N_30818);
and U38700 (N_38700,N_32291,N_31762);
xor U38701 (N_38701,N_30452,N_33777);
nor U38702 (N_38702,N_30965,N_34415);
and U38703 (N_38703,N_30793,N_34243);
nand U38704 (N_38704,N_30876,N_32807);
or U38705 (N_38705,N_31376,N_31170);
and U38706 (N_38706,N_32901,N_33495);
or U38707 (N_38707,N_30478,N_31900);
or U38708 (N_38708,N_34253,N_31637);
and U38709 (N_38709,N_31723,N_32304);
and U38710 (N_38710,N_33914,N_32139);
nand U38711 (N_38711,N_31334,N_34588);
nand U38712 (N_38712,N_32002,N_34307);
nor U38713 (N_38713,N_31184,N_33891);
nand U38714 (N_38714,N_33692,N_30807);
nor U38715 (N_38715,N_32734,N_31044);
or U38716 (N_38716,N_30214,N_31481);
xor U38717 (N_38717,N_33915,N_34429);
xnor U38718 (N_38718,N_32694,N_30277);
nor U38719 (N_38719,N_33125,N_34391);
nor U38720 (N_38720,N_33125,N_34333);
or U38721 (N_38721,N_31216,N_32465);
or U38722 (N_38722,N_34998,N_31755);
nor U38723 (N_38723,N_30518,N_32589);
nand U38724 (N_38724,N_30486,N_34398);
nor U38725 (N_38725,N_32430,N_30381);
nand U38726 (N_38726,N_32596,N_32778);
and U38727 (N_38727,N_31535,N_30422);
nand U38728 (N_38728,N_31864,N_30659);
nor U38729 (N_38729,N_31370,N_33294);
nand U38730 (N_38730,N_32062,N_31410);
or U38731 (N_38731,N_34835,N_31320);
and U38732 (N_38732,N_31023,N_30298);
nor U38733 (N_38733,N_33656,N_34397);
xor U38734 (N_38734,N_31726,N_31792);
and U38735 (N_38735,N_32518,N_32673);
nor U38736 (N_38736,N_34136,N_33053);
nand U38737 (N_38737,N_33698,N_31406);
nand U38738 (N_38738,N_32538,N_31235);
or U38739 (N_38739,N_31040,N_34395);
or U38740 (N_38740,N_34729,N_30818);
nand U38741 (N_38741,N_34703,N_34496);
xnor U38742 (N_38742,N_34830,N_34532);
nor U38743 (N_38743,N_33799,N_31493);
nand U38744 (N_38744,N_31889,N_33276);
nand U38745 (N_38745,N_32806,N_33697);
and U38746 (N_38746,N_34712,N_32909);
nand U38747 (N_38747,N_32647,N_32840);
nor U38748 (N_38748,N_30363,N_34325);
or U38749 (N_38749,N_34750,N_30557);
nor U38750 (N_38750,N_32169,N_33591);
and U38751 (N_38751,N_30232,N_32437);
nor U38752 (N_38752,N_30175,N_30571);
nor U38753 (N_38753,N_33677,N_30963);
nor U38754 (N_38754,N_33297,N_31473);
nor U38755 (N_38755,N_30143,N_32994);
nand U38756 (N_38756,N_34073,N_34855);
nor U38757 (N_38757,N_32264,N_32472);
and U38758 (N_38758,N_32996,N_34906);
xor U38759 (N_38759,N_31976,N_32618);
and U38760 (N_38760,N_31062,N_32168);
nand U38761 (N_38761,N_30755,N_34607);
and U38762 (N_38762,N_30737,N_31375);
nor U38763 (N_38763,N_30044,N_31338);
and U38764 (N_38764,N_31932,N_33667);
nor U38765 (N_38765,N_30927,N_31596);
xor U38766 (N_38766,N_34362,N_31275);
nand U38767 (N_38767,N_31353,N_32460);
xnor U38768 (N_38768,N_34974,N_32559);
nor U38769 (N_38769,N_31023,N_33653);
and U38770 (N_38770,N_32861,N_32896);
nor U38771 (N_38771,N_34028,N_31089);
nor U38772 (N_38772,N_33894,N_31078);
xnor U38773 (N_38773,N_32432,N_33342);
and U38774 (N_38774,N_33168,N_31284);
nor U38775 (N_38775,N_33979,N_32108);
or U38776 (N_38776,N_34679,N_31038);
nand U38777 (N_38777,N_33172,N_31708);
or U38778 (N_38778,N_30311,N_31167);
or U38779 (N_38779,N_31561,N_33731);
xnor U38780 (N_38780,N_32805,N_32540);
or U38781 (N_38781,N_31213,N_31900);
or U38782 (N_38782,N_31202,N_31268);
and U38783 (N_38783,N_33910,N_34573);
and U38784 (N_38784,N_32671,N_30610);
xnor U38785 (N_38785,N_32177,N_33454);
and U38786 (N_38786,N_33018,N_31624);
and U38787 (N_38787,N_30781,N_32196);
and U38788 (N_38788,N_34625,N_30034);
nor U38789 (N_38789,N_31884,N_34838);
and U38790 (N_38790,N_33652,N_30357);
and U38791 (N_38791,N_34357,N_32862);
and U38792 (N_38792,N_33366,N_33051);
or U38793 (N_38793,N_34017,N_31664);
nor U38794 (N_38794,N_31709,N_31770);
nor U38795 (N_38795,N_30029,N_32237);
nor U38796 (N_38796,N_32856,N_34538);
nor U38797 (N_38797,N_30119,N_31166);
and U38798 (N_38798,N_31209,N_31273);
nor U38799 (N_38799,N_33992,N_34266);
nor U38800 (N_38800,N_32934,N_31817);
or U38801 (N_38801,N_31297,N_30439);
nand U38802 (N_38802,N_33434,N_34012);
or U38803 (N_38803,N_34817,N_31162);
nor U38804 (N_38804,N_31497,N_32075);
and U38805 (N_38805,N_30373,N_32447);
or U38806 (N_38806,N_31082,N_33455);
nor U38807 (N_38807,N_34212,N_32000);
and U38808 (N_38808,N_34114,N_34030);
nand U38809 (N_38809,N_32106,N_34234);
nor U38810 (N_38810,N_33863,N_31779);
xnor U38811 (N_38811,N_32466,N_32549);
nand U38812 (N_38812,N_32744,N_33005);
and U38813 (N_38813,N_31927,N_30169);
nand U38814 (N_38814,N_30323,N_31182);
nand U38815 (N_38815,N_30249,N_31136);
nor U38816 (N_38816,N_34433,N_32064);
nand U38817 (N_38817,N_34758,N_34909);
and U38818 (N_38818,N_34315,N_33854);
or U38819 (N_38819,N_30268,N_34666);
and U38820 (N_38820,N_31069,N_30940);
nor U38821 (N_38821,N_30471,N_34170);
xor U38822 (N_38822,N_34055,N_30684);
nand U38823 (N_38823,N_31288,N_30738);
nor U38824 (N_38824,N_32861,N_33288);
nand U38825 (N_38825,N_31784,N_31292);
and U38826 (N_38826,N_30847,N_34477);
or U38827 (N_38827,N_32089,N_32908);
or U38828 (N_38828,N_32794,N_32630);
and U38829 (N_38829,N_30370,N_32087);
and U38830 (N_38830,N_33621,N_30920);
nor U38831 (N_38831,N_33448,N_34299);
or U38832 (N_38832,N_34574,N_34228);
nor U38833 (N_38833,N_30679,N_30148);
or U38834 (N_38834,N_30165,N_30320);
or U38835 (N_38835,N_30508,N_33461);
nor U38836 (N_38836,N_32166,N_34353);
or U38837 (N_38837,N_34621,N_31919);
nor U38838 (N_38838,N_30173,N_30482);
and U38839 (N_38839,N_30512,N_34047);
and U38840 (N_38840,N_34769,N_34730);
and U38841 (N_38841,N_34349,N_31977);
xnor U38842 (N_38842,N_33613,N_33216);
nand U38843 (N_38843,N_33234,N_30562);
xor U38844 (N_38844,N_33666,N_32701);
nor U38845 (N_38845,N_32924,N_30768);
nand U38846 (N_38846,N_32231,N_34693);
nand U38847 (N_38847,N_34378,N_33784);
nor U38848 (N_38848,N_34383,N_31432);
nand U38849 (N_38849,N_33010,N_31547);
or U38850 (N_38850,N_31737,N_34435);
and U38851 (N_38851,N_32128,N_33552);
nand U38852 (N_38852,N_30297,N_33536);
and U38853 (N_38853,N_31882,N_33416);
or U38854 (N_38854,N_32452,N_30079);
nor U38855 (N_38855,N_30495,N_30659);
or U38856 (N_38856,N_32800,N_34576);
and U38857 (N_38857,N_32193,N_31625);
or U38858 (N_38858,N_32601,N_30349);
nor U38859 (N_38859,N_30802,N_31038);
and U38860 (N_38860,N_34442,N_31963);
or U38861 (N_38861,N_34418,N_34318);
nor U38862 (N_38862,N_33586,N_34273);
and U38863 (N_38863,N_31530,N_34444);
nor U38864 (N_38864,N_31606,N_30953);
xnor U38865 (N_38865,N_34595,N_33809);
and U38866 (N_38866,N_32541,N_34886);
and U38867 (N_38867,N_31183,N_31094);
and U38868 (N_38868,N_31597,N_34695);
nor U38869 (N_38869,N_34351,N_32523);
nor U38870 (N_38870,N_31574,N_30792);
and U38871 (N_38871,N_33181,N_30419);
or U38872 (N_38872,N_31544,N_33168);
nor U38873 (N_38873,N_32869,N_32290);
or U38874 (N_38874,N_34399,N_30723);
or U38875 (N_38875,N_34001,N_33836);
xor U38876 (N_38876,N_33720,N_34667);
xor U38877 (N_38877,N_31923,N_30151);
nand U38878 (N_38878,N_33088,N_30859);
and U38879 (N_38879,N_30277,N_31412);
and U38880 (N_38880,N_32816,N_30778);
nand U38881 (N_38881,N_33553,N_34831);
or U38882 (N_38882,N_30284,N_30328);
xnor U38883 (N_38883,N_34371,N_34547);
nor U38884 (N_38884,N_31607,N_34996);
xnor U38885 (N_38885,N_34852,N_32623);
nor U38886 (N_38886,N_32995,N_32346);
xor U38887 (N_38887,N_34471,N_31939);
and U38888 (N_38888,N_33269,N_33319);
nor U38889 (N_38889,N_30411,N_30191);
or U38890 (N_38890,N_30139,N_31531);
xor U38891 (N_38891,N_30947,N_30049);
xor U38892 (N_38892,N_34643,N_31999);
nand U38893 (N_38893,N_31321,N_30132);
nor U38894 (N_38894,N_32404,N_30285);
xnor U38895 (N_38895,N_32787,N_34109);
nand U38896 (N_38896,N_31763,N_33771);
xor U38897 (N_38897,N_33686,N_33597);
or U38898 (N_38898,N_34966,N_30576);
nand U38899 (N_38899,N_30410,N_33923);
nor U38900 (N_38900,N_32337,N_33958);
or U38901 (N_38901,N_30744,N_32817);
nor U38902 (N_38902,N_33597,N_32259);
xor U38903 (N_38903,N_31940,N_30312);
nand U38904 (N_38904,N_32482,N_33951);
or U38905 (N_38905,N_31464,N_33534);
nor U38906 (N_38906,N_31817,N_34065);
and U38907 (N_38907,N_33429,N_34392);
nor U38908 (N_38908,N_30542,N_31206);
nor U38909 (N_38909,N_31671,N_32431);
or U38910 (N_38910,N_30725,N_34988);
or U38911 (N_38911,N_33567,N_32352);
nor U38912 (N_38912,N_34816,N_30553);
nand U38913 (N_38913,N_34456,N_32954);
xnor U38914 (N_38914,N_30629,N_31368);
xnor U38915 (N_38915,N_30767,N_33251);
or U38916 (N_38916,N_32943,N_33913);
xnor U38917 (N_38917,N_30712,N_32191);
nand U38918 (N_38918,N_33864,N_34886);
nor U38919 (N_38919,N_30981,N_30454);
xor U38920 (N_38920,N_34655,N_33905);
nand U38921 (N_38921,N_33909,N_32097);
nand U38922 (N_38922,N_31418,N_31905);
nor U38923 (N_38923,N_32022,N_33905);
nor U38924 (N_38924,N_32775,N_34997);
nand U38925 (N_38925,N_32873,N_33847);
or U38926 (N_38926,N_33874,N_31176);
nand U38927 (N_38927,N_30084,N_33869);
xor U38928 (N_38928,N_34364,N_30767);
xnor U38929 (N_38929,N_33813,N_31692);
and U38930 (N_38930,N_32339,N_33474);
nand U38931 (N_38931,N_32435,N_30608);
or U38932 (N_38932,N_31328,N_31285);
and U38933 (N_38933,N_30590,N_33543);
nor U38934 (N_38934,N_31471,N_30887);
or U38935 (N_38935,N_34383,N_32942);
or U38936 (N_38936,N_30187,N_30630);
or U38937 (N_38937,N_30244,N_34044);
and U38938 (N_38938,N_33507,N_34996);
nor U38939 (N_38939,N_30069,N_32402);
nand U38940 (N_38940,N_32708,N_34404);
or U38941 (N_38941,N_33068,N_33513);
nand U38942 (N_38942,N_30883,N_34761);
nor U38943 (N_38943,N_34936,N_33853);
nor U38944 (N_38944,N_30774,N_34585);
xor U38945 (N_38945,N_33205,N_34401);
nand U38946 (N_38946,N_32482,N_30156);
nand U38947 (N_38947,N_30900,N_32695);
or U38948 (N_38948,N_33737,N_31001);
nor U38949 (N_38949,N_31153,N_32277);
nor U38950 (N_38950,N_30396,N_34316);
or U38951 (N_38951,N_34029,N_31722);
or U38952 (N_38952,N_33421,N_30699);
and U38953 (N_38953,N_31598,N_31337);
xor U38954 (N_38954,N_34913,N_31415);
or U38955 (N_38955,N_34511,N_33590);
nand U38956 (N_38956,N_32282,N_33686);
nor U38957 (N_38957,N_32079,N_30558);
xor U38958 (N_38958,N_31105,N_31436);
and U38959 (N_38959,N_33137,N_33011);
nand U38960 (N_38960,N_30611,N_31341);
nor U38961 (N_38961,N_30125,N_31833);
nor U38962 (N_38962,N_34821,N_34113);
and U38963 (N_38963,N_30188,N_34656);
nor U38964 (N_38964,N_34916,N_32149);
or U38965 (N_38965,N_31462,N_32530);
or U38966 (N_38966,N_34326,N_30087);
or U38967 (N_38967,N_32223,N_34044);
and U38968 (N_38968,N_33973,N_31010);
xnor U38969 (N_38969,N_33337,N_31746);
nor U38970 (N_38970,N_33865,N_32496);
and U38971 (N_38971,N_30106,N_33508);
nand U38972 (N_38972,N_32095,N_32610);
and U38973 (N_38973,N_31084,N_32493);
nor U38974 (N_38974,N_30481,N_33345);
and U38975 (N_38975,N_33625,N_33039);
nand U38976 (N_38976,N_33500,N_30535);
and U38977 (N_38977,N_30317,N_34904);
nand U38978 (N_38978,N_33587,N_30577);
nand U38979 (N_38979,N_30769,N_34640);
and U38980 (N_38980,N_34190,N_33983);
nand U38981 (N_38981,N_30646,N_32753);
and U38982 (N_38982,N_34046,N_33977);
and U38983 (N_38983,N_31038,N_32488);
and U38984 (N_38984,N_30820,N_34497);
or U38985 (N_38985,N_32851,N_33435);
and U38986 (N_38986,N_34068,N_34505);
xor U38987 (N_38987,N_31507,N_31733);
and U38988 (N_38988,N_32796,N_33505);
and U38989 (N_38989,N_34172,N_30581);
nand U38990 (N_38990,N_32569,N_30612);
or U38991 (N_38991,N_34791,N_34149);
or U38992 (N_38992,N_33313,N_30916);
or U38993 (N_38993,N_30468,N_32721);
or U38994 (N_38994,N_34986,N_31094);
nor U38995 (N_38995,N_33861,N_30413);
and U38996 (N_38996,N_30000,N_34228);
nor U38997 (N_38997,N_31074,N_34295);
nor U38998 (N_38998,N_30044,N_34946);
nor U38999 (N_38999,N_33805,N_34786);
and U39000 (N_39000,N_32874,N_34145);
and U39001 (N_39001,N_30813,N_32750);
and U39002 (N_39002,N_33862,N_34448);
nand U39003 (N_39003,N_34976,N_30806);
xnor U39004 (N_39004,N_32037,N_31488);
nand U39005 (N_39005,N_34433,N_31458);
xnor U39006 (N_39006,N_32712,N_33492);
nor U39007 (N_39007,N_33218,N_30804);
nor U39008 (N_39008,N_30466,N_30749);
and U39009 (N_39009,N_30497,N_30244);
or U39010 (N_39010,N_31072,N_34926);
nand U39011 (N_39011,N_33439,N_33705);
and U39012 (N_39012,N_34613,N_30299);
or U39013 (N_39013,N_33205,N_30621);
or U39014 (N_39014,N_31849,N_32757);
xor U39015 (N_39015,N_30384,N_30638);
and U39016 (N_39016,N_34777,N_31811);
nand U39017 (N_39017,N_33475,N_31062);
nor U39018 (N_39018,N_30376,N_30415);
and U39019 (N_39019,N_32835,N_30593);
nand U39020 (N_39020,N_34908,N_31933);
nor U39021 (N_39021,N_33730,N_30806);
nor U39022 (N_39022,N_34124,N_33022);
nor U39023 (N_39023,N_34154,N_32809);
or U39024 (N_39024,N_34585,N_33020);
or U39025 (N_39025,N_30237,N_31655);
or U39026 (N_39026,N_30493,N_32773);
nor U39027 (N_39027,N_34513,N_31085);
xor U39028 (N_39028,N_31926,N_34330);
nor U39029 (N_39029,N_31368,N_32414);
nand U39030 (N_39030,N_34355,N_31413);
nor U39031 (N_39031,N_33469,N_34717);
xor U39032 (N_39032,N_33697,N_33194);
and U39033 (N_39033,N_34476,N_31536);
and U39034 (N_39034,N_34095,N_32951);
nor U39035 (N_39035,N_32542,N_30205);
and U39036 (N_39036,N_30906,N_33691);
nand U39037 (N_39037,N_31233,N_31379);
or U39038 (N_39038,N_32412,N_31606);
or U39039 (N_39039,N_34727,N_31665);
and U39040 (N_39040,N_34580,N_31497);
and U39041 (N_39041,N_30034,N_34150);
and U39042 (N_39042,N_30243,N_33473);
or U39043 (N_39043,N_30676,N_31201);
nand U39044 (N_39044,N_30979,N_32936);
nor U39045 (N_39045,N_33293,N_32935);
and U39046 (N_39046,N_32960,N_31520);
nand U39047 (N_39047,N_34577,N_30828);
and U39048 (N_39048,N_31913,N_34149);
nor U39049 (N_39049,N_32081,N_31028);
nand U39050 (N_39050,N_33798,N_33707);
nor U39051 (N_39051,N_33468,N_31198);
nor U39052 (N_39052,N_31453,N_30149);
or U39053 (N_39053,N_32610,N_31190);
xor U39054 (N_39054,N_34049,N_34039);
nand U39055 (N_39055,N_34505,N_32408);
or U39056 (N_39056,N_32648,N_30144);
nor U39057 (N_39057,N_31460,N_34793);
nand U39058 (N_39058,N_30168,N_33552);
nand U39059 (N_39059,N_34895,N_33186);
nand U39060 (N_39060,N_31662,N_34846);
or U39061 (N_39061,N_32695,N_34048);
or U39062 (N_39062,N_34694,N_31731);
or U39063 (N_39063,N_30921,N_30895);
nor U39064 (N_39064,N_33597,N_31846);
and U39065 (N_39065,N_33352,N_30669);
or U39066 (N_39066,N_30875,N_31891);
nand U39067 (N_39067,N_30163,N_31452);
and U39068 (N_39068,N_33696,N_31638);
or U39069 (N_39069,N_31552,N_31846);
or U39070 (N_39070,N_33322,N_31056);
nor U39071 (N_39071,N_32050,N_32880);
nand U39072 (N_39072,N_33749,N_34476);
and U39073 (N_39073,N_32793,N_33449);
or U39074 (N_39074,N_33375,N_31353);
nor U39075 (N_39075,N_34390,N_31698);
and U39076 (N_39076,N_30605,N_34015);
and U39077 (N_39077,N_31027,N_30294);
nand U39078 (N_39078,N_32673,N_31545);
and U39079 (N_39079,N_32767,N_30461);
and U39080 (N_39080,N_32299,N_32384);
and U39081 (N_39081,N_30207,N_32903);
and U39082 (N_39082,N_32798,N_32478);
nor U39083 (N_39083,N_30292,N_31725);
and U39084 (N_39084,N_31896,N_33079);
nand U39085 (N_39085,N_33961,N_33841);
and U39086 (N_39086,N_32103,N_33668);
nand U39087 (N_39087,N_34350,N_32278);
or U39088 (N_39088,N_31510,N_31431);
nand U39089 (N_39089,N_34146,N_32378);
or U39090 (N_39090,N_31799,N_30764);
nand U39091 (N_39091,N_33830,N_34636);
nand U39092 (N_39092,N_33085,N_34358);
nor U39093 (N_39093,N_34740,N_30348);
and U39094 (N_39094,N_30706,N_31017);
and U39095 (N_39095,N_30763,N_32555);
xnor U39096 (N_39096,N_32986,N_31256);
or U39097 (N_39097,N_34122,N_34092);
or U39098 (N_39098,N_34775,N_31127);
and U39099 (N_39099,N_30366,N_34610);
and U39100 (N_39100,N_34919,N_33505);
and U39101 (N_39101,N_34967,N_31459);
nand U39102 (N_39102,N_32589,N_32399);
xnor U39103 (N_39103,N_31780,N_32716);
or U39104 (N_39104,N_30709,N_31516);
and U39105 (N_39105,N_30476,N_33396);
and U39106 (N_39106,N_34063,N_32983);
nand U39107 (N_39107,N_31435,N_31806);
nor U39108 (N_39108,N_32615,N_31346);
nor U39109 (N_39109,N_32165,N_31395);
or U39110 (N_39110,N_33248,N_31603);
nor U39111 (N_39111,N_30926,N_34679);
xnor U39112 (N_39112,N_32380,N_32858);
nand U39113 (N_39113,N_32793,N_33471);
or U39114 (N_39114,N_33976,N_32873);
nor U39115 (N_39115,N_34965,N_32204);
nor U39116 (N_39116,N_31517,N_34982);
and U39117 (N_39117,N_34286,N_32937);
nor U39118 (N_39118,N_32870,N_31351);
or U39119 (N_39119,N_30130,N_30531);
and U39120 (N_39120,N_33411,N_32509);
or U39121 (N_39121,N_34094,N_34376);
xor U39122 (N_39122,N_34939,N_32538);
nand U39123 (N_39123,N_33123,N_33000);
and U39124 (N_39124,N_34394,N_31301);
or U39125 (N_39125,N_34463,N_34736);
and U39126 (N_39126,N_32436,N_30978);
or U39127 (N_39127,N_32274,N_32287);
xor U39128 (N_39128,N_31847,N_34933);
nor U39129 (N_39129,N_30286,N_32855);
or U39130 (N_39130,N_30240,N_31005);
and U39131 (N_39131,N_33289,N_32897);
and U39132 (N_39132,N_30559,N_32337);
nor U39133 (N_39133,N_34814,N_32002);
and U39134 (N_39134,N_31726,N_32816);
and U39135 (N_39135,N_31274,N_33347);
and U39136 (N_39136,N_31148,N_33982);
nand U39137 (N_39137,N_31193,N_34211);
nand U39138 (N_39138,N_31682,N_32007);
or U39139 (N_39139,N_32639,N_31942);
nand U39140 (N_39140,N_30388,N_32675);
nand U39141 (N_39141,N_32756,N_34227);
nand U39142 (N_39142,N_33458,N_30803);
nand U39143 (N_39143,N_31184,N_34452);
xnor U39144 (N_39144,N_34092,N_30515);
nor U39145 (N_39145,N_33496,N_31805);
and U39146 (N_39146,N_34344,N_33851);
and U39147 (N_39147,N_33877,N_32408);
nand U39148 (N_39148,N_32750,N_31663);
nand U39149 (N_39149,N_32682,N_30997);
xnor U39150 (N_39150,N_34288,N_30707);
nand U39151 (N_39151,N_30022,N_33658);
and U39152 (N_39152,N_30988,N_30534);
nand U39153 (N_39153,N_31672,N_30599);
and U39154 (N_39154,N_31597,N_32031);
or U39155 (N_39155,N_33455,N_34595);
and U39156 (N_39156,N_32119,N_31089);
nor U39157 (N_39157,N_32079,N_30023);
nor U39158 (N_39158,N_30994,N_32713);
nor U39159 (N_39159,N_34702,N_32686);
nor U39160 (N_39160,N_31600,N_32624);
nand U39161 (N_39161,N_32392,N_30419);
or U39162 (N_39162,N_32462,N_32189);
xnor U39163 (N_39163,N_30274,N_31431);
nand U39164 (N_39164,N_34234,N_31978);
or U39165 (N_39165,N_31669,N_31057);
or U39166 (N_39166,N_33476,N_33307);
xor U39167 (N_39167,N_31398,N_34300);
or U39168 (N_39168,N_30668,N_30151);
and U39169 (N_39169,N_32300,N_32215);
or U39170 (N_39170,N_30093,N_34342);
or U39171 (N_39171,N_33940,N_30841);
nand U39172 (N_39172,N_33265,N_33884);
nand U39173 (N_39173,N_30199,N_31842);
nor U39174 (N_39174,N_30138,N_31384);
and U39175 (N_39175,N_34788,N_34597);
and U39176 (N_39176,N_32076,N_32188);
nand U39177 (N_39177,N_30163,N_33931);
nor U39178 (N_39178,N_33612,N_34329);
nand U39179 (N_39179,N_32258,N_33877);
nand U39180 (N_39180,N_32929,N_33921);
xor U39181 (N_39181,N_34839,N_31553);
or U39182 (N_39182,N_32122,N_33079);
nor U39183 (N_39183,N_31696,N_33206);
and U39184 (N_39184,N_32755,N_34616);
nor U39185 (N_39185,N_34776,N_31209);
or U39186 (N_39186,N_32392,N_32958);
nand U39187 (N_39187,N_33712,N_34621);
and U39188 (N_39188,N_31302,N_34211);
nor U39189 (N_39189,N_32633,N_31658);
or U39190 (N_39190,N_34243,N_33876);
nand U39191 (N_39191,N_30391,N_31516);
nand U39192 (N_39192,N_31902,N_33876);
nor U39193 (N_39193,N_34566,N_33399);
nor U39194 (N_39194,N_32450,N_34011);
nand U39195 (N_39195,N_33889,N_32199);
nand U39196 (N_39196,N_33887,N_31560);
xnor U39197 (N_39197,N_32849,N_33052);
and U39198 (N_39198,N_31056,N_31636);
and U39199 (N_39199,N_30147,N_32391);
and U39200 (N_39200,N_33967,N_33904);
nor U39201 (N_39201,N_30783,N_31909);
xnor U39202 (N_39202,N_30880,N_34878);
or U39203 (N_39203,N_31685,N_34120);
nand U39204 (N_39204,N_34031,N_32734);
and U39205 (N_39205,N_33306,N_32156);
nand U39206 (N_39206,N_34784,N_31388);
and U39207 (N_39207,N_34946,N_31859);
nor U39208 (N_39208,N_30195,N_34404);
nand U39209 (N_39209,N_32827,N_33582);
or U39210 (N_39210,N_31959,N_31963);
xor U39211 (N_39211,N_32915,N_31136);
and U39212 (N_39212,N_34604,N_34531);
nor U39213 (N_39213,N_30508,N_33428);
xor U39214 (N_39214,N_33882,N_31657);
and U39215 (N_39215,N_30909,N_32670);
nand U39216 (N_39216,N_32654,N_33398);
or U39217 (N_39217,N_30971,N_31125);
and U39218 (N_39218,N_34461,N_30747);
and U39219 (N_39219,N_33610,N_30264);
and U39220 (N_39220,N_30558,N_31748);
or U39221 (N_39221,N_33771,N_32242);
nor U39222 (N_39222,N_33848,N_32528);
nor U39223 (N_39223,N_31132,N_30562);
nor U39224 (N_39224,N_33328,N_33465);
or U39225 (N_39225,N_30054,N_30044);
or U39226 (N_39226,N_32661,N_33717);
and U39227 (N_39227,N_30648,N_32915);
nand U39228 (N_39228,N_31914,N_34249);
or U39229 (N_39229,N_31978,N_33074);
and U39230 (N_39230,N_31788,N_30859);
and U39231 (N_39231,N_33723,N_31577);
and U39232 (N_39232,N_31463,N_34895);
nor U39233 (N_39233,N_30987,N_30319);
nand U39234 (N_39234,N_34795,N_31389);
nand U39235 (N_39235,N_32565,N_31696);
nor U39236 (N_39236,N_32783,N_33901);
nor U39237 (N_39237,N_32677,N_31257);
xnor U39238 (N_39238,N_30256,N_30049);
and U39239 (N_39239,N_33230,N_30663);
or U39240 (N_39240,N_32823,N_31313);
nand U39241 (N_39241,N_34539,N_34523);
nand U39242 (N_39242,N_31731,N_33804);
and U39243 (N_39243,N_31439,N_34039);
or U39244 (N_39244,N_30414,N_31528);
nor U39245 (N_39245,N_33745,N_30817);
xnor U39246 (N_39246,N_34932,N_30581);
nor U39247 (N_39247,N_33815,N_33161);
nand U39248 (N_39248,N_30551,N_32728);
and U39249 (N_39249,N_30167,N_34745);
or U39250 (N_39250,N_31346,N_33647);
or U39251 (N_39251,N_34835,N_34089);
or U39252 (N_39252,N_34275,N_34495);
and U39253 (N_39253,N_32612,N_31634);
xnor U39254 (N_39254,N_32507,N_32146);
nor U39255 (N_39255,N_30226,N_31510);
and U39256 (N_39256,N_31365,N_32428);
nand U39257 (N_39257,N_31360,N_32609);
nor U39258 (N_39258,N_31155,N_30237);
nand U39259 (N_39259,N_30363,N_34570);
nand U39260 (N_39260,N_34916,N_34164);
and U39261 (N_39261,N_32097,N_34501);
and U39262 (N_39262,N_33070,N_34763);
xor U39263 (N_39263,N_31078,N_32152);
xnor U39264 (N_39264,N_30142,N_30922);
and U39265 (N_39265,N_30250,N_31917);
xnor U39266 (N_39266,N_31270,N_34309);
or U39267 (N_39267,N_31189,N_31748);
or U39268 (N_39268,N_34129,N_34498);
nand U39269 (N_39269,N_31647,N_32716);
and U39270 (N_39270,N_32210,N_33935);
nand U39271 (N_39271,N_34794,N_31269);
nand U39272 (N_39272,N_30196,N_34433);
nor U39273 (N_39273,N_34923,N_31969);
nor U39274 (N_39274,N_31820,N_31653);
nand U39275 (N_39275,N_31333,N_32185);
or U39276 (N_39276,N_34999,N_30818);
nor U39277 (N_39277,N_32851,N_32664);
nand U39278 (N_39278,N_30236,N_30289);
nor U39279 (N_39279,N_34527,N_33699);
and U39280 (N_39280,N_31579,N_32756);
or U39281 (N_39281,N_33702,N_33049);
and U39282 (N_39282,N_33971,N_30856);
or U39283 (N_39283,N_31840,N_30517);
xnor U39284 (N_39284,N_34407,N_32031);
or U39285 (N_39285,N_31939,N_30986);
or U39286 (N_39286,N_34060,N_30605);
and U39287 (N_39287,N_30066,N_31062);
nand U39288 (N_39288,N_32693,N_30917);
or U39289 (N_39289,N_34692,N_32204);
and U39290 (N_39290,N_32684,N_33745);
and U39291 (N_39291,N_30867,N_34841);
and U39292 (N_39292,N_32399,N_32329);
nand U39293 (N_39293,N_30730,N_33826);
or U39294 (N_39294,N_32861,N_30626);
nand U39295 (N_39295,N_31675,N_31478);
or U39296 (N_39296,N_32846,N_30768);
and U39297 (N_39297,N_33212,N_30595);
xnor U39298 (N_39298,N_33061,N_32027);
nand U39299 (N_39299,N_31822,N_31420);
nand U39300 (N_39300,N_34192,N_30240);
or U39301 (N_39301,N_32224,N_30529);
nor U39302 (N_39302,N_31076,N_32193);
xnor U39303 (N_39303,N_33331,N_32458);
or U39304 (N_39304,N_31929,N_31253);
xnor U39305 (N_39305,N_33297,N_31083);
nor U39306 (N_39306,N_31638,N_31155);
or U39307 (N_39307,N_32739,N_30330);
and U39308 (N_39308,N_30055,N_30407);
and U39309 (N_39309,N_32464,N_33811);
nand U39310 (N_39310,N_33848,N_33624);
nand U39311 (N_39311,N_34923,N_30704);
nand U39312 (N_39312,N_30262,N_34578);
xor U39313 (N_39313,N_30661,N_31898);
xnor U39314 (N_39314,N_33163,N_30152);
nand U39315 (N_39315,N_32483,N_34754);
nand U39316 (N_39316,N_31917,N_31665);
or U39317 (N_39317,N_30075,N_32786);
xnor U39318 (N_39318,N_30544,N_32097);
xnor U39319 (N_39319,N_33179,N_31773);
nand U39320 (N_39320,N_32697,N_31342);
nand U39321 (N_39321,N_33937,N_33708);
or U39322 (N_39322,N_31693,N_34154);
xor U39323 (N_39323,N_31064,N_34424);
nor U39324 (N_39324,N_32401,N_34011);
nand U39325 (N_39325,N_31206,N_31382);
nor U39326 (N_39326,N_31642,N_32953);
xor U39327 (N_39327,N_30354,N_32100);
nand U39328 (N_39328,N_31426,N_31201);
xnor U39329 (N_39329,N_33853,N_31754);
and U39330 (N_39330,N_34176,N_31002);
xor U39331 (N_39331,N_31915,N_30057);
nor U39332 (N_39332,N_30849,N_31693);
or U39333 (N_39333,N_32949,N_32721);
or U39334 (N_39334,N_31209,N_32255);
nor U39335 (N_39335,N_33637,N_34745);
or U39336 (N_39336,N_32926,N_31272);
nor U39337 (N_39337,N_33385,N_34653);
xnor U39338 (N_39338,N_32918,N_31838);
nand U39339 (N_39339,N_32398,N_34467);
and U39340 (N_39340,N_33882,N_30014);
or U39341 (N_39341,N_31550,N_34240);
or U39342 (N_39342,N_33385,N_33823);
nand U39343 (N_39343,N_32869,N_32301);
nand U39344 (N_39344,N_34325,N_30913);
or U39345 (N_39345,N_34775,N_30743);
nand U39346 (N_39346,N_31422,N_33207);
and U39347 (N_39347,N_34859,N_31376);
or U39348 (N_39348,N_31640,N_32459);
xor U39349 (N_39349,N_34275,N_33326);
and U39350 (N_39350,N_32552,N_32222);
and U39351 (N_39351,N_31119,N_31883);
nand U39352 (N_39352,N_34817,N_34717);
or U39353 (N_39353,N_31593,N_33848);
and U39354 (N_39354,N_34070,N_32569);
nor U39355 (N_39355,N_34127,N_31601);
or U39356 (N_39356,N_32477,N_34005);
and U39357 (N_39357,N_32860,N_31083);
nor U39358 (N_39358,N_31848,N_30129);
or U39359 (N_39359,N_31249,N_30821);
or U39360 (N_39360,N_34280,N_33141);
nand U39361 (N_39361,N_32839,N_32900);
and U39362 (N_39362,N_33923,N_30948);
or U39363 (N_39363,N_34197,N_30336);
and U39364 (N_39364,N_32081,N_30540);
or U39365 (N_39365,N_31051,N_31315);
or U39366 (N_39366,N_30894,N_33308);
and U39367 (N_39367,N_33496,N_34596);
and U39368 (N_39368,N_30145,N_33528);
nand U39369 (N_39369,N_30583,N_33757);
and U39370 (N_39370,N_34000,N_33305);
nor U39371 (N_39371,N_34451,N_33158);
and U39372 (N_39372,N_33254,N_31283);
and U39373 (N_39373,N_31646,N_30155);
xor U39374 (N_39374,N_33706,N_30149);
nor U39375 (N_39375,N_33564,N_33224);
and U39376 (N_39376,N_31270,N_30538);
nor U39377 (N_39377,N_33931,N_32921);
and U39378 (N_39378,N_34779,N_34123);
nand U39379 (N_39379,N_34664,N_30310);
and U39380 (N_39380,N_34356,N_32451);
nor U39381 (N_39381,N_32953,N_34387);
and U39382 (N_39382,N_34445,N_33757);
nor U39383 (N_39383,N_34652,N_33953);
xnor U39384 (N_39384,N_30759,N_30405);
nand U39385 (N_39385,N_31920,N_34230);
nor U39386 (N_39386,N_33203,N_30862);
nor U39387 (N_39387,N_33781,N_33614);
or U39388 (N_39388,N_30875,N_33244);
and U39389 (N_39389,N_34280,N_30952);
nand U39390 (N_39390,N_32105,N_31443);
or U39391 (N_39391,N_31335,N_34260);
xnor U39392 (N_39392,N_34518,N_33344);
nor U39393 (N_39393,N_33311,N_34226);
nor U39394 (N_39394,N_31300,N_32990);
xor U39395 (N_39395,N_33684,N_34494);
or U39396 (N_39396,N_30275,N_30427);
xor U39397 (N_39397,N_30758,N_32710);
xnor U39398 (N_39398,N_34487,N_31078);
xor U39399 (N_39399,N_30406,N_30074);
or U39400 (N_39400,N_30936,N_32894);
xnor U39401 (N_39401,N_32320,N_34506);
xor U39402 (N_39402,N_33289,N_33425);
nor U39403 (N_39403,N_34359,N_32086);
nand U39404 (N_39404,N_31556,N_31727);
and U39405 (N_39405,N_33741,N_34444);
or U39406 (N_39406,N_32977,N_31930);
nand U39407 (N_39407,N_34702,N_32853);
or U39408 (N_39408,N_30178,N_32014);
nor U39409 (N_39409,N_30799,N_30680);
nor U39410 (N_39410,N_34654,N_32951);
xnor U39411 (N_39411,N_30092,N_30357);
or U39412 (N_39412,N_33938,N_33460);
nand U39413 (N_39413,N_31882,N_32470);
nand U39414 (N_39414,N_30113,N_34979);
nor U39415 (N_39415,N_33657,N_33656);
nor U39416 (N_39416,N_34227,N_32980);
nor U39417 (N_39417,N_31125,N_34689);
xor U39418 (N_39418,N_34064,N_31928);
or U39419 (N_39419,N_31615,N_34283);
or U39420 (N_39420,N_33687,N_31709);
and U39421 (N_39421,N_32150,N_32381);
nor U39422 (N_39422,N_31255,N_30674);
or U39423 (N_39423,N_31738,N_32700);
or U39424 (N_39424,N_32762,N_31115);
and U39425 (N_39425,N_30711,N_31592);
nor U39426 (N_39426,N_32035,N_32601);
and U39427 (N_39427,N_31570,N_33808);
or U39428 (N_39428,N_32123,N_32655);
and U39429 (N_39429,N_32782,N_34305);
nand U39430 (N_39430,N_30047,N_33040);
xnor U39431 (N_39431,N_31654,N_30408);
nor U39432 (N_39432,N_31529,N_32221);
nor U39433 (N_39433,N_32289,N_31277);
or U39434 (N_39434,N_30986,N_34180);
nor U39435 (N_39435,N_30040,N_34434);
and U39436 (N_39436,N_33984,N_31785);
or U39437 (N_39437,N_33519,N_34502);
or U39438 (N_39438,N_34093,N_32146);
xnor U39439 (N_39439,N_30306,N_30900);
and U39440 (N_39440,N_30591,N_33736);
and U39441 (N_39441,N_31384,N_32510);
and U39442 (N_39442,N_32728,N_31622);
or U39443 (N_39443,N_34062,N_32084);
xnor U39444 (N_39444,N_32587,N_30043);
or U39445 (N_39445,N_34789,N_33664);
and U39446 (N_39446,N_34824,N_33946);
nor U39447 (N_39447,N_31012,N_32224);
nand U39448 (N_39448,N_33018,N_31649);
xnor U39449 (N_39449,N_31718,N_34364);
xnor U39450 (N_39450,N_33864,N_31734);
nand U39451 (N_39451,N_32294,N_32779);
nor U39452 (N_39452,N_32639,N_32790);
or U39453 (N_39453,N_31821,N_32610);
and U39454 (N_39454,N_34292,N_31907);
or U39455 (N_39455,N_33420,N_33232);
and U39456 (N_39456,N_33637,N_33915);
nor U39457 (N_39457,N_31736,N_33758);
xnor U39458 (N_39458,N_33111,N_33731);
nor U39459 (N_39459,N_30210,N_34102);
nor U39460 (N_39460,N_32588,N_31285);
or U39461 (N_39461,N_34251,N_32609);
and U39462 (N_39462,N_32140,N_31260);
or U39463 (N_39463,N_33869,N_30349);
or U39464 (N_39464,N_34371,N_31365);
xnor U39465 (N_39465,N_32476,N_30495);
nand U39466 (N_39466,N_32520,N_30217);
or U39467 (N_39467,N_31041,N_32356);
nor U39468 (N_39468,N_32217,N_31226);
and U39469 (N_39469,N_33203,N_31392);
or U39470 (N_39470,N_31378,N_32161);
or U39471 (N_39471,N_31506,N_30719);
nor U39472 (N_39472,N_33974,N_30893);
nor U39473 (N_39473,N_32789,N_32694);
nand U39474 (N_39474,N_31410,N_30627);
and U39475 (N_39475,N_34674,N_33501);
nor U39476 (N_39476,N_30269,N_34403);
and U39477 (N_39477,N_34255,N_33003);
or U39478 (N_39478,N_34467,N_33969);
and U39479 (N_39479,N_30080,N_34629);
and U39480 (N_39480,N_30038,N_34300);
and U39481 (N_39481,N_31621,N_30279);
or U39482 (N_39482,N_30886,N_33063);
nor U39483 (N_39483,N_32754,N_33808);
nor U39484 (N_39484,N_31530,N_32937);
and U39485 (N_39485,N_33229,N_30880);
nor U39486 (N_39486,N_32952,N_31743);
nand U39487 (N_39487,N_30018,N_33011);
and U39488 (N_39488,N_30094,N_32191);
nor U39489 (N_39489,N_34003,N_34032);
or U39490 (N_39490,N_31865,N_33585);
nand U39491 (N_39491,N_33264,N_33680);
or U39492 (N_39492,N_30333,N_33305);
and U39493 (N_39493,N_34442,N_31233);
and U39494 (N_39494,N_32905,N_30244);
nand U39495 (N_39495,N_31414,N_30746);
nor U39496 (N_39496,N_33877,N_34076);
xnor U39497 (N_39497,N_33529,N_32537);
nand U39498 (N_39498,N_30383,N_30204);
or U39499 (N_39499,N_34681,N_32828);
nand U39500 (N_39500,N_32435,N_31599);
nor U39501 (N_39501,N_33134,N_32618);
nand U39502 (N_39502,N_32351,N_34682);
nand U39503 (N_39503,N_30196,N_34482);
nor U39504 (N_39504,N_31838,N_31796);
nand U39505 (N_39505,N_33674,N_32450);
or U39506 (N_39506,N_31308,N_33754);
and U39507 (N_39507,N_34237,N_30869);
nand U39508 (N_39508,N_34196,N_31034);
or U39509 (N_39509,N_31788,N_33256);
nand U39510 (N_39510,N_33791,N_32416);
nand U39511 (N_39511,N_31167,N_30651);
nor U39512 (N_39512,N_32026,N_34207);
nor U39513 (N_39513,N_33156,N_31910);
and U39514 (N_39514,N_34221,N_32536);
nand U39515 (N_39515,N_34772,N_30855);
nand U39516 (N_39516,N_31528,N_31982);
xnor U39517 (N_39517,N_33979,N_30930);
nand U39518 (N_39518,N_33738,N_32512);
and U39519 (N_39519,N_30366,N_34259);
nor U39520 (N_39520,N_31883,N_33216);
or U39521 (N_39521,N_31987,N_31151);
and U39522 (N_39522,N_31312,N_30481);
nand U39523 (N_39523,N_32012,N_31457);
and U39524 (N_39524,N_31147,N_30959);
nand U39525 (N_39525,N_31299,N_34447);
nand U39526 (N_39526,N_33671,N_32821);
or U39527 (N_39527,N_31422,N_32119);
nor U39528 (N_39528,N_33771,N_31184);
nand U39529 (N_39529,N_32226,N_32091);
or U39530 (N_39530,N_34979,N_33429);
or U39531 (N_39531,N_34147,N_30500);
nor U39532 (N_39532,N_33345,N_30259);
or U39533 (N_39533,N_32711,N_33832);
and U39534 (N_39534,N_34919,N_30613);
or U39535 (N_39535,N_34440,N_32121);
or U39536 (N_39536,N_32158,N_30769);
nor U39537 (N_39537,N_34583,N_31868);
xor U39538 (N_39538,N_34135,N_30783);
nor U39539 (N_39539,N_30507,N_34157);
nand U39540 (N_39540,N_32103,N_30993);
xor U39541 (N_39541,N_30905,N_32819);
nand U39542 (N_39542,N_33321,N_30277);
xor U39543 (N_39543,N_34712,N_30194);
or U39544 (N_39544,N_34039,N_32532);
nand U39545 (N_39545,N_30949,N_30769);
nand U39546 (N_39546,N_30840,N_30205);
nand U39547 (N_39547,N_32649,N_32820);
and U39548 (N_39548,N_32910,N_33270);
xnor U39549 (N_39549,N_33636,N_33787);
nand U39550 (N_39550,N_30529,N_31791);
or U39551 (N_39551,N_30084,N_33288);
nand U39552 (N_39552,N_31260,N_31850);
nor U39553 (N_39553,N_31417,N_31317);
nor U39554 (N_39554,N_34648,N_32329);
and U39555 (N_39555,N_31769,N_30213);
or U39556 (N_39556,N_33271,N_32960);
and U39557 (N_39557,N_30418,N_33978);
xnor U39558 (N_39558,N_33794,N_34575);
or U39559 (N_39559,N_32987,N_34902);
or U39560 (N_39560,N_32963,N_33025);
or U39561 (N_39561,N_31934,N_31134);
nand U39562 (N_39562,N_32378,N_31288);
or U39563 (N_39563,N_31797,N_30238);
and U39564 (N_39564,N_34357,N_30148);
and U39565 (N_39565,N_31585,N_34571);
or U39566 (N_39566,N_32149,N_33408);
or U39567 (N_39567,N_33632,N_34020);
and U39568 (N_39568,N_30432,N_33740);
nor U39569 (N_39569,N_31625,N_31565);
or U39570 (N_39570,N_33124,N_34456);
nor U39571 (N_39571,N_31254,N_31064);
or U39572 (N_39572,N_33896,N_32102);
nand U39573 (N_39573,N_32240,N_32981);
and U39574 (N_39574,N_34578,N_30280);
or U39575 (N_39575,N_32558,N_33906);
and U39576 (N_39576,N_33925,N_33900);
nand U39577 (N_39577,N_32522,N_31962);
or U39578 (N_39578,N_34951,N_33692);
or U39579 (N_39579,N_34258,N_33959);
xnor U39580 (N_39580,N_31753,N_32364);
or U39581 (N_39581,N_30918,N_31829);
xnor U39582 (N_39582,N_31303,N_32049);
nor U39583 (N_39583,N_31934,N_32626);
nand U39584 (N_39584,N_33586,N_34557);
nor U39585 (N_39585,N_32230,N_33761);
xor U39586 (N_39586,N_34498,N_30461);
xor U39587 (N_39587,N_34594,N_31606);
nand U39588 (N_39588,N_32413,N_32195);
and U39589 (N_39589,N_31151,N_32542);
nand U39590 (N_39590,N_34725,N_33597);
or U39591 (N_39591,N_32369,N_34445);
and U39592 (N_39592,N_32554,N_32474);
or U39593 (N_39593,N_32647,N_30692);
xnor U39594 (N_39594,N_33119,N_32908);
or U39595 (N_39595,N_34534,N_34258);
and U39596 (N_39596,N_32995,N_31792);
nand U39597 (N_39597,N_34956,N_33581);
nand U39598 (N_39598,N_33969,N_30222);
or U39599 (N_39599,N_30608,N_30693);
and U39600 (N_39600,N_32795,N_33232);
and U39601 (N_39601,N_33758,N_31991);
or U39602 (N_39602,N_31273,N_31892);
nand U39603 (N_39603,N_34644,N_34628);
and U39604 (N_39604,N_34047,N_30755);
or U39605 (N_39605,N_31925,N_34846);
or U39606 (N_39606,N_32637,N_32821);
and U39607 (N_39607,N_31458,N_33599);
or U39608 (N_39608,N_31285,N_30437);
or U39609 (N_39609,N_34377,N_34470);
nand U39610 (N_39610,N_34290,N_32497);
or U39611 (N_39611,N_30647,N_31253);
and U39612 (N_39612,N_30585,N_31831);
nand U39613 (N_39613,N_34176,N_32665);
nor U39614 (N_39614,N_31305,N_32325);
nor U39615 (N_39615,N_31519,N_30414);
and U39616 (N_39616,N_34838,N_30718);
nand U39617 (N_39617,N_33087,N_31455);
nand U39618 (N_39618,N_30120,N_30306);
or U39619 (N_39619,N_33548,N_30098);
nor U39620 (N_39620,N_32568,N_32510);
nor U39621 (N_39621,N_33744,N_33373);
and U39622 (N_39622,N_34761,N_30128);
or U39623 (N_39623,N_31893,N_33254);
and U39624 (N_39624,N_32784,N_34031);
xor U39625 (N_39625,N_34244,N_32385);
nand U39626 (N_39626,N_34328,N_32453);
or U39627 (N_39627,N_31964,N_31682);
nand U39628 (N_39628,N_33426,N_31914);
and U39629 (N_39629,N_30851,N_32485);
xnor U39630 (N_39630,N_31822,N_33766);
or U39631 (N_39631,N_30810,N_30035);
nand U39632 (N_39632,N_32285,N_34666);
nor U39633 (N_39633,N_33795,N_31874);
nand U39634 (N_39634,N_34560,N_34641);
nand U39635 (N_39635,N_33314,N_34940);
nor U39636 (N_39636,N_31186,N_31266);
and U39637 (N_39637,N_33865,N_34089);
nor U39638 (N_39638,N_32640,N_31110);
nor U39639 (N_39639,N_30349,N_30122);
and U39640 (N_39640,N_33442,N_32623);
or U39641 (N_39641,N_30687,N_33011);
nand U39642 (N_39642,N_32349,N_31897);
nand U39643 (N_39643,N_33351,N_34094);
or U39644 (N_39644,N_32728,N_33574);
or U39645 (N_39645,N_31953,N_33562);
nor U39646 (N_39646,N_31889,N_34422);
nand U39647 (N_39647,N_32871,N_30161);
nor U39648 (N_39648,N_31448,N_32438);
nand U39649 (N_39649,N_31785,N_33914);
and U39650 (N_39650,N_31746,N_33584);
nand U39651 (N_39651,N_32738,N_33205);
nand U39652 (N_39652,N_30206,N_31199);
nand U39653 (N_39653,N_31344,N_34963);
and U39654 (N_39654,N_31707,N_33691);
nand U39655 (N_39655,N_30801,N_32143);
nand U39656 (N_39656,N_34060,N_30652);
nor U39657 (N_39657,N_31767,N_30120);
or U39658 (N_39658,N_30577,N_34900);
nand U39659 (N_39659,N_31752,N_30592);
or U39660 (N_39660,N_33687,N_31046);
nor U39661 (N_39661,N_33980,N_31409);
and U39662 (N_39662,N_32199,N_33356);
nand U39663 (N_39663,N_34463,N_30698);
nand U39664 (N_39664,N_34209,N_32576);
xnor U39665 (N_39665,N_30427,N_30842);
or U39666 (N_39666,N_30966,N_34066);
nor U39667 (N_39667,N_31446,N_31628);
nand U39668 (N_39668,N_30061,N_32663);
and U39669 (N_39669,N_34378,N_32534);
nand U39670 (N_39670,N_34030,N_31574);
or U39671 (N_39671,N_33393,N_32649);
and U39672 (N_39672,N_32625,N_34786);
nand U39673 (N_39673,N_33791,N_34187);
nand U39674 (N_39674,N_30122,N_33295);
or U39675 (N_39675,N_33076,N_31301);
nor U39676 (N_39676,N_34098,N_34200);
or U39677 (N_39677,N_30602,N_34827);
and U39678 (N_39678,N_34284,N_34373);
and U39679 (N_39679,N_34568,N_33909);
nor U39680 (N_39680,N_33936,N_32265);
nor U39681 (N_39681,N_31954,N_31779);
or U39682 (N_39682,N_30326,N_32734);
or U39683 (N_39683,N_31917,N_32941);
or U39684 (N_39684,N_31188,N_30481);
and U39685 (N_39685,N_32610,N_33421);
or U39686 (N_39686,N_31954,N_30995);
or U39687 (N_39687,N_31996,N_31012);
or U39688 (N_39688,N_33066,N_33336);
and U39689 (N_39689,N_32422,N_34705);
and U39690 (N_39690,N_30177,N_34977);
and U39691 (N_39691,N_34141,N_31217);
xnor U39692 (N_39692,N_30500,N_32340);
nor U39693 (N_39693,N_34011,N_34374);
nand U39694 (N_39694,N_31088,N_34492);
nor U39695 (N_39695,N_31451,N_30477);
xnor U39696 (N_39696,N_33066,N_31390);
nand U39697 (N_39697,N_30804,N_32087);
nor U39698 (N_39698,N_32397,N_31750);
and U39699 (N_39699,N_34077,N_34350);
nand U39700 (N_39700,N_31821,N_33611);
and U39701 (N_39701,N_32913,N_34992);
and U39702 (N_39702,N_33711,N_33358);
and U39703 (N_39703,N_30440,N_34038);
xnor U39704 (N_39704,N_33159,N_32694);
nor U39705 (N_39705,N_31483,N_32551);
and U39706 (N_39706,N_32798,N_34849);
nor U39707 (N_39707,N_32853,N_32701);
or U39708 (N_39708,N_31061,N_32994);
and U39709 (N_39709,N_33025,N_34031);
and U39710 (N_39710,N_31962,N_31115);
nand U39711 (N_39711,N_30630,N_30060);
nor U39712 (N_39712,N_33448,N_32004);
xnor U39713 (N_39713,N_32595,N_31002);
nand U39714 (N_39714,N_31204,N_31605);
and U39715 (N_39715,N_33065,N_33315);
nand U39716 (N_39716,N_33583,N_31525);
or U39717 (N_39717,N_32864,N_31058);
nor U39718 (N_39718,N_31255,N_32021);
nand U39719 (N_39719,N_34439,N_31482);
nand U39720 (N_39720,N_34030,N_31724);
nor U39721 (N_39721,N_32833,N_32699);
or U39722 (N_39722,N_31148,N_31066);
xnor U39723 (N_39723,N_32037,N_32767);
or U39724 (N_39724,N_34168,N_32698);
and U39725 (N_39725,N_33236,N_32037);
and U39726 (N_39726,N_31150,N_34533);
nor U39727 (N_39727,N_31293,N_33962);
nor U39728 (N_39728,N_34242,N_33500);
nor U39729 (N_39729,N_30997,N_33744);
xor U39730 (N_39730,N_32802,N_33141);
nand U39731 (N_39731,N_30905,N_31897);
and U39732 (N_39732,N_31242,N_31274);
nand U39733 (N_39733,N_31546,N_34781);
and U39734 (N_39734,N_33805,N_30821);
xnor U39735 (N_39735,N_33593,N_30670);
nor U39736 (N_39736,N_31721,N_34994);
nor U39737 (N_39737,N_31787,N_34418);
or U39738 (N_39738,N_32144,N_33063);
nand U39739 (N_39739,N_31232,N_31143);
and U39740 (N_39740,N_30232,N_31853);
nor U39741 (N_39741,N_30851,N_34320);
nor U39742 (N_39742,N_33455,N_34816);
and U39743 (N_39743,N_30364,N_30731);
and U39744 (N_39744,N_32569,N_31368);
and U39745 (N_39745,N_31639,N_31811);
and U39746 (N_39746,N_33135,N_33874);
nand U39747 (N_39747,N_33710,N_32776);
nor U39748 (N_39748,N_31353,N_30031);
or U39749 (N_39749,N_31632,N_31576);
or U39750 (N_39750,N_30132,N_31547);
nand U39751 (N_39751,N_33613,N_34542);
and U39752 (N_39752,N_32994,N_33930);
nor U39753 (N_39753,N_32513,N_33831);
xnor U39754 (N_39754,N_34750,N_30792);
and U39755 (N_39755,N_31374,N_33730);
and U39756 (N_39756,N_34316,N_30998);
nand U39757 (N_39757,N_30054,N_34215);
and U39758 (N_39758,N_34927,N_31565);
or U39759 (N_39759,N_34766,N_33433);
nand U39760 (N_39760,N_32304,N_31706);
or U39761 (N_39761,N_31298,N_34596);
and U39762 (N_39762,N_30625,N_33783);
nor U39763 (N_39763,N_32518,N_33433);
nor U39764 (N_39764,N_31386,N_31132);
nor U39765 (N_39765,N_34185,N_31570);
nand U39766 (N_39766,N_32058,N_34281);
nor U39767 (N_39767,N_33978,N_34896);
nor U39768 (N_39768,N_33206,N_32705);
or U39769 (N_39769,N_34929,N_34140);
xnor U39770 (N_39770,N_33487,N_31815);
xor U39771 (N_39771,N_30085,N_31962);
or U39772 (N_39772,N_30361,N_32532);
nor U39773 (N_39773,N_31875,N_34120);
or U39774 (N_39774,N_33069,N_30035);
and U39775 (N_39775,N_32955,N_32186);
and U39776 (N_39776,N_33698,N_33941);
and U39777 (N_39777,N_33850,N_33810);
nor U39778 (N_39778,N_33215,N_31327);
nand U39779 (N_39779,N_34052,N_31449);
or U39780 (N_39780,N_32131,N_30704);
or U39781 (N_39781,N_33807,N_31409);
xor U39782 (N_39782,N_30573,N_32386);
and U39783 (N_39783,N_32031,N_31217);
nor U39784 (N_39784,N_31271,N_31678);
nand U39785 (N_39785,N_31148,N_30455);
nand U39786 (N_39786,N_34431,N_32741);
or U39787 (N_39787,N_33599,N_32815);
and U39788 (N_39788,N_33750,N_30449);
nor U39789 (N_39789,N_30049,N_34566);
or U39790 (N_39790,N_32278,N_32352);
and U39791 (N_39791,N_30708,N_32139);
nor U39792 (N_39792,N_31283,N_34085);
nand U39793 (N_39793,N_32897,N_32337);
nor U39794 (N_39794,N_31233,N_30424);
and U39795 (N_39795,N_34364,N_31055);
and U39796 (N_39796,N_32799,N_30376);
nand U39797 (N_39797,N_32343,N_30502);
nand U39798 (N_39798,N_32185,N_30819);
or U39799 (N_39799,N_32962,N_31521);
nand U39800 (N_39800,N_34107,N_33493);
and U39801 (N_39801,N_32951,N_34954);
or U39802 (N_39802,N_32936,N_33596);
xor U39803 (N_39803,N_31846,N_34489);
nand U39804 (N_39804,N_34208,N_34027);
or U39805 (N_39805,N_31076,N_32645);
nand U39806 (N_39806,N_31256,N_32429);
xnor U39807 (N_39807,N_34533,N_30005);
nor U39808 (N_39808,N_34453,N_30304);
nor U39809 (N_39809,N_33211,N_32652);
or U39810 (N_39810,N_33310,N_32282);
and U39811 (N_39811,N_34754,N_33155);
nand U39812 (N_39812,N_30298,N_32688);
or U39813 (N_39813,N_31701,N_33703);
nand U39814 (N_39814,N_33560,N_34613);
nand U39815 (N_39815,N_31046,N_32086);
and U39816 (N_39816,N_32054,N_31990);
xnor U39817 (N_39817,N_30542,N_34010);
nand U39818 (N_39818,N_30370,N_32563);
xor U39819 (N_39819,N_30946,N_33878);
or U39820 (N_39820,N_32151,N_30763);
nand U39821 (N_39821,N_33644,N_32177);
or U39822 (N_39822,N_33885,N_32352);
nor U39823 (N_39823,N_31027,N_31774);
nor U39824 (N_39824,N_30748,N_30645);
or U39825 (N_39825,N_32674,N_33131);
and U39826 (N_39826,N_33353,N_34044);
and U39827 (N_39827,N_30655,N_31843);
nor U39828 (N_39828,N_31789,N_31937);
and U39829 (N_39829,N_32825,N_30285);
nand U39830 (N_39830,N_34385,N_34492);
nand U39831 (N_39831,N_32016,N_30250);
or U39832 (N_39832,N_32530,N_31490);
or U39833 (N_39833,N_31683,N_34085);
xnor U39834 (N_39834,N_34520,N_31028);
and U39835 (N_39835,N_32299,N_32464);
and U39836 (N_39836,N_30356,N_34835);
or U39837 (N_39837,N_31522,N_34631);
nor U39838 (N_39838,N_31252,N_31475);
or U39839 (N_39839,N_32129,N_34712);
or U39840 (N_39840,N_30450,N_30352);
xnor U39841 (N_39841,N_30743,N_34715);
or U39842 (N_39842,N_34393,N_31513);
or U39843 (N_39843,N_34697,N_34072);
or U39844 (N_39844,N_30673,N_34986);
and U39845 (N_39845,N_34812,N_33951);
nand U39846 (N_39846,N_32763,N_32368);
nand U39847 (N_39847,N_30045,N_31389);
xor U39848 (N_39848,N_31882,N_30530);
nor U39849 (N_39849,N_32874,N_34195);
nand U39850 (N_39850,N_33230,N_30605);
xor U39851 (N_39851,N_33218,N_33171);
nand U39852 (N_39852,N_33105,N_32930);
or U39853 (N_39853,N_31071,N_33996);
and U39854 (N_39854,N_34831,N_32050);
nor U39855 (N_39855,N_32807,N_31238);
or U39856 (N_39856,N_31795,N_31925);
nor U39857 (N_39857,N_31732,N_33779);
and U39858 (N_39858,N_32840,N_33802);
nor U39859 (N_39859,N_33871,N_32183);
or U39860 (N_39860,N_31146,N_34638);
and U39861 (N_39861,N_31833,N_31582);
xor U39862 (N_39862,N_34950,N_30656);
nor U39863 (N_39863,N_34980,N_32903);
and U39864 (N_39864,N_33803,N_30774);
nand U39865 (N_39865,N_33044,N_32792);
nand U39866 (N_39866,N_30151,N_33418);
nand U39867 (N_39867,N_33125,N_32501);
and U39868 (N_39868,N_30077,N_33235);
or U39869 (N_39869,N_31253,N_33128);
nor U39870 (N_39870,N_30078,N_34065);
and U39871 (N_39871,N_34144,N_33847);
and U39872 (N_39872,N_33539,N_33212);
nor U39873 (N_39873,N_33444,N_31912);
nor U39874 (N_39874,N_30356,N_33449);
or U39875 (N_39875,N_33181,N_34884);
nor U39876 (N_39876,N_32970,N_31188);
and U39877 (N_39877,N_32193,N_34543);
or U39878 (N_39878,N_31097,N_32083);
nand U39879 (N_39879,N_31677,N_32024);
and U39880 (N_39880,N_32679,N_32682);
or U39881 (N_39881,N_33220,N_32345);
nand U39882 (N_39882,N_31714,N_31913);
nand U39883 (N_39883,N_33515,N_31522);
nand U39884 (N_39884,N_30472,N_32485);
nand U39885 (N_39885,N_32780,N_33222);
and U39886 (N_39886,N_34811,N_31742);
or U39887 (N_39887,N_31190,N_32315);
and U39888 (N_39888,N_31435,N_31962);
and U39889 (N_39889,N_34312,N_33662);
nand U39890 (N_39890,N_31853,N_31783);
nor U39891 (N_39891,N_33569,N_33143);
and U39892 (N_39892,N_33076,N_31795);
or U39893 (N_39893,N_34402,N_32155);
and U39894 (N_39894,N_31606,N_33097);
or U39895 (N_39895,N_30068,N_32666);
nor U39896 (N_39896,N_30928,N_34591);
nand U39897 (N_39897,N_33696,N_33974);
and U39898 (N_39898,N_31423,N_31653);
or U39899 (N_39899,N_34914,N_30550);
nand U39900 (N_39900,N_32055,N_30890);
and U39901 (N_39901,N_32203,N_32546);
or U39902 (N_39902,N_34696,N_32378);
nor U39903 (N_39903,N_33244,N_32457);
xnor U39904 (N_39904,N_30323,N_34264);
nor U39905 (N_39905,N_31008,N_30498);
xnor U39906 (N_39906,N_30682,N_31149);
and U39907 (N_39907,N_32278,N_30710);
and U39908 (N_39908,N_30050,N_34871);
nor U39909 (N_39909,N_34108,N_34337);
or U39910 (N_39910,N_34591,N_33757);
xor U39911 (N_39911,N_34274,N_30869);
and U39912 (N_39912,N_31185,N_30628);
nand U39913 (N_39913,N_30424,N_33056);
and U39914 (N_39914,N_31998,N_33598);
or U39915 (N_39915,N_34534,N_34578);
nand U39916 (N_39916,N_32660,N_31638);
nor U39917 (N_39917,N_33327,N_31551);
and U39918 (N_39918,N_32283,N_30957);
or U39919 (N_39919,N_34623,N_30968);
xnor U39920 (N_39920,N_30567,N_30677);
xnor U39921 (N_39921,N_33628,N_32945);
or U39922 (N_39922,N_34831,N_34956);
and U39923 (N_39923,N_34647,N_30738);
or U39924 (N_39924,N_33738,N_31263);
nand U39925 (N_39925,N_33004,N_33928);
or U39926 (N_39926,N_32295,N_34057);
nand U39927 (N_39927,N_32409,N_30451);
and U39928 (N_39928,N_33313,N_33280);
or U39929 (N_39929,N_31127,N_33400);
nand U39930 (N_39930,N_34635,N_33924);
or U39931 (N_39931,N_31139,N_31266);
nor U39932 (N_39932,N_34343,N_30582);
nor U39933 (N_39933,N_34674,N_31600);
nand U39934 (N_39934,N_33401,N_33497);
and U39935 (N_39935,N_30825,N_33884);
and U39936 (N_39936,N_30248,N_34656);
nor U39937 (N_39937,N_30663,N_34401);
and U39938 (N_39938,N_32821,N_34424);
or U39939 (N_39939,N_32732,N_32638);
nand U39940 (N_39940,N_32533,N_30644);
nand U39941 (N_39941,N_31811,N_32593);
nor U39942 (N_39942,N_32000,N_31254);
and U39943 (N_39943,N_31048,N_33820);
nand U39944 (N_39944,N_31127,N_34723);
and U39945 (N_39945,N_32776,N_30646);
nor U39946 (N_39946,N_30365,N_31971);
or U39947 (N_39947,N_33604,N_30235);
xor U39948 (N_39948,N_32757,N_32727);
xor U39949 (N_39949,N_30963,N_31423);
xor U39950 (N_39950,N_30157,N_31670);
or U39951 (N_39951,N_31600,N_34041);
nor U39952 (N_39952,N_32121,N_33295);
nand U39953 (N_39953,N_30352,N_32832);
nor U39954 (N_39954,N_30909,N_33271);
nor U39955 (N_39955,N_30146,N_33129);
or U39956 (N_39956,N_34666,N_30308);
nand U39957 (N_39957,N_30294,N_31161);
nand U39958 (N_39958,N_34038,N_31759);
and U39959 (N_39959,N_33512,N_32544);
nor U39960 (N_39960,N_33193,N_30778);
nand U39961 (N_39961,N_31161,N_34471);
nand U39962 (N_39962,N_33116,N_34502);
and U39963 (N_39963,N_32559,N_34220);
nor U39964 (N_39964,N_30984,N_33034);
nand U39965 (N_39965,N_34360,N_32460);
or U39966 (N_39966,N_34362,N_32548);
or U39967 (N_39967,N_34009,N_31202);
nand U39968 (N_39968,N_30021,N_33269);
nor U39969 (N_39969,N_31977,N_30787);
nor U39970 (N_39970,N_32888,N_32079);
nand U39971 (N_39971,N_32214,N_31213);
nor U39972 (N_39972,N_30993,N_31548);
and U39973 (N_39973,N_32836,N_34512);
nand U39974 (N_39974,N_32619,N_32394);
nand U39975 (N_39975,N_32944,N_30526);
nor U39976 (N_39976,N_33628,N_33204);
xor U39977 (N_39977,N_34666,N_30159);
or U39978 (N_39978,N_30299,N_34930);
and U39979 (N_39979,N_32541,N_31681);
and U39980 (N_39980,N_33973,N_33098);
nand U39981 (N_39981,N_30734,N_32678);
and U39982 (N_39982,N_34674,N_32225);
and U39983 (N_39983,N_33781,N_30292);
nand U39984 (N_39984,N_30582,N_32400);
or U39985 (N_39985,N_33174,N_33122);
nor U39986 (N_39986,N_34876,N_34610);
and U39987 (N_39987,N_33115,N_31687);
nand U39988 (N_39988,N_34947,N_31818);
nand U39989 (N_39989,N_34023,N_31616);
nor U39990 (N_39990,N_30194,N_30555);
and U39991 (N_39991,N_32846,N_30985);
and U39992 (N_39992,N_34628,N_30338);
nor U39993 (N_39993,N_33833,N_31470);
nand U39994 (N_39994,N_31756,N_33492);
nor U39995 (N_39995,N_34884,N_31336);
nor U39996 (N_39996,N_33432,N_30022);
nor U39997 (N_39997,N_30692,N_30127);
nor U39998 (N_39998,N_31702,N_31091);
and U39999 (N_39999,N_33409,N_30035);
xnor U40000 (N_40000,N_38753,N_39456);
nand U40001 (N_40001,N_36779,N_39419);
or U40002 (N_40002,N_37965,N_35910);
or U40003 (N_40003,N_38198,N_35329);
nand U40004 (N_40004,N_37885,N_35141);
nand U40005 (N_40005,N_35229,N_38965);
nor U40006 (N_40006,N_38031,N_35855);
xnor U40007 (N_40007,N_35864,N_37998);
or U40008 (N_40008,N_35734,N_39748);
and U40009 (N_40009,N_36632,N_39780);
and U40010 (N_40010,N_39195,N_38448);
xnor U40011 (N_40011,N_39186,N_36511);
nor U40012 (N_40012,N_37544,N_37235);
or U40013 (N_40013,N_35072,N_35677);
nor U40014 (N_40014,N_35820,N_37204);
nor U40015 (N_40015,N_39513,N_35196);
nand U40016 (N_40016,N_36650,N_37445);
and U40017 (N_40017,N_39343,N_36372);
or U40018 (N_40018,N_36721,N_39175);
nor U40019 (N_40019,N_37761,N_38558);
nand U40020 (N_40020,N_39486,N_37663);
nor U40021 (N_40021,N_38065,N_39709);
nand U40022 (N_40022,N_37936,N_37193);
xor U40023 (N_40023,N_36738,N_37304);
nor U40024 (N_40024,N_38902,N_37215);
nor U40025 (N_40025,N_39638,N_38266);
xor U40026 (N_40026,N_37924,N_38102);
or U40027 (N_40027,N_38204,N_38899);
or U40028 (N_40028,N_37608,N_35756);
or U40029 (N_40029,N_36853,N_36197);
and U40030 (N_40030,N_38919,N_35180);
and U40031 (N_40031,N_37670,N_39432);
or U40032 (N_40032,N_38110,N_39968);
nand U40033 (N_40033,N_38386,N_37653);
and U40034 (N_40034,N_36232,N_38949);
xor U40035 (N_40035,N_35256,N_37527);
and U40036 (N_40036,N_37941,N_36841);
nand U40037 (N_40037,N_38005,N_35553);
or U40038 (N_40038,N_36868,N_37805);
nor U40039 (N_40039,N_37351,N_36183);
nor U40040 (N_40040,N_39753,N_35304);
xnor U40041 (N_40041,N_39276,N_36475);
and U40042 (N_40042,N_35242,N_38347);
or U40043 (N_40043,N_35411,N_35981);
and U40044 (N_40044,N_37757,N_39037);
nand U40045 (N_40045,N_36058,N_39939);
nor U40046 (N_40046,N_36393,N_35453);
nor U40047 (N_40047,N_35599,N_37562);
nand U40048 (N_40048,N_36057,N_39352);
and U40049 (N_40049,N_37706,N_39291);
or U40050 (N_40050,N_37514,N_39478);
nor U40051 (N_40051,N_35047,N_35994);
and U40052 (N_40052,N_36077,N_36992);
nor U40053 (N_40053,N_39153,N_39068);
or U40054 (N_40054,N_39604,N_37388);
and U40055 (N_40055,N_39878,N_35851);
nor U40056 (N_40056,N_35414,N_37600);
nor U40057 (N_40057,N_37389,N_36777);
xnor U40058 (N_40058,N_38549,N_37901);
or U40059 (N_40059,N_35446,N_36244);
nor U40060 (N_40060,N_39913,N_39231);
and U40061 (N_40061,N_35257,N_35381);
or U40062 (N_40062,N_39362,N_39140);
or U40063 (N_40063,N_35836,N_38015);
or U40064 (N_40064,N_38686,N_35771);
or U40065 (N_40065,N_35829,N_39090);
xor U40066 (N_40066,N_38675,N_37201);
nand U40067 (N_40067,N_39577,N_39468);
or U40068 (N_40068,N_38539,N_37289);
and U40069 (N_40069,N_35164,N_36881);
nor U40070 (N_40070,N_35117,N_38837);
and U40071 (N_40071,N_39514,N_38817);
xnor U40072 (N_40072,N_38037,N_37371);
nor U40073 (N_40073,N_35083,N_39793);
and U40074 (N_40074,N_35785,N_36949);
or U40075 (N_40075,N_36552,N_39387);
or U40076 (N_40076,N_39644,N_36678);
or U40077 (N_40077,N_37742,N_35236);
and U40078 (N_40078,N_39457,N_37962);
or U40079 (N_40079,N_36256,N_35189);
or U40080 (N_40080,N_38116,N_35584);
and U40081 (N_40081,N_36640,N_36139);
nor U40082 (N_40082,N_37881,N_37124);
nor U40083 (N_40083,N_35374,N_39842);
or U40084 (N_40084,N_35992,N_35560);
nor U40085 (N_40085,N_37749,N_36609);
nand U40086 (N_40086,N_35642,N_36491);
or U40087 (N_40087,N_36285,N_36998);
nor U40088 (N_40088,N_35922,N_35426);
or U40089 (N_40089,N_39379,N_35106);
nor U40090 (N_40090,N_37430,N_39081);
nor U40091 (N_40091,N_38107,N_37584);
nor U40092 (N_40092,N_37700,N_38618);
nor U40093 (N_40093,N_39716,N_39874);
nor U40094 (N_40094,N_36110,N_38332);
xnor U40095 (N_40095,N_38134,N_36108);
and U40096 (N_40096,N_35863,N_39070);
or U40097 (N_40097,N_37348,N_39377);
nand U40098 (N_40098,N_35755,N_38971);
nand U40099 (N_40099,N_37482,N_39242);
nor U40100 (N_40100,N_35975,N_36990);
or U40101 (N_40101,N_38123,N_36870);
nand U40102 (N_40102,N_38795,N_37084);
nand U40103 (N_40103,N_39161,N_37104);
or U40104 (N_40104,N_39394,N_37303);
nor U40105 (N_40105,N_38727,N_37766);
and U40106 (N_40106,N_37362,N_39662);
and U40107 (N_40107,N_39006,N_37080);
or U40108 (N_40108,N_36905,N_35684);
or U40109 (N_40109,N_37202,N_39307);
and U40110 (N_40110,N_38423,N_37739);
and U40111 (N_40111,N_38540,N_37571);
and U40112 (N_40112,N_36846,N_38158);
and U40113 (N_40113,N_38024,N_37787);
or U40114 (N_40114,N_37100,N_39616);
nand U40115 (N_40115,N_39687,N_38950);
nor U40116 (N_40116,N_35669,N_37838);
nand U40117 (N_40117,N_36874,N_35693);
and U40118 (N_40118,N_36278,N_37411);
and U40119 (N_40119,N_36324,N_39071);
nand U40120 (N_40120,N_35650,N_38963);
nand U40121 (N_40121,N_39091,N_39851);
or U40122 (N_40122,N_37230,N_39578);
nand U40123 (N_40123,N_37576,N_38997);
nor U40124 (N_40124,N_37790,N_37505);
and U40125 (N_40125,N_38062,N_36843);
nor U40126 (N_40126,N_37341,N_35935);
nor U40127 (N_40127,N_39283,N_37909);
nand U40128 (N_40128,N_37454,N_37317);
nand U40129 (N_40129,N_37444,N_37532);
nand U40130 (N_40130,N_38688,N_37218);
or U40131 (N_40131,N_36923,N_38537);
and U40132 (N_40132,N_36961,N_36298);
nand U40133 (N_40133,N_36249,N_36999);
or U40134 (N_40134,N_38479,N_37840);
and U40135 (N_40135,N_37123,N_35744);
nor U40136 (N_40136,N_35831,N_38330);
nand U40137 (N_40137,N_39656,N_36595);
and U40138 (N_40138,N_36798,N_38086);
or U40139 (N_40139,N_37814,N_39522);
and U40140 (N_40140,N_39477,N_39686);
nor U40141 (N_40141,N_35574,N_38509);
and U40142 (N_40142,N_38691,N_36412);
nor U40143 (N_40143,N_35258,N_36492);
nand U40144 (N_40144,N_37067,N_38040);
and U40145 (N_40145,N_37301,N_39722);
or U40146 (N_40146,N_36011,N_39765);
xnor U40147 (N_40147,N_35228,N_38981);
or U40148 (N_40148,N_38173,N_39712);
xor U40149 (N_40149,N_38326,N_37117);
nor U40150 (N_40150,N_36126,N_38584);
nand U40151 (N_40151,N_35046,N_37643);
and U40152 (N_40152,N_35812,N_39932);
or U40153 (N_40153,N_39378,N_37113);
nand U40154 (N_40154,N_37287,N_37929);
and U40155 (N_40155,N_38576,N_37645);
or U40156 (N_40156,N_35240,N_35463);
nor U40157 (N_40157,N_39399,N_36432);
nand U40158 (N_40158,N_37631,N_37709);
nand U40159 (N_40159,N_37073,N_38682);
and U40160 (N_40160,N_36358,N_35770);
and U40161 (N_40161,N_36171,N_39627);
or U40162 (N_40162,N_37183,N_38029);
or U40163 (N_40163,N_36226,N_39224);
and U40164 (N_40164,N_39326,N_38181);
nand U40165 (N_40165,N_38099,N_35491);
and U40166 (N_40166,N_38671,N_38853);
or U40167 (N_40167,N_36234,N_39773);
nor U40168 (N_40168,N_36699,N_39052);
xnor U40169 (N_40169,N_35275,N_36043);
and U40170 (N_40170,N_39087,N_38349);
or U40171 (N_40171,N_38418,N_37078);
and U40172 (N_40172,N_39946,N_37164);
xnor U40173 (N_40173,N_39436,N_39476);
and U40174 (N_40174,N_39936,N_36378);
and U40175 (N_40175,N_36837,N_38334);
nor U40176 (N_40176,N_36858,N_36896);
and U40177 (N_40177,N_35389,N_39763);
nor U40178 (N_40178,N_38186,N_37774);
nand U40179 (N_40179,N_38398,N_38737);
nand U40180 (N_40180,N_36113,N_38866);
nand U40181 (N_40181,N_35551,N_38410);
nand U40182 (N_40182,N_35134,N_39758);
nor U40183 (N_40183,N_38259,N_39919);
or U40184 (N_40184,N_36112,N_37199);
nor U40185 (N_40185,N_35472,N_37788);
or U40186 (N_40186,N_35621,N_37336);
and U40187 (N_40187,N_36296,N_38694);
nand U40188 (N_40188,N_39511,N_36490);
xor U40189 (N_40189,N_36463,N_38786);
nand U40190 (N_40190,N_39809,N_39413);
nand U40191 (N_40191,N_39770,N_39023);
nand U40192 (N_40192,N_36729,N_35522);
xnor U40193 (N_40193,N_36302,N_39924);
and U40194 (N_40194,N_35948,N_39097);
nand U40195 (N_40195,N_36444,N_38904);
nor U40196 (N_40196,N_38275,N_35231);
xnor U40197 (N_40197,N_38032,N_37300);
and U40198 (N_40198,N_38747,N_36439);
nand U40199 (N_40199,N_36505,N_38705);
and U40200 (N_40200,N_39059,N_39044);
or U40201 (N_40201,N_38909,N_39222);
and U40202 (N_40202,N_38052,N_39426);
or U40203 (N_40203,N_38288,N_36227);
and U40204 (N_40204,N_37768,N_38480);
or U40205 (N_40205,N_37171,N_36394);
and U40206 (N_40206,N_35663,N_36670);
nand U40207 (N_40207,N_38660,N_36158);
nand U40208 (N_40208,N_35489,N_39049);
or U40209 (N_40209,N_35243,N_35919);
or U40210 (N_40210,N_37405,N_35154);
and U40211 (N_40211,N_35286,N_36268);
xor U40212 (N_40212,N_38486,N_38121);
and U40213 (N_40213,N_38443,N_36293);
nor U40214 (N_40214,N_37770,N_37903);
nand U40215 (N_40215,N_36816,N_37234);
and U40216 (N_40216,N_35865,N_39746);
nand U40217 (N_40217,N_38583,N_37627);
nand U40218 (N_40218,N_35958,N_37721);
and U40219 (N_40219,N_35912,N_35531);
nor U40220 (N_40220,N_39949,N_36387);
nand U40221 (N_40221,N_37189,N_37604);
or U40222 (N_40222,N_39796,N_39263);
xor U40223 (N_40223,N_36196,N_37145);
and U40224 (N_40224,N_37119,N_35273);
and U40225 (N_40225,N_39385,N_38006);
or U40226 (N_40226,N_35097,N_35401);
and U40227 (N_40227,N_39527,N_36287);
nor U40228 (N_40228,N_39050,N_36917);
nor U40229 (N_40229,N_35719,N_39095);
nor U40230 (N_40230,N_39256,N_36718);
nand U40231 (N_40231,N_36177,N_36562);
or U40232 (N_40232,N_39459,N_38255);
xnor U40233 (N_40233,N_38523,N_35708);
nand U40234 (N_40234,N_37826,N_38744);
nor U40235 (N_40235,N_38044,N_35034);
and U40236 (N_40236,N_39189,N_37718);
and U40237 (N_40237,N_36485,N_37421);
nor U40238 (N_40238,N_35456,N_39560);
nor U40239 (N_40239,N_35547,N_35316);
nand U40240 (N_40240,N_36031,N_38828);
xor U40241 (N_40241,N_37539,N_38177);
or U40242 (N_40242,N_39568,N_35730);
nand U40243 (N_40243,N_37652,N_38436);
and U40244 (N_40244,N_39009,N_37834);
and U40245 (N_40245,N_37188,N_38638);
nor U40246 (N_40246,N_35932,N_35440);
and U40247 (N_40247,N_36713,N_38724);
xnor U40248 (N_40248,N_38802,N_39659);
nand U40249 (N_40249,N_38194,N_38193);
nor U40250 (N_40250,N_39458,N_36789);
nor U40251 (N_40251,N_37040,N_37244);
or U40252 (N_40252,N_38308,N_38388);
nand U40253 (N_40253,N_36345,N_39103);
nand U40254 (N_40254,N_39930,N_35872);
or U40255 (N_40255,N_39469,N_35956);
nor U40256 (N_40256,N_39681,N_35007);
or U40257 (N_40257,N_39393,N_38946);
nand U40258 (N_40258,N_37907,N_35077);
nand U40259 (N_40259,N_38515,N_38336);
and U40260 (N_40260,N_35048,N_35419);
nor U40261 (N_40261,N_39641,N_39795);
nor U40262 (N_40262,N_35351,N_38372);
nor U40263 (N_40263,N_36689,N_38770);
nor U40264 (N_40264,N_36450,N_39265);
or U40265 (N_40265,N_37007,N_39160);
and U40266 (N_40266,N_39859,N_36742);
or U40267 (N_40267,N_38556,N_35585);
nand U40268 (N_40268,N_39027,N_37856);
or U40269 (N_40269,N_35568,N_35962);
or U40270 (N_40270,N_35937,N_38568);
and U40271 (N_40271,N_35542,N_35695);
and U40272 (N_40272,N_36851,N_35783);
nand U40273 (N_40273,N_37485,N_38835);
and U40274 (N_40274,N_38395,N_39807);
xnor U40275 (N_40275,N_37333,N_35073);
nand U40276 (N_40276,N_37589,N_35210);
nor U40277 (N_40277,N_37549,N_37793);
and U40278 (N_40278,N_36022,N_36190);
or U40279 (N_40279,N_39646,N_37459);
nor U40280 (N_40280,N_37177,N_37972);
and U40281 (N_40281,N_39933,N_35029);
nor U40282 (N_40282,N_39489,N_36238);
nor U40283 (N_40283,N_36532,N_39618);
and U40284 (N_40284,N_36431,N_36591);
or U40285 (N_40285,N_38662,N_36514);
and U40286 (N_40286,N_35887,N_36447);
nor U40287 (N_40287,N_39916,N_38360);
xor U40288 (N_40288,N_38111,N_39319);
or U40289 (N_40289,N_36026,N_38041);
nor U40290 (N_40290,N_35646,N_36557);
nor U40291 (N_40291,N_39496,N_39002);
nand U40292 (N_40292,N_36411,N_37484);
nand U40293 (N_40293,N_36107,N_36782);
nor U40294 (N_40294,N_39204,N_35685);
nor U40295 (N_40295,N_36835,N_38416);
xor U40296 (N_40296,N_35746,N_36817);
nand U40297 (N_40297,N_36985,N_38818);
or U40298 (N_40298,N_38068,N_36109);
nor U40299 (N_40299,N_36243,N_35010);
nand U40300 (N_40300,N_37120,N_37845);
nor U40301 (N_40301,N_35717,N_35881);
nor U40302 (N_40302,N_38728,N_35690);
nor U40303 (N_40303,N_37537,N_38254);
nand U40304 (N_40304,N_39806,N_36312);
or U40305 (N_40305,N_35457,N_35654);
or U40306 (N_40306,N_35715,N_35063);
nand U40307 (N_40307,N_35628,N_35019);
and U40308 (N_40308,N_36796,N_36198);
or U40309 (N_40309,N_38734,N_38518);
and U40310 (N_40310,N_36279,N_39462);
or U40311 (N_40311,N_39512,N_35823);
or U40312 (N_40312,N_39934,N_38516);
nand U40313 (N_40313,N_35671,N_36034);
nand U40314 (N_40314,N_36928,N_37051);
nand U40315 (N_40315,N_38830,N_37474);
or U40316 (N_40316,N_37667,N_35689);
nand U40317 (N_40317,N_38054,N_37010);
nand U40318 (N_40318,N_35078,N_39072);
nor U40319 (N_40319,N_38884,N_39988);
nand U40320 (N_40320,N_39048,N_37071);
and U40321 (N_40321,N_38187,N_38408);
nand U40322 (N_40322,N_37391,N_38176);
xor U40323 (N_40323,N_39275,N_35718);
and U40324 (N_40324,N_39182,N_35040);
nor U40325 (N_40325,N_39232,N_38806);
and U40326 (N_40326,N_39159,N_37919);
and U40327 (N_40327,N_37436,N_36346);
and U40328 (N_40328,N_35699,N_37566);
nand U40329 (N_40329,N_35873,N_35899);
nor U40330 (N_40330,N_35622,N_36397);
nand U40331 (N_40331,N_37516,N_36828);
or U40332 (N_40332,N_39952,N_35536);
or U40333 (N_40333,N_36307,N_38419);
or U40334 (N_40334,N_38613,N_39270);
nand U40335 (N_40335,N_38138,N_36160);
nand U40336 (N_40336,N_39840,N_37775);
xnor U40337 (N_40337,N_36960,N_39607);
nor U40338 (N_40338,N_37806,N_38461);
and U40339 (N_40339,N_35697,N_38468);
nor U40340 (N_40340,N_38021,N_38458);
and U40341 (N_40341,N_38536,N_38180);
nand U40342 (N_40342,N_35939,N_36887);
or U40343 (N_40343,N_37184,N_38983);
xnor U40344 (N_40344,N_37355,N_36461);
and U40345 (N_40345,N_35687,N_36771);
nor U40346 (N_40346,N_36458,N_36213);
nor U40347 (N_40347,N_36506,N_39609);
and U40348 (N_40348,N_36130,N_39284);
or U40349 (N_40349,N_39693,N_37112);
nand U40350 (N_40350,N_39020,N_37050);
or U40351 (N_40351,N_37061,N_37324);
nand U40352 (N_40352,N_39749,N_36649);
nor U40353 (N_40353,N_35452,N_35371);
and U40354 (N_40354,N_35345,N_36630);
nand U40355 (N_40355,N_35090,N_36087);
nor U40356 (N_40356,N_36168,N_36179);
nand U40357 (N_40357,N_35777,N_38766);
nand U40358 (N_40358,N_36820,N_38738);
nand U40359 (N_40359,N_39948,N_37918);
nand U40360 (N_40360,N_35348,N_38757);
nor U40361 (N_40361,N_36061,N_35601);
and U40362 (N_40362,N_35195,N_38894);
or U40363 (N_40363,N_37846,N_37708);
nand U40364 (N_40364,N_37085,N_37012);
nand U40365 (N_40365,N_38311,N_36755);
nor U40366 (N_40366,N_39595,N_36683);
or U40367 (N_40367,N_36446,N_36013);
nor U40368 (N_40368,N_36628,N_39925);
or U40369 (N_40369,N_36053,N_36062);
nor U40370 (N_40370,N_37990,N_35184);
nor U40371 (N_40371,N_35808,N_36954);
and U40372 (N_40372,N_35590,N_35576);
or U40373 (N_40373,N_35619,N_36250);
xnor U40374 (N_40374,N_39254,N_36042);
nand U40375 (N_40375,N_39813,N_39248);
nor U40376 (N_40376,N_39332,N_37837);
or U40377 (N_40377,N_35447,N_37847);
nor U40378 (N_40378,N_38577,N_39983);
xor U40379 (N_40379,N_35918,N_36472);
nor U40380 (N_40380,N_36739,N_39530);
and U40381 (N_40381,N_35884,N_37981);
and U40382 (N_40382,N_35750,N_38522);
nand U40383 (N_40383,N_35121,N_36629);
or U40384 (N_40384,N_35431,N_35165);
and U40385 (N_40385,N_38834,N_38790);
nor U40386 (N_40386,N_38714,N_39093);
nor U40387 (N_40387,N_36111,N_35636);
and U40388 (N_40388,N_36512,N_35878);
and U40389 (N_40389,N_39785,N_37857);
nor U40390 (N_40390,N_37418,N_39033);
and U40391 (N_40391,N_35665,N_39778);
or U40392 (N_40392,N_37951,N_38531);
or U40393 (N_40393,N_36059,N_36300);
xor U40394 (N_40394,N_36323,N_36242);
nand U40395 (N_40395,N_39771,N_38217);
nor U40396 (N_40396,N_37028,N_37613);
nand U40397 (N_40397,N_37471,N_39541);
nand U40398 (N_40398,N_35728,N_35496);
nor U40399 (N_40399,N_35144,N_37035);
nand U40400 (N_40400,N_35995,N_35786);
nor U40401 (N_40401,N_35486,N_39757);
or U40402 (N_40402,N_36714,N_38424);
or U40403 (N_40403,N_37704,N_38491);
and U40404 (N_40404,N_37994,N_36748);
nand U40405 (N_40405,N_38513,N_37633);
nor U40406 (N_40406,N_36152,N_37536);
nand U40407 (N_40407,N_35260,N_37580);
and U40408 (N_40408,N_37947,N_36487);
or U40409 (N_40409,N_39228,N_35942);
nand U40410 (N_40410,N_39185,N_37223);
and U40411 (N_40411,N_38269,N_36981);
nor U40412 (N_40412,N_38721,N_35483);
xnor U40413 (N_40413,N_35434,N_35330);
and U40414 (N_40414,N_36143,N_38357);
or U40415 (N_40415,N_36994,N_35269);
or U40416 (N_40416,N_35527,N_38609);
and U40417 (N_40417,N_36658,N_35834);
nor U40418 (N_40418,N_37390,N_36003);
nand U40419 (N_40419,N_36124,N_38890);
nor U40420 (N_40420,N_35960,N_38677);
nand U40421 (N_40421,N_36855,N_39928);
and U40422 (N_40422,N_37394,N_38067);
or U40423 (N_40423,N_38078,N_39045);
xnor U40424 (N_40424,N_35006,N_35500);
and U40425 (N_40425,N_38455,N_35779);
nand U40426 (N_40426,N_37809,N_37386);
nand U40427 (N_40427,N_39398,N_39582);
or U40428 (N_40428,N_35811,N_35732);
nand U40429 (N_40429,N_38122,N_36806);
xor U40430 (N_40430,N_35766,N_35058);
or U40431 (N_40431,N_37187,N_36894);
or U40432 (N_40432,N_36586,N_38179);
nand U40433 (N_40433,N_37158,N_37447);
or U40434 (N_40434,N_38597,N_39938);
and U40435 (N_40435,N_35679,N_37374);
xor U40436 (N_40436,N_36661,N_35475);
nor U40437 (N_40437,N_38081,N_39623);
and U40438 (N_40438,N_39479,N_36045);
nand U40439 (N_40439,N_39835,N_37313);
nor U40440 (N_40440,N_37132,N_35603);
or U40441 (N_40441,N_38743,N_37554);
and U40442 (N_40442,N_37298,N_35296);
and U40443 (N_40443,N_35694,N_37945);
nand U40444 (N_40444,N_38773,N_39881);
nor U40445 (N_40445,N_36409,N_39480);
or U40446 (N_40446,N_35041,N_35629);
nor U40447 (N_40447,N_35420,N_37958);
and U40448 (N_40448,N_37329,N_39098);
nor U40449 (N_40449,N_35798,N_35492);
and U40450 (N_40450,N_35407,N_37480);
or U40451 (N_40451,N_38628,N_39244);
and U40452 (N_40452,N_35614,N_39839);
or U40453 (N_40453,N_37200,N_37760);
and U40454 (N_40454,N_39294,N_38846);
nand U40455 (N_40455,N_38857,N_36078);
or U40456 (N_40456,N_35305,N_38341);
nor U40457 (N_40457,N_37377,N_38881);
and U40458 (N_40458,N_36496,N_38075);
nand U40459 (N_40459,N_39931,N_39207);
or U40460 (N_40460,N_35290,N_36639);
and U40461 (N_40461,N_38257,N_38156);
and U40462 (N_40462,N_39581,N_38670);
and U40463 (N_40463,N_37062,N_35516);
xnor U40464 (N_40464,N_38990,N_36740);
nand U40465 (N_40465,N_36737,N_39664);
xnor U40466 (N_40466,N_35810,N_36838);
nor U40467 (N_40467,N_39154,N_39978);
or U40468 (N_40468,N_36856,N_37282);
and U40469 (N_40469,N_37555,N_37038);
xor U40470 (N_40470,N_38563,N_37872);
nor U40471 (N_40471,N_37109,N_35340);
or U40472 (N_40472,N_37398,N_36906);
nor U40473 (N_40473,N_39801,N_36593);
nor U40474 (N_40474,N_39943,N_39761);
nand U40475 (N_40475,N_37603,N_35176);
nor U40476 (N_40476,N_35157,N_37949);
nor U40477 (N_40477,N_39505,N_36615);
nand U40478 (N_40478,N_37136,N_38886);
and U40479 (N_40479,N_37861,N_39826);
or U40480 (N_40480,N_39137,N_36473);
and U40481 (N_40481,N_39502,N_35448);
nor U40482 (N_40482,N_39293,N_36029);
nand U40483 (N_40483,N_38637,N_35030);
or U40484 (N_40484,N_38742,N_37649);
nand U40485 (N_40485,N_35026,N_38559);
nor U40486 (N_40486,N_39483,N_37696);
and U40487 (N_40487,N_39877,N_36947);
xor U40488 (N_40488,N_36276,N_37494);
nand U40489 (N_40489,N_35495,N_36823);
nand U40490 (N_40490,N_35169,N_36958);
or U40491 (N_40491,N_39316,N_39836);
and U40492 (N_40492,N_39860,N_38279);
nand U40493 (N_40493,N_39374,N_37294);
nor U40494 (N_40494,N_35039,N_38298);
or U40495 (N_40495,N_38244,N_36653);
nor U40496 (N_40496,N_36877,N_35898);
nor U40497 (N_40497,N_36437,N_38202);
and U40498 (N_40498,N_38891,N_39668);
or U40499 (N_40499,N_37605,N_39285);
nor U40500 (N_40500,N_39351,N_35354);
and U40501 (N_40501,N_38236,N_38604);
and U40502 (N_40502,N_39309,N_36317);
nand U40503 (N_40503,N_36021,N_35792);
xnor U40504 (N_40504,N_39756,N_37185);
or U40505 (N_40505,N_36944,N_39868);
and U40506 (N_40506,N_39911,N_38520);
or U40507 (N_40507,N_36373,N_36971);
xnor U40508 (N_40508,N_35916,N_36481);
nor U40509 (N_40509,N_38463,N_35989);
nand U40510 (N_40510,N_36395,N_38264);
and U40511 (N_40511,N_39241,N_35990);
and U40512 (N_40512,N_35913,N_38028);
and U40513 (N_40513,N_37508,N_39051);
nor U40514 (N_40514,N_38726,N_38166);
nand U40515 (N_40515,N_39471,N_39754);
and U40516 (N_40516,N_38702,N_38013);
or U40517 (N_40517,N_38689,N_37732);
nor U40518 (N_40518,N_36647,N_37433);
and U40519 (N_40519,N_38009,N_36784);
and U40520 (N_40520,N_36340,N_39674);
xor U40521 (N_40521,N_39906,N_37481);
or U40522 (N_40522,N_35643,N_39148);
xor U40523 (N_40523,N_35714,N_39202);
nand U40524 (N_40524,N_36704,N_36263);
nor U40525 (N_40525,N_35763,N_38221);
or U40526 (N_40526,N_38844,N_39180);
nand U40527 (N_40527,N_37672,N_39976);
xnor U40528 (N_40528,N_35634,N_39015);
or U40529 (N_40529,N_38046,N_36741);
nand U40530 (N_40530,N_36028,N_38203);
or U40531 (N_40531,N_36533,N_38150);
xnor U40532 (N_40532,N_35901,N_35565);
nand U40533 (N_40533,N_39660,N_35692);
nand U40534 (N_40534,N_35828,N_39714);
xnor U40535 (N_40535,N_36840,N_36854);
and U40536 (N_40536,N_36023,N_38145);
nor U40537 (N_40537,N_39114,N_35882);
and U40538 (N_40538,N_39369,N_39448);
or U40539 (N_40539,N_38370,N_35721);
nor U40540 (N_40540,N_35682,N_37843);
nand U40541 (N_40541,N_35367,N_38319);
and U40542 (N_40542,N_37404,N_35856);
nor U40543 (N_40543,N_39308,N_38389);
nand U40544 (N_40544,N_39318,N_35592);
xnor U40545 (N_40545,N_37916,N_38807);
xnor U40546 (N_40546,N_35065,N_39696);
nand U40547 (N_40547,N_37824,N_37399);
and U40548 (N_40548,N_39022,N_35436);
or U40549 (N_40549,N_39080,N_35344);
nor U40550 (N_40550,N_37288,N_38998);
and U40551 (N_40551,N_37651,N_35888);
and U40552 (N_40552,N_38557,N_37064);
or U40553 (N_40553,N_36495,N_36539);
nor U40554 (N_40554,N_37626,N_35894);
nor U40555 (N_40555,N_37882,N_37915);
xnor U40556 (N_40556,N_35148,N_36459);
nand U40557 (N_40557,N_35111,N_36984);
and U40558 (N_40558,N_38752,N_35709);
nor U40559 (N_40559,N_38605,N_36092);
and U40560 (N_40560,N_35379,N_37648);
xnor U40561 (N_40561,N_38631,N_39593);
nand U40562 (N_40562,N_36553,N_39628);
nor U40563 (N_40563,N_35661,N_35464);
or U40564 (N_40564,N_38865,N_37607);
nor U40565 (N_40565,N_37069,N_35541);
nor U40566 (N_40566,N_38083,N_39173);
and U40567 (N_40567,N_39260,N_36938);
or U40568 (N_40568,N_36477,N_39854);
nand U40569 (N_40569,N_39129,N_39852);
nand U40570 (N_40570,N_37906,N_35042);
nand U40571 (N_40571,N_35548,N_36036);
or U40572 (N_40572,N_39314,N_38362);
or U40573 (N_40573,N_35772,N_37299);
nand U40574 (N_40574,N_35247,N_39955);
or U40575 (N_40575,N_38126,N_36930);
nor U40576 (N_40576,N_35926,N_39895);
or U40577 (N_40577,N_35691,N_39133);
nor U40578 (N_40578,N_35889,N_35526);
nor U40579 (N_40579,N_38528,N_35775);
nand U40580 (N_40580,N_36150,N_36685);
nand U40581 (N_40581,N_37895,N_38146);
or U40582 (N_40582,N_35571,N_36725);
nand U40583 (N_40583,N_39727,N_38049);
nor U40584 (N_40584,N_39531,N_38142);
or U40585 (N_40585,N_39838,N_36385);
xnor U40586 (N_40586,N_37720,N_37877);
nor U40587 (N_40587,N_35156,N_39481);
xor U40588 (N_40588,N_39554,N_38252);
xor U40589 (N_40589,N_35241,N_36155);
nor U40590 (N_40590,N_38188,N_39981);
nand U40591 (N_40591,N_35789,N_37034);
xnor U40592 (N_40592,N_36237,N_39450);
nor U40593 (N_40593,N_38979,N_36519);
or U40594 (N_40594,N_38190,N_39384);
and U40595 (N_40595,N_37961,N_37922);
or U40596 (N_40596,N_37440,N_39350);
nand U40597 (N_40597,N_37046,N_39893);
nand U40598 (N_40598,N_38771,N_38383);
and U40599 (N_40599,N_38928,N_36265);
nor U40600 (N_40600,N_37570,N_39675);
or U40601 (N_40601,N_37468,N_35386);
and U40602 (N_40602,N_38938,N_37754);
nand U40603 (N_40603,N_37638,N_39191);
or U40604 (N_40604,N_39794,N_37364);
xnor U40605 (N_40605,N_36436,N_39297);
nand U40606 (N_40606,N_39225,N_36055);
and U40607 (N_40607,N_39252,N_38120);
nand U40608 (N_40608,N_37940,N_38566);
and U40609 (N_40609,N_39329,N_38701);
nand U40610 (N_40610,N_39152,N_38160);
nor U40611 (N_40611,N_38096,N_39742);
and U40612 (N_40612,N_37206,N_38722);
xor U40613 (N_40613,N_37462,N_38995);
and U40614 (N_40614,N_36859,N_38353);
or U40615 (N_40615,N_35736,N_39069);
nand U40616 (N_40616,N_39372,N_38841);
and U40617 (N_40617,N_36831,N_36405);
or U40618 (N_40618,N_36063,N_35723);
nor U40619 (N_40619,N_39029,N_36066);
and U40620 (N_40620,N_36270,N_35549);
xor U40621 (N_40621,N_35218,N_35444);
nand U40622 (N_40622,N_36507,N_39171);
nor U40623 (N_40623,N_36698,N_39543);
and U40624 (N_40624,N_35712,N_36788);
nand U40625 (N_40625,N_37782,N_35649);
and U40626 (N_40626,N_36778,N_37509);
and U40627 (N_40627,N_37661,N_36845);
xnor U40628 (N_40628,N_36486,N_39649);
nand U40629 (N_40629,N_35883,N_35767);
nor U40630 (N_40630,N_39219,N_39891);
xor U40631 (N_40631,N_38492,N_35455);
or U40632 (N_40632,N_37928,N_38839);
xor U40633 (N_40633,N_39181,N_37680);
and U40634 (N_40634,N_38809,N_37041);
and U40635 (N_40635,N_37252,N_39608);
nand U40636 (N_40636,N_37488,N_39589);
nor U40637 (N_40637,N_36955,N_38680);
or U40638 (N_40638,N_37347,N_36371);
nor U40639 (N_40639,N_35979,N_38501);
nor U40640 (N_40640,N_37455,N_38407);
and U40641 (N_40641,N_36973,N_39677);
or U40642 (N_40642,N_36451,N_37261);
and U40643 (N_40643,N_37673,N_39017);
nand U40644 (N_40644,N_37068,N_38088);
nand U40645 (N_40645,N_38474,N_38810);
nor U40646 (N_40646,N_37000,N_37889);
or U40647 (N_40647,N_35337,N_36319);
xnor U40648 (N_40648,N_39603,N_35617);
nand U40649 (N_40649,N_39897,N_37569);
nand U40650 (N_40650,N_39972,N_35627);
nor U40651 (N_40651,N_35611,N_36556);
nor U40652 (N_40652,N_37683,N_35416);
or U40653 (N_40653,N_37344,N_38579);
nor U40654 (N_40654,N_36797,N_37350);
nand U40655 (N_40655,N_38027,N_35155);
or U40656 (N_40656,N_39873,N_38483);
nor U40657 (N_40657,N_39333,N_38606);
and U40658 (N_40658,N_36880,N_37515);
or U40659 (N_40659,N_35825,N_37968);
nor U40660 (N_40660,N_35101,N_35320);
or U40661 (N_40661,N_35091,N_35118);
and U40662 (N_40662,N_36618,N_39869);
nor U40663 (N_40663,N_37305,N_37609);
and U40664 (N_40664,N_37955,N_38452);
nand U40665 (N_40665,N_36580,N_39900);
or U40666 (N_40666,N_37987,N_36251);
nor U40667 (N_40667,N_38033,N_39940);
nor U40668 (N_40668,N_35835,N_36619);
and U40669 (N_40669,N_36608,N_36776);
or U40670 (N_40670,N_37491,N_36239);
nor U40671 (N_40671,N_36138,N_35869);
nand U40672 (N_40672,N_37726,N_37884);
and U40673 (N_40673,N_35350,N_37182);
and U40674 (N_40674,N_39493,N_37151);
nor U40675 (N_40675,N_37599,N_38933);
and U40676 (N_40676,N_35623,N_39238);
and U40677 (N_40677,N_35647,N_38673);
nor U40678 (N_40678,N_36216,N_36343);
and U40679 (N_40679,N_38053,N_38199);
and U40680 (N_40680,N_39909,N_39518);
or U40681 (N_40681,N_39340,N_39962);
nor U40682 (N_40682,N_39950,N_39600);
and U40683 (N_40683,N_38898,N_38706);
nand U40684 (N_40684,N_39509,N_36662);
nand U40685 (N_40685,N_39035,N_37339);
nand U40686 (N_40686,N_35754,N_38948);
nor U40687 (N_40687,N_37747,N_39269);
nand U40688 (N_40688,N_38213,N_39447);
nand U40689 (N_40689,N_37475,N_35146);
nor U40690 (N_40690,N_35529,N_36717);
and U40691 (N_40691,N_36009,N_39574);
nand U40692 (N_40692,N_35280,N_35822);
nand U40693 (N_40693,N_39184,N_36732);
and U40694 (N_40694,N_36240,N_35322);
nor U40695 (N_40695,N_37785,N_39845);
or U40696 (N_40696,N_37851,N_39408);
nor U40697 (N_40697,N_35264,N_37135);
and U40698 (N_40698,N_38535,N_39960);
and U40699 (N_40699,N_38079,N_38413);
and U40700 (N_40700,N_37976,N_37671);
or U40701 (N_40701,N_37559,N_38476);
or U40702 (N_40702,N_38935,N_36513);
nand U40703 (N_40703,N_37143,N_39289);
or U40704 (N_40704,N_38824,N_39657);
nor U40705 (N_40705,N_38625,N_38498);
nand U40706 (N_40706,N_37635,N_38849);
nand U40707 (N_40707,N_35086,N_35996);
and U40708 (N_40708,N_38402,N_39392);
or U40709 (N_40709,N_36939,N_36136);
xnor U40710 (N_40710,N_37490,N_36211);
or U40711 (N_40711,N_36997,N_36176);
nor U40712 (N_40712,N_38860,N_36368);
nand U40713 (N_40713,N_38709,N_37912);
and U40714 (N_40714,N_36675,N_38404);
xnor U40715 (N_40715,N_37357,N_37281);
or U40716 (N_40716,N_35982,N_36032);
nand U40717 (N_40717,N_35587,N_37866);
and U40718 (N_40718,N_35387,N_38913);
nor U40719 (N_40719,N_38635,N_35469);
nand U40720 (N_40720,N_38784,N_38861);
nor U40721 (N_40721,N_39233,N_38366);
or U40722 (N_40722,N_39213,N_35844);
or U40723 (N_40723,N_39357,N_37056);
and U40724 (N_40724,N_36898,N_35487);
nand U40725 (N_40725,N_35235,N_37796);
nand U40726 (N_40726,N_37013,N_35022);
and U40727 (N_40727,N_35084,N_38945);
nor U40728 (N_40728,N_39557,N_38712);
nor U40729 (N_40729,N_39491,N_39170);
and U40730 (N_40730,N_35009,N_38090);
nand U40731 (N_40731,N_35914,N_35740);
xnor U40732 (N_40732,N_39435,N_38124);
nand U40733 (N_40733,N_39075,N_37533);
nor U40734 (N_40734,N_38101,N_39421);
and U40735 (N_40735,N_37959,N_37110);
or U40736 (N_40736,N_35702,N_35398);
nand U40737 (N_40737,N_37469,N_39100);
or U40738 (N_40738,N_37096,N_37059);
or U40739 (N_40739,N_39115,N_38183);
nand U40740 (N_40740,N_38970,N_35412);
xnor U40741 (N_40741,N_35075,N_37550);
nand U40742 (N_40742,N_38430,N_36941);
or U40743 (N_40743,N_38554,N_37783);
nor U40744 (N_40744,N_39798,N_38328);
and U40745 (N_40745,N_39279,N_36151);
nand U40746 (N_40746,N_38663,N_39703);
nor U40747 (N_40747,N_39719,N_38533);
and U40748 (N_40748,N_35251,N_39074);
nor U40749 (N_40749,N_37413,N_39440);
or U40750 (N_40750,N_35589,N_39253);
or U40751 (N_40751,N_35974,N_36805);
and U40752 (N_40752,N_39396,N_36201);
nor U40753 (N_40753,N_36406,N_39032);
nor U40754 (N_40754,N_37385,N_36728);
nand U40755 (N_40755,N_39391,N_38787);
or U40756 (N_40756,N_37558,N_36535);
nand U40757 (N_40757,N_37737,N_36086);
or U40758 (N_40758,N_39145,N_39847);
nand U40759 (N_40759,N_35624,N_39910);
and U40760 (N_40760,N_36581,N_39151);
and U40761 (N_40761,N_37717,N_35521);
or U40762 (N_40762,N_37254,N_38442);
xnor U40763 (N_40763,N_37746,N_39532);
and U40764 (N_40764,N_39036,N_35246);
or U40765 (N_40765,N_39439,N_38265);
and U40766 (N_40766,N_39915,N_38612);
and U40767 (N_40767,N_37727,N_38035);
nand U40768 (N_40768,N_36824,N_39846);
and U40769 (N_40769,N_36688,N_35225);
nor U40770 (N_40770,N_36030,N_36563);
nor U40771 (N_40771,N_36585,N_37320);
and U40772 (N_40772,N_37037,N_36510);
or U40773 (N_40773,N_35860,N_38794);
or U40774 (N_40774,N_37776,N_35802);
nand U40775 (N_40775,N_37973,N_36094);
or U40776 (N_40776,N_36518,N_39963);
xnor U40777 (N_40777,N_37380,N_39510);
nor U40778 (N_40778,N_37896,N_38621);
or U40779 (N_40779,N_36365,N_39808);
and U40780 (N_40780,N_37054,N_37157);
and U40781 (N_40781,N_39484,N_36832);
or U40782 (N_40782,N_37573,N_36515);
or U40783 (N_40783,N_38918,N_36566);
or U40784 (N_40784,N_35339,N_38996);
or U40785 (N_40785,N_37507,N_37030);
nand U40786 (N_40786,N_36957,N_36555);
nand U40787 (N_40787,N_35674,N_38655);
nand U40788 (N_40788,N_37194,N_38434);
nor U40789 (N_40789,N_35907,N_35570);
nand U40790 (N_40790,N_36230,N_35816);
nand U40791 (N_40791,N_38004,N_36974);
nor U40792 (N_40792,N_37343,N_37913);
nor U40793 (N_40793,N_36564,N_37950);
xor U40794 (N_40794,N_38415,N_35093);
or U40795 (N_40795,N_38297,N_37106);
and U40796 (N_40796,N_35274,N_39633);
and U40797 (N_40797,N_39237,N_35207);
and U40798 (N_40798,N_36720,N_35814);
and U40799 (N_40799,N_35089,N_39596);
nor U40800 (N_40800,N_36258,N_38547);
nor U40801 (N_40801,N_39084,N_39474);
and U40802 (N_40802,N_36715,N_35250);
xor U40803 (N_40803,N_39054,N_36174);
or U40804 (N_40804,N_35900,N_38924);
nor U40805 (N_40805,N_38292,N_35462);
and U40806 (N_40806,N_39134,N_39652);
or U40807 (N_40807,N_39167,N_39550);
nor U40808 (N_40808,N_35375,N_36790);
nor U40809 (N_40809,N_39800,N_35890);
nor U40810 (N_40810,N_37302,N_35920);
or U40811 (N_40811,N_38708,N_35027);
and U40812 (N_40812,N_38085,N_38781);
nor U40813 (N_40813,N_38651,N_37590);
or U40814 (N_40814,N_38304,N_39896);
or U40815 (N_40815,N_35216,N_37690);
and U40816 (N_40816,N_36453,N_37277);
or U40817 (N_40817,N_38674,N_38154);
and U40818 (N_40818,N_39739,N_37065);
nor U40819 (N_40819,N_36117,N_39572);
nor U40820 (N_40820,N_35466,N_36399);
or U40821 (N_40821,N_38832,N_35227);
xnor U40822 (N_40822,N_37108,N_35711);
or U40823 (N_40823,N_39176,N_36599);
nand U40824 (N_40824,N_35102,N_35613);
xnor U40825 (N_40825,N_36587,N_38230);
or U40826 (N_40826,N_37620,N_37166);
nand U40827 (N_40827,N_37331,N_35896);
and U40828 (N_40828,N_35353,N_39546);
or U40829 (N_40829,N_38163,N_39941);
and U40830 (N_40830,N_37196,N_35604);
nor U40831 (N_40831,N_38622,N_36137);
and U40832 (N_40832,N_36246,N_38109);
or U40833 (N_40833,N_37619,N_39544);
or U40834 (N_40834,N_36148,N_36700);
nor U40835 (N_40835,N_37771,N_37087);
nor U40836 (N_40836,N_39113,N_36541);
xor U40837 (N_40837,N_37142,N_35945);
or U40838 (N_40838,N_36104,N_37162);
or U40839 (N_40839,N_39953,N_38741);
and U40840 (N_40840,N_35530,N_38503);
and U40841 (N_40841,N_37926,N_35435);
nand U40842 (N_40842,N_39131,N_39206);
xor U40843 (N_40843,N_39201,N_37777);
or U40844 (N_40844,N_38457,N_36803);
or U40845 (N_40845,N_38586,N_37297);
and U40846 (N_40846,N_38337,N_35722);
nor U40847 (N_40847,N_38984,N_37974);
and U40848 (N_40848,N_39655,N_37964);
and U40849 (N_40849,N_35673,N_35382);
nor U40850 (N_40850,N_35088,N_39682);
and U40851 (N_40851,N_35965,N_37246);
nor U40852 (N_40852,N_38363,N_38344);
and U40853 (N_40853,N_39508,N_37406);
nand U40854 (N_40854,N_38381,N_39556);
nand U40855 (N_40855,N_37773,N_35033);
nor U40856 (N_40856,N_36048,N_39516);
xor U40857 (N_40857,N_35023,N_35513);
or U40858 (N_40858,N_35204,N_35037);
xnor U40859 (N_40859,N_35532,N_35174);
or U40860 (N_40860,N_36056,N_38544);
and U40861 (N_40861,N_37253,N_37992);
xnor U40862 (N_40862,N_36015,N_37072);
and U40863 (N_40863,N_38560,N_38943);
and U40864 (N_40864,N_39487,N_35705);
or U40865 (N_40865,N_37323,N_39908);
nor U40866 (N_40866,N_35332,N_38218);
and U40867 (N_40867,N_36710,N_38490);
and U40868 (N_40868,N_39443,N_35265);
and U40869 (N_40869,N_39349,N_38369);
nor U40870 (N_40870,N_35535,N_35610);
or U40871 (N_40871,N_35707,N_37551);
nor U40872 (N_40872,N_36849,N_37552);
nor U40873 (N_40873,N_36864,N_35197);
or U40874 (N_40874,N_38189,N_36951);
and U40875 (N_40875,N_38934,N_38669);
nor U40876 (N_40876,N_38338,N_38007);
nor U40877 (N_40877,N_36830,N_38901);
and U40878 (N_40878,N_39982,N_36702);
nand U40879 (N_40879,N_37219,N_39884);
or U40880 (N_40880,N_35186,N_35580);
nand U40881 (N_40881,N_39814,N_37102);
and U40882 (N_40882,N_39268,N_39957);
and U40883 (N_40883,N_39583,N_38797);
nor U40884 (N_40884,N_39315,N_35769);
and U40885 (N_40885,N_38848,N_35991);
and U40886 (N_40886,N_38825,N_35404);
nor U40887 (N_40887,N_35237,N_39812);
or U40888 (N_40888,N_38594,N_38952);
nand U40889 (N_40889,N_36968,N_37844);
nand U40890 (N_40890,N_39220,N_39288);
nor U40891 (N_40891,N_38885,N_37815);
and U40892 (N_40892,N_39929,N_39467);
or U40893 (N_40893,N_37954,N_36758);
or U40894 (N_40894,N_36425,N_37988);
and U40895 (N_40895,N_39680,N_39102);
or U40896 (N_40896,N_38070,N_38852);
and U40897 (N_40897,N_38331,N_37160);
and U40898 (N_40898,N_39292,N_36041);
nor U40899 (N_40899,N_38593,N_36331);
nor U40900 (N_40900,N_38128,N_35335);
and U40901 (N_40901,N_36652,N_37174);
nand U40902 (N_40902,N_37216,N_37004);
nor U40903 (N_40903,N_36660,N_36132);
and U40904 (N_40904,N_39843,N_39885);
and U40905 (N_40905,N_39500,N_38619);
xnor U40906 (N_40906,N_36284,N_39987);
xnor U40907 (N_40907,N_37353,N_38445);
nor U40908 (N_40908,N_36223,N_35145);
nor U40909 (N_40909,N_37914,N_35333);
xor U40910 (N_40910,N_38723,N_36785);
xnor U40911 (N_40911,N_39364,N_37526);
or U40912 (N_40912,N_38999,N_39112);
nand U40913 (N_40913,N_39298,N_38211);
and U40914 (N_40914,N_38106,N_35151);
nand U40915 (N_40915,N_37039,N_35842);
nand U40916 (N_40916,N_36222,N_37137);
or U40917 (N_40917,N_37236,N_36362);
nand U40918 (N_40918,N_39555,N_37725);
and U40919 (N_40919,N_37332,N_38466);
nor U40920 (N_40920,N_36091,N_39030);
or U40921 (N_40921,N_36597,N_36388);
nand U40922 (N_40922,N_35946,N_36082);
or U40923 (N_40923,N_39547,N_38778);
xnor U40924 (N_40924,N_37931,N_37093);
and U40925 (N_40925,N_35909,N_36808);
xor U40926 (N_40926,N_37147,N_35281);
nor U40927 (N_40927,N_38358,N_35866);
or U40928 (N_40928,N_37827,N_37702);
and U40929 (N_40929,N_39648,N_35774);
and U40930 (N_40930,N_35804,N_35940);
and U40931 (N_40931,N_39971,N_36192);
and U40932 (N_40932,N_38532,N_36904);
and U40933 (N_40933,N_38469,N_36191);
and U40934 (N_40934,N_37890,N_38432);
and U40935 (N_40935,N_38073,N_37695);
nor U40936 (N_40936,N_39679,N_37986);
and U40937 (N_40937,N_38962,N_37434);
nor U40938 (N_40938,N_38958,N_35268);
xnor U40939 (N_40939,N_35626,N_39788);
nor U40940 (N_40940,N_38683,N_35113);
xor U40941 (N_40941,N_38939,N_37634);
and U40942 (N_40942,N_39460,N_39395);
nand U40943 (N_40943,N_36301,N_39523);
xor U40944 (N_40944,N_35607,N_37543);
xor U40945 (N_40945,N_38080,N_35185);
nor U40946 (N_40946,N_37862,N_36188);
or U40947 (N_40947,N_38284,N_35068);
nand U40948 (N_40948,N_39833,N_38322);
nand U40949 (N_40949,N_35349,N_35360);
nand U40950 (N_40950,N_39642,N_38439);
nor U40951 (N_40951,N_39515,N_36900);
nand U40952 (N_40952,N_35837,N_35409);
nand U40953 (N_40953,N_37659,N_38143);
nand U40954 (N_40954,N_35861,N_36719);
nor U40955 (N_40955,N_38889,N_37676);
or U40956 (N_40956,N_39494,N_37593);
nand U40957 (N_40957,N_38310,N_36099);
nand U40958 (N_40958,N_35212,N_35546);
nor U40959 (N_40959,N_39848,N_37874);
or U40960 (N_40960,N_36382,N_37522);
or U40961 (N_40961,N_37260,N_35506);
nor U40962 (N_40962,N_35713,N_37750);
and U40963 (N_40963,N_35393,N_38878);
or U40964 (N_40964,N_38247,N_35205);
xnor U40965 (N_40965,N_38050,N_39614);
nor U40966 (N_40966,N_39871,N_35929);
nor U40967 (N_40967,N_36161,N_39822);
nand U40968 (N_40968,N_36149,N_38412);
or U40969 (N_40969,N_35641,N_35343);
nand U40970 (N_40970,N_35092,N_39127);
nand U40971 (N_40971,N_36722,N_37740);
nor U40972 (N_40972,N_35978,N_39031);
nand U40973 (N_40973,N_38530,N_37003);
nand U40974 (N_40974,N_38327,N_38703);
or U40975 (N_40975,N_35519,N_38226);
nor U40976 (N_40976,N_38930,N_36210);
and U40977 (N_40977,N_36389,N_37836);
nand U40978 (N_40978,N_36297,N_35159);
nand U40979 (N_40979,N_39262,N_38076);
nor U40980 (N_40980,N_36907,N_39569);
nand U40981 (N_40981,N_37807,N_38800);
nor U40982 (N_40982,N_35875,N_36848);
xor U40983 (N_40983,N_39143,N_37169);
nor U40984 (N_40984,N_38294,N_36892);
or U40985 (N_40985,N_38152,N_36663);
or U40986 (N_40986,N_35983,N_39082);
nand U40987 (N_40987,N_38258,N_39376);
and U40988 (N_40988,N_36865,N_35988);
and U40989 (N_40989,N_38379,N_37991);
nor U40990 (N_40990,N_37257,N_35594);
or U40991 (N_40991,N_37052,N_35973);
nand U40992 (N_40992,N_37574,N_37255);
nor U40993 (N_40993,N_39046,N_39816);
and U40994 (N_40994,N_37057,N_35969);
and U40995 (N_40995,N_37818,N_36337);
nand U40996 (N_40996,N_39466,N_39083);
nand U40997 (N_40997,N_38289,N_37049);
or U40998 (N_40998,N_39615,N_35168);
and U40999 (N_40999,N_36381,N_38196);
nand U41000 (N_41000,N_36332,N_39077);
nor U41001 (N_41001,N_37891,N_35954);
and U41002 (N_41002,N_37212,N_37220);
and U41003 (N_41003,N_38681,N_37181);
xnor U41004 (N_41004,N_39287,N_36972);
and U41005 (N_41005,N_35163,N_38527);
and U41006 (N_41006,N_39139,N_39996);
nor U41007 (N_41007,N_35016,N_39879);
or U41008 (N_41008,N_38325,N_37799);
nor U41009 (N_41009,N_35279,N_35729);
and U41010 (N_41010,N_39565,N_35095);
nor U41011 (N_41011,N_35934,N_38792);
or U41012 (N_41012,N_35302,N_35538);
nor U41013 (N_41013,N_37439,N_35291);
nor U41014 (N_41014,N_35893,N_38664);
xor U41015 (N_41015,N_38201,N_37628);
and U41016 (N_41016,N_37152,N_37479);
or U41017 (N_41017,N_39517,N_36768);
xnor U41018 (N_41018,N_38271,N_38936);
nor U41019 (N_41019,N_38697,N_39060);
and U41020 (N_41020,N_38667,N_37476);
nor U41021 (N_41021,N_38858,N_37415);
or U41022 (N_41022,N_36919,N_36144);
and U41023 (N_41023,N_35399,N_36522);
and U41024 (N_41024,N_37731,N_37295);
and U41025 (N_41025,N_39498,N_37178);
and U41026 (N_41026,N_37452,N_37443);
xnor U41027 (N_41027,N_38059,N_36834);
nor U41028 (N_41028,N_35081,N_35806);
nand U41029 (N_41029,N_37267,N_39886);
nor U41030 (N_41030,N_39043,N_39956);
or U41031 (N_41031,N_36286,N_37728);
nand U41032 (N_41032,N_39061,N_35943);
nor U41033 (N_41033,N_39373,N_36369);
nor U41034 (N_41034,N_39872,N_36690);
and U41035 (N_41035,N_39864,N_37249);
nor U41036 (N_41036,N_35752,N_37111);
and U41037 (N_41037,N_39306,N_38855);
or U41038 (N_41038,N_36731,N_39830);
nor U41039 (N_41039,N_35787,N_36936);
or U41040 (N_41040,N_39506,N_39013);
nand U41041 (N_41041,N_36948,N_39912);
nand U41042 (N_41042,N_39942,N_37089);
or U41043 (N_41043,N_38863,N_39358);
or U41044 (N_41044,N_36166,N_37666);
and U41045 (N_41045,N_37917,N_39882);
and U41046 (N_41046,N_35100,N_38197);
nor U41047 (N_41047,N_37904,N_39475);
nor U41048 (N_41048,N_37553,N_39470);
xnor U41049 (N_41049,N_39094,N_35087);
nor U41050 (N_41050,N_38799,N_38698);
or U41051 (N_41051,N_39804,N_35266);
nand U41052 (N_41052,N_36814,N_35429);
and U41053 (N_41053,N_38497,N_35559);
and U41054 (N_41054,N_38060,N_38534);
nand U41055 (N_41055,N_39168,N_38329);
nand U41056 (N_41056,N_35206,N_39899);
nand U41057 (N_41057,N_38003,N_35011);
and U41058 (N_41058,N_36786,N_35045);
xor U41059 (N_41059,N_37602,N_36330);
nand U41060 (N_41060,N_39718,N_37311);
xor U41061 (N_41061,N_36402,N_35867);
nand U41062 (N_41062,N_38069,N_36430);
xnor U41063 (N_41063,N_37133,N_38801);
or U41064 (N_41064,N_36612,N_37944);
and U41065 (N_41065,N_37711,N_35562);
and U41066 (N_41066,N_39740,N_38610);
or U41067 (N_41067,N_36520,N_38856);
and U41068 (N_41068,N_39923,N_39365);
nand U41069 (N_41069,N_39637,N_36484);
nor U41070 (N_41070,N_36355,N_39575);
nor U41071 (N_41071,N_39705,N_39926);
or U41072 (N_41072,N_39867,N_37330);
and U41073 (N_41073,N_39330,N_37420);
nor U41074 (N_41074,N_35377,N_38253);
xnor U41075 (N_41075,N_39750,N_38882);
nand U41076 (N_41076,N_37138,N_36600);
and U41077 (N_41077,N_39461,N_36525);
or U41078 (N_41078,N_36528,N_38862);
nand U41079 (N_41079,N_38393,N_39602);
nand U41080 (N_41080,N_36545,N_35421);
nand U41081 (N_41081,N_38926,N_37828);
and U41082 (N_41082,N_38135,N_35366);
or U41083 (N_41083,N_37208,N_38012);
xor U41084 (N_41084,N_37753,N_38763);
nand U41085 (N_41085,N_36804,N_39643);
or U41086 (N_41086,N_39247,N_35832);
and U41087 (N_41087,N_39592,N_37451);
nand U41088 (N_41088,N_38966,N_36352);
nand U41089 (N_41089,N_39217,N_35748);
nand U41090 (N_41090,N_39922,N_38133);
or U41091 (N_41091,N_39055,N_35971);
nor U41092 (N_41092,N_36872,N_35652);
or U41093 (N_41093,N_39999,N_38627);
or U41094 (N_41094,N_38967,N_39625);
nand U41095 (N_41095,N_38750,N_36509);
and U41096 (N_41096,N_36233,N_39295);
nand U41097 (N_41097,N_38151,N_36756);
nor U41098 (N_41098,N_39296,N_36083);
nor U41099 (N_41099,N_39729,N_37501);
and U41100 (N_41100,N_36733,N_38493);
xor U41101 (N_41101,N_35064,N_35445);
or U41102 (N_41102,N_35451,N_38223);
and U41103 (N_41103,N_37293,N_37980);
and U41104 (N_41104,N_39904,N_37763);
or U41105 (N_41105,N_36765,N_38346);
or U41106 (N_41106,N_35005,N_35254);
or U41107 (N_41107,N_38564,N_37092);
nand U41108 (N_41108,N_36878,N_35479);
xor U41109 (N_41109,N_36980,N_35651);
nand U41110 (N_41110,N_35957,N_35733);
and U41111 (N_41111,N_37383,N_36979);
nor U41112 (N_41112,N_38268,N_35788);
or U41113 (N_41113,N_37248,N_37026);
nand U41114 (N_41114,N_35949,N_35400);
nor U41115 (N_41115,N_36257,N_36554);
nand U41116 (N_41116,N_38045,N_39631);
nor U41117 (N_41117,N_36578,N_38428);
and U41118 (N_41118,N_35494,N_39147);
xor U41119 (N_41119,N_37486,N_38182);
nor U41120 (N_41120,N_38238,N_35923);
and U41121 (N_41121,N_37762,N_38927);
nand U41122 (N_41122,N_37900,N_39218);
nor U41123 (N_41123,N_36952,N_38459);
nand U41124 (N_41124,N_36129,N_36572);
nor U41125 (N_41125,N_37168,N_36857);
or U41126 (N_41126,N_37376,N_35182);
or U41127 (N_41127,N_39747,N_36468);
nand U41128 (N_41128,N_39697,N_39335);
xor U41129 (N_41129,N_37167,N_37131);
and U41130 (N_41130,N_36908,N_38731);
nand U41131 (N_41131,N_37247,N_35321);
nand U41132 (N_41132,N_36375,N_35085);
nor U41133 (N_41133,N_35028,N_38504);
and U41134 (N_41134,N_35328,N_38782);
nor U41135 (N_41135,N_36157,N_38237);
xnor U41136 (N_41136,N_38499,N_37179);
nor U41137 (N_41137,N_37345,N_37899);
or U41138 (N_41138,N_35490,N_39118);
nand U41139 (N_41139,N_35478,N_39520);
nor U41140 (N_41140,N_35395,N_37765);
nand U41141 (N_41141,N_38008,N_37063);
and U41142 (N_41142,N_37614,N_36342);
xor U41143 (N_41143,N_38167,N_38352);
and U41144 (N_41144,N_36559,N_37978);
or U41145 (N_41145,N_37400,N_36068);
nand U41146 (N_41146,N_36781,N_39799);
nor U41147 (N_41147,N_37741,N_37198);
or U41148 (N_41148,N_36754,N_36277);
or U41149 (N_41149,N_39540,N_36634);
nand U41150 (N_41150,N_39117,N_37340);
and U41151 (N_41151,N_38178,N_35104);
or U41152 (N_41152,N_37328,N_36114);
or U41153 (N_41153,N_39053,N_39203);
nor U41154 (N_41154,N_38058,N_35778);
and U41155 (N_41155,N_38214,N_37019);
nand U41156 (N_41156,N_37920,N_37647);
or U41157 (N_41157,N_39451,N_37854);
or U41158 (N_41158,N_37587,N_38961);
nor U41159 (N_41159,N_38581,N_38877);
xor U41160 (N_41160,N_37759,N_39588);
xnor U41161 (N_41161,N_38569,N_36886);
or U41162 (N_41162,N_37733,N_37513);
nor U41163 (N_41163,N_35015,N_39047);
xnor U41164 (N_41164,N_38232,N_36575);
and U41165 (N_41165,N_39691,N_37665);
or U41166 (N_41166,N_35512,N_37617);
nor U41167 (N_41167,N_37784,N_39755);
nor U41168 (N_41168,N_38220,N_37971);
or U41169 (N_41169,N_39164,N_35417);
nor U41170 (N_41170,N_39078,N_37203);
nand U41171 (N_41171,N_39193,N_36521);
and U41172 (N_41172,N_35768,N_35050);
and U41173 (N_41173,N_38780,N_38788);
or U41174 (N_41174,N_37465,N_38986);
and U41175 (N_41175,N_35550,N_39503);
nand U41176 (N_41176,N_37266,N_38973);
nor U41177 (N_41177,N_38018,N_36657);
and U41178 (N_41178,N_37227,N_35352);
and U41179 (N_41179,N_37456,N_37118);
and U41180 (N_41180,N_37048,N_35612);
or U41181 (N_41181,N_38982,N_38729);
and U41182 (N_41182,N_36185,N_39710);
xnor U41183 (N_41183,N_38785,N_35128);
and U41184 (N_41184,N_35249,N_37441);
nor U41185 (N_41185,N_35032,N_36869);
or U41186 (N_41186,N_36033,N_39415);
and U41187 (N_41187,N_39038,N_36548);
nor U41188 (N_41188,N_39752,N_37523);
nand U41189 (N_41189,N_36020,N_39717);
nand U41190 (N_41190,N_36707,N_35653);
or U41191 (N_41191,N_36433,N_36396);
and U41192 (N_41192,N_38312,N_39424);
and U41193 (N_41193,N_36311,N_36523);
xnor U41194 (N_41194,N_35933,N_38654);
xnor U41195 (N_41195,N_39834,N_38917);
nand U41196 (N_41196,N_35892,N_37588);
nor U41197 (N_41197,N_37032,N_35303);
and U41198 (N_41198,N_36386,N_36254);
nand U41199 (N_41199,N_39007,N_39135);
nand U41200 (N_41200,N_36611,N_35021);
or U41201 (N_41201,N_39827,N_38444);
or U41202 (N_41202,N_36423,N_38879);
nand U41203 (N_41203,N_39345,N_35403);
and U41204 (N_41204,N_35796,N_38758);
nor U41205 (N_41205,N_35660,N_35481);
xnor U41206 (N_41206,N_38417,N_36882);
nand U41207 (N_41207,N_39695,N_35797);
and U41208 (N_41208,N_37825,N_37982);
and U41209 (N_41209,N_37156,N_39651);
nand U41210 (N_41210,N_39359,N_39772);
or U41211 (N_41211,N_39101,N_36200);
nor U41212 (N_41212,N_35600,N_39767);
nor U41213 (N_41213,N_39810,N_39629);
nor U41214 (N_41214,N_37417,N_37276);
or U41215 (N_41215,N_38473,N_39632);
nand U41216 (N_41216,N_39671,N_35428);
and U41217 (N_41217,N_36862,N_37625);
nand U41218 (N_41218,N_38596,N_35342);
or U41219 (N_41219,N_39702,N_39323);
and U41220 (N_41220,N_38922,N_36408);
nand U41221 (N_41221,N_38603,N_35760);
and U41222 (N_41222,N_38991,N_38148);
or U41223 (N_41223,N_38507,N_39549);
nor U41224 (N_41224,N_38589,N_35248);
or U41225 (N_41225,N_35306,N_37556);
nand U41226 (N_41226,N_39802,N_37542);
nor U41227 (N_41227,N_36189,N_38633);
nor U41228 (N_41228,N_39640,N_36912);
or U41229 (N_41229,N_38285,N_38478);
or U41230 (N_41230,N_35807,N_36531);
nor U41231 (N_41231,N_35586,N_35018);
nor U41232 (N_41232,N_37363,N_39235);
nor U41233 (N_41233,N_36730,N_37714);
and U41234 (N_41234,N_38382,N_39545);
or U41235 (N_41235,N_38514,N_39249);
and U41236 (N_41236,N_36426,N_38871);
nor U41237 (N_41237,N_38429,N_36792);
xor U41238 (N_41238,N_36264,N_38477);
or U41239 (N_41239,N_35985,N_37029);
and U41240 (N_41240,N_37801,N_36706);
nand U41241 (N_41241,N_37623,N_39427);
and U41242 (N_41242,N_38302,N_39774);
nor U41243 (N_41243,N_36051,N_39828);
nor U41244 (N_41244,N_39188,N_36121);
and U41245 (N_41245,N_38433,N_35906);
or U41246 (N_41246,N_39420,N_36594);
nor U41247 (N_41247,N_37499,N_37531);
or U41248 (N_41248,N_38157,N_38117);
and U41249 (N_41249,N_39278,N_38296);
nor U41250 (N_41250,N_38010,N_39529);
or U41251 (N_41251,N_36054,N_38321);
and U41252 (N_41252,N_37239,N_36404);
or U41253 (N_41253,N_36916,N_36601);
or U41254 (N_41254,N_35357,N_36344);
nand U41255 (N_41255,N_35024,N_36418);
and U41256 (N_41256,N_39542,N_39402);
nand U41257 (N_41257,N_38131,N_39149);
and U41258 (N_41258,N_39437,N_36267);
or U41259 (N_41259,N_36527,N_37472);
and U41260 (N_41260,N_37506,N_39425);
nor U41261 (N_41261,N_37654,N_36592);
nor U41262 (N_41262,N_36076,N_39803);
or U41263 (N_41263,N_36291,N_35917);
nand U41264 (N_41264,N_36550,N_36536);
nand U41265 (N_41265,N_37817,N_37150);
and U41266 (N_41266,N_36866,N_36407);
and U41267 (N_41267,N_35346,N_38215);
and U41268 (N_41268,N_38391,N_39903);
nand U41269 (N_41269,N_39116,N_39348);
nor U41270 (N_41270,N_36901,N_36454);
or U41271 (N_41271,N_36321,N_36773);
or U41272 (N_41272,N_37373,N_37939);
and U41273 (N_41273,N_35631,N_39528);
nand U41274 (N_41274,N_38629,N_36701);
nor U41275 (N_41275,N_35301,N_35666);
and U41276 (N_41276,N_36579,N_37778);
xnor U41277 (N_41277,N_38912,N_37833);
and U41278 (N_41278,N_39239,N_39272);
or U41279 (N_41279,N_35126,N_38164);
and U41280 (N_41280,N_35502,N_35239);
and U41281 (N_41281,N_37756,N_35199);
or U41282 (N_41282,N_39199,N_35655);
nor U41283 (N_41283,N_37639,N_36379);
or U41284 (N_41284,N_38426,N_38260);
nand U41285 (N_41285,N_36703,N_37031);
and U41286 (N_41286,N_37707,N_39088);
nor U41287 (N_41287,N_38646,N_37612);
and U41288 (N_41288,N_39781,N_36852);
and U41289 (N_41289,N_37424,N_35388);
nor U41290 (N_41290,N_35468,N_37848);
or U41291 (N_41291,N_39210,N_37053);
xnor U41292 (N_41292,N_39277,N_35976);
nand U41293 (N_41293,N_37091,N_38210);
nand U41294 (N_41294,N_37270,N_37461);
nor U41295 (N_41295,N_37372,N_37207);
nand U41296 (N_41296,N_35071,N_37905);
nor U41297 (N_41297,N_37797,N_37878);
nand U41298 (N_41298,N_37910,N_38411);
nor U41299 (N_41299,N_38307,N_35511);
nand U41300 (N_41300,N_38896,N_37879);
nand U41301 (N_41301,N_36793,N_35805);
nand U41302 (N_41302,N_38409,N_36673);
xnor U41303 (N_41303,N_39346,N_35132);
nor U41304 (N_41304,N_37898,N_36354);
nor U41305 (N_41305,N_38812,N_36534);
xnor U41306 (N_41306,N_37975,N_36927);
nor U41307 (N_41307,N_36895,N_35394);
nor U41308 (N_41308,N_35569,N_37274);
nor U41309 (N_41309,N_35220,N_39108);
or U41310 (N_41310,N_39907,N_38136);
nor U41311 (N_41311,N_36248,N_36829);
nand U41312 (N_41312,N_39267,N_39737);
nor U41313 (N_41313,N_37165,N_35477);
and U41314 (N_41314,N_38643,N_39617);
nand U41315 (N_41315,N_38047,N_38019);
or U41316 (N_41316,N_36314,N_35931);
xor U41317 (N_41317,N_35025,N_35984);
nand U41318 (N_41318,N_37835,N_37205);
nor U41319 (N_41319,N_37027,N_39920);
or U41320 (N_41320,N_36976,N_35193);
nor U41321 (N_41321,N_39676,N_36676);
nand U41322 (N_41322,N_36810,N_38091);
nand U41323 (N_41323,N_36260,N_36255);
xor U41324 (N_41324,N_38207,N_38573);
and U41325 (N_41325,N_35977,N_36175);
or U41326 (N_41326,N_36146,N_35602);
or U41327 (N_41327,N_39573,N_35753);
and U41328 (N_41328,N_36826,N_36236);
and U41329 (N_41329,N_35208,N_39079);
or U41330 (N_41330,N_38923,N_37864);
and U41331 (N_41331,N_38805,N_39856);
nor U41332 (N_41332,N_39429,N_37592);
and U41333 (N_41333,N_35418,N_38301);
nor U41334 (N_41334,N_37015,N_37791);
nand U41335 (N_41335,N_37908,N_38462);
or U41336 (N_41336,N_39155,N_37375);
nor U41337 (N_41337,N_36967,N_38350);
or U41338 (N_41338,N_38036,N_35287);
nor U41339 (N_41339,N_35582,N_38869);
and U41340 (N_41340,N_36133,N_35848);
nand U41341 (N_41341,N_37969,N_37598);
and U41342 (N_41342,N_39974,N_36850);
or U41343 (N_41343,N_36606,N_36089);
xor U41344 (N_41344,N_38570,N_38840);
or U41345 (N_41345,N_35686,N_36452);
nor U41346 (N_41346,N_35821,N_35501);
and U41347 (N_41347,N_36813,N_38114);
nand U41348 (N_41348,N_38639,N_39634);
or U41349 (N_41349,N_37280,N_35618);
nor U41350 (N_41350,N_36208,N_39688);
xor U41351 (N_41351,N_36266,N_37076);
and U41352 (N_41352,N_35336,N_37860);
or U41353 (N_41353,N_38071,N_36364);
and U41354 (N_41354,N_37577,N_35911);
and U41355 (N_41355,N_38064,N_38113);
nor U41356 (N_41356,N_36497,N_39775);
nand U41357 (N_41357,N_39177,N_38261);
nand U41358 (N_41358,N_37957,N_37688);
nand U41359 (N_41359,N_39694,N_38947);
and U41360 (N_41360,N_35743,N_39000);
nor U41361 (N_41361,N_38500,N_37960);
nand U41362 (N_41362,N_36019,N_38072);
nand U41363 (N_41363,N_35564,N_35588);
and U41364 (N_41364,N_39331,N_36924);
and U41365 (N_41365,N_35966,N_35368);
or U41366 (N_41366,N_35630,N_39024);
nand U41367 (N_41367,N_37743,N_37226);
nor U41368 (N_41368,N_36376,N_38333);
xnor U41369 (N_41369,N_37923,N_36123);
or U41370 (N_41370,N_38431,N_39163);
and U41371 (N_41371,N_39417,N_36162);
and U41372 (N_41372,N_35859,N_39887);
nor U41373 (N_41373,N_35737,N_39741);
nand U41374 (N_41374,N_36780,N_36122);
and U41375 (N_41375,N_36006,N_35422);
or U41376 (N_41376,N_39211,N_36100);
and U41377 (N_41377,N_35928,N_35739);
nor U41378 (N_41378,N_36039,N_35471);
or U41379 (N_41379,N_38482,N_35773);
nand U41380 (N_41380,N_39076,N_35179);
nand U41381 (N_41381,N_38676,N_36684);
and U41382 (N_41382,N_35510,N_38195);
and U41383 (N_41383,N_35903,N_37460);
or U41384 (N_41384,N_39311,N_39106);
nor U41385 (N_41385,N_36427,N_37744);
xor U41386 (N_41386,N_35784,N_38403);
nand U41387 (N_41387,N_35238,N_37921);
nand U41388 (N_41388,N_35107,N_38836);
nor U41389 (N_41389,N_38969,N_39488);
nor U41390 (N_41390,N_39042,N_35656);
or U41391 (N_41391,N_38281,N_37819);
nand U41392 (N_41392,N_37495,N_39334);
xor U41393 (N_41393,N_35742,N_35698);
xor U41394 (N_41394,N_37594,N_38228);
and U41395 (N_41395,N_37098,N_36203);
nor U41396 (N_41396,N_39504,N_37927);
or U41397 (N_41397,N_38920,N_39305);
or U41398 (N_41398,N_36010,N_36131);
or U41399 (N_41399,N_36604,N_36449);
nor U41400 (N_41400,N_36479,N_35066);
or U41401 (N_41401,N_37225,N_39606);
nand U41402 (N_41402,N_36281,N_35070);
nor U41403 (N_41403,N_36995,N_36392);
nor U41404 (N_41404,N_37107,N_39354);
or U41405 (N_41405,N_38880,N_37883);
nor U41406 (N_41406,N_38615,N_39434);
or U41407 (N_41407,N_38614,N_35334);
or U41408 (N_41408,N_39105,N_36476);
xnor U41409 (N_41409,N_37769,N_35038);
nor U41410 (N_41410,N_35192,N_35941);
nor U41411 (N_41411,N_35904,N_39526);
xnor U41412 (N_41412,N_38191,N_36642);
or U41413 (N_41413,N_37804,N_37510);
xnor U41414 (N_41414,N_39338,N_38470);
or U41415 (N_41415,N_36377,N_38567);
nor U41416 (N_41416,N_36049,N_39062);
or U41417 (N_41417,N_39132,N_35214);
or U41418 (N_41418,N_38502,N_38875);
nor U41419 (N_41419,N_36524,N_39563);
or U41420 (N_41420,N_39138,N_38206);
nand U41421 (N_41421,N_36403,N_37214);
nor U41422 (N_41422,N_37370,N_35410);
and U41423 (N_41423,N_37984,N_39700);
nor U41424 (N_41424,N_35644,N_38730);
and U41425 (N_41425,N_38348,N_36456);
nor U41426 (N_41426,N_39726,N_38066);
nor U41427 (N_41427,N_35593,N_38475);
nand U41428 (N_41428,N_35232,N_36558);
and U41429 (N_41429,N_36989,N_38777);
nand U41430 (N_41430,N_35049,N_35298);
or U41431 (N_41431,N_37487,N_35142);
and U41432 (N_41432,N_36614,N_38587);
or U41433 (N_41433,N_39945,N_35004);
nor U41434 (N_41434,N_38762,N_37699);
nand U41435 (N_41435,N_37572,N_36460);
and U41436 (N_41436,N_36384,N_39403);
or U41437 (N_41437,N_38980,N_39018);
or U41438 (N_41438,N_36709,N_39111);
nor U41439 (N_41439,N_38921,N_38942);
and U41440 (N_41440,N_38887,N_35879);
nand U41441 (N_41441,N_38916,N_36470);
nand U41442 (N_41442,N_38042,N_37319);
nand U41443 (N_41443,N_35776,N_39157);
nand U41444 (N_41444,N_39464,N_38303);
nand U41445 (N_41445,N_38873,N_35595);
and U41446 (N_41446,N_36480,N_37467);
nor U41447 (N_41447,N_39552,N_39551);
and U41448 (N_41448,N_37095,N_37423);
or U41449 (N_41449,N_39388,N_35523);
nor U41450 (N_41450,N_38335,N_38546);
nand U41451 (N_41451,N_35020,N_37520);
nor U41452 (N_41452,N_38324,N_39012);
nand U41453 (N_41453,N_37977,N_38808);
nand U41454 (N_41454,N_37687,N_37875);
and U41455 (N_41455,N_38165,N_39875);
and U41456 (N_41456,N_38964,N_38666);
nand U41457 (N_41457,N_38263,N_36410);
and U41458 (N_41458,N_36348,N_35122);
xor U41459 (N_41459,N_36932,N_35520);
nand U41460 (N_41460,N_35749,N_37701);
or U41461 (N_41461,N_38907,N_39599);
or U41462 (N_41462,N_36800,N_37310);
or U41463 (N_41463,N_38847,N_35967);
and U41464 (N_41464,N_35498,N_39257);
and U41465 (N_41465,N_36664,N_39172);
xor U41466 (N_41466,N_37664,N_35953);
nand U41467 (N_41467,N_37335,N_35318);
and U41468 (N_41468,N_39322,N_38815);
nand U41469 (N_41469,N_36526,N_37116);
nand U41470 (N_41470,N_39921,N_37650);
nand U41471 (N_41471,N_39339,N_39985);
and U41472 (N_41472,N_39654,N_35219);
nand U41473 (N_41473,N_37524,N_39914);
nor U41474 (N_41474,N_38578,N_39713);
or U41475 (N_41475,N_36180,N_35637);
nand U41476 (N_41476,N_38026,N_38864);
nor U41477 (N_41477,N_38900,N_36613);
and U41478 (N_41478,N_35099,N_39961);
nand U41479 (N_41479,N_39905,N_38030);
or U41480 (N_41480,N_39226,N_37781);
xor U41481 (N_41481,N_36547,N_38082);
and U41482 (N_41482,N_35745,N_35525);
nor U41483 (N_41483,N_37859,N_37892);
xnor U41484 (N_41484,N_37611,N_35190);
nor U41485 (N_41485,N_37309,N_35508);
xnor U41486 (N_41486,N_36421,N_39817);
or U41487 (N_41487,N_39610,N_38385);
or U41488 (N_41488,N_39724,N_38449);
nor U41489 (N_41489,N_35131,N_37568);
or U41490 (N_41490,N_39011,N_37764);
xnor U41491 (N_41491,N_35376,N_36991);
nor U41492 (N_41492,N_39274,N_37642);
nor U41493 (N_41493,N_39245,N_37989);
or U41494 (N_41494,N_37621,N_37518);
nand U41495 (N_41495,N_38590,N_37264);
nor U41496 (N_41496,N_36821,N_38993);
and U41497 (N_41497,N_36902,N_36060);
or U41498 (N_41498,N_36088,N_37047);
nor U41499 (N_41499,N_38524,N_38425);
nand U41500 (N_41500,N_36891,N_36598);
nor U41501 (N_41501,N_35017,N_36380);
or U41502 (N_41502,N_39375,N_36889);
and U41503 (N_41503,N_36819,N_35963);
nor U41504 (N_41504,N_35672,N_35458);
xnor U41505 (N_41505,N_39123,N_36206);
and U41506 (N_41506,N_39993,N_37956);
and U41507 (N_41507,N_35925,N_38823);
xor U41508 (N_41508,N_37564,N_37464);
nor U41509 (N_41509,N_39178,N_38234);
nand U41510 (N_41510,N_38978,N_38575);
nand U41511 (N_41511,N_37055,N_38870);
nand U41512 (N_41512,N_37378,N_36897);
and U41513 (N_41513,N_35314,N_36390);
or U41514 (N_41514,N_39973,N_36313);
nand U41515 (N_41515,N_37795,N_39647);
nor U41516 (N_41516,N_38687,N_39769);
and U41517 (N_41517,N_35300,N_37172);
and U41518 (N_41518,N_35657,N_38316);
and U41519 (N_41519,N_36977,N_37449);
nor U41520 (N_41520,N_38243,N_35224);
nand U41521 (N_41521,N_39183,N_35211);
nand U41522 (N_41522,N_38001,N_37349);
nor U41523 (N_41523,N_39128,N_35710);
or U41524 (N_41524,N_35271,N_35670);
xor U41525 (N_41525,N_36935,N_38634);
and U41526 (N_41526,N_37993,N_39980);
nand U41527 (N_41527,N_36325,N_36212);
xnor U41528 (N_41528,N_36186,N_39944);
xor U41529 (N_41529,N_35166,N_38095);
nand U41530 (N_41530,N_39585,N_38868);
or U41531 (N_41531,N_35947,N_36329);
nand U41532 (N_41532,N_35908,N_38506);
xnor U41533 (N_41533,N_39984,N_36825);
xnor U41534 (N_41534,N_38291,N_36860);
and U41535 (N_41535,N_39670,N_37382);
nand U41536 (N_41536,N_37002,N_37141);
or U41537 (N_41537,N_35150,N_38118);
xnor U41538 (N_41538,N_38246,N_37099);
nor U41539 (N_41539,N_35897,N_37849);
or U41540 (N_41540,N_38820,N_38314);
and U41541 (N_41541,N_36488,N_35380);
nor U41542 (N_41542,N_37458,N_35461);
nor U41543 (N_41543,N_36584,N_37839);
and U41544 (N_41544,N_37367,N_38168);
nor U41545 (N_41545,N_35668,N_37710);
and U41546 (N_41546,N_36745,N_37222);
nand U41547 (N_41547,N_38910,N_36966);
and U41548 (N_41548,N_37422,N_38719);
or U41549 (N_41549,N_39411,N_37630);
and U41550 (N_41550,N_39766,N_35299);
or U41551 (N_41551,N_38172,N_38775);
nor U41552 (N_41552,N_37703,N_36757);
xor U41553 (N_41553,N_37129,N_36272);
nor U41554 (N_41554,N_37272,N_37070);
nand U41555 (N_41555,N_36622,N_38427);
nand U41556 (N_41556,N_36391,N_37540);
or U41557 (N_41557,N_39414,N_36761);
or U41558 (N_41558,N_36669,N_37365);
nand U41559 (N_41559,N_36316,N_39158);
xor U41560 (N_41560,N_38355,N_38754);
and U41561 (N_41561,N_35524,N_39156);
nor U41562 (N_41562,N_38672,N_37712);
nand U41563 (N_41563,N_37497,N_36116);
nand U41564 (N_41564,N_38574,N_39003);
or U41565 (N_41565,N_38783,N_39431);
and U41566 (N_41566,N_38611,N_35579);
nor U41567 (N_41567,N_36214,N_36920);
nand U41568 (N_41568,N_36283,N_35517);
xor U41569 (N_41569,N_38022,N_37886);
nor U41570 (N_41570,N_36457,N_36235);
nand U41571 (N_41571,N_37005,N_38283);
nor U41572 (N_41572,N_39865,N_36753);
and U41573 (N_41573,N_38313,N_35082);
nor U41574 (N_41574,N_36681,N_37758);
nor U41575 (N_41575,N_35288,N_36680);
nand U41576 (N_41576,N_39347,N_37705);
or U41577 (N_41577,N_38941,N_36929);
nor U41578 (N_41578,N_36164,N_37397);
and U41579 (N_41579,N_36750,N_39209);
or U41580 (N_41580,N_39473,N_36493);
nor U41581 (N_41581,N_36950,N_37887);
xor U41582 (N_41582,N_39969,N_36273);
nand U41583 (N_41583,N_36434,N_36693);
and U41584 (N_41584,N_37816,N_38813);
nor U41585 (N_41585,N_38231,N_39597);
nor U41586 (N_41586,N_35849,N_37629);
nor U41587 (N_41587,N_39673,N_35683);
or U41588 (N_41588,N_36946,N_37477);
nand U41589 (N_41589,N_35751,N_37263);
nor U41590 (N_41590,N_36570,N_38955);
and U41591 (N_41591,N_38693,N_37407);
nor U41592 (N_41592,N_37873,N_39259);
and U41593 (N_41593,N_39300,N_36299);
nand U41594 (N_41594,N_39937,N_38209);
or U41595 (N_41595,N_37393,N_37610);
nor U41596 (N_41596,N_39214,N_38055);
nor U41597 (N_41597,N_36668,N_37036);
nor U41598 (N_41598,N_39892,N_38827);
and U41599 (N_41599,N_39321,N_38717);
xnor U41600 (N_41600,N_38906,N_39958);
nand U41601 (N_41601,N_38772,N_35704);
and U41602 (N_41602,N_39580,N_35841);
nor U41603 (N_41603,N_35793,N_39355);
or U41604 (N_41604,N_36140,N_39954);
nand U41605 (N_41605,N_38240,N_36469);
nand U41606 (N_41606,N_38764,N_36621);
or U41607 (N_41607,N_38224,N_38940);
and U41608 (N_41608,N_36290,N_37601);
or U41609 (N_41609,N_39782,N_38384);
xor U41610 (N_41610,N_39630,N_39760);
or U41611 (N_41611,N_35474,N_39663);
nand U41612 (N_41612,N_39708,N_37525);
nand U41613 (N_41613,N_36616,N_37948);
and U41614 (N_41614,N_39041,N_38000);
nand U41615 (N_41615,N_39704,N_37426);
or U41616 (N_41616,N_37803,N_37694);
nand U41617 (N_41617,N_39832,N_37125);
or U41618 (N_41618,N_35129,N_35936);
or U41619 (N_41619,N_38467,N_35226);
and U41620 (N_41620,N_36571,N_36795);
xnor U41621 (N_41621,N_37946,N_36659);
nand U41622 (N_41622,N_39979,N_37618);
nor U41623 (N_41623,N_38098,N_36752);
nor U41624 (N_41624,N_38585,N_37970);
nand U41625 (N_41625,N_35120,N_39998);
and U41626 (N_41626,N_39197,N_35833);
nand U41627 (N_41627,N_39064,N_37863);
xor U41628 (N_41628,N_36383,N_35980);
nand U41629 (N_41629,N_37159,N_38239);
nand U41630 (N_41630,N_39564,N_38225);
and U41631 (N_41631,N_37735,N_35103);
nand U41632 (N_41632,N_38831,N_37597);
nand U41633 (N_41633,N_39715,N_35359);
and U41634 (N_41634,N_39720,N_39337);
nor U41635 (N_41635,N_37698,N_35167);
nand U41636 (N_41636,N_39198,N_39611);
nand U41637 (N_41637,N_37871,N_38658);
nand U41638 (N_41638,N_39888,N_36147);
xor U41639 (N_41639,N_35152,N_37730);
nand U41640 (N_41640,N_38620,N_35961);
or U41641 (N_41641,N_37256,N_39635);
nor U41642 (N_41642,N_37284,N_37530);
and U41643 (N_41643,N_36288,N_36241);
xor U41644 (N_41644,N_37736,N_39250);
or U41645 (N_41645,N_36885,N_38796);
nand U41646 (N_41646,N_37767,N_35096);
and U41647 (N_41647,N_37115,N_35261);
and U41648 (N_41648,N_38833,N_38854);
nand U41649 (N_41649,N_37258,N_38380);
nand U41650 (N_41650,N_37269,N_38174);
and U41651 (N_41651,N_35645,N_39786);
nand U41652 (N_41652,N_36959,N_36686);
nor U41653 (N_41653,N_38161,N_37243);
nor U41654 (N_41654,N_39302,N_39751);
or U41655 (N_41655,N_38739,N_37213);
or U41656 (N_41656,N_38751,N_39236);
nor U41657 (N_41657,N_37802,N_35794);
xnor U41658 (N_41658,N_37996,N_38440);
or U41659 (N_41659,N_36398,N_38915);
and U41660 (N_41660,N_38414,N_36445);
or U41661 (N_41661,N_35383,N_37779);
and U41662 (N_41662,N_35130,N_38051);
nor U41663 (N_41663,N_38720,N_36093);
or U41664 (N_41664,N_37853,N_36202);
nor U41665 (N_41665,N_36666,N_36050);
or U41666 (N_41666,N_36549,N_36128);
or U41667 (N_41667,N_37163,N_39501);
and U41668 (N_41668,N_36749,N_39363);
or U41669 (N_41669,N_37231,N_38811);
nor U41670 (N_41670,N_36726,N_37446);
nand U41671 (N_41671,N_39566,N_35408);
or U41672 (N_41672,N_38399,N_38465);
nand U41673 (N_41673,N_37483,N_37811);
or U41674 (N_41674,N_36489,N_38435);
or U41675 (N_41675,N_39519,N_38104);
nor U41676 (N_41676,N_37346,N_39733);
nor U41677 (N_41677,N_37217,N_39004);
or U41678 (N_41678,N_39538,N_35648);
nor U41679 (N_41679,N_36336,N_35606);
and U41680 (N_41680,N_38147,N_35554);
and U41681 (N_41681,N_38274,N_39261);
nand U41682 (N_41682,N_36542,N_37271);
and U41683 (N_41683,N_38450,N_37641);
nand U41684 (N_41684,N_38488,N_35460);
and U41685 (N_41685,N_37327,N_35136);
or U41686 (N_41686,N_35056,N_36356);
nor U41687 (N_41687,N_37858,N_36289);
nand U41688 (N_41688,N_39404,N_36428);
or U41689 (N_41689,N_36005,N_36764);
nor U41690 (N_41690,N_37682,N_36746);
and U41691 (N_41691,N_38821,N_35390);
and U41692 (N_41692,N_37999,N_36787);
and U41693 (N_41693,N_38888,N_36734);
nand U41694 (N_41694,N_38339,N_35116);
nor U41695 (N_41695,N_35635,N_37153);
xnor U41696 (N_41696,N_38375,N_35054);
or U41697 (N_41697,N_36098,N_39281);
and U41698 (N_41698,N_38159,N_38700);
or U41699 (N_41699,N_39390,N_36627);
or U41700 (N_41700,N_37615,N_37438);
and U41701 (N_41701,N_36772,N_36573);
nor U41702 (N_41702,N_37334,N_38867);
nand U41703 (N_41703,N_39124,N_37808);
or U41704 (N_41704,N_37997,N_39590);
nand U41705 (N_41705,N_36401,N_39085);
and U41706 (N_41706,N_38850,N_39438);
or U41707 (N_41707,N_39870,N_37148);
or U41708 (N_41708,N_37541,N_35764);
or U41709 (N_41709,N_37358,N_36001);
nor U41710 (N_41710,N_39858,N_37691);
and U41711 (N_41711,N_38601,N_35223);
xor U41712 (N_41712,N_37755,N_38108);
nor U41713 (N_41713,N_39683,N_39935);
nor U41714 (N_41714,N_39039,N_37130);
nor U41715 (N_41715,N_35780,N_35544);
and U41716 (N_41716,N_39366,N_39965);
nor U41717 (N_41717,N_38511,N_38299);
or U41718 (N_41718,N_39576,N_35430);
and U41719 (N_41719,N_39407,N_37001);
nand U41720 (N_41720,N_36253,N_35938);
or U41721 (N_41721,N_38039,N_38565);
or U41722 (N_41722,N_38732,N_36170);
or U41723 (N_41723,N_38793,N_35175);
nand U41724 (N_41724,N_38323,N_37428);
nor U41725 (N_41725,N_36105,N_39057);
or U41726 (N_41726,N_39258,N_38859);
nand U41727 (N_41727,N_38400,N_35688);
and U41728 (N_41728,N_38130,N_38774);
or U41729 (N_41729,N_37616,N_38367);
nand U41730 (N_41730,N_36794,N_35370);
or U41731 (N_41731,N_36516,N_37493);
xor U41732 (N_41732,N_37596,N_36435);
nor U41733 (N_41733,N_38819,N_38273);
nand U41734 (N_41734,N_38679,N_37354);
xnor U41735 (N_41735,N_38084,N_35509);
and U41736 (N_41736,N_38555,N_38267);
nor U41737 (N_41737,N_35905,N_39521);
nor U41738 (N_41738,N_37952,N_37496);
or U41739 (N_41739,N_35790,N_39725);
xor U41740 (N_41740,N_37752,N_36081);
nand U41741 (N_41741,N_36103,N_36351);
or U41742 (N_41742,N_36863,N_36502);
and U41743 (N_41743,N_36903,N_39166);
xor U41744 (N_41744,N_39689,N_37009);
nand U41745 (N_41745,N_36873,N_36893);
nor U41746 (N_41746,N_39304,N_39622);
or U41747 (N_41747,N_35706,N_37127);
nand U41748 (N_41748,N_37979,N_35877);
or U41749 (N_41749,N_38845,N_37075);
nor U41750 (N_41750,N_37392,N_39146);
nand U41751 (N_41751,N_38592,N_35608);
nand U41752 (N_41752,N_39889,N_37155);
or U41753 (N_41753,N_37425,N_36762);
and U41754 (N_41754,N_37893,N_39762);
nand U41755 (N_41755,N_36219,N_37855);
and U41756 (N_41756,N_39661,N_35405);
nand U41757 (N_41757,N_39453,N_36271);
or U41758 (N_41758,N_36926,N_36292);
nor U41759 (N_41759,N_35173,N_36827);
xor U41760 (N_41760,N_36815,N_37128);
xor U41761 (N_41761,N_35215,N_37268);
xor U41762 (N_41762,N_35217,N_39658);
xnor U41763 (N_41763,N_37224,N_37315);
nor U41764 (N_41764,N_37238,N_38127);
and U41765 (N_41765,N_38485,N_38767);
and U41766 (N_41766,N_35449,N_39016);
or U41767 (N_41767,N_38804,N_35640);
or U41768 (N_41768,N_35098,N_36644);
nand U41769 (N_41769,N_36018,N_39405);
nor U41770 (N_41770,N_38883,N_38749);
xor U41771 (N_41771,N_36357,N_36228);
or U41772 (N_41772,N_36070,N_35036);
xnor U41773 (N_41773,N_37241,N_38144);
nand U41774 (N_41774,N_39571,N_35222);
and U41775 (N_41775,N_38368,N_37938);
nor U41776 (N_41776,N_37450,N_35504);
and U41777 (N_41777,N_38139,N_38438);
and U41778 (N_41778,N_37582,N_36341);
or U41779 (N_41779,N_39196,N_36096);
nor U41780 (N_41780,N_39723,N_37934);
and U41781 (N_41781,N_39562,N_36691);
xor U41782 (N_41782,N_37937,N_38170);
nor U41783 (N_41783,N_37232,N_38526);
and U41784 (N_41784,N_37876,N_37692);
xor U41785 (N_41785,N_36163,N_35315);
or U41786 (N_41786,N_35609,N_36142);
or U41787 (N_41787,N_37668,N_38242);
and U41788 (N_41788,N_35438,N_35364);
nor U41789 (N_41789,N_39790,N_38892);
nor U41790 (N_41790,N_35277,N_36607);
nor U41791 (N_41791,N_35213,N_35819);
nand U41792 (N_41792,N_38093,N_37008);
and U41793 (N_41793,N_37575,N_39797);
or U41794 (N_41794,N_39898,N_37563);
nand U41795 (N_41795,N_39205,N_37356);
nor U41796 (N_41796,N_37175,N_35874);
xor U41797 (N_41797,N_37024,N_35326);
or U41798 (N_41798,N_36156,N_36429);
or U41799 (N_41799,N_36079,N_37431);
or U41800 (N_41800,N_39619,N_35986);
nor U41801 (N_41801,N_37176,N_38038);
nand U41802 (N_41802,N_35055,N_36145);
or U41803 (N_41803,N_37800,N_38496);
or U41804 (N_41804,N_37669,N_36925);
or U41805 (N_41805,N_37786,N_35035);
or U41806 (N_41806,N_37813,N_36909);
nor U41807 (N_41807,N_39805,N_35060);
or U41808 (N_41808,N_35292,N_39829);
or U41809 (N_41809,N_39119,N_38256);
xnor U41810 (N_41810,N_37251,N_38571);
or U41811 (N_41811,N_36589,N_39418);
nor U41812 (N_41812,N_36209,N_39861);
or U41813 (N_41813,N_37387,N_37723);
nor U41814 (N_41814,N_36303,N_36913);
and U41815 (N_41815,N_39997,N_35373);
nor U41816 (N_41816,N_36215,N_39192);
nand U41817 (N_41817,N_35800,N_38599);
and U41818 (N_41818,N_39028,N_38077);
and U41819 (N_41819,N_38460,N_35338);
nand U41820 (N_41820,N_37995,N_38644);
nand U41821 (N_41821,N_35726,N_39692);
nand U41822 (N_41822,N_36478,N_39964);
or U41823 (N_41823,N_35633,N_38545);
nand U41824 (N_41824,N_37240,N_35680);
and U41825 (N_41825,N_38318,N_39150);
nor U41826 (N_41826,N_38641,N_38125);
nor U41827 (N_41827,N_37831,N_37585);
or U41828 (N_41828,N_37935,N_35397);
or U41829 (N_41829,N_35858,N_39792);
xnor U41830 (N_41830,N_39975,N_36711);
and U41831 (N_41831,N_36983,N_38624);
nor U41832 (N_41832,N_38422,N_39299);
nand U41833 (N_41833,N_38718,N_39567);
xor U41834 (N_41834,N_37674,N_36743);
xor U41835 (N_41835,N_37591,N_39092);
nand U41836 (N_41836,N_35309,N_35639);
nor U41837 (N_41837,N_35845,N_39533);
nand U41838 (N_41838,N_39065,N_36335);
and U41839 (N_41839,N_38011,N_37985);
nor U41840 (N_41840,N_38765,N_38392);
nand U41841 (N_41841,N_36247,N_36310);
xnor U41842 (N_41842,N_38582,N_39234);
or U41843 (N_41843,N_39579,N_39371);
nand U41844 (N_41844,N_35310,N_37081);
or U41845 (N_41845,N_36875,N_37228);
nor U41846 (N_41846,N_35267,N_37017);
and U41847 (N_41847,N_37279,N_35465);
and U41848 (N_41848,N_38711,N_38636);
nand U41849 (N_41849,N_35731,N_39266);
or U41850 (N_41850,N_38171,N_36448);
xnor U41851 (N_41851,N_39731,N_38897);
nand U41852 (N_41852,N_39672,N_39040);
nand U41853 (N_41853,N_37190,N_35002);
nand U41854 (N_41854,N_35801,N_37021);
and U41855 (N_41855,N_36027,N_38387);
or U41856 (N_41856,N_39187,N_38607);
nor U41857 (N_41857,N_39853,N_35124);
nor U41858 (N_41858,N_39310,N_38061);
xor U41859 (N_41859,N_35282,N_35703);
or U41860 (N_41860,N_36899,N_35885);
and U41861 (N_41861,N_38175,N_36295);
nand U41862 (N_41862,N_38760,N_37545);
nand U41863 (N_41863,N_35365,N_39216);
nand U41864 (N_41864,N_35557,N_35427);
nor U41865 (N_41865,N_38315,N_38249);
and U41866 (N_41866,N_38512,N_36304);
nand U41867 (N_41867,N_35484,N_36414);
nand U41868 (N_41868,N_36165,N_38378);
xnor U41869 (N_41869,N_37250,N_39142);
or U41870 (N_41870,N_36546,N_35043);
nand U41871 (N_41871,N_35625,N_39089);
and U41872 (N_41872,N_35003,N_35272);
xnor U41873 (N_41873,N_38716,N_37022);
and U41874 (N_41874,N_35194,N_39823);
nand U41875 (N_41875,N_35094,N_35577);
nor U41876 (N_41876,N_38956,N_36065);
or U41877 (N_41877,N_38025,N_36280);
nor U41878 (N_41878,N_37379,N_35423);
or U41879 (N_41879,N_39344,N_37401);
and U41880 (N_41880,N_36000,N_37014);
and U41881 (N_41881,N_38481,N_36467);
nor U41882 (N_41882,N_38598,N_38974);
and U41883 (N_41883,N_36193,N_39844);
nand U41884 (N_41884,N_37275,N_35720);
nand U41885 (N_41885,N_38272,N_36173);
xnor U41886 (N_41886,N_36017,N_37963);
nand U41887 (N_41887,N_37521,N_38056);
nor U41888 (N_41888,N_37870,N_35997);
nand U41889 (N_41889,N_36134,N_35930);
and U41890 (N_41890,N_37595,N_36441);
nor U41891 (N_41891,N_36118,N_39650);
nor U41892 (N_41892,N_38735,N_35507);
and U41893 (N_41893,N_35951,N_35127);
nor U41894 (N_41894,N_35295,N_38895);
nand U41895 (N_41895,N_39824,N_38623);
xor U41896 (N_41896,N_38994,N_36424);
nor U41897 (N_41897,N_36665,N_35158);
nor U41898 (N_41898,N_38872,N_39820);
nor U41899 (N_41899,N_35758,N_37850);
nor U41900 (N_41900,N_38456,N_38162);
nand U41901 (N_41901,N_35276,N_36530);
nor U41902 (N_41902,N_39465,N_38200);
or U41903 (N_41903,N_37448,N_37242);
or U41904 (N_41904,N_35284,N_38548);
and U41905 (N_41905,N_36471,N_37565);
nand U41906 (N_41906,N_36465,N_38100);
nor U41907 (N_41907,N_39894,N_36347);
xnor U41908 (N_41908,N_35597,N_36736);
xnor U41909 (N_41909,N_38280,N_39613);
nor U41910 (N_41910,N_35701,N_35915);
and U41911 (N_41911,N_36551,N_38287);
nor U41912 (N_41912,N_39190,N_36225);
nand U41913 (N_41913,N_37902,N_39073);
or U41914 (N_41914,N_35762,N_36982);
and U41915 (N_41915,N_36818,N_38972);
and U41916 (N_41916,N_36809,N_35791);
nor U41917 (N_41917,N_39730,N_37504);
nand U41918 (N_41918,N_39764,N_38925);
nand U41919 (N_41919,N_37655,N_35757);
and U41920 (N_41920,N_35470,N_38270);
nand U41921 (N_41921,N_38489,N_37414);
nor U41922 (N_41922,N_39584,N_35355);
nand U41923 (N_41923,N_38699,N_38521);
and U41924 (N_41924,N_36540,N_35188);
and U41925 (N_41925,N_36933,N_38112);
nor U41926 (N_41926,N_37547,N_38608);
xnor U41927 (N_41927,N_36141,N_39698);
nor U41928 (N_41928,N_39594,N_39524);
nor U41929 (N_41929,N_37579,N_37312);
nor U41930 (N_41930,N_39855,N_36442);
nor U41931 (N_41931,N_37473,N_39495);
nor U41932 (N_41932,N_35662,N_35181);
xor U41933 (N_41933,N_38446,N_39994);
xnor U41934 (N_41934,N_39428,N_36876);
xor U41935 (N_41935,N_35696,N_37018);
or U41936 (N_41936,N_36327,N_38276);
nor U41937 (N_41937,N_39890,N_37581);
nor U41938 (N_41938,N_36567,N_35183);
nand U41939 (N_41939,N_37546,N_38371);
xnor U41940 (N_41940,N_36366,N_37637);
nor U41941 (N_41941,N_36004,N_35839);
or U41942 (N_41942,N_37812,N_38087);
nor U41943 (N_41943,N_35678,N_39107);
or U41944 (N_41944,N_37097,N_36724);
or U41945 (N_41945,N_39255,N_35605);
xor U41946 (N_41946,N_37492,N_39317);
or U41947 (N_41947,N_38944,N_35543);
or U41948 (N_41948,N_35170,N_38149);
nor U41949 (N_41949,N_37221,N_35384);
or U41950 (N_41950,N_38954,N_38550);
nor U41951 (N_41951,N_36440,N_39636);
xnor U41952 (N_41952,N_36360,N_38977);
and U41953 (N_41953,N_36400,N_37489);
nor U41954 (N_41954,N_39821,N_35485);
nand U41955 (N_41955,N_39735,N_36194);
nand U41956 (N_41956,N_37114,N_38132);
nand U41957 (N_41957,N_37646,N_39227);
xnor U41958 (N_41958,N_37321,N_37025);
and U41959 (N_41959,N_39721,N_36646);
nor U41960 (N_41960,N_35347,N_36318);
nand U41961 (N_41961,N_39063,N_37466);
or U41962 (N_41962,N_39966,N_37006);
or U41963 (N_41963,N_37967,N_37210);
or U41964 (N_41964,N_37149,N_38057);
nor U41965 (N_41965,N_39883,N_39342);
nor U41966 (N_41966,N_38219,N_36207);
and U41967 (N_41967,N_37868,N_35061);
or U41968 (N_41968,N_37416,N_35902);
nor U41969 (N_41969,N_36044,N_36500);
nand U41970 (N_41970,N_35133,N_37326);
nor U41971 (N_41971,N_37503,N_36154);
and U41972 (N_41972,N_36931,N_37058);
nand U41973 (N_41973,N_39380,N_36097);
nor U41974 (N_41974,N_39406,N_39301);
nor U41975 (N_41975,N_39463,N_36775);
or U41976 (N_41976,N_37237,N_37693);
nand U41977 (N_41977,N_37192,N_36978);
or U41978 (N_41978,N_35993,N_39109);
or U41979 (N_41979,N_37079,N_39422);
or U41980 (N_41980,N_36014,N_38129);
nand U41981 (N_41981,N_35846,N_38632);
nor U41982 (N_41982,N_36052,N_36603);
or U41983 (N_41983,N_36760,N_35297);
nand U41984 (N_41984,N_38192,N_37020);
xnor U41985 (N_41985,N_36582,N_36626);
or U41986 (N_41986,N_36822,N_36072);
or U41987 (N_41987,N_36723,N_38851);
and U41988 (N_41988,N_37535,N_39472);
nand U41989 (N_41989,N_38951,N_35294);
or U41990 (N_41990,N_36274,N_39223);
and U41991 (N_41991,N_36986,N_37722);
and U41992 (N_41992,N_35857,N_39086);
nand U41993 (N_41993,N_39862,N_35924);
nand U41994 (N_41994,N_36633,N_36884);
nor U41995 (N_41995,N_38668,N_35135);
and U41996 (N_41996,N_37229,N_37314);
and U41997 (N_41997,N_36269,N_35450);
and U41998 (N_41998,N_39818,N_38115);
nand U41999 (N_41999,N_36937,N_38227);
or U42000 (N_42000,N_37173,N_37822);
nand U42001 (N_42001,N_39684,N_36333);
and U42002 (N_42002,N_37798,N_35724);
nand U42003 (N_42003,N_35847,N_39970);
nand U42004 (N_42004,N_35341,N_37724);
xor U42005 (N_42005,N_39454,N_38293);
and U42006 (N_42006,N_39014,N_36282);
nor U42007 (N_42007,N_39110,N_38505);
xor U42008 (N_42008,N_36956,N_35200);
or U42009 (N_42009,N_35402,N_36940);
xor U42010 (N_42010,N_38649,N_39121);
xnor U42011 (N_42011,N_35591,N_36416);
and U42012 (N_42012,N_36922,N_38769);
or U42013 (N_42013,N_35533,N_36075);
and U42014 (N_42014,N_35840,N_37366);
or U42015 (N_42015,N_39525,N_37478);
nand U42016 (N_42016,N_38212,N_35782);
nor U42017 (N_42017,N_39612,N_37751);
nand U42018 (N_42018,N_35664,N_37789);
nand U42019 (N_42019,N_36801,N_37409);
nand U42020 (N_42020,N_35059,N_39312);
nand U42021 (N_42021,N_39539,N_38245);
or U42022 (N_42022,N_35443,N_39485);
and U42023 (N_42023,N_39548,N_36695);
or U42024 (N_42024,N_35850,N_36883);
xor U42025 (N_42025,N_38988,N_37195);
or U42026 (N_42026,N_37657,N_37719);
or U42027 (N_42027,N_37306,N_35817);
nor U42028 (N_42028,N_38519,N_35761);
nor U42029 (N_42029,N_36610,N_36417);
nor U42030 (N_42030,N_38074,N_36259);
xor U42031 (N_42031,N_35203,N_38137);
or U42032 (N_42032,N_39290,N_35392);
nand U42033 (N_42033,N_39430,N_35147);
or U42034 (N_42034,N_36969,N_38975);
nor U42035 (N_42035,N_38931,N_37402);
and U42036 (N_42036,N_39370,N_39598);
or U42037 (N_42037,N_36455,N_36623);
or U42038 (N_42038,N_38377,N_37262);
or U42039 (N_42039,N_37519,N_35441);
nand U42040 (N_42040,N_36261,N_37832);
nand U42041 (N_42041,N_38103,N_35583);
and U42042 (N_42042,N_38903,N_36635);
and U42043 (N_42043,N_36667,N_36574);
or U42044 (N_42044,N_38097,N_38745);
nand U42045 (N_42045,N_39353,N_39591);
and U42046 (N_42046,N_39441,N_39745);
and U42047 (N_42047,N_35378,N_38650);
nand U42048 (N_42048,N_39200,N_35480);
or U42049 (N_42049,N_39067,N_39857);
and U42050 (N_42050,N_38390,N_39685);
xnor U42051 (N_42051,N_37066,N_35454);
xor U42052 (N_42052,N_35781,N_35172);
or U42053 (N_42053,N_38776,N_35658);
xor U42054 (N_42054,N_37561,N_38725);
nand U42055 (N_42055,N_36178,N_35534);
or U42056 (N_42056,N_35119,N_36696);
nor U42057 (N_42057,N_37897,N_36008);
or U42058 (N_42058,N_36221,N_38089);
nor U42059 (N_42059,N_39141,N_36964);
xnor U42060 (N_42060,N_39776,N_39768);
and U42061 (N_42061,N_36422,N_38262);
and U42062 (N_42062,N_36624,N_39605);
nor U42063 (N_42063,N_37395,N_37429);
nor U42064 (N_42064,N_37622,N_39208);
nor U42065 (N_42065,N_36204,N_39120);
nor U42066 (N_42066,N_37209,N_38653);
or U42067 (N_42067,N_37869,N_38987);
and U42068 (N_42068,N_35311,N_35558);
and U42069 (N_42069,N_35361,N_37074);
and U42070 (N_42070,N_37583,N_35391);
nor U42071 (N_42071,N_38704,N_36231);
nor U42072 (N_42072,N_39328,N_38286);
and U42073 (N_42073,N_38048,N_39831);
nor U42074 (N_42074,N_35439,N_39010);
and U42075 (N_42075,N_37419,N_38908);
or U42076 (N_42076,N_36182,N_37660);
and U42077 (N_42077,N_36565,N_35171);
nand U42078 (N_42078,N_39779,N_39019);
xnor U42079 (N_42079,N_36708,N_37161);
nand U42080 (N_42080,N_37044,N_37738);
nand U42081 (N_42081,N_36769,N_35202);
or U42082 (N_42082,N_35868,N_36367);
or U42083 (N_42083,N_35285,N_37180);
or U42084 (N_42084,N_36965,N_38696);
or U42085 (N_42085,N_37083,N_38816);
or U42086 (N_42086,N_38543,N_35818);
or U42087 (N_42087,N_36620,N_37245);
nor U42088 (N_42088,N_36774,N_37932);
xor U42089 (N_42089,N_39959,N_35413);
nor U42090 (N_42090,N_35125,N_38517);
nor U42091 (N_42091,N_35001,N_37170);
nor U42092 (N_42092,N_38756,N_36517);
and U42093 (N_42093,N_35062,N_37273);
nor U42094 (N_42094,N_36687,N_37453);
and U42095 (N_42095,N_35675,N_38248);
nor U42096 (N_42096,N_39162,N_36415);
nand U42097 (N_42097,N_38937,N_38759);
and U42098 (N_42098,N_35795,N_35312);
and U42099 (N_42099,N_35944,N_39825);
nor U42100 (N_42100,N_39445,N_37442);
and U42101 (N_42101,N_35123,N_35563);
nor U42102 (N_42102,N_39416,N_39743);
or U42103 (N_42103,N_38661,N_37865);
and U42104 (N_42104,N_38205,N_38216);
nand U42105 (N_42105,N_35528,N_37342);
or U42106 (N_42106,N_37632,N_35014);
nor U42107 (N_42107,N_36220,N_35473);
and U42108 (N_42108,N_35245,N_36671);
nor U42109 (N_42109,N_38305,N_37512);
and U42110 (N_42110,N_35555,N_36656);
or U42111 (N_42111,N_39212,N_36694);
nor U42112 (N_42112,N_39789,N_39811);
nand U42113 (N_42113,N_35459,N_37560);
nand U42114 (N_42114,N_38561,N_37772);
or U42115 (N_42115,N_37841,N_37359);
or U42116 (N_42116,N_35153,N_36538);
or U42117 (N_42117,N_36504,N_37259);
nand U42118 (N_42118,N_38405,N_36474);
nand U42119 (N_42119,N_37285,N_37567);
nor U42120 (N_42120,N_35659,N_39005);
or U42121 (N_42121,N_37140,N_35044);
xor U42122 (N_42122,N_38169,N_36945);
and U42123 (N_42123,N_37678,N_38359);
or U42124 (N_42124,N_38652,N_35149);
or U42125 (N_42125,N_37930,N_35765);
nor U42126 (N_42126,N_37644,N_35886);
or U42127 (N_42127,N_36322,N_36590);
or U42128 (N_42128,N_37211,N_39678);
and U42129 (N_42129,N_37684,N_37748);
nand U42130 (N_42130,N_36349,N_38235);
nand U42131 (N_42131,N_36561,N_39784);
and U42132 (N_42132,N_39243,N_36759);
nand U42133 (N_42133,N_39707,N_39452);
nor U42134 (N_42134,N_38647,N_36638);
xnor U42135 (N_42135,N_37911,N_35008);
nor U42136 (N_42136,N_36172,N_36879);
nand U42137 (N_42137,N_39144,N_38317);
and U42138 (N_42138,N_35115,N_35244);
and U42139 (N_42139,N_39444,N_39320);
and U42140 (N_42140,N_35700,N_38451);
nand U42141 (N_42141,N_37307,N_35324);
nand U42142 (N_42142,N_38184,N_37606);
nor U42143 (N_42143,N_39901,N_35537);
nor U42144 (N_42144,N_36125,N_39787);
or U42145 (N_42145,N_38510,N_38365);
xor U42146 (N_42146,N_38300,N_38600);
nand U42147 (N_42147,N_35667,N_36914);
nor U42148 (N_42148,N_36074,N_35747);
xor U42149 (N_42149,N_39229,N_38929);
or U42150 (N_42150,N_39433,N_38376);
xnor U42151 (N_42151,N_36024,N_35880);
or U42152 (N_42152,N_36963,N_37384);
nor U42153 (N_42153,N_35308,N_37322);
nor U42154 (N_42154,N_35278,N_36106);
or U42155 (N_42155,N_35253,N_35013);
nor U42156 (N_42156,N_38141,N_37042);
nand U42157 (N_42157,N_37470,N_35252);
and U42158 (N_42158,N_35307,N_37154);
nand U42159 (N_42159,N_39008,N_39356);
nand U42160 (N_42160,N_35505,N_36438);
nor U42161 (N_42161,N_38562,N_35363);
and U42162 (N_42162,N_39951,N_38630);
nand U42163 (N_42163,N_39389,N_39361);
or U42164 (N_42164,N_39174,N_37432);
nor U42165 (N_42165,N_38740,N_39221);
nor U42166 (N_42166,N_36326,N_35843);
nand U42167 (N_42167,N_38340,N_35499);
and U42168 (N_42168,N_39381,N_36943);
and U42169 (N_42169,N_38580,N_37337);
nor U42170 (N_42170,N_37144,N_38695);
nor U42171 (N_42171,N_39446,N_36464);
nand U42172 (N_42172,N_36338,N_35057);
nor U42173 (N_42173,N_39918,N_38684);
nand U42174 (N_42174,N_38989,N_38495);
nor U42175 (N_42175,N_35854,N_35545);
or U42176 (N_42176,N_38447,N_39561);
and U42177 (N_42177,N_39645,N_35293);
or U42178 (N_42178,N_37498,N_36370);
or U42179 (N_42179,N_35138,N_38976);
nor U42180 (N_42180,N_38768,N_38553);
xnor U42181 (N_42181,N_35433,N_39759);
and U42182 (N_42182,N_39412,N_37338);
nor U42183 (N_42183,N_36890,N_39711);
or U42184 (N_42184,N_39706,N_38595);
xor U42185 (N_42185,N_36921,N_36361);
nor U42186 (N_42186,N_39026,N_38789);
and U42187 (N_42187,N_36655,N_38755);
or U42188 (N_42188,N_39699,N_36217);
or U42189 (N_42189,N_35567,N_35968);
or U42190 (N_42190,N_39482,N_36812);
xnor U42191 (N_42191,N_37290,N_39977);
and U42192 (N_42192,N_37983,N_38932);
nand U42193 (N_42193,N_39455,N_35741);
or U42194 (N_42194,N_36084,N_35827);
nor U42195 (N_42195,N_38733,N_39667);
or U42196 (N_42196,N_36420,N_36712);
or U42197 (N_42197,N_37122,N_36374);
nand U42198 (N_42198,N_37082,N_37830);
nand U42199 (N_42199,N_35362,N_35230);
nand U42200 (N_42200,N_39025,N_38016);
and U42201 (N_42201,N_39327,N_36328);
nand U42202 (N_42202,N_38282,N_36135);
nand U42203 (N_42203,N_36482,N_37308);
xnor U42204 (N_42204,N_36218,N_37457);
xnor U42205 (N_42205,N_37677,N_38278);
and U42206 (N_42206,N_39639,N_38572);
nand U42207 (N_42207,N_39586,N_39866);
or U42208 (N_42208,N_37381,N_36679);
nor U42209 (N_42209,N_38829,N_37823);
and U42210 (N_42210,N_38953,N_35815);
or U42211 (N_42211,N_38119,N_39991);
xnor U42212 (N_42212,N_37435,N_35809);
and U42213 (N_42213,N_38155,N_36791);
or U42214 (N_42214,N_39559,N_39442);
nand U42215 (N_42215,N_38251,N_36836);
xor U42216 (N_42216,N_39165,N_36915);
nor U42217 (N_42217,N_37191,N_36320);
nor U42218 (N_42218,N_39368,N_39497);
nor U42219 (N_42219,N_39492,N_39215);
or U42220 (N_42220,N_36224,N_38472);
and U42221 (N_42221,N_37578,N_39056);
and U42222 (N_42222,N_36631,N_38968);
and U42223 (N_42223,N_39669,N_39690);
and U42224 (N_42224,N_39849,N_37427);
nor U42225 (N_42225,N_38017,N_35178);
nor U42226 (N_42226,N_36334,N_39570);
nand U42227 (N_42227,N_38406,N_38542);
and U42228 (N_42228,N_36245,N_37094);
nand U42229 (N_42229,N_37729,N_39360);
xor U42230 (N_42230,N_39125,N_39280);
and U42231 (N_42231,N_36102,N_36988);
xnor U42232 (N_42232,N_35177,N_37283);
nand U42233 (N_42233,N_37502,N_35725);
nor U42234 (N_42234,N_38959,N_36727);
nor U42235 (N_42235,N_35514,N_37713);
nor U42236 (N_42236,N_37640,N_38656);
or U42237 (N_42237,N_37966,N_39876);
and U42238 (N_42238,N_38229,N_35853);
and U42239 (N_42239,N_36844,N_35112);
nor U42240 (N_42240,N_39791,N_36637);
nor U42241 (N_42241,N_36262,N_38208);
nor U42242 (N_42242,N_39880,N_35488);
or U42243 (N_42243,N_36716,N_35561);
and U42244 (N_42244,N_35160,N_36252);
xnor U42245 (N_42245,N_38874,N_39096);
nand U42246 (N_42246,N_39537,N_39246);
nand U42247 (N_42247,N_37134,N_39286);
nand U42248 (N_42248,N_39744,N_38105);
xnor U42249 (N_42249,N_35283,N_35325);
nand U42250 (N_42250,N_39194,N_39535);
and U42251 (N_42251,N_38233,N_38525);
and U42252 (N_42252,N_38487,N_35000);
or U42253 (N_42253,N_36617,N_35270);
nand U42254 (N_42254,N_37286,N_36942);
nor U42255 (N_42255,N_38957,N_38692);
and U42256 (N_42256,N_35255,N_36993);
nand U42257 (N_42257,N_39728,N_37517);
or U42258 (N_42258,N_38893,N_35425);
or U42259 (N_42259,N_39507,N_39989);
or U42260 (N_42260,N_37103,N_35735);
nor U42261 (N_42261,N_35467,N_35201);
nor U42262 (N_42262,N_36002,N_39130);
or U42263 (N_42263,N_36996,N_36962);
or U42264 (N_42264,N_38309,N_37016);
and U42265 (N_42265,N_36672,N_37360);
nor U42266 (N_42266,N_35862,N_39850);
nor U42267 (N_42267,N_37511,N_35596);
nand U42268 (N_42268,N_38551,N_39325);
or U42269 (N_42269,N_37557,N_37662);
or U42270 (N_42270,N_35069,N_37410);
nand U42271 (N_42271,N_36038,N_39986);
nor U42272 (N_42272,N_38373,N_37888);
or U42273 (N_42273,N_35676,N_35620);
and U42274 (N_42274,N_38023,N_37403);
nor U42275 (N_42275,N_35076,N_37586);
nor U42276 (N_42276,N_37685,N_36115);
nand U42277 (N_42277,N_35051,N_36833);
or U42278 (N_42278,N_36543,N_35955);
xor U42279 (N_42279,N_37636,N_35209);
or U42280 (N_42280,N_35871,N_38985);
and U42281 (N_42281,N_39927,N_35358);
and U42282 (N_42282,N_35615,N_35109);
or U42283 (N_42283,N_36466,N_37011);
or U42284 (N_42284,N_37894,N_39324);
nand U42285 (N_42285,N_36413,N_39553);
xor U42286 (N_42286,N_35108,N_38063);
nand U42287 (N_42287,N_38648,N_38779);
nand U42288 (N_42288,N_38354,N_37943);
or U42289 (N_42289,N_39734,N_36766);
nand U42290 (N_42290,N_36641,N_36783);
and U42291 (N_42291,N_39534,N_36159);
or U42292 (N_42292,N_39499,N_39126);
nor U42293 (N_42293,N_38992,N_37500);
and U42294 (N_42294,N_35262,N_37369);
xor U42295 (N_42295,N_35891,N_38715);
nor U42296 (N_42296,N_36498,N_38092);
nand U42297 (N_42297,N_36503,N_36802);
nand U42298 (N_42298,N_39034,N_35137);
or U42299 (N_42299,N_38748,N_36588);
nor U42300 (N_42300,N_35759,N_35573);
nand U42301 (N_42301,N_35575,N_39665);
and U42302 (N_42302,N_39666,N_35493);
nor U42303 (N_42303,N_39490,N_36953);
and U42304 (N_42304,N_37715,N_37697);
and U42305 (N_42305,N_38374,N_35139);
or U42306 (N_42306,N_39601,N_35803);
xnor U42307 (N_42307,N_38657,N_39777);
or U42308 (N_42308,N_38437,N_37658);
and U42309 (N_42309,N_35616,N_37933);
xnor U42310 (N_42310,N_35959,N_36153);
and U42311 (N_42311,N_39271,N_39653);
or U42312 (N_42312,N_36187,N_36569);
or U42313 (N_42313,N_38645,N_37043);
or U42314 (N_42314,N_35313,N_36970);
nor U42315 (N_42315,N_37656,N_38351);
nor U42316 (N_42316,N_36596,N_36025);
nand U42317 (N_42317,N_37197,N_35826);
xor U42318 (N_42318,N_38640,N_37810);
or U42319 (N_42319,N_37045,N_36645);
nand U42320 (N_42320,N_35503,N_37408);
nor U42321 (N_42321,N_39397,N_36643);
nand U42322 (N_42322,N_36167,N_37101);
nand U42323 (N_42323,N_35638,N_37352);
or U42324 (N_42324,N_36537,N_36443);
and U42325 (N_42325,N_35681,N_37679);
xnor U42326 (N_42326,N_35442,N_35110);
or U42327 (N_42327,N_38616,N_38277);
nor U42328 (N_42328,N_37088,N_36744);
and U42329 (N_42329,N_38014,N_36807);
or U42330 (N_42330,N_39341,N_36918);
or U42331 (N_42331,N_36636,N_35053);
nand U42332 (N_42332,N_38761,N_37534);
xor U42333 (N_42333,N_36007,N_35432);
and U42334 (N_42334,N_38690,N_36294);
xnor U42335 (N_42335,N_37538,N_35187);
or U42336 (N_42336,N_38454,N_36308);
nand U42337 (N_42337,N_39336,N_35162);
and U42338 (N_42338,N_35327,N_36071);
nand U42339 (N_42339,N_36697,N_37396);
or U42340 (N_42340,N_36169,N_36839);
or U42341 (N_42341,N_36871,N_39066);
nor U42342 (N_42342,N_38529,N_36195);
nand U42343 (N_42343,N_36747,N_35921);
xor U42344 (N_42344,N_37105,N_37689);
and U42345 (N_42345,N_36040,N_36095);
or U42346 (N_42346,N_37842,N_36751);
xor U42347 (N_42347,N_36577,N_36767);
nor U42348 (N_42348,N_38707,N_39621);
or U42349 (N_42349,N_39967,N_37316);
or U42350 (N_42350,N_35406,N_37529);
or U42351 (N_42351,N_37829,N_36350);
xor U42352 (N_42352,N_38002,N_36847);
or U42353 (N_42353,N_37794,N_39251);
xnor U42354 (N_42354,N_38791,N_39902);
and U42355 (N_42355,N_36544,N_36205);
nand U42356 (N_42356,N_39783,N_35552);
nand U42357 (N_42357,N_35950,N_35539);
nand U42358 (N_42358,N_37716,N_38250);
or U42359 (N_42359,N_39587,N_35813);
or U42360 (N_42360,N_36127,N_37186);
or U42361 (N_42361,N_36037,N_36911);
nor U42362 (N_42362,N_37146,N_38665);
xor U42363 (N_42363,N_39449,N_38464);
nor U42364 (N_42364,N_38678,N_38642);
nor U42365 (N_42365,N_36625,N_35482);
or U42366 (N_42366,N_36085,N_36499);
or U42367 (N_42367,N_39558,N_37686);
or U42368 (N_42368,N_36339,N_38401);
xor U42369 (N_42369,N_37780,N_35114);
xnor U42370 (N_42370,N_36305,N_36568);
or U42371 (N_42371,N_35233,N_35476);
and U42372 (N_42372,N_38659,N_38343);
nor U42373 (N_42373,N_36046,N_36605);
xor U42374 (N_42374,N_36090,N_39136);
and U42375 (N_42375,N_36529,N_38911);
nand U42376 (N_42376,N_35727,N_38905);
and U42377 (N_42377,N_38043,N_37318);
nand U42378 (N_42378,N_38222,N_39104);
nand U42379 (N_42379,N_39819,N_36080);
nand U42380 (N_42380,N_35998,N_38822);
or U42381 (N_42381,N_36067,N_35927);
or U42382 (N_42382,N_37925,N_36583);
and U42383 (N_42383,N_36419,N_37121);
or U42384 (N_42384,N_39410,N_36120);
or U42385 (N_42385,N_38617,N_38342);
or U42386 (N_42386,N_37548,N_36229);
nor U42387 (N_42387,N_38710,N_38356);
xnor U42388 (N_42388,N_39264,N_39409);
xnor U42389 (N_42389,N_36842,N_37368);
xnor U42390 (N_42390,N_35259,N_36677);
and U42391 (N_42391,N_37077,N_38306);
nand U42392 (N_42392,N_36064,N_35970);
and U42393 (N_42393,N_35396,N_38602);
and U42394 (N_42394,N_37792,N_35632);
xnor U42395 (N_42395,N_38626,N_37278);
and U42396 (N_42396,N_38484,N_39701);
nor U42397 (N_42397,N_38538,N_36888);
nor U42398 (N_42398,N_35437,N_38397);
nor U42399 (N_42399,N_36735,N_39001);
nor U42400 (N_42400,N_35518,N_35198);
or U42401 (N_42401,N_36651,N_36867);
or U42402 (N_42402,N_38153,N_37361);
and U42403 (N_42403,N_35572,N_35372);
or U42404 (N_42404,N_39240,N_38876);
or U42405 (N_42405,N_36576,N_36692);
and U42406 (N_42406,N_35738,N_37942);
nor U42407 (N_42407,N_35263,N_38494);
xnor U42408 (N_42408,N_37437,N_38453);
nor U42409 (N_42409,N_39122,N_36483);
and U42410 (N_42410,N_36674,N_39099);
nor U42411 (N_42411,N_36910,N_36353);
xnor U42412 (N_42412,N_37060,N_36012);
nand U42413 (N_42413,N_39303,N_37265);
nand U42414 (N_42414,N_37681,N_38814);
and U42415 (N_42415,N_38290,N_39863);
nor U42416 (N_42416,N_38798,N_38843);
nand U42417 (N_42417,N_39273,N_37880);
xnor U42418 (N_42418,N_35331,N_35319);
and U42419 (N_42419,N_35317,N_37292);
nor U42420 (N_42420,N_35987,N_39624);
nor U42421 (N_42421,N_38960,N_35895);
xor U42422 (N_42422,N_39990,N_38914);
and U42423 (N_42423,N_35964,N_37233);
nor U42424 (N_42424,N_35067,N_39282);
and U42425 (N_42425,N_35852,N_36494);
nand U42426 (N_42426,N_38746,N_37139);
and U42427 (N_42427,N_36560,N_35012);
and U42428 (N_42428,N_38471,N_36363);
nand U42429 (N_42429,N_36016,N_38541);
nand U42430 (N_42430,N_36654,N_38588);
xor U42431 (N_42431,N_38094,N_35581);
nor U42432 (N_42432,N_35221,N_35052);
or U42433 (N_42433,N_36101,N_37820);
nor U42434 (N_42434,N_35598,N_35234);
nand U42435 (N_42435,N_39230,N_39021);
nor U42436 (N_42436,N_37090,N_38320);
and U42437 (N_42437,N_35385,N_35140);
and U42438 (N_42438,N_35424,N_38394);
or U42439 (N_42439,N_38441,N_36682);
nor U42440 (N_42440,N_36602,N_36987);
nor U42441 (N_42441,N_39058,N_35870);
nand U42442 (N_42442,N_38396,N_36934);
or U42443 (N_42443,N_38295,N_38713);
xor U42444 (N_42444,N_36073,N_39736);
nand U42445 (N_42445,N_36309,N_36799);
nand U42446 (N_42446,N_38034,N_39367);
nor U42447 (N_42447,N_36315,N_37745);
or U42448 (N_42448,N_39992,N_39423);
nand U42449 (N_42449,N_39815,N_35999);
and U42450 (N_42450,N_35079,N_39995);
and U42451 (N_42451,N_39947,N_35838);
nor U42452 (N_42452,N_36861,N_38736);
nor U42453 (N_42453,N_35972,N_35105);
nor U42454 (N_42454,N_36181,N_35540);
nand U42455 (N_42455,N_38345,N_37086);
and U42456 (N_42456,N_37852,N_38803);
nand U42457 (N_42457,N_37821,N_35824);
or U42458 (N_42458,N_37675,N_35566);
and U42459 (N_42459,N_36199,N_39536);
and U42460 (N_42460,N_36035,N_36184);
nand U42461 (N_42461,N_37953,N_38826);
xor U42462 (N_42462,N_35191,N_35830);
nor U42463 (N_42463,N_39841,N_39626);
nand U42464 (N_42464,N_35080,N_35716);
nand U42465 (N_42465,N_35876,N_35515);
nor U42466 (N_42466,N_38020,N_37463);
nand U42467 (N_42467,N_37296,N_35369);
and U42468 (N_42468,N_37624,N_39400);
nor U42469 (N_42469,N_35415,N_36770);
nor U42470 (N_42470,N_35799,N_36306);
or U42471 (N_42471,N_39732,N_37033);
and U42472 (N_42472,N_36359,N_39620);
nor U42473 (N_42473,N_36811,N_35578);
nor U42474 (N_42474,N_39382,N_35952);
nand U42475 (N_42475,N_36462,N_36705);
or U42476 (N_42476,N_39837,N_36275);
nor U42477 (N_42477,N_36069,N_39383);
nand U42478 (N_42478,N_38364,N_35323);
xor U42479 (N_42479,N_35161,N_38361);
nor U42480 (N_42480,N_37023,N_39401);
or U42481 (N_42481,N_37126,N_35074);
xor U42482 (N_42482,N_35556,N_38420);
nand U42483 (N_42483,N_35289,N_38552);
and U42484 (N_42484,N_38508,N_36763);
and U42485 (N_42485,N_36119,N_37412);
nor U42486 (N_42486,N_35143,N_37734);
nor U42487 (N_42487,N_38185,N_37528);
nand U42488 (N_42488,N_38842,N_36975);
nor U42489 (N_42489,N_36047,N_38140);
nor U42490 (N_42490,N_37867,N_35356);
nand U42491 (N_42491,N_39179,N_39313);
or U42492 (N_42492,N_38241,N_39738);
or U42493 (N_42493,N_39386,N_35031);
or U42494 (N_42494,N_36501,N_38838);
or U42495 (N_42495,N_35497,N_39169);
and U42496 (N_42496,N_38685,N_38421);
xor U42497 (N_42497,N_37291,N_37325);
and U42498 (N_42498,N_38591,N_36508);
and U42499 (N_42499,N_36648,N_39917);
nand U42500 (N_42500,N_35000,N_39182);
or U42501 (N_42501,N_37654,N_37210);
nor U42502 (N_42502,N_36678,N_35892);
and U42503 (N_42503,N_38969,N_37591);
or U42504 (N_42504,N_39696,N_37748);
xor U42505 (N_42505,N_38427,N_39595);
nor U42506 (N_42506,N_38251,N_37902);
nor U42507 (N_42507,N_38256,N_37192);
or U42508 (N_42508,N_39113,N_38112);
nor U42509 (N_42509,N_35463,N_39382);
or U42510 (N_42510,N_39881,N_35622);
nand U42511 (N_42511,N_37053,N_38905);
xnor U42512 (N_42512,N_36353,N_36309);
nor U42513 (N_42513,N_39237,N_37852);
and U42514 (N_42514,N_36662,N_35768);
nor U42515 (N_42515,N_38477,N_35861);
or U42516 (N_42516,N_36036,N_35437);
or U42517 (N_42517,N_35126,N_39130);
xor U42518 (N_42518,N_37515,N_37127);
or U42519 (N_42519,N_36781,N_38477);
and U42520 (N_42520,N_37107,N_37719);
nand U42521 (N_42521,N_38102,N_36820);
xnor U42522 (N_42522,N_38667,N_38875);
or U42523 (N_42523,N_37687,N_38244);
nor U42524 (N_42524,N_36456,N_35394);
nor U42525 (N_42525,N_39030,N_36811);
or U42526 (N_42526,N_35102,N_37731);
or U42527 (N_42527,N_39673,N_35354);
and U42528 (N_42528,N_36512,N_37333);
or U42529 (N_42529,N_36863,N_39947);
nor U42530 (N_42530,N_39121,N_35595);
and U42531 (N_42531,N_37082,N_37663);
nor U42532 (N_42532,N_38759,N_36872);
or U42533 (N_42533,N_39322,N_35304);
xnor U42534 (N_42534,N_35038,N_36539);
nand U42535 (N_42535,N_36459,N_35088);
nor U42536 (N_42536,N_39626,N_36601);
and U42537 (N_42537,N_39276,N_35098);
xor U42538 (N_42538,N_37658,N_37185);
and U42539 (N_42539,N_39262,N_37006);
and U42540 (N_42540,N_38766,N_36320);
xnor U42541 (N_42541,N_38869,N_35485);
or U42542 (N_42542,N_35442,N_38126);
and U42543 (N_42543,N_36629,N_39843);
xor U42544 (N_42544,N_37135,N_39538);
nand U42545 (N_42545,N_37114,N_35356);
or U42546 (N_42546,N_35263,N_39149);
and U42547 (N_42547,N_39523,N_37309);
or U42548 (N_42548,N_35655,N_35982);
nor U42549 (N_42549,N_39726,N_35589);
nor U42550 (N_42550,N_35737,N_37189);
or U42551 (N_42551,N_39856,N_36406);
nor U42552 (N_42552,N_38783,N_35299);
xor U42553 (N_42553,N_35068,N_35179);
and U42554 (N_42554,N_39014,N_36417);
and U42555 (N_42555,N_39109,N_39586);
nor U42556 (N_42556,N_39191,N_39391);
or U42557 (N_42557,N_36387,N_38320);
xnor U42558 (N_42558,N_38742,N_35623);
nor U42559 (N_42559,N_38142,N_39445);
nand U42560 (N_42560,N_39431,N_36793);
nor U42561 (N_42561,N_36033,N_38041);
nand U42562 (N_42562,N_36068,N_35577);
nand U42563 (N_42563,N_35827,N_38138);
and U42564 (N_42564,N_36326,N_38703);
nor U42565 (N_42565,N_38724,N_38420);
nand U42566 (N_42566,N_37771,N_39962);
nor U42567 (N_42567,N_37419,N_39783);
or U42568 (N_42568,N_36147,N_36459);
nor U42569 (N_42569,N_38118,N_36544);
and U42570 (N_42570,N_37447,N_35178);
nand U42571 (N_42571,N_35285,N_39719);
nor U42572 (N_42572,N_36805,N_39828);
and U42573 (N_42573,N_35197,N_37836);
nor U42574 (N_42574,N_36514,N_36758);
nand U42575 (N_42575,N_38875,N_38642);
nor U42576 (N_42576,N_37046,N_37909);
nand U42577 (N_42577,N_39382,N_38125);
nor U42578 (N_42578,N_39595,N_39124);
nor U42579 (N_42579,N_36736,N_38783);
nand U42580 (N_42580,N_36290,N_36471);
nor U42581 (N_42581,N_35886,N_38149);
xor U42582 (N_42582,N_37462,N_38209);
and U42583 (N_42583,N_35296,N_37143);
and U42584 (N_42584,N_38499,N_38762);
xnor U42585 (N_42585,N_36914,N_39313);
nand U42586 (N_42586,N_37371,N_37269);
or U42587 (N_42587,N_38999,N_38090);
or U42588 (N_42588,N_36193,N_39392);
or U42589 (N_42589,N_37095,N_35700);
nor U42590 (N_42590,N_38209,N_36165);
nor U42591 (N_42591,N_36055,N_37148);
or U42592 (N_42592,N_38788,N_38491);
and U42593 (N_42593,N_39936,N_36027);
and U42594 (N_42594,N_37351,N_35769);
nor U42595 (N_42595,N_39593,N_39731);
nor U42596 (N_42596,N_35513,N_35729);
nor U42597 (N_42597,N_36474,N_39621);
nor U42598 (N_42598,N_39536,N_37660);
nor U42599 (N_42599,N_36247,N_39494);
or U42600 (N_42600,N_39031,N_39240);
nor U42601 (N_42601,N_36294,N_39295);
nor U42602 (N_42602,N_38805,N_36867);
or U42603 (N_42603,N_35930,N_38328);
nand U42604 (N_42604,N_38948,N_37279);
nand U42605 (N_42605,N_37524,N_38342);
and U42606 (N_42606,N_35981,N_35204);
nand U42607 (N_42607,N_36640,N_38612);
or U42608 (N_42608,N_35266,N_38344);
xor U42609 (N_42609,N_37244,N_35743);
or U42610 (N_42610,N_36841,N_35807);
nor U42611 (N_42611,N_39947,N_35353);
and U42612 (N_42612,N_38008,N_37242);
nor U42613 (N_42613,N_39125,N_39262);
nand U42614 (N_42614,N_39003,N_36191);
and U42615 (N_42615,N_39577,N_36932);
and U42616 (N_42616,N_38329,N_36917);
xnor U42617 (N_42617,N_36095,N_36000);
and U42618 (N_42618,N_39981,N_35946);
or U42619 (N_42619,N_37336,N_36502);
or U42620 (N_42620,N_36040,N_37636);
and U42621 (N_42621,N_39939,N_36396);
or U42622 (N_42622,N_38763,N_37543);
and U42623 (N_42623,N_37397,N_36577);
nor U42624 (N_42624,N_38397,N_39864);
and U42625 (N_42625,N_35998,N_38094);
or U42626 (N_42626,N_35252,N_38654);
or U42627 (N_42627,N_37143,N_38842);
xor U42628 (N_42628,N_39329,N_38865);
or U42629 (N_42629,N_39852,N_38744);
or U42630 (N_42630,N_39601,N_35958);
xnor U42631 (N_42631,N_38756,N_37422);
or U42632 (N_42632,N_35405,N_38677);
nor U42633 (N_42633,N_37229,N_36100);
or U42634 (N_42634,N_39768,N_35947);
nand U42635 (N_42635,N_37960,N_37545);
nand U42636 (N_42636,N_35293,N_37835);
and U42637 (N_42637,N_38953,N_35505);
or U42638 (N_42638,N_39108,N_37533);
and U42639 (N_42639,N_37039,N_35424);
or U42640 (N_42640,N_37922,N_38532);
nor U42641 (N_42641,N_37010,N_38603);
nor U42642 (N_42642,N_39770,N_37504);
xor U42643 (N_42643,N_35146,N_37148);
nand U42644 (N_42644,N_37374,N_35447);
and U42645 (N_42645,N_39762,N_39974);
and U42646 (N_42646,N_38553,N_37076);
nand U42647 (N_42647,N_39488,N_36333);
nor U42648 (N_42648,N_39833,N_38694);
nand U42649 (N_42649,N_36016,N_37552);
nand U42650 (N_42650,N_38857,N_35760);
or U42651 (N_42651,N_35953,N_35362);
nor U42652 (N_42652,N_37305,N_39306);
and U42653 (N_42653,N_38851,N_37883);
xnor U42654 (N_42654,N_36524,N_39026);
xnor U42655 (N_42655,N_35543,N_39054);
nand U42656 (N_42656,N_37593,N_37924);
xor U42657 (N_42657,N_35816,N_36234);
xor U42658 (N_42658,N_36233,N_38661);
or U42659 (N_42659,N_37334,N_39677);
nor U42660 (N_42660,N_37159,N_35740);
nand U42661 (N_42661,N_36359,N_36474);
and U42662 (N_42662,N_36297,N_35449);
and U42663 (N_42663,N_38840,N_35340);
xnor U42664 (N_42664,N_37276,N_39148);
xor U42665 (N_42665,N_38205,N_39751);
and U42666 (N_42666,N_35762,N_35617);
nand U42667 (N_42667,N_39125,N_39784);
nand U42668 (N_42668,N_36488,N_39162);
nor U42669 (N_42669,N_39113,N_35630);
nand U42670 (N_42670,N_37952,N_37472);
nand U42671 (N_42671,N_35551,N_35477);
nor U42672 (N_42672,N_36992,N_37934);
nor U42673 (N_42673,N_35993,N_37637);
nor U42674 (N_42674,N_36981,N_38141);
or U42675 (N_42675,N_39191,N_38476);
nand U42676 (N_42676,N_37285,N_35475);
nand U42677 (N_42677,N_39554,N_39295);
nor U42678 (N_42678,N_35864,N_36647);
and U42679 (N_42679,N_39800,N_37861);
xnor U42680 (N_42680,N_39040,N_38968);
nor U42681 (N_42681,N_39632,N_35174);
and U42682 (N_42682,N_39854,N_38790);
or U42683 (N_42683,N_38555,N_35294);
xnor U42684 (N_42684,N_38652,N_35114);
or U42685 (N_42685,N_39139,N_36397);
and U42686 (N_42686,N_35218,N_38003);
or U42687 (N_42687,N_38337,N_38066);
xnor U42688 (N_42688,N_37752,N_38087);
or U42689 (N_42689,N_35466,N_36791);
and U42690 (N_42690,N_35589,N_36398);
and U42691 (N_42691,N_38949,N_38957);
nor U42692 (N_42692,N_35378,N_36431);
xor U42693 (N_42693,N_37958,N_36041);
or U42694 (N_42694,N_37007,N_38046);
or U42695 (N_42695,N_36176,N_36144);
and U42696 (N_42696,N_37603,N_39483);
nor U42697 (N_42697,N_36651,N_36661);
nor U42698 (N_42698,N_39025,N_36310);
nor U42699 (N_42699,N_35220,N_36488);
and U42700 (N_42700,N_38601,N_39070);
nand U42701 (N_42701,N_38755,N_39130);
nand U42702 (N_42702,N_35139,N_39265);
nand U42703 (N_42703,N_38501,N_38129);
or U42704 (N_42704,N_37875,N_36854);
and U42705 (N_42705,N_37278,N_38835);
or U42706 (N_42706,N_37208,N_39409);
and U42707 (N_42707,N_36576,N_38633);
nand U42708 (N_42708,N_35379,N_39037);
nor U42709 (N_42709,N_35094,N_39734);
or U42710 (N_42710,N_39067,N_38138);
and U42711 (N_42711,N_36173,N_35708);
and U42712 (N_42712,N_38633,N_38199);
or U42713 (N_42713,N_38862,N_36124);
nor U42714 (N_42714,N_36094,N_39925);
nand U42715 (N_42715,N_39585,N_36533);
nand U42716 (N_42716,N_37128,N_38236);
or U42717 (N_42717,N_39590,N_38544);
nor U42718 (N_42718,N_37066,N_39021);
nand U42719 (N_42719,N_38080,N_36087);
or U42720 (N_42720,N_37099,N_36114);
or U42721 (N_42721,N_36796,N_36618);
or U42722 (N_42722,N_39538,N_35193);
or U42723 (N_42723,N_35222,N_35258);
and U42724 (N_42724,N_39402,N_37186);
nand U42725 (N_42725,N_39900,N_37537);
nor U42726 (N_42726,N_35448,N_36661);
and U42727 (N_42727,N_37882,N_38259);
and U42728 (N_42728,N_36539,N_37165);
nor U42729 (N_42729,N_37567,N_38717);
xnor U42730 (N_42730,N_36414,N_39438);
and U42731 (N_42731,N_37679,N_36157);
nand U42732 (N_42732,N_39248,N_35268);
or U42733 (N_42733,N_37347,N_37225);
or U42734 (N_42734,N_35076,N_38597);
and U42735 (N_42735,N_37028,N_39510);
and U42736 (N_42736,N_39738,N_38249);
or U42737 (N_42737,N_38291,N_39119);
and U42738 (N_42738,N_36727,N_37914);
nor U42739 (N_42739,N_38374,N_37678);
nand U42740 (N_42740,N_36653,N_36602);
nand U42741 (N_42741,N_39441,N_38403);
or U42742 (N_42742,N_37181,N_36982);
or U42743 (N_42743,N_37602,N_39734);
and U42744 (N_42744,N_37463,N_35880);
nor U42745 (N_42745,N_37872,N_36081);
or U42746 (N_42746,N_35304,N_35683);
nand U42747 (N_42747,N_35969,N_38987);
or U42748 (N_42748,N_37046,N_37092);
and U42749 (N_42749,N_38954,N_35128);
nor U42750 (N_42750,N_35306,N_37935);
and U42751 (N_42751,N_35892,N_39371);
and U42752 (N_42752,N_37975,N_36792);
xor U42753 (N_42753,N_39342,N_35788);
nor U42754 (N_42754,N_39404,N_38504);
nor U42755 (N_42755,N_39315,N_36572);
nor U42756 (N_42756,N_37535,N_37197);
nand U42757 (N_42757,N_37264,N_36627);
or U42758 (N_42758,N_37504,N_38213);
and U42759 (N_42759,N_37577,N_35958);
or U42760 (N_42760,N_37905,N_35723);
xor U42761 (N_42761,N_37411,N_36134);
or U42762 (N_42762,N_38508,N_36950);
or U42763 (N_42763,N_36150,N_38272);
and U42764 (N_42764,N_38129,N_38025);
or U42765 (N_42765,N_35906,N_38925);
nor U42766 (N_42766,N_35546,N_39010);
xor U42767 (N_42767,N_38865,N_36080);
nor U42768 (N_42768,N_38668,N_35508);
nor U42769 (N_42769,N_35967,N_39885);
and U42770 (N_42770,N_38240,N_38773);
xnor U42771 (N_42771,N_39660,N_35872);
or U42772 (N_42772,N_37899,N_37386);
and U42773 (N_42773,N_37651,N_36086);
xnor U42774 (N_42774,N_35496,N_35835);
and U42775 (N_42775,N_37783,N_38047);
and U42776 (N_42776,N_39239,N_39830);
or U42777 (N_42777,N_38187,N_38998);
nand U42778 (N_42778,N_38003,N_39294);
nor U42779 (N_42779,N_35182,N_39160);
and U42780 (N_42780,N_35085,N_37725);
or U42781 (N_42781,N_35719,N_38416);
nor U42782 (N_42782,N_35677,N_39359);
nand U42783 (N_42783,N_39244,N_38480);
xnor U42784 (N_42784,N_35302,N_39347);
or U42785 (N_42785,N_37984,N_36574);
and U42786 (N_42786,N_36242,N_35129);
xor U42787 (N_42787,N_36291,N_38003);
and U42788 (N_42788,N_38010,N_37240);
nand U42789 (N_42789,N_39779,N_37075);
xnor U42790 (N_42790,N_35944,N_37901);
nand U42791 (N_42791,N_38198,N_38243);
or U42792 (N_42792,N_36363,N_35616);
and U42793 (N_42793,N_38136,N_37421);
and U42794 (N_42794,N_35317,N_37112);
nand U42795 (N_42795,N_36022,N_36650);
and U42796 (N_42796,N_35976,N_36227);
or U42797 (N_42797,N_38102,N_36615);
or U42798 (N_42798,N_37930,N_39800);
xor U42799 (N_42799,N_35058,N_38244);
or U42800 (N_42800,N_39490,N_36260);
nand U42801 (N_42801,N_36168,N_36353);
and U42802 (N_42802,N_35519,N_38231);
and U42803 (N_42803,N_39548,N_36162);
nand U42804 (N_42804,N_36716,N_39468);
xor U42805 (N_42805,N_39720,N_39496);
or U42806 (N_42806,N_36457,N_35274);
and U42807 (N_42807,N_39837,N_37073);
and U42808 (N_42808,N_35996,N_38558);
nor U42809 (N_42809,N_36140,N_39614);
or U42810 (N_42810,N_36791,N_35258);
or U42811 (N_42811,N_38314,N_37305);
nand U42812 (N_42812,N_37075,N_35875);
nor U42813 (N_42813,N_35675,N_38306);
xnor U42814 (N_42814,N_38359,N_35664);
or U42815 (N_42815,N_36662,N_36124);
nand U42816 (N_42816,N_35540,N_36959);
or U42817 (N_42817,N_35817,N_36236);
or U42818 (N_42818,N_36091,N_36150);
nand U42819 (N_42819,N_39741,N_38055);
xnor U42820 (N_42820,N_37029,N_36037);
and U42821 (N_42821,N_36038,N_38647);
or U42822 (N_42822,N_38563,N_36210);
nor U42823 (N_42823,N_35056,N_39255);
or U42824 (N_42824,N_37316,N_38622);
nor U42825 (N_42825,N_38969,N_37378);
or U42826 (N_42826,N_39679,N_36259);
nand U42827 (N_42827,N_38855,N_37862);
and U42828 (N_42828,N_38717,N_36477);
nor U42829 (N_42829,N_38254,N_38659);
nor U42830 (N_42830,N_35888,N_38761);
nor U42831 (N_42831,N_38160,N_38739);
and U42832 (N_42832,N_37840,N_35870);
or U42833 (N_42833,N_38103,N_35926);
xnor U42834 (N_42834,N_39831,N_38409);
nand U42835 (N_42835,N_39610,N_35372);
nor U42836 (N_42836,N_36352,N_37397);
and U42837 (N_42837,N_35773,N_37687);
or U42838 (N_42838,N_39487,N_35731);
nor U42839 (N_42839,N_37517,N_37042);
nor U42840 (N_42840,N_39802,N_36008);
or U42841 (N_42841,N_35021,N_38942);
nor U42842 (N_42842,N_39965,N_35375);
nor U42843 (N_42843,N_38225,N_38549);
nand U42844 (N_42844,N_39999,N_36777);
and U42845 (N_42845,N_38145,N_36393);
nor U42846 (N_42846,N_39560,N_38654);
nand U42847 (N_42847,N_36767,N_35047);
and U42848 (N_42848,N_37981,N_39731);
nand U42849 (N_42849,N_36034,N_36161);
and U42850 (N_42850,N_37569,N_37536);
nor U42851 (N_42851,N_35672,N_39402);
nand U42852 (N_42852,N_35891,N_39479);
and U42853 (N_42853,N_37347,N_37389);
nand U42854 (N_42854,N_38639,N_37925);
or U42855 (N_42855,N_38269,N_36045);
nand U42856 (N_42856,N_37771,N_35222);
nand U42857 (N_42857,N_36370,N_39880);
nor U42858 (N_42858,N_35080,N_37271);
nor U42859 (N_42859,N_37146,N_38859);
nand U42860 (N_42860,N_39132,N_37516);
nor U42861 (N_42861,N_39217,N_39197);
nand U42862 (N_42862,N_35647,N_36070);
and U42863 (N_42863,N_37483,N_38912);
xor U42864 (N_42864,N_36870,N_35050);
or U42865 (N_42865,N_39495,N_36269);
and U42866 (N_42866,N_38541,N_37970);
nor U42867 (N_42867,N_38583,N_35185);
or U42868 (N_42868,N_39005,N_39877);
or U42869 (N_42869,N_36229,N_38986);
or U42870 (N_42870,N_37454,N_35857);
nor U42871 (N_42871,N_39361,N_36689);
and U42872 (N_42872,N_35766,N_35684);
nand U42873 (N_42873,N_38204,N_39318);
nand U42874 (N_42874,N_39008,N_39127);
nand U42875 (N_42875,N_38357,N_39350);
or U42876 (N_42876,N_37331,N_38026);
and U42877 (N_42877,N_35090,N_35225);
nand U42878 (N_42878,N_35774,N_35671);
and U42879 (N_42879,N_38251,N_37098);
and U42880 (N_42880,N_37477,N_35003);
and U42881 (N_42881,N_37725,N_38082);
or U42882 (N_42882,N_37821,N_39928);
nand U42883 (N_42883,N_39173,N_37783);
nand U42884 (N_42884,N_39037,N_39354);
xor U42885 (N_42885,N_36029,N_39263);
nor U42886 (N_42886,N_35199,N_37794);
nor U42887 (N_42887,N_39545,N_35042);
and U42888 (N_42888,N_35540,N_38659);
nand U42889 (N_42889,N_36825,N_35232);
and U42890 (N_42890,N_38870,N_39234);
or U42891 (N_42891,N_36639,N_35932);
or U42892 (N_42892,N_39222,N_35560);
nor U42893 (N_42893,N_35776,N_35470);
or U42894 (N_42894,N_36170,N_39462);
xor U42895 (N_42895,N_35546,N_35017);
nand U42896 (N_42896,N_38199,N_38331);
nand U42897 (N_42897,N_35081,N_36339);
nor U42898 (N_42898,N_36627,N_36393);
nor U42899 (N_42899,N_37841,N_37302);
nand U42900 (N_42900,N_36818,N_38068);
and U42901 (N_42901,N_37259,N_35870);
and U42902 (N_42902,N_37125,N_35792);
nor U42903 (N_42903,N_35102,N_37170);
nor U42904 (N_42904,N_36593,N_35858);
nor U42905 (N_42905,N_38748,N_36865);
or U42906 (N_42906,N_36667,N_35170);
and U42907 (N_42907,N_39706,N_39359);
xor U42908 (N_42908,N_37406,N_38896);
and U42909 (N_42909,N_36921,N_38051);
nor U42910 (N_42910,N_35778,N_35069);
or U42911 (N_42911,N_38453,N_36611);
or U42912 (N_42912,N_38465,N_39021);
and U42913 (N_42913,N_37054,N_35669);
and U42914 (N_42914,N_39524,N_35773);
nor U42915 (N_42915,N_38109,N_37837);
and U42916 (N_42916,N_39816,N_35583);
nand U42917 (N_42917,N_37517,N_39089);
xnor U42918 (N_42918,N_37009,N_37012);
nor U42919 (N_42919,N_35965,N_36427);
nor U42920 (N_42920,N_35307,N_36820);
or U42921 (N_42921,N_39475,N_37037);
nand U42922 (N_42922,N_35533,N_35176);
nand U42923 (N_42923,N_36452,N_35607);
nor U42924 (N_42924,N_39874,N_37133);
xnor U42925 (N_42925,N_36104,N_37727);
nor U42926 (N_42926,N_36956,N_38121);
xnor U42927 (N_42927,N_38051,N_37433);
nor U42928 (N_42928,N_37034,N_39043);
and U42929 (N_42929,N_38214,N_38896);
or U42930 (N_42930,N_35098,N_35746);
or U42931 (N_42931,N_36880,N_36248);
nor U42932 (N_42932,N_35849,N_36090);
and U42933 (N_42933,N_37381,N_38232);
nand U42934 (N_42934,N_38969,N_35773);
nor U42935 (N_42935,N_39444,N_37068);
or U42936 (N_42936,N_38997,N_37442);
or U42937 (N_42937,N_36397,N_37257);
and U42938 (N_42938,N_35231,N_37238);
and U42939 (N_42939,N_39045,N_37563);
nor U42940 (N_42940,N_36724,N_38011);
or U42941 (N_42941,N_37444,N_36932);
nand U42942 (N_42942,N_39814,N_37535);
nand U42943 (N_42943,N_38197,N_36720);
and U42944 (N_42944,N_38392,N_37995);
and U42945 (N_42945,N_38367,N_38569);
or U42946 (N_42946,N_37526,N_39386);
and U42947 (N_42947,N_39387,N_39137);
xor U42948 (N_42948,N_38137,N_39678);
nor U42949 (N_42949,N_35717,N_37768);
xnor U42950 (N_42950,N_36781,N_38862);
nand U42951 (N_42951,N_36848,N_38944);
and U42952 (N_42952,N_38411,N_35811);
nand U42953 (N_42953,N_38957,N_37354);
nor U42954 (N_42954,N_39851,N_39408);
and U42955 (N_42955,N_38488,N_35150);
and U42956 (N_42956,N_38467,N_37148);
or U42957 (N_42957,N_39724,N_36894);
and U42958 (N_42958,N_38417,N_39040);
and U42959 (N_42959,N_36298,N_35290);
or U42960 (N_42960,N_37630,N_39987);
nand U42961 (N_42961,N_38175,N_35384);
nor U42962 (N_42962,N_37192,N_36003);
xnor U42963 (N_42963,N_35071,N_35542);
xnor U42964 (N_42964,N_39386,N_38187);
and U42965 (N_42965,N_39283,N_38603);
or U42966 (N_42966,N_35355,N_35762);
and U42967 (N_42967,N_35800,N_37189);
or U42968 (N_42968,N_37091,N_37378);
nand U42969 (N_42969,N_38355,N_38493);
and U42970 (N_42970,N_38545,N_39391);
and U42971 (N_42971,N_35994,N_35798);
and U42972 (N_42972,N_35594,N_37407);
nor U42973 (N_42973,N_37521,N_35062);
nor U42974 (N_42974,N_36878,N_35574);
and U42975 (N_42975,N_37960,N_35043);
xor U42976 (N_42976,N_35426,N_38639);
nor U42977 (N_42977,N_36761,N_38320);
or U42978 (N_42978,N_35469,N_37859);
or U42979 (N_42979,N_38231,N_36052);
or U42980 (N_42980,N_39589,N_37880);
and U42981 (N_42981,N_36091,N_38210);
nand U42982 (N_42982,N_35143,N_35083);
nand U42983 (N_42983,N_38440,N_36045);
xnor U42984 (N_42984,N_37043,N_38052);
nand U42985 (N_42985,N_37937,N_35961);
nor U42986 (N_42986,N_38098,N_37710);
and U42987 (N_42987,N_39032,N_35899);
or U42988 (N_42988,N_36076,N_39065);
nor U42989 (N_42989,N_36742,N_38890);
nor U42990 (N_42990,N_39992,N_39919);
xor U42991 (N_42991,N_38371,N_36938);
nand U42992 (N_42992,N_37580,N_38696);
or U42993 (N_42993,N_38347,N_38219);
or U42994 (N_42994,N_39337,N_39822);
and U42995 (N_42995,N_37190,N_39923);
xor U42996 (N_42996,N_38438,N_38007);
and U42997 (N_42997,N_36905,N_38809);
nor U42998 (N_42998,N_36167,N_35536);
xor U42999 (N_42999,N_35734,N_37118);
or U43000 (N_43000,N_39025,N_37107);
or U43001 (N_43001,N_38930,N_36940);
nor U43002 (N_43002,N_39828,N_36269);
xor U43003 (N_43003,N_35977,N_39167);
and U43004 (N_43004,N_38564,N_39693);
and U43005 (N_43005,N_39940,N_36422);
xnor U43006 (N_43006,N_37025,N_39248);
nand U43007 (N_43007,N_39680,N_37573);
nand U43008 (N_43008,N_36217,N_37125);
nand U43009 (N_43009,N_37869,N_35942);
or U43010 (N_43010,N_37706,N_39186);
or U43011 (N_43011,N_36865,N_37007);
nor U43012 (N_43012,N_38258,N_37264);
or U43013 (N_43013,N_38546,N_36806);
nand U43014 (N_43014,N_39180,N_39703);
and U43015 (N_43015,N_38887,N_35081);
and U43016 (N_43016,N_36732,N_35789);
nand U43017 (N_43017,N_35130,N_39458);
or U43018 (N_43018,N_37531,N_36799);
nor U43019 (N_43019,N_39770,N_39691);
and U43020 (N_43020,N_38708,N_35156);
or U43021 (N_43021,N_35077,N_38579);
or U43022 (N_43022,N_39778,N_38271);
nand U43023 (N_43023,N_39272,N_37319);
nor U43024 (N_43024,N_36653,N_35971);
and U43025 (N_43025,N_36947,N_38362);
nor U43026 (N_43026,N_39059,N_35674);
nor U43027 (N_43027,N_35248,N_35011);
and U43028 (N_43028,N_35971,N_36058);
xnor U43029 (N_43029,N_37742,N_39536);
or U43030 (N_43030,N_39111,N_38857);
or U43031 (N_43031,N_39669,N_39076);
nand U43032 (N_43032,N_38071,N_35046);
and U43033 (N_43033,N_38385,N_37164);
xor U43034 (N_43034,N_36799,N_35772);
or U43035 (N_43035,N_36968,N_35329);
or U43036 (N_43036,N_37406,N_35902);
nor U43037 (N_43037,N_36907,N_38143);
nor U43038 (N_43038,N_35583,N_36352);
nor U43039 (N_43039,N_35416,N_35630);
or U43040 (N_43040,N_39708,N_37947);
nor U43041 (N_43041,N_38593,N_37403);
or U43042 (N_43042,N_36222,N_35631);
nand U43043 (N_43043,N_35817,N_39045);
nand U43044 (N_43044,N_36581,N_35865);
and U43045 (N_43045,N_36151,N_39491);
nor U43046 (N_43046,N_36118,N_35282);
or U43047 (N_43047,N_39069,N_37494);
or U43048 (N_43048,N_36454,N_38744);
nand U43049 (N_43049,N_35517,N_36393);
nor U43050 (N_43050,N_35493,N_38452);
nand U43051 (N_43051,N_37846,N_37352);
or U43052 (N_43052,N_39858,N_36475);
nand U43053 (N_43053,N_39314,N_36314);
nand U43054 (N_43054,N_39072,N_37201);
nor U43055 (N_43055,N_36077,N_35119);
nor U43056 (N_43056,N_36058,N_37841);
nor U43057 (N_43057,N_38868,N_38702);
nand U43058 (N_43058,N_38946,N_36890);
and U43059 (N_43059,N_35870,N_38077);
nor U43060 (N_43060,N_35524,N_37782);
nand U43061 (N_43061,N_36208,N_35816);
nand U43062 (N_43062,N_38200,N_35134);
and U43063 (N_43063,N_35375,N_38887);
or U43064 (N_43064,N_38675,N_38730);
xnor U43065 (N_43065,N_37702,N_38700);
or U43066 (N_43066,N_38855,N_37578);
xnor U43067 (N_43067,N_38011,N_36763);
nor U43068 (N_43068,N_38227,N_39274);
nand U43069 (N_43069,N_38991,N_35895);
nand U43070 (N_43070,N_37804,N_37952);
or U43071 (N_43071,N_35136,N_36946);
or U43072 (N_43072,N_37874,N_38344);
or U43073 (N_43073,N_39836,N_37631);
nand U43074 (N_43074,N_39784,N_38912);
nor U43075 (N_43075,N_38429,N_38836);
and U43076 (N_43076,N_39911,N_36191);
and U43077 (N_43077,N_36128,N_38931);
nand U43078 (N_43078,N_36259,N_38213);
nand U43079 (N_43079,N_38744,N_38838);
or U43080 (N_43080,N_38305,N_38941);
and U43081 (N_43081,N_39593,N_36428);
nand U43082 (N_43082,N_35409,N_39371);
and U43083 (N_43083,N_37821,N_38302);
nand U43084 (N_43084,N_37379,N_39763);
and U43085 (N_43085,N_35163,N_36654);
and U43086 (N_43086,N_38853,N_39830);
nor U43087 (N_43087,N_35023,N_35634);
nor U43088 (N_43088,N_39068,N_37991);
nor U43089 (N_43089,N_35920,N_37134);
nor U43090 (N_43090,N_37345,N_37424);
or U43091 (N_43091,N_36260,N_38798);
nand U43092 (N_43092,N_39069,N_37159);
and U43093 (N_43093,N_37081,N_36090);
and U43094 (N_43094,N_37390,N_37293);
nand U43095 (N_43095,N_37171,N_35109);
nand U43096 (N_43096,N_36463,N_36645);
nor U43097 (N_43097,N_39800,N_35247);
nand U43098 (N_43098,N_38604,N_37089);
xor U43099 (N_43099,N_39506,N_37282);
or U43100 (N_43100,N_39281,N_36821);
nand U43101 (N_43101,N_36459,N_36754);
xnor U43102 (N_43102,N_39317,N_38958);
and U43103 (N_43103,N_37580,N_38257);
or U43104 (N_43104,N_39727,N_36995);
and U43105 (N_43105,N_37018,N_36589);
or U43106 (N_43106,N_37442,N_37411);
or U43107 (N_43107,N_35073,N_39819);
nor U43108 (N_43108,N_36101,N_35892);
and U43109 (N_43109,N_38724,N_37951);
and U43110 (N_43110,N_35319,N_35945);
and U43111 (N_43111,N_39191,N_36902);
or U43112 (N_43112,N_35219,N_37561);
and U43113 (N_43113,N_38553,N_36325);
xnor U43114 (N_43114,N_38486,N_35988);
nor U43115 (N_43115,N_37578,N_37240);
nand U43116 (N_43116,N_39043,N_37770);
and U43117 (N_43117,N_35634,N_37993);
nand U43118 (N_43118,N_39738,N_38113);
and U43119 (N_43119,N_37196,N_39587);
nand U43120 (N_43120,N_37440,N_36880);
xnor U43121 (N_43121,N_38342,N_36567);
nor U43122 (N_43122,N_39579,N_35533);
nor U43123 (N_43123,N_35629,N_35114);
nor U43124 (N_43124,N_38429,N_37217);
xnor U43125 (N_43125,N_37725,N_37925);
and U43126 (N_43126,N_37190,N_37249);
nor U43127 (N_43127,N_36004,N_39320);
or U43128 (N_43128,N_35373,N_36640);
nand U43129 (N_43129,N_35191,N_37189);
or U43130 (N_43130,N_35885,N_38415);
or U43131 (N_43131,N_36004,N_35099);
and U43132 (N_43132,N_35897,N_39951);
nand U43133 (N_43133,N_39911,N_39302);
nor U43134 (N_43134,N_36200,N_38812);
or U43135 (N_43135,N_39992,N_38778);
nand U43136 (N_43136,N_37652,N_35953);
nor U43137 (N_43137,N_39015,N_38301);
nand U43138 (N_43138,N_37216,N_37762);
nand U43139 (N_43139,N_38718,N_39622);
and U43140 (N_43140,N_36488,N_36721);
nor U43141 (N_43141,N_38988,N_35179);
xnor U43142 (N_43142,N_36262,N_39933);
nor U43143 (N_43143,N_35386,N_35696);
or U43144 (N_43144,N_38411,N_35044);
and U43145 (N_43145,N_39935,N_38622);
and U43146 (N_43146,N_36996,N_36836);
and U43147 (N_43147,N_35865,N_37845);
nor U43148 (N_43148,N_37206,N_36088);
or U43149 (N_43149,N_37158,N_35421);
nor U43150 (N_43150,N_37127,N_35982);
and U43151 (N_43151,N_37295,N_39450);
nor U43152 (N_43152,N_35552,N_38780);
or U43153 (N_43153,N_38099,N_39475);
or U43154 (N_43154,N_39724,N_36501);
and U43155 (N_43155,N_35715,N_36051);
nand U43156 (N_43156,N_35811,N_35709);
xnor U43157 (N_43157,N_35992,N_35419);
and U43158 (N_43158,N_37642,N_39586);
xor U43159 (N_43159,N_35872,N_39342);
nand U43160 (N_43160,N_39081,N_37590);
and U43161 (N_43161,N_39499,N_36067);
or U43162 (N_43162,N_36710,N_39364);
or U43163 (N_43163,N_39910,N_38972);
and U43164 (N_43164,N_39522,N_37220);
nand U43165 (N_43165,N_39116,N_37484);
nor U43166 (N_43166,N_36668,N_35758);
nor U43167 (N_43167,N_35540,N_38066);
nand U43168 (N_43168,N_38239,N_35477);
xor U43169 (N_43169,N_37116,N_39260);
nor U43170 (N_43170,N_35228,N_37332);
and U43171 (N_43171,N_37713,N_36489);
nor U43172 (N_43172,N_37275,N_39831);
and U43173 (N_43173,N_35051,N_37786);
nor U43174 (N_43174,N_39849,N_39111);
nand U43175 (N_43175,N_39715,N_39256);
xor U43176 (N_43176,N_37534,N_37350);
or U43177 (N_43177,N_39152,N_38064);
and U43178 (N_43178,N_35521,N_37765);
nor U43179 (N_43179,N_35735,N_35339);
or U43180 (N_43180,N_35057,N_38758);
or U43181 (N_43181,N_36841,N_38878);
and U43182 (N_43182,N_38338,N_37180);
nand U43183 (N_43183,N_39897,N_38960);
nor U43184 (N_43184,N_39159,N_36656);
or U43185 (N_43185,N_35178,N_36059);
xnor U43186 (N_43186,N_37824,N_37817);
xnor U43187 (N_43187,N_39472,N_35531);
or U43188 (N_43188,N_38811,N_37202);
or U43189 (N_43189,N_39585,N_36719);
nand U43190 (N_43190,N_35572,N_39872);
and U43191 (N_43191,N_37842,N_37111);
xor U43192 (N_43192,N_38794,N_37283);
nor U43193 (N_43193,N_36995,N_37026);
nand U43194 (N_43194,N_39877,N_35705);
or U43195 (N_43195,N_38067,N_37978);
and U43196 (N_43196,N_38349,N_37017);
nand U43197 (N_43197,N_35834,N_37911);
nand U43198 (N_43198,N_38966,N_35917);
nor U43199 (N_43199,N_39910,N_38668);
or U43200 (N_43200,N_39593,N_38212);
or U43201 (N_43201,N_38968,N_38257);
nand U43202 (N_43202,N_35077,N_35340);
or U43203 (N_43203,N_37418,N_35991);
xor U43204 (N_43204,N_39541,N_37761);
or U43205 (N_43205,N_38371,N_39747);
and U43206 (N_43206,N_37088,N_35175);
nand U43207 (N_43207,N_37636,N_36893);
nor U43208 (N_43208,N_38768,N_37171);
nor U43209 (N_43209,N_35267,N_37249);
nand U43210 (N_43210,N_36244,N_37745);
nand U43211 (N_43211,N_38303,N_37778);
nor U43212 (N_43212,N_39688,N_39632);
and U43213 (N_43213,N_37905,N_38658);
nor U43214 (N_43214,N_37298,N_39340);
nor U43215 (N_43215,N_36802,N_37353);
or U43216 (N_43216,N_35047,N_38125);
and U43217 (N_43217,N_37922,N_37616);
nor U43218 (N_43218,N_39395,N_37197);
nor U43219 (N_43219,N_39148,N_36871);
and U43220 (N_43220,N_38537,N_36520);
nor U43221 (N_43221,N_35284,N_35954);
or U43222 (N_43222,N_38388,N_36083);
or U43223 (N_43223,N_35839,N_37135);
and U43224 (N_43224,N_35196,N_38709);
nand U43225 (N_43225,N_39554,N_36867);
nor U43226 (N_43226,N_39314,N_35890);
and U43227 (N_43227,N_39261,N_36785);
or U43228 (N_43228,N_36196,N_39898);
or U43229 (N_43229,N_39840,N_39936);
and U43230 (N_43230,N_39391,N_36759);
nor U43231 (N_43231,N_39348,N_39579);
nand U43232 (N_43232,N_35961,N_36114);
nand U43233 (N_43233,N_37547,N_39919);
nand U43234 (N_43234,N_35053,N_36540);
or U43235 (N_43235,N_39112,N_38381);
nand U43236 (N_43236,N_38244,N_38891);
nor U43237 (N_43237,N_37509,N_38222);
nand U43238 (N_43238,N_36866,N_39754);
nor U43239 (N_43239,N_35058,N_36581);
or U43240 (N_43240,N_36850,N_38021);
or U43241 (N_43241,N_35261,N_35231);
nor U43242 (N_43242,N_37995,N_36132);
xor U43243 (N_43243,N_37455,N_38758);
nand U43244 (N_43244,N_37872,N_38059);
nand U43245 (N_43245,N_35417,N_38484);
xor U43246 (N_43246,N_37779,N_38973);
and U43247 (N_43247,N_35124,N_37827);
or U43248 (N_43248,N_39354,N_37049);
and U43249 (N_43249,N_36572,N_39121);
or U43250 (N_43250,N_38839,N_38250);
and U43251 (N_43251,N_38517,N_38604);
nor U43252 (N_43252,N_35278,N_36222);
or U43253 (N_43253,N_36577,N_38103);
nor U43254 (N_43254,N_36982,N_37646);
nor U43255 (N_43255,N_35660,N_38696);
nor U43256 (N_43256,N_38164,N_36419);
and U43257 (N_43257,N_39791,N_35848);
and U43258 (N_43258,N_37803,N_39561);
nand U43259 (N_43259,N_36250,N_37460);
xor U43260 (N_43260,N_36956,N_39519);
or U43261 (N_43261,N_35506,N_38294);
nor U43262 (N_43262,N_36802,N_35776);
nand U43263 (N_43263,N_38430,N_39424);
and U43264 (N_43264,N_35147,N_37315);
nor U43265 (N_43265,N_36580,N_38775);
or U43266 (N_43266,N_37117,N_38822);
and U43267 (N_43267,N_36042,N_35500);
or U43268 (N_43268,N_37230,N_38403);
nand U43269 (N_43269,N_36081,N_35611);
nand U43270 (N_43270,N_38786,N_39434);
nand U43271 (N_43271,N_38717,N_39667);
or U43272 (N_43272,N_38270,N_39886);
and U43273 (N_43273,N_35356,N_38612);
nand U43274 (N_43274,N_38674,N_39146);
or U43275 (N_43275,N_35838,N_39169);
or U43276 (N_43276,N_38834,N_35440);
nand U43277 (N_43277,N_35203,N_39257);
nand U43278 (N_43278,N_38672,N_38109);
nor U43279 (N_43279,N_36416,N_36681);
and U43280 (N_43280,N_37918,N_37431);
nor U43281 (N_43281,N_39452,N_39126);
or U43282 (N_43282,N_38621,N_37666);
nor U43283 (N_43283,N_38127,N_37367);
and U43284 (N_43284,N_38754,N_37418);
nor U43285 (N_43285,N_39976,N_35763);
nor U43286 (N_43286,N_35204,N_36170);
nand U43287 (N_43287,N_37974,N_39009);
nand U43288 (N_43288,N_35538,N_36602);
nand U43289 (N_43289,N_38995,N_39214);
and U43290 (N_43290,N_37462,N_39548);
and U43291 (N_43291,N_35179,N_38646);
or U43292 (N_43292,N_39736,N_37941);
nand U43293 (N_43293,N_38116,N_35429);
nand U43294 (N_43294,N_35403,N_35708);
or U43295 (N_43295,N_35512,N_36471);
and U43296 (N_43296,N_39193,N_36395);
xnor U43297 (N_43297,N_35265,N_35495);
or U43298 (N_43298,N_38332,N_38245);
nand U43299 (N_43299,N_38783,N_38359);
or U43300 (N_43300,N_38444,N_36145);
and U43301 (N_43301,N_38615,N_36521);
and U43302 (N_43302,N_38291,N_37669);
xor U43303 (N_43303,N_38204,N_35120);
nor U43304 (N_43304,N_39523,N_35933);
or U43305 (N_43305,N_39111,N_38777);
and U43306 (N_43306,N_38936,N_36035);
and U43307 (N_43307,N_37405,N_36792);
nor U43308 (N_43308,N_37946,N_38698);
nand U43309 (N_43309,N_35021,N_35870);
and U43310 (N_43310,N_38400,N_38286);
and U43311 (N_43311,N_38923,N_36963);
nor U43312 (N_43312,N_37731,N_39088);
or U43313 (N_43313,N_38681,N_39934);
and U43314 (N_43314,N_39253,N_37519);
and U43315 (N_43315,N_39173,N_38630);
nand U43316 (N_43316,N_38671,N_37776);
nand U43317 (N_43317,N_36481,N_38552);
or U43318 (N_43318,N_36482,N_39777);
xnor U43319 (N_43319,N_38834,N_37438);
nor U43320 (N_43320,N_38923,N_35695);
xnor U43321 (N_43321,N_38780,N_35484);
or U43322 (N_43322,N_36214,N_35124);
nor U43323 (N_43323,N_37793,N_37991);
nor U43324 (N_43324,N_37181,N_37961);
and U43325 (N_43325,N_35261,N_35612);
nand U43326 (N_43326,N_36783,N_36607);
nand U43327 (N_43327,N_37541,N_35563);
nor U43328 (N_43328,N_38806,N_39937);
nand U43329 (N_43329,N_36263,N_36210);
or U43330 (N_43330,N_36699,N_36523);
and U43331 (N_43331,N_38892,N_36005);
or U43332 (N_43332,N_35872,N_36710);
and U43333 (N_43333,N_36487,N_39913);
xnor U43334 (N_43334,N_35729,N_38699);
or U43335 (N_43335,N_37451,N_35287);
nor U43336 (N_43336,N_36018,N_37623);
or U43337 (N_43337,N_35467,N_38817);
or U43338 (N_43338,N_35124,N_39372);
nand U43339 (N_43339,N_35852,N_38542);
and U43340 (N_43340,N_38871,N_38833);
or U43341 (N_43341,N_38915,N_37783);
or U43342 (N_43342,N_38774,N_36672);
nor U43343 (N_43343,N_36213,N_37078);
or U43344 (N_43344,N_36670,N_39867);
or U43345 (N_43345,N_35103,N_35775);
or U43346 (N_43346,N_38165,N_35694);
or U43347 (N_43347,N_36045,N_38364);
or U43348 (N_43348,N_36532,N_37250);
nand U43349 (N_43349,N_38063,N_37002);
nor U43350 (N_43350,N_37177,N_38809);
and U43351 (N_43351,N_38553,N_36007);
or U43352 (N_43352,N_35540,N_39305);
or U43353 (N_43353,N_39062,N_35533);
or U43354 (N_43354,N_37311,N_36905);
nand U43355 (N_43355,N_36961,N_38814);
or U43356 (N_43356,N_37240,N_35525);
xor U43357 (N_43357,N_38857,N_35851);
nor U43358 (N_43358,N_36721,N_37820);
xnor U43359 (N_43359,N_38362,N_35154);
or U43360 (N_43360,N_39875,N_37551);
nor U43361 (N_43361,N_38031,N_36402);
nor U43362 (N_43362,N_37526,N_39111);
nor U43363 (N_43363,N_38570,N_35845);
nor U43364 (N_43364,N_35182,N_35138);
or U43365 (N_43365,N_39458,N_36109);
nand U43366 (N_43366,N_36428,N_36624);
and U43367 (N_43367,N_39880,N_39177);
nand U43368 (N_43368,N_39551,N_38148);
and U43369 (N_43369,N_38292,N_36616);
or U43370 (N_43370,N_36474,N_39829);
nand U43371 (N_43371,N_36070,N_38370);
nor U43372 (N_43372,N_37338,N_39183);
nor U43373 (N_43373,N_38834,N_39740);
nand U43374 (N_43374,N_38277,N_36517);
nor U43375 (N_43375,N_39078,N_38481);
and U43376 (N_43376,N_39309,N_38229);
nor U43377 (N_43377,N_38864,N_37386);
nand U43378 (N_43378,N_39202,N_38482);
nand U43379 (N_43379,N_35761,N_37049);
or U43380 (N_43380,N_36967,N_36435);
or U43381 (N_43381,N_38421,N_38207);
nand U43382 (N_43382,N_35894,N_36631);
nand U43383 (N_43383,N_35210,N_35815);
and U43384 (N_43384,N_35326,N_37968);
nand U43385 (N_43385,N_36849,N_38840);
nor U43386 (N_43386,N_37212,N_39651);
nand U43387 (N_43387,N_39168,N_37828);
or U43388 (N_43388,N_36112,N_38129);
nand U43389 (N_43389,N_36804,N_36612);
and U43390 (N_43390,N_39098,N_35515);
or U43391 (N_43391,N_37308,N_36277);
xor U43392 (N_43392,N_39878,N_35743);
nor U43393 (N_43393,N_37407,N_39263);
or U43394 (N_43394,N_38958,N_38497);
nor U43395 (N_43395,N_35845,N_36769);
and U43396 (N_43396,N_36580,N_39778);
nand U43397 (N_43397,N_37222,N_37591);
and U43398 (N_43398,N_38764,N_38010);
or U43399 (N_43399,N_38112,N_38110);
nand U43400 (N_43400,N_39695,N_35659);
nor U43401 (N_43401,N_36694,N_39790);
or U43402 (N_43402,N_35276,N_39882);
nand U43403 (N_43403,N_35745,N_39793);
nor U43404 (N_43404,N_39274,N_38599);
and U43405 (N_43405,N_35470,N_37867);
or U43406 (N_43406,N_39535,N_37244);
or U43407 (N_43407,N_35695,N_39669);
xnor U43408 (N_43408,N_37237,N_35256);
and U43409 (N_43409,N_36478,N_38562);
xor U43410 (N_43410,N_38423,N_39186);
and U43411 (N_43411,N_36454,N_39501);
xnor U43412 (N_43412,N_36192,N_38118);
nand U43413 (N_43413,N_36695,N_35289);
and U43414 (N_43414,N_38804,N_37568);
or U43415 (N_43415,N_38843,N_36636);
nand U43416 (N_43416,N_37659,N_35525);
or U43417 (N_43417,N_38925,N_35880);
and U43418 (N_43418,N_39013,N_38699);
and U43419 (N_43419,N_39478,N_39793);
and U43420 (N_43420,N_35131,N_36929);
nand U43421 (N_43421,N_37525,N_35954);
nand U43422 (N_43422,N_38672,N_39122);
nor U43423 (N_43423,N_38137,N_39301);
or U43424 (N_43424,N_37933,N_36246);
xor U43425 (N_43425,N_37912,N_36034);
or U43426 (N_43426,N_35501,N_38948);
or U43427 (N_43427,N_35364,N_36998);
and U43428 (N_43428,N_38130,N_39598);
xor U43429 (N_43429,N_38668,N_37496);
xor U43430 (N_43430,N_38042,N_38611);
nand U43431 (N_43431,N_38719,N_38376);
nor U43432 (N_43432,N_37000,N_36112);
xnor U43433 (N_43433,N_36567,N_35846);
or U43434 (N_43434,N_35252,N_39429);
xnor U43435 (N_43435,N_36177,N_36033);
or U43436 (N_43436,N_36830,N_38692);
or U43437 (N_43437,N_38566,N_39614);
xor U43438 (N_43438,N_36834,N_38382);
and U43439 (N_43439,N_38740,N_35562);
and U43440 (N_43440,N_39896,N_39096);
and U43441 (N_43441,N_37314,N_38011);
xor U43442 (N_43442,N_38961,N_39232);
and U43443 (N_43443,N_38424,N_38146);
nand U43444 (N_43444,N_37204,N_37788);
or U43445 (N_43445,N_38405,N_36482);
nor U43446 (N_43446,N_38666,N_37142);
xnor U43447 (N_43447,N_37882,N_39782);
nand U43448 (N_43448,N_38090,N_35610);
and U43449 (N_43449,N_38780,N_38606);
and U43450 (N_43450,N_35123,N_37157);
xor U43451 (N_43451,N_37998,N_38515);
xor U43452 (N_43452,N_35552,N_37119);
and U43453 (N_43453,N_37470,N_36039);
xnor U43454 (N_43454,N_38049,N_36651);
nor U43455 (N_43455,N_35797,N_37661);
and U43456 (N_43456,N_37275,N_35092);
xnor U43457 (N_43457,N_36420,N_38901);
and U43458 (N_43458,N_35551,N_36369);
nand U43459 (N_43459,N_35953,N_38145);
or U43460 (N_43460,N_36043,N_36811);
or U43461 (N_43461,N_37160,N_39856);
or U43462 (N_43462,N_36372,N_36179);
and U43463 (N_43463,N_37099,N_37231);
or U43464 (N_43464,N_39332,N_37050);
or U43465 (N_43465,N_36069,N_35722);
and U43466 (N_43466,N_35100,N_37483);
xnor U43467 (N_43467,N_39996,N_38892);
nand U43468 (N_43468,N_39871,N_38313);
and U43469 (N_43469,N_38505,N_36458);
or U43470 (N_43470,N_38605,N_37924);
or U43471 (N_43471,N_37322,N_35201);
or U43472 (N_43472,N_37148,N_38101);
or U43473 (N_43473,N_37547,N_39042);
and U43474 (N_43474,N_37920,N_36248);
and U43475 (N_43475,N_35424,N_39744);
nor U43476 (N_43476,N_37734,N_38546);
and U43477 (N_43477,N_35984,N_36299);
nor U43478 (N_43478,N_36789,N_37807);
and U43479 (N_43479,N_37757,N_39812);
or U43480 (N_43480,N_38822,N_37174);
or U43481 (N_43481,N_37022,N_37984);
xor U43482 (N_43482,N_36552,N_35441);
nor U43483 (N_43483,N_35974,N_36974);
or U43484 (N_43484,N_36634,N_38608);
nand U43485 (N_43485,N_38140,N_36273);
or U43486 (N_43486,N_38529,N_38457);
or U43487 (N_43487,N_39386,N_37677);
nor U43488 (N_43488,N_37996,N_37938);
and U43489 (N_43489,N_38922,N_36777);
and U43490 (N_43490,N_35314,N_38823);
and U43491 (N_43491,N_37173,N_35843);
nor U43492 (N_43492,N_36156,N_36404);
or U43493 (N_43493,N_39087,N_36907);
nand U43494 (N_43494,N_36829,N_39260);
or U43495 (N_43495,N_38783,N_37725);
nor U43496 (N_43496,N_39155,N_38858);
nor U43497 (N_43497,N_39618,N_39149);
or U43498 (N_43498,N_38038,N_36867);
and U43499 (N_43499,N_38918,N_36103);
or U43500 (N_43500,N_38297,N_38120);
nand U43501 (N_43501,N_36183,N_36844);
nor U43502 (N_43502,N_37059,N_38672);
nor U43503 (N_43503,N_37200,N_39111);
nor U43504 (N_43504,N_37223,N_37110);
nor U43505 (N_43505,N_36177,N_39943);
nor U43506 (N_43506,N_36905,N_39009);
or U43507 (N_43507,N_39703,N_35441);
and U43508 (N_43508,N_36670,N_35843);
nand U43509 (N_43509,N_35621,N_36722);
nand U43510 (N_43510,N_39467,N_39479);
nand U43511 (N_43511,N_36861,N_37490);
nor U43512 (N_43512,N_36275,N_38211);
or U43513 (N_43513,N_36518,N_38474);
xor U43514 (N_43514,N_35442,N_35142);
nor U43515 (N_43515,N_39216,N_38039);
or U43516 (N_43516,N_38774,N_37163);
and U43517 (N_43517,N_35482,N_38716);
and U43518 (N_43518,N_36341,N_38373);
or U43519 (N_43519,N_39310,N_37987);
and U43520 (N_43520,N_35978,N_39766);
xor U43521 (N_43521,N_39169,N_37323);
or U43522 (N_43522,N_38052,N_39769);
and U43523 (N_43523,N_38579,N_37448);
nor U43524 (N_43524,N_39589,N_38614);
xnor U43525 (N_43525,N_37142,N_35973);
nor U43526 (N_43526,N_35350,N_39270);
or U43527 (N_43527,N_39603,N_38032);
nor U43528 (N_43528,N_39346,N_38314);
nand U43529 (N_43529,N_35243,N_35307);
nand U43530 (N_43530,N_38857,N_38419);
and U43531 (N_43531,N_37298,N_35062);
nand U43532 (N_43532,N_36485,N_37838);
nor U43533 (N_43533,N_37313,N_36371);
or U43534 (N_43534,N_39401,N_38085);
and U43535 (N_43535,N_39952,N_36691);
nor U43536 (N_43536,N_38952,N_37044);
and U43537 (N_43537,N_36616,N_36676);
nor U43538 (N_43538,N_37008,N_35417);
nor U43539 (N_43539,N_36142,N_38040);
nor U43540 (N_43540,N_37607,N_37203);
nor U43541 (N_43541,N_38209,N_36235);
and U43542 (N_43542,N_39856,N_37455);
nor U43543 (N_43543,N_35187,N_35792);
nor U43544 (N_43544,N_36105,N_38740);
and U43545 (N_43545,N_38139,N_36524);
nor U43546 (N_43546,N_37254,N_35769);
xor U43547 (N_43547,N_37511,N_39306);
nor U43548 (N_43548,N_39010,N_39033);
and U43549 (N_43549,N_35847,N_35425);
xnor U43550 (N_43550,N_38637,N_36318);
or U43551 (N_43551,N_35882,N_38387);
or U43552 (N_43552,N_36668,N_36448);
nand U43553 (N_43553,N_37252,N_38929);
xnor U43554 (N_43554,N_37509,N_35797);
or U43555 (N_43555,N_37678,N_36459);
nand U43556 (N_43556,N_36722,N_37492);
or U43557 (N_43557,N_38753,N_36225);
or U43558 (N_43558,N_37572,N_38115);
nand U43559 (N_43559,N_36706,N_35816);
nand U43560 (N_43560,N_36403,N_38606);
and U43561 (N_43561,N_39551,N_35221);
xnor U43562 (N_43562,N_38516,N_38292);
xor U43563 (N_43563,N_38149,N_36470);
nor U43564 (N_43564,N_36384,N_37994);
and U43565 (N_43565,N_35419,N_35554);
nand U43566 (N_43566,N_35681,N_39319);
and U43567 (N_43567,N_37792,N_37950);
xor U43568 (N_43568,N_36914,N_35374);
nand U43569 (N_43569,N_38533,N_38349);
and U43570 (N_43570,N_36161,N_39395);
and U43571 (N_43571,N_35952,N_37850);
or U43572 (N_43572,N_36767,N_37415);
nor U43573 (N_43573,N_39968,N_38327);
nand U43574 (N_43574,N_38410,N_39904);
or U43575 (N_43575,N_39836,N_38193);
or U43576 (N_43576,N_38312,N_35545);
or U43577 (N_43577,N_37017,N_39138);
nand U43578 (N_43578,N_38405,N_39248);
nor U43579 (N_43579,N_36755,N_39528);
and U43580 (N_43580,N_36634,N_37705);
nand U43581 (N_43581,N_35701,N_35433);
nand U43582 (N_43582,N_39971,N_37875);
nand U43583 (N_43583,N_35859,N_39326);
xor U43584 (N_43584,N_37229,N_39180);
nor U43585 (N_43585,N_39463,N_35901);
or U43586 (N_43586,N_37654,N_38831);
and U43587 (N_43587,N_38937,N_37159);
and U43588 (N_43588,N_39159,N_39216);
nor U43589 (N_43589,N_37724,N_38582);
nand U43590 (N_43590,N_38355,N_39042);
and U43591 (N_43591,N_35989,N_39367);
nor U43592 (N_43592,N_39869,N_36222);
or U43593 (N_43593,N_38349,N_39970);
xnor U43594 (N_43594,N_36633,N_36645);
or U43595 (N_43595,N_37455,N_36440);
nand U43596 (N_43596,N_35356,N_38606);
xnor U43597 (N_43597,N_38304,N_38641);
and U43598 (N_43598,N_36539,N_37092);
nand U43599 (N_43599,N_36379,N_38951);
nand U43600 (N_43600,N_36343,N_35077);
nor U43601 (N_43601,N_39674,N_36043);
or U43602 (N_43602,N_35487,N_37324);
nor U43603 (N_43603,N_36966,N_38358);
and U43604 (N_43604,N_39405,N_36903);
nand U43605 (N_43605,N_35937,N_38112);
nor U43606 (N_43606,N_36999,N_35922);
xor U43607 (N_43607,N_37879,N_39995);
and U43608 (N_43608,N_38423,N_39883);
xnor U43609 (N_43609,N_39058,N_37398);
nor U43610 (N_43610,N_38942,N_37470);
nand U43611 (N_43611,N_38756,N_35300);
or U43612 (N_43612,N_36126,N_36901);
or U43613 (N_43613,N_39746,N_39098);
or U43614 (N_43614,N_38711,N_36351);
or U43615 (N_43615,N_36023,N_39048);
nor U43616 (N_43616,N_35313,N_38784);
nand U43617 (N_43617,N_38374,N_36342);
nor U43618 (N_43618,N_35117,N_35661);
nor U43619 (N_43619,N_39012,N_35490);
nand U43620 (N_43620,N_35073,N_35026);
and U43621 (N_43621,N_35713,N_39467);
and U43622 (N_43622,N_38768,N_38048);
nor U43623 (N_43623,N_39593,N_38215);
nor U43624 (N_43624,N_38866,N_39958);
nand U43625 (N_43625,N_36133,N_35275);
nand U43626 (N_43626,N_38887,N_37764);
and U43627 (N_43627,N_38965,N_36004);
xor U43628 (N_43628,N_37835,N_37405);
nor U43629 (N_43629,N_39229,N_37745);
or U43630 (N_43630,N_37736,N_37025);
nor U43631 (N_43631,N_37342,N_38529);
and U43632 (N_43632,N_35141,N_36978);
or U43633 (N_43633,N_37833,N_36244);
nand U43634 (N_43634,N_35310,N_39851);
and U43635 (N_43635,N_36181,N_36019);
and U43636 (N_43636,N_39086,N_37164);
or U43637 (N_43637,N_35321,N_35330);
nor U43638 (N_43638,N_37459,N_36348);
and U43639 (N_43639,N_39450,N_35234);
or U43640 (N_43640,N_37629,N_36614);
xor U43641 (N_43641,N_37264,N_39115);
nor U43642 (N_43642,N_38336,N_39732);
nor U43643 (N_43643,N_35419,N_37519);
nand U43644 (N_43644,N_35829,N_35554);
nand U43645 (N_43645,N_38277,N_39768);
nor U43646 (N_43646,N_35735,N_38386);
or U43647 (N_43647,N_38280,N_36307);
nand U43648 (N_43648,N_38772,N_35446);
and U43649 (N_43649,N_35159,N_38838);
nor U43650 (N_43650,N_39573,N_36278);
nor U43651 (N_43651,N_39080,N_37609);
xnor U43652 (N_43652,N_36447,N_39467);
nand U43653 (N_43653,N_37528,N_35645);
or U43654 (N_43654,N_38975,N_36574);
nand U43655 (N_43655,N_36024,N_38685);
and U43656 (N_43656,N_38684,N_37222);
xnor U43657 (N_43657,N_35595,N_36838);
and U43658 (N_43658,N_37021,N_38811);
xor U43659 (N_43659,N_37165,N_36250);
nand U43660 (N_43660,N_36661,N_38970);
or U43661 (N_43661,N_35458,N_38448);
nor U43662 (N_43662,N_37166,N_35437);
and U43663 (N_43663,N_37378,N_37092);
nand U43664 (N_43664,N_35886,N_37470);
nor U43665 (N_43665,N_38929,N_38898);
nand U43666 (N_43666,N_36063,N_35027);
or U43667 (N_43667,N_37433,N_36368);
and U43668 (N_43668,N_36389,N_35204);
and U43669 (N_43669,N_38911,N_36631);
or U43670 (N_43670,N_37205,N_35431);
or U43671 (N_43671,N_38009,N_38031);
nor U43672 (N_43672,N_39105,N_35537);
nor U43673 (N_43673,N_35253,N_38129);
and U43674 (N_43674,N_35764,N_37820);
nand U43675 (N_43675,N_39876,N_37822);
and U43676 (N_43676,N_36358,N_39425);
and U43677 (N_43677,N_37287,N_39086);
or U43678 (N_43678,N_37390,N_38983);
or U43679 (N_43679,N_37027,N_38617);
nand U43680 (N_43680,N_35744,N_38532);
nor U43681 (N_43681,N_35510,N_39407);
nor U43682 (N_43682,N_37382,N_37936);
nand U43683 (N_43683,N_38456,N_35913);
nor U43684 (N_43684,N_39581,N_37010);
nand U43685 (N_43685,N_38917,N_35030);
nand U43686 (N_43686,N_35828,N_37189);
xnor U43687 (N_43687,N_38100,N_39594);
nand U43688 (N_43688,N_37284,N_35735);
nor U43689 (N_43689,N_39563,N_38722);
and U43690 (N_43690,N_38425,N_38588);
nand U43691 (N_43691,N_36364,N_37456);
and U43692 (N_43692,N_35370,N_39934);
and U43693 (N_43693,N_36575,N_36157);
or U43694 (N_43694,N_38758,N_36373);
nand U43695 (N_43695,N_36593,N_38501);
and U43696 (N_43696,N_39033,N_37205);
nand U43697 (N_43697,N_38118,N_38864);
nor U43698 (N_43698,N_36858,N_39889);
nor U43699 (N_43699,N_35855,N_38212);
and U43700 (N_43700,N_35404,N_35000);
nand U43701 (N_43701,N_35246,N_39726);
or U43702 (N_43702,N_36269,N_39248);
nand U43703 (N_43703,N_36129,N_38072);
or U43704 (N_43704,N_38236,N_35307);
or U43705 (N_43705,N_35735,N_36261);
nand U43706 (N_43706,N_39605,N_36024);
or U43707 (N_43707,N_39635,N_39264);
nor U43708 (N_43708,N_38417,N_35818);
and U43709 (N_43709,N_35282,N_38967);
nand U43710 (N_43710,N_37410,N_39831);
xnor U43711 (N_43711,N_39619,N_37797);
nor U43712 (N_43712,N_37150,N_37227);
nor U43713 (N_43713,N_38758,N_39296);
nand U43714 (N_43714,N_36016,N_35672);
nor U43715 (N_43715,N_37034,N_38267);
xor U43716 (N_43716,N_36123,N_39768);
nor U43717 (N_43717,N_36507,N_39016);
nand U43718 (N_43718,N_37540,N_37715);
nor U43719 (N_43719,N_38638,N_37145);
or U43720 (N_43720,N_39225,N_39592);
nand U43721 (N_43721,N_37312,N_38762);
or U43722 (N_43722,N_37166,N_35445);
nor U43723 (N_43723,N_35548,N_38165);
or U43724 (N_43724,N_36697,N_36799);
nor U43725 (N_43725,N_39510,N_38331);
xor U43726 (N_43726,N_38163,N_37888);
or U43727 (N_43727,N_38924,N_35298);
nand U43728 (N_43728,N_38893,N_35514);
or U43729 (N_43729,N_36782,N_36229);
nor U43730 (N_43730,N_39947,N_35221);
nor U43731 (N_43731,N_35910,N_37184);
nand U43732 (N_43732,N_39897,N_36253);
and U43733 (N_43733,N_37980,N_39370);
or U43734 (N_43734,N_35162,N_39837);
and U43735 (N_43735,N_37767,N_35106);
or U43736 (N_43736,N_36896,N_38879);
and U43737 (N_43737,N_37012,N_38650);
xor U43738 (N_43738,N_39067,N_36787);
nand U43739 (N_43739,N_38321,N_38623);
and U43740 (N_43740,N_37600,N_37503);
and U43741 (N_43741,N_35999,N_38488);
nand U43742 (N_43742,N_38176,N_38275);
or U43743 (N_43743,N_36121,N_38682);
and U43744 (N_43744,N_38787,N_36754);
nor U43745 (N_43745,N_35798,N_38096);
nand U43746 (N_43746,N_39406,N_35185);
nor U43747 (N_43747,N_36550,N_35392);
or U43748 (N_43748,N_35502,N_35105);
nor U43749 (N_43749,N_36143,N_37051);
and U43750 (N_43750,N_37826,N_37776);
nand U43751 (N_43751,N_35284,N_36233);
or U43752 (N_43752,N_39819,N_35782);
nor U43753 (N_43753,N_35561,N_35304);
and U43754 (N_43754,N_36766,N_38628);
xor U43755 (N_43755,N_39655,N_36917);
nor U43756 (N_43756,N_35467,N_35833);
nand U43757 (N_43757,N_38212,N_38166);
nand U43758 (N_43758,N_36235,N_36632);
or U43759 (N_43759,N_38183,N_38331);
or U43760 (N_43760,N_37464,N_35101);
and U43761 (N_43761,N_39333,N_37270);
nor U43762 (N_43762,N_35916,N_36790);
and U43763 (N_43763,N_37265,N_39870);
or U43764 (N_43764,N_37167,N_35116);
and U43765 (N_43765,N_39094,N_35742);
nand U43766 (N_43766,N_39774,N_35098);
or U43767 (N_43767,N_38073,N_35948);
nand U43768 (N_43768,N_38220,N_37672);
and U43769 (N_43769,N_38454,N_39873);
nor U43770 (N_43770,N_36734,N_35598);
or U43771 (N_43771,N_36207,N_36201);
and U43772 (N_43772,N_39911,N_37107);
nor U43773 (N_43773,N_39888,N_38641);
or U43774 (N_43774,N_39155,N_38112);
or U43775 (N_43775,N_39214,N_35373);
and U43776 (N_43776,N_35555,N_35277);
xor U43777 (N_43777,N_36194,N_37107);
nor U43778 (N_43778,N_39182,N_35435);
and U43779 (N_43779,N_38503,N_35165);
nand U43780 (N_43780,N_35062,N_38384);
nor U43781 (N_43781,N_39910,N_37656);
nor U43782 (N_43782,N_39216,N_36173);
and U43783 (N_43783,N_37743,N_38473);
nand U43784 (N_43784,N_36807,N_39968);
and U43785 (N_43785,N_38976,N_39776);
and U43786 (N_43786,N_35459,N_39884);
nand U43787 (N_43787,N_35064,N_36581);
xnor U43788 (N_43788,N_37471,N_36728);
or U43789 (N_43789,N_36091,N_36451);
nand U43790 (N_43790,N_38123,N_37989);
and U43791 (N_43791,N_39485,N_37061);
nor U43792 (N_43792,N_35763,N_35860);
nor U43793 (N_43793,N_36362,N_35534);
nand U43794 (N_43794,N_38868,N_36783);
and U43795 (N_43795,N_37257,N_38099);
nand U43796 (N_43796,N_35415,N_35706);
or U43797 (N_43797,N_36207,N_36923);
nand U43798 (N_43798,N_37407,N_37003);
or U43799 (N_43799,N_38181,N_35074);
nand U43800 (N_43800,N_35434,N_35625);
nand U43801 (N_43801,N_37617,N_35335);
or U43802 (N_43802,N_37380,N_39601);
nand U43803 (N_43803,N_37958,N_39903);
nor U43804 (N_43804,N_35646,N_35876);
and U43805 (N_43805,N_37310,N_37201);
nor U43806 (N_43806,N_35990,N_37739);
or U43807 (N_43807,N_39697,N_37683);
nor U43808 (N_43808,N_35046,N_39020);
and U43809 (N_43809,N_36639,N_38293);
and U43810 (N_43810,N_35834,N_35176);
xnor U43811 (N_43811,N_38162,N_39512);
nand U43812 (N_43812,N_38272,N_35051);
or U43813 (N_43813,N_35586,N_37825);
or U43814 (N_43814,N_38442,N_37927);
or U43815 (N_43815,N_36438,N_37550);
nand U43816 (N_43816,N_36060,N_35825);
nand U43817 (N_43817,N_39757,N_36831);
and U43818 (N_43818,N_35891,N_39575);
or U43819 (N_43819,N_35855,N_36593);
nand U43820 (N_43820,N_35346,N_37523);
xnor U43821 (N_43821,N_38036,N_35121);
nand U43822 (N_43822,N_39534,N_38548);
nor U43823 (N_43823,N_37157,N_35543);
and U43824 (N_43824,N_36060,N_38686);
nor U43825 (N_43825,N_38660,N_38518);
xnor U43826 (N_43826,N_37125,N_37654);
and U43827 (N_43827,N_37611,N_35292);
or U43828 (N_43828,N_37780,N_39774);
and U43829 (N_43829,N_35770,N_39016);
and U43830 (N_43830,N_36245,N_36333);
or U43831 (N_43831,N_35263,N_37403);
nor U43832 (N_43832,N_37409,N_37506);
or U43833 (N_43833,N_35300,N_37561);
nand U43834 (N_43834,N_37836,N_38718);
nand U43835 (N_43835,N_38716,N_39160);
nand U43836 (N_43836,N_38718,N_37633);
xnor U43837 (N_43837,N_37084,N_38753);
and U43838 (N_43838,N_38101,N_39263);
or U43839 (N_43839,N_39143,N_35173);
nand U43840 (N_43840,N_36511,N_37429);
and U43841 (N_43841,N_37127,N_35316);
nand U43842 (N_43842,N_38422,N_35289);
nand U43843 (N_43843,N_38587,N_39229);
nand U43844 (N_43844,N_39037,N_35970);
nand U43845 (N_43845,N_35812,N_35909);
or U43846 (N_43846,N_35526,N_37684);
nand U43847 (N_43847,N_39421,N_39592);
or U43848 (N_43848,N_37292,N_39634);
and U43849 (N_43849,N_35104,N_36990);
xnor U43850 (N_43850,N_36450,N_37388);
and U43851 (N_43851,N_37562,N_36376);
and U43852 (N_43852,N_39517,N_36880);
nand U43853 (N_43853,N_35989,N_37083);
and U43854 (N_43854,N_37923,N_38673);
and U43855 (N_43855,N_35772,N_35288);
nand U43856 (N_43856,N_37351,N_36609);
or U43857 (N_43857,N_37923,N_38889);
and U43858 (N_43858,N_37948,N_39180);
and U43859 (N_43859,N_38773,N_38241);
nand U43860 (N_43860,N_36196,N_36432);
nor U43861 (N_43861,N_39627,N_39120);
xnor U43862 (N_43862,N_36702,N_36595);
nor U43863 (N_43863,N_39387,N_35188);
and U43864 (N_43864,N_36472,N_36642);
nor U43865 (N_43865,N_35426,N_39594);
xor U43866 (N_43866,N_36848,N_35566);
nand U43867 (N_43867,N_39221,N_37118);
nand U43868 (N_43868,N_36702,N_39582);
nand U43869 (N_43869,N_38799,N_39652);
xor U43870 (N_43870,N_36738,N_38911);
nand U43871 (N_43871,N_37883,N_39954);
or U43872 (N_43872,N_37924,N_35160);
and U43873 (N_43873,N_38234,N_39777);
nand U43874 (N_43874,N_36275,N_35710);
or U43875 (N_43875,N_38622,N_35237);
nand U43876 (N_43876,N_35479,N_38194);
xnor U43877 (N_43877,N_38929,N_39670);
or U43878 (N_43878,N_38062,N_37273);
and U43879 (N_43879,N_36643,N_35740);
and U43880 (N_43880,N_35667,N_36453);
or U43881 (N_43881,N_35731,N_37121);
and U43882 (N_43882,N_39361,N_36496);
nor U43883 (N_43883,N_39112,N_39327);
nand U43884 (N_43884,N_35987,N_38520);
and U43885 (N_43885,N_39380,N_35067);
nor U43886 (N_43886,N_35379,N_38303);
or U43887 (N_43887,N_38070,N_37431);
and U43888 (N_43888,N_35691,N_36790);
or U43889 (N_43889,N_39728,N_38867);
or U43890 (N_43890,N_36690,N_36288);
and U43891 (N_43891,N_35912,N_38912);
nor U43892 (N_43892,N_37910,N_36023);
nor U43893 (N_43893,N_36100,N_38617);
nor U43894 (N_43894,N_35331,N_38824);
nand U43895 (N_43895,N_37156,N_38747);
and U43896 (N_43896,N_36165,N_38087);
or U43897 (N_43897,N_37144,N_37220);
nand U43898 (N_43898,N_39870,N_36990);
and U43899 (N_43899,N_35754,N_37849);
nand U43900 (N_43900,N_35605,N_38674);
and U43901 (N_43901,N_39847,N_39676);
nor U43902 (N_43902,N_35189,N_36996);
and U43903 (N_43903,N_39246,N_35555);
nand U43904 (N_43904,N_37518,N_36103);
nor U43905 (N_43905,N_36776,N_37570);
and U43906 (N_43906,N_35889,N_38344);
and U43907 (N_43907,N_36919,N_36012);
or U43908 (N_43908,N_37937,N_35149);
and U43909 (N_43909,N_39924,N_39707);
nand U43910 (N_43910,N_39479,N_37805);
xor U43911 (N_43911,N_35213,N_37185);
nor U43912 (N_43912,N_37178,N_35031);
and U43913 (N_43913,N_38325,N_36165);
nor U43914 (N_43914,N_38699,N_38963);
xnor U43915 (N_43915,N_39167,N_36889);
and U43916 (N_43916,N_39338,N_37052);
or U43917 (N_43917,N_36671,N_38879);
and U43918 (N_43918,N_36646,N_39040);
xor U43919 (N_43919,N_37649,N_37257);
nor U43920 (N_43920,N_37623,N_36719);
xnor U43921 (N_43921,N_38371,N_38949);
or U43922 (N_43922,N_37203,N_35869);
and U43923 (N_43923,N_36843,N_37745);
nor U43924 (N_43924,N_37623,N_38020);
and U43925 (N_43925,N_37460,N_35328);
nand U43926 (N_43926,N_35619,N_39195);
or U43927 (N_43927,N_36631,N_36853);
nand U43928 (N_43928,N_35916,N_39758);
nand U43929 (N_43929,N_35811,N_37094);
xnor U43930 (N_43930,N_35400,N_38977);
xnor U43931 (N_43931,N_38373,N_35997);
nand U43932 (N_43932,N_38590,N_35853);
or U43933 (N_43933,N_39135,N_38957);
nand U43934 (N_43934,N_38078,N_38143);
and U43935 (N_43935,N_39583,N_36720);
or U43936 (N_43936,N_38663,N_37139);
nor U43937 (N_43937,N_36876,N_37204);
nor U43938 (N_43938,N_39602,N_38591);
and U43939 (N_43939,N_35353,N_39485);
nand U43940 (N_43940,N_37461,N_37956);
nor U43941 (N_43941,N_35318,N_37802);
nor U43942 (N_43942,N_35950,N_35006);
or U43943 (N_43943,N_39725,N_39740);
nor U43944 (N_43944,N_38754,N_38604);
nor U43945 (N_43945,N_35487,N_39247);
or U43946 (N_43946,N_36628,N_36257);
nor U43947 (N_43947,N_36469,N_35535);
or U43948 (N_43948,N_37409,N_35589);
or U43949 (N_43949,N_37922,N_35171);
nor U43950 (N_43950,N_37838,N_36185);
nand U43951 (N_43951,N_39082,N_38486);
nor U43952 (N_43952,N_36688,N_35382);
xor U43953 (N_43953,N_38037,N_38009);
nand U43954 (N_43954,N_39919,N_36879);
or U43955 (N_43955,N_37948,N_38671);
or U43956 (N_43956,N_39405,N_38330);
nand U43957 (N_43957,N_36214,N_36317);
xnor U43958 (N_43958,N_37585,N_38566);
or U43959 (N_43959,N_39813,N_35285);
nor U43960 (N_43960,N_39179,N_39351);
and U43961 (N_43961,N_39450,N_35030);
nand U43962 (N_43962,N_35503,N_35109);
and U43963 (N_43963,N_37393,N_39411);
or U43964 (N_43964,N_36294,N_35690);
or U43965 (N_43965,N_37327,N_38855);
or U43966 (N_43966,N_39872,N_38488);
and U43967 (N_43967,N_37086,N_38484);
nand U43968 (N_43968,N_39565,N_36720);
nand U43969 (N_43969,N_38536,N_39365);
nand U43970 (N_43970,N_38638,N_37977);
or U43971 (N_43971,N_39119,N_37205);
or U43972 (N_43972,N_38964,N_36982);
or U43973 (N_43973,N_38375,N_36597);
nand U43974 (N_43974,N_36024,N_36765);
and U43975 (N_43975,N_35778,N_39487);
or U43976 (N_43976,N_35285,N_38752);
and U43977 (N_43977,N_35052,N_35770);
nor U43978 (N_43978,N_39414,N_38340);
or U43979 (N_43979,N_37151,N_36525);
or U43980 (N_43980,N_39092,N_37855);
or U43981 (N_43981,N_37423,N_35829);
nor U43982 (N_43982,N_37985,N_35517);
or U43983 (N_43983,N_37491,N_38235);
and U43984 (N_43984,N_35381,N_39502);
and U43985 (N_43985,N_37302,N_38593);
or U43986 (N_43986,N_35210,N_37377);
xnor U43987 (N_43987,N_35636,N_38930);
nand U43988 (N_43988,N_36748,N_35388);
and U43989 (N_43989,N_36895,N_36109);
xor U43990 (N_43990,N_39625,N_36151);
xnor U43991 (N_43991,N_38352,N_39034);
nand U43992 (N_43992,N_36439,N_39084);
or U43993 (N_43993,N_38028,N_36636);
nand U43994 (N_43994,N_36571,N_38058);
nor U43995 (N_43995,N_35126,N_37941);
and U43996 (N_43996,N_36161,N_39429);
or U43997 (N_43997,N_35560,N_37155);
xor U43998 (N_43998,N_39027,N_36369);
and U43999 (N_43999,N_35780,N_35839);
or U44000 (N_44000,N_39303,N_36876);
nor U44001 (N_44001,N_37697,N_37410);
nor U44002 (N_44002,N_35599,N_37520);
nand U44003 (N_44003,N_35180,N_38547);
and U44004 (N_44004,N_38262,N_35241);
or U44005 (N_44005,N_36259,N_37135);
or U44006 (N_44006,N_39878,N_38311);
or U44007 (N_44007,N_35953,N_39418);
nor U44008 (N_44008,N_39447,N_36306);
nor U44009 (N_44009,N_37079,N_36165);
or U44010 (N_44010,N_37619,N_39640);
and U44011 (N_44011,N_36474,N_36944);
nand U44012 (N_44012,N_38840,N_38370);
or U44013 (N_44013,N_36631,N_36957);
and U44014 (N_44014,N_36389,N_37979);
nand U44015 (N_44015,N_39144,N_36029);
and U44016 (N_44016,N_35863,N_36173);
and U44017 (N_44017,N_37706,N_38294);
and U44018 (N_44018,N_36804,N_37349);
nor U44019 (N_44019,N_37833,N_36892);
or U44020 (N_44020,N_39685,N_39995);
nor U44021 (N_44021,N_38921,N_35851);
and U44022 (N_44022,N_37660,N_39470);
or U44023 (N_44023,N_35767,N_37476);
nor U44024 (N_44024,N_38883,N_39604);
and U44025 (N_44025,N_38840,N_39233);
and U44026 (N_44026,N_35358,N_35003);
and U44027 (N_44027,N_37501,N_36653);
nor U44028 (N_44028,N_36976,N_35363);
nand U44029 (N_44029,N_39310,N_38891);
nand U44030 (N_44030,N_37282,N_36394);
nor U44031 (N_44031,N_38271,N_38655);
or U44032 (N_44032,N_35466,N_39611);
nor U44033 (N_44033,N_38923,N_39225);
xor U44034 (N_44034,N_39105,N_37464);
xnor U44035 (N_44035,N_36486,N_37271);
nor U44036 (N_44036,N_38442,N_37337);
or U44037 (N_44037,N_37902,N_35924);
and U44038 (N_44038,N_35283,N_36754);
or U44039 (N_44039,N_38198,N_35039);
and U44040 (N_44040,N_35265,N_36206);
nand U44041 (N_44041,N_38976,N_39572);
xor U44042 (N_44042,N_39060,N_36639);
xor U44043 (N_44043,N_37216,N_35538);
and U44044 (N_44044,N_35918,N_37572);
or U44045 (N_44045,N_36893,N_36307);
xnor U44046 (N_44046,N_39720,N_36150);
or U44047 (N_44047,N_35896,N_37016);
nand U44048 (N_44048,N_37806,N_39373);
xnor U44049 (N_44049,N_39099,N_38597);
nor U44050 (N_44050,N_38659,N_37490);
nand U44051 (N_44051,N_39357,N_37642);
and U44052 (N_44052,N_38344,N_39128);
or U44053 (N_44053,N_38297,N_36460);
nor U44054 (N_44054,N_36423,N_35541);
nor U44055 (N_44055,N_37642,N_36822);
or U44056 (N_44056,N_36007,N_37949);
nor U44057 (N_44057,N_39830,N_38842);
nand U44058 (N_44058,N_37374,N_35317);
or U44059 (N_44059,N_39022,N_39075);
nand U44060 (N_44060,N_35800,N_38811);
nor U44061 (N_44061,N_38444,N_39714);
nor U44062 (N_44062,N_37159,N_38431);
xor U44063 (N_44063,N_35250,N_35721);
xor U44064 (N_44064,N_35975,N_35476);
and U44065 (N_44065,N_36321,N_35449);
nor U44066 (N_44066,N_38483,N_36331);
xnor U44067 (N_44067,N_36277,N_38555);
nor U44068 (N_44068,N_39760,N_38024);
and U44069 (N_44069,N_37435,N_37834);
or U44070 (N_44070,N_39401,N_35538);
or U44071 (N_44071,N_39055,N_36710);
and U44072 (N_44072,N_35988,N_39397);
or U44073 (N_44073,N_35978,N_35676);
and U44074 (N_44074,N_39039,N_37507);
nor U44075 (N_44075,N_37777,N_37966);
nor U44076 (N_44076,N_37119,N_39607);
nor U44077 (N_44077,N_39981,N_39182);
nor U44078 (N_44078,N_37228,N_39937);
nor U44079 (N_44079,N_36160,N_36865);
or U44080 (N_44080,N_36917,N_35011);
nor U44081 (N_44081,N_37372,N_37099);
or U44082 (N_44082,N_37464,N_35150);
and U44083 (N_44083,N_37882,N_35788);
nand U44084 (N_44084,N_35866,N_38789);
xor U44085 (N_44085,N_37405,N_38725);
nor U44086 (N_44086,N_36162,N_39914);
nor U44087 (N_44087,N_37918,N_35944);
and U44088 (N_44088,N_37249,N_38497);
or U44089 (N_44089,N_35400,N_39979);
or U44090 (N_44090,N_38228,N_39699);
and U44091 (N_44091,N_36576,N_39328);
nor U44092 (N_44092,N_37531,N_36303);
or U44093 (N_44093,N_36920,N_37059);
nor U44094 (N_44094,N_36391,N_36237);
or U44095 (N_44095,N_37871,N_39870);
and U44096 (N_44096,N_38188,N_35326);
nand U44097 (N_44097,N_39060,N_36287);
nor U44098 (N_44098,N_38552,N_35324);
and U44099 (N_44099,N_37623,N_38162);
nor U44100 (N_44100,N_37697,N_38826);
nand U44101 (N_44101,N_35001,N_39446);
xor U44102 (N_44102,N_38047,N_35329);
nand U44103 (N_44103,N_37781,N_35881);
and U44104 (N_44104,N_39128,N_37373);
or U44105 (N_44105,N_35320,N_38398);
or U44106 (N_44106,N_35150,N_36327);
nand U44107 (N_44107,N_37536,N_36030);
nand U44108 (N_44108,N_35191,N_38605);
nand U44109 (N_44109,N_38388,N_39169);
or U44110 (N_44110,N_39885,N_37280);
nor U44111 (N_44111,N_38525,N_37285);
xor U44112 (N_44112,N_35736,N_35510);
or U44113 (N_44113,N_36097,N_37222);
and U44114 (N_44114,N_37777,N_39383);
nand U44115 (N_44115,N_35125,N_35932);
nand U44116 (N_44116,N_38443,N_36794);
xor U44117 (N_44117,N_37990,N_39435);
or U44118 (N_44118,N_37629,N_39964);
or U44119 (N_44119,N_35149,N_38943);
nand U44120 (N_44120,N_36894,N_39527);
or U44121 (N_44121,N_37109,N_37546);
nor U44122 (N_44122,N_38265,N_37326);
nand U44123 (N_44123,N_37441,N_35454);
or U44124 (N_44124,N_39921,N_38387);
nor U44125 (N_44125,N_37959,N_35920);
nor U44126 (N_44126,N_39572,N_35355);
or U44127 (N_44127,N_37372,N_39963);
nand U44128 (N_44128,N_38679,N_38946);
or U44129 (N_44129,N_35231,N_36174);
nor U44130 (N_44130,N_37208,N_39419);
nand U44131 (N_44131,N_36873,N_39474);
or U44132 (N_44132,N_38770,N_37540);
nor U44133 (N_44133,N_39823,N_36866);
or U44134 (N_44134,N_37713,N_35304);
and U44135 (N_44135,N_39615,N_38925);
nor U44136 (N_44136,N_37292,N_37761);
and U44137 (N_44137,N_35123,N_35446);
nand U44138 (N_44138,N_35573,N_39412);
and U44139 (N_44139,N_39416,N_37976);
xnor U44140 (N_44140,N_37744,N_38149);
xor U44141 (N_44141,N_35904,N_39811);
or U44142 (N_44142,N_37322,N_38069);
or U44143 (N_44143,N_38892,N_35004);
or U44144 (N_44144,N_35952,N_35523);
nand U44145 (N_44145,N_35457,N_36984);
or U44146 (N_44146,N_39279,N_35391);
and U44147 (N_44147,N_36160,N_38457);
nand U44148 (N_44148,N_39285,N_35440);
nor U44149 (N_44149,N_37768,N_35570);
and U44150 (N_44150,N_39866,N_36383);
nor U44151 (N_44151,N_38391,N_38828);
xor U44152 (N_44152,N_35277,N_39728);
and U44153 (N_44153,N_36185,N_37358);
nand U44154 (N_44154,N_36301,N_35012);
and U44155 (N_44155,N_36096,N_36621);
nand U44156 (N_44156,N_37792,N_38534);
nand U44157 (N_44157,N_37113,N_38449);
nor U44158 (N_44158,N_38489,N_39271);
and U44159 (N_44159,N_37856,N_38585);
nand U44160 (N_44160,N_39709,N_36497);
xnor U44161 (N_44161,N_37428,N_35646);
nor U44162 (N_44162,N_38199,N_38016);
nand U44163 (N_44163,N_38701,N_37343);
nor U44164 (N_44164,N_39090,N_35201);
or U44165 (N_44165,N_36701,N_36272);
nor U44166 (N_44166,N_36398,N_38955);
nor U44167 (N_44167,N_39925,N_39030);
nor U44168 (N_44168,N_36346,N_37101);
nand U44169 (N_44169,N_39738,N_35387);
nand U44170 (N_44170,N_37641,N_35089);
and U44171 (N_44171,N_39954,N_37991);
nor U44172 (N_44172,N_39112,N_37350);
nor U44173 (N_44173,N_35972,N_36772);
and U44174 (N_44174,N_37889,N_36504);
nor U44175 (N_44175,N_36649,N_35507);
and U44176 (N_44176,N_37063,N_36303);
nor U44177 (N_44177,N_37474,N_39113);
and U44178 (N_44178,N_37809,N_35534);
nand U44179 (N_44179,N_35671,N_39836);
or U44180 (N_44180,N_36230,N_38184);
nand U44181 (N_44181,N_38199,N_35198);
and U44182 (N_44182,N_35474,N_36583);
xor U44183 (N_44183,N_35654,N_38266);
and U44184 (N_44184,N_37482,N_38175);
nor U44185 (N_44185,N_37189,N_36546);
and U44186 (N_44186,N_39705,N_36603);
or U44187 (N_44187,N_38367,N_38262);
nor U44188 (N_44188,N_38379,N_36581);
or U44189 (N_44189,N_36401,N_38968);
and U44190 (N_44190,N_39207,N_39695);
and U44191 (N_44191,N_38227,N_36762);
and U44192 (N_44192,N_35614,N_36545);
nor U44193 (N_44193,N_39206,N_39307);
or U44194 (N_44194,N_39569,N_39563);
or U44195 (N_44195,N_39641,N_37772);
or U44196 (N_44196,N_38549,N_38459);
xnor U44197 (N_44197,N_35709,N_38375);
nor U44198 (N_44198,N_36817,N_37418);
or U44199 (N_44199,N_38724,N_38367);
and U44200 (N_44200,N_35632,N_39543);
xnor U44201 (N_44201,N_37255,N_37620);
nand U44202 (N_44202,N_38694,N_38870);
nor U44203 (N_44203,N_36577,N_39912);
nor U44204 (N_44204,N_39807,N_35671);
or U44205 (N_44205,N_36288,N_37589);
nand U44206 (N_44206,N_39893,N_35262);
or U44207 (N_44207,N_38161,N_37666);
or U44208 (N_44208,N_35266,N_38334);
or U44209 (N_44209,N_38604,N_38627);
nand U44210 (N_44210,N_35474,N_39830);
nor U44211 (N_44211,N_38652,N_36413);
nor U44212 (N_44212,N_39867,N_39784);
or U44213 (N_44213,N_38861,N_35447);
and U44214 (N_44214,N_36467,N_39922);
nor U44215 (N_44215,N_39074,N_36917);
and U44216 (N_44216,N_39662,N_35662);
or U44217 (N_44217,N_37878,N_35677);
and U44218 (N_44218,N_38228,N_37246);
nand U44219 (N_44219,N_36171,N_36060);
and U44220 (N_44220,N_35863,N_37077);
nand U44221 (N_44221,N_38489,N_38800);
nand U44222 (N_44222,N_37897,N_37103);
or U44223 (N_44223,N_39995,N_38955);
nor U44224 (N_44224,N_39326,N_39810);
xnor U44225 (N_44225,N_38269,N_37117);
and U44226 (N_44226,N_36775,N_37123);
or U44227 (N_44227,N_37288,N_38422);
and U44228 (N_44228,N_37953,N_39829);
or U44229 (N_44229,N_36705,N_36506);
or U44230 (N_44230,N_35175,N_37175);
nor U44231 (N_44231,N_35666,N_39496);
and U44232 (N_44232,N_36525,N_38893);
or U44233 (N_44233,N_35745,N_37974);
nand U44234 (N_44234,N_38356,N_38544);
and U44235 (N_44235,N_37024,N_36052);
and U44236 (N_44236,N_37907,N_35980);
or U44237 (N_44237,N_38521,N_38135);
and U44238 (N_44238,N_36298,N_37546);
xor U44239 (N_44239,N_38155,N_37508);
nand U44240 (N_44240,N_39269,N_36606);
or U44241 (N_44241,N_37861,N_37509);
nand U44242 (N_44242,N_39658,N_36935);
nand U44243 (N_44243,N_38990,N_39850);
or U44244 (N_44244,N_38932,N_36492);
nor U44245 (N_44245,N_38215,N_38675);
or U44246 (N_44246,N_37436,N_39667);
nor U44247 (N_44247,N_39891,N_37244);
xnor U44248 (N_44248,N_36581,N_37113);
nand U44249 (N_44249,N_36626,N_38850);
and U44250 (N_44250,N_37060,N_37748);
nand U44251 (N_44251,N_38073,N_36679);
and U44252 (N_44252,N_35713,N_36816);
or U44253 (N_44253,N_35513,N_38025);
nor U44254 (N_44254,N_37820,N_37682);
or U44255 (N_44255,N_36117,N_35449);
nand U44256 (N_44256,N_39668,N_36352);
nand U44257 (N_44257,N_36348,N_37372);
and U44258 (N_44258,N_39506,N_38040);
xnor U44259 (N_44259,N_35267,N_38496);
nand U44260 (N_44260,N_39817,N_35464);
nand U44261 (N_44261,N_36884,N_35860);
and U44262 (N_44262,N_39016,N_35797);
or U44263 (N_44263,N_37379,N_39929);
nand U44264 (N_44264,N_37490,N_36579);
nand U44265 (N_44265,N_38773,N_38725);
nor U44266 (N_44266,N_39119,N_37984);
nor U44267 (N_44267,N_39630,N_38493);
or U44268 (N_44268,N_38402,N_36238);
or U44269 (N_44269,N_39391,N_36865);
nand U44270 (N_44270,N_38903,N_36795);
nand U44271 (N_44271,N_38477,N_38687);
nor U44272 (N_44272,N_38862,N_36400);
nor U44273 (N_44273,N_38869,N_37659);
and U44274 (N_44274,N_39135,N_38617);
nand U44275 (N_44275,N_37227,N_36799);
or U44276 (N_44276,N_36168,N_37828);
and U44277 (N_44277,N_37830,N_38326);
and U44278 (N_44278,N_39040,N_35447);
nor U44279 (N_44279,N_38309,N_37342);
and U44280 (N_44280,N_35581,N_36362);
nand U44281 (N_44281,N_39861,N_37601);
nand U44282 (N_44282,N_39664,N_36465);
or U44283 (N_44283,N_35863,N_36494);
nand U44284 (N_44284,N_38975,N_36286);
xnor U44285 (N_44285,N_39770,N_35148);
nand U44286 (N_44286,N_35673,N_37836);
and U44287 (N_44287,N_35890,N_39007);
nor U44288 (N_44288,N_37163,N_39488);
nand U44289 (N_44289,N_36352,N_36092);
nand U44290 (N_44290,N_38466,N_37736);
xor U44291 (N_44291,N_35573,N_35328);
xor U44292 (N_44292,N_36875,N_39082);
nor U44293 (N_44293,N_39936,N_35441);
and U44294 (N_44294,N_35521,N_38238);
and U44295 (N_44295,N_35209,N_39644);
and U44296 (N_44296,N_37551,N_37603);
and U44297 (N_44297,N_39528,N_39284);
and U44298 (N_44298,N_38193,N_35582);
and U44299 (N_44299,N_35042,N_39550);
nand U44300 (N_44300,N_37402,N_39879);
and U44301 (N_44301,N_35766,N_36299);
or U44302 (N_44302,N_39792,N_35788);
or U44303 (N_44303,N_39096,N_38577);
or U44304 (N_44304,N_36490,N_35135);
and U44305 (N_44305,N_37632,N_35937);
xor U44306 (N_44306,N_35419,N_36893);
nor U44307 (N_44307,N_36854,N_39446);
nor U44308 (N_44308,N_39281,N_39492);
nor U44309 (N_44309,N_35623,N_38888);
xor U44310 (N_44310,N_35448,N_35223);
or U44311 (N_44311,N_35919,N_38456);
nor U44312 (N_44312,N_37498,N_37935);
or U44313 (N_44313,N_36060,N_38334);
and U44314 (N_44314,N_38538,N_39055);
nand U44315 (N_44315,N_37642,N_39991);
nor U44316 (N_44316,N_37423,N_38541);
nand U44317 (N_44317,N_39431,N_35527);
nor U44318 (N_44318,N_36739,N_39960);
or U44319 (N_44319,N_39907,N_36976);
xor U44320 (N_44320,N_38701,N_35973);
and U44321 (N_44321,N_35645,N_37828);
or U44322 (N_44322,N_39873,N_39163);
or U44323 (N_44323,N_38536,N_35724);
and U44324 (N_44324,N_35010,N_35463);
or U44325 (N_44325,N_39591,N_35713);
nand U44326 (N_44326,N_38246,N_39558);
and U44327 (N_44327,N_38178,N_36643);
nor U44328 (N_44328,N_39482,N_36354);
nand U44329 (N_44329,N_37270,N_35357);
and U44330 (N_44330,N_39186,N_38438);
xnor U44331 (N_44331,N_38934,N_36201);
or U44332 (N_44332,N_37609,N_36139);
nand U44333 (N_44333,N_38631,N_36427);
and U44334 (N_44334,N_36268,N_39250);
nor U44335 (N_44335,N_36089,N_35299);
or U44336 (N_44336,N_35812,N_35714);
nand U44337 (N_44337,N_37336,N_35726);
nand U44338 (N_44338,N_36134,N_36387);
and U44339 (N_44339,N_35086,N_37702);
or U44340 (N_44340,N_38126,N_39580);
nand U44341 (N_44341,N_39436,N_36737);
nor U44342 (N_44342,N_35914,N_36271);
nand U44343 (N_44343,N_37970,N_35747);
and U44344 (N_44344,N_35922,N_37395);
and U44345 (N_44345,N_35935,N_39526);
nor U44346 (N_44346,N_36522,N_36751);
nand U44347 (N_44347,N_37245,N_36627);
nand U44348 (N_44348,N_39010,N_37665);
or U44349 (N_44349,N_36974,N_39895);
nor U44350 (N_44350,N_38741,N_35721);
or U44351 (N_44351,N_38750,N_35112);
xor U44352 (N_44352,N_37975,N_36361);
or U44353 (N_44353,N_36203,N_36449);
and U44354 (N_44354,N_37312,N_38177);
and U44355 (N_44355,N_36575,N_39096);
or U44356 (N_44356,N_37351,N_39530);
nand U44357 (N_44357,N_38637,N_36310);
nand U44358 (N_44358,N_36302,N_36033);
xor U44359 (N_44359,N_36904,N_38194);
nor U44360 (N_44360,N_39753,N_37901);
and U44361 (N_44361,N_37936,N_37994);
nand U44362 (N_44362,N_35897,N_35088);
and U44363 (N_44363,N_36260,N_39806);
xor U44364 (N_44364,N_38448,N_38627);
nor U44365 (N_44365,N_38270,N_35509);
and U44366 (N_44366,N_39046,N_39973);
nor U44367 (N_44367,N_35990,N_39382);
nand U44368 (N_44368,N_36495,N_36140);
nor U44369 (N_44369,N_39242,N_38343);
and U44370 (N_44370,N_36872,N_38857);
xor U44371 (N_44371,N_38798,N_36714);
or U44372 (N_44372,N_38273,N_39141);
nand U44373 (N_44373,N_37432,N_36196);
and U44374 (N_44374,N_35941,N_36433);
nor U44375 (N_44375,N_36527,N_37750);
xor U44376 (N_44376,N_39765,N_38829);
or U44377 (N_44377,N_37783,N_35137);
and U44378 (N_44378,N_38676,N_37168);
nand U44379 (N_44379,N_37759,N_37831);
nor U44380 (N_44380,N_38049,N_35650);
or U44381 (N_44381,N_35963,N_36994);
xnor U44382 (N_44382,N_38131,N_37897);
and U44383 (N_44383,N_35749,N_39471);
xnor U44384 (N_44384,N_39819,N_35414);
or U44385 (N_44385,N_35410,N_36740);
nand U44386 (N_44386,N_35038,N_37448);
or U44387 (N_44387,N_36593,N_37516);
and U44388 (N_44388,N_36041,N_37194);
and U44389 (N_44389,N_35379,N_38601);
nand U44390 (N_44390,N_36834,N_35830);
and U44391 (N_44391,N_39091,N_36798);
and U44392 (N_44392,N_38501,N_39160);
and U44393 (N_44393,N_36184,N_38009);
nand U44394 (N_44394,N_38855,N_35136);
or U44395 (N_44395,N_38489,N_37282);
nor U44396 (N_44396,N_38795,N_39903);
or U44397 (N_44397,N_38184,N_39036);
and U44398 (N_44398,N_36057,N_36718);
and U44399 (N_44399,N_35222,N_39060);
nand U44400 (N_44400,N_38475,N_39981);
nand U44401 (N_44401,N_38008,N_37475);
and U44402 (N_44402,N_38195,N_36836);
or U44403 (N_44403,N_37430,N_36601);
nand U44404 (N_44404,N_39532,N_38376);
nand U44405 (N_44405,N_37358,N_35295);
xnor U44406 (N_44406,N_37253,N_38066);
and U44407 (N_44407,N_36454,N_39365);
and U44408 (N_44408,N_36455,N_36353);
xor U44409 (N_44409,N_37204,N_36846);
or U44410 (N_44410,N_39751,N_35010);
and U44411 (N_44411,N_39607,N_39569);
or U44412 (N_44412,N_39862,N_38867);
or U44413 (N_44413,N_38120,N_38597);
and U44414 (N_44414,N_38774,N_38974);
nor U44415 (N_44415,N_38370,N_37467);
or U44416 (N_44416,N_35326,N_37971);
or U44417 (N_44417,N_35892,N_36275);
nand U44418 (N_44418,N_39970,N_39466);
nor U44419 (N_44419,N_38603,N_38633);
or U44420 (N_44420,N_38671,N_38022);
or U44421 (N_44421,N_39679,N_35540);
or U44422 (N_44422,N_37886,N_39882);
and U44423 (N_44423,N_36687,N_39847);
xor U44424 (N_44424,N_39369,N_38099);
and U44425 (N_44425,N_35120,N_38141);
nand U44426 (N_44426,N_35781,N_38968);
nor U44427 (N_44427,N_37737,N_39548);
nor U44428 (N_44428,N_38544,N_37657);
or U44429 (N_44429,N_39561,N_38661);
nor U44430 (N_44430,N_36597,N_39192);
nand U44431 (N_44431,N_39064,N_38303);
nand U44432 (N_44432,N_39344,N_37750);
nor U44433 (N_44433,N_35478,N_36056);
or U44434 (N_44434,N_38121,N_39445);
nor U44435 (N_44435,N_35739,N_39854);
nor U44436 (N_44436,N_39040,N_38748);
xor U44437 (N_44437,N_37322,N_35311);
and U44438 (N_44438,N_37807,N_37306);
nand U44439 (N_44439,N_38243,N_38570);
and U44440 (N_44440,N_38170,N_35820);
and U44441 (N_44441,N_38111,N_36254);
and U44442 (N_44442,N_38297,N_36850);
nand U44443 (N_44443,N_36746,N_37004);
nand U44444 (N_44444,N_35126,N_39068);
xor U44445 (N_44445,N_35904,N_37747);
nor U44446 (N_44446,N_36379,N_35917);
nand U44447 (N_44447,N_38469,N_37499);
or U44448 (N_44448,N_35556,N_39217);
nor U44449 (N_44449,N_36696,N_38978);
nor U44450 (N_44450,N_37503,N_37096);
nor U44451 (N_44451,N_37216,N_38305);
nor U44452 (N_44452,N_36935,N_39739);
nor U44453 (N_44453,N_36387,N_35775);
and U44454 (N_44454,N_36295,N_36988);
and U44455 (N_44455,N_38243,N_36209);
and U44456 (N_44456,N_39285,N_36289);
nand U44457 (N_44457,N_39654,N_35387);
nand U44458 (N_44458,N_35589,N_36163);
nor U44459 (N_44459,N_38059,N_38869);
or U44460 (N_44460,N_39560,N_39531);
nor U44461 (N_44461,N_37240,N_35926);
and U44462 (N_44462,N_37320,N_38880);
nor U44463 (N_44463,N_35208,N_38706);
and U44464 (N_44464,N_35340,N_35419);
nand U44465 (N_44465,N_35479,N_36730);
nor U44466 (N_44466,N_38085,N_36130);
or U44467 (N_44467,N_38365,N_36971);
nand U44468 (N_44468,N_35508,N_37567);
or U44469 (N_44469,N_36405,N_39545);
and U44470 (N_44470,N_37533,N_36253);
or U44471 (N_44471,N_39700,N_36204);
nor U44472 (N_44472,N_36211,N_35925);
or U44473 (N_44473,N_39785,N_37471);
or U44474 (N_44474,N_38098,N_39425);
nand U44475 (N_44475,N_37306,N_36414);
nor U44476 (N_44476,N_35981,N_35775);
nand U44477 (N_44477,N_36571,N_35135);
xnor U44478 (N_44478,N_36755,N_39838);
nand U44479 (N_44479,N_39707,N_36686);
nor U44480 (N_44480,N_36687,N_36466);
xor U44481 (N_44481,N_37182,N_36799);
or U44482 (N_44482,N_35244,N_37275);
or U44483 (N_44483,N_35211,N_38848);
nand U44484 (N_44484,N_39682,N_37456);
or U44485 (N_44485,N_39564,N_35116);
nor U44486 (N_44486,N_37779,N_35680);
nor U44487 (N_44487,N_37075,N_37507);
and U44488 (N_44488,N_37882,N_37326);
and U44489 (N_44489,N_38857,N_38058);
or U44490 (N_44490,N_39455,N_38351);
and U44491 (N_44491,N_38183,N_39656);
xor U44492 (N_44492,N_37123,N_36709);
or U44493 (N_44493,N_36768,N_36632);
xor U44494 (N_44494,N_35826,N_37229);
nor U44495 (N_44495,N_35175,N_36699);
nor U44496 (N_44496,N_38140,N_39175);
or U44497 (N_44497,N_37923,N_39547);
and U44498 (N_44498,N_35923,N_35523);
or U44499 (N_44499,N_35468,N_37823);
and U44500 (N_44500,N_39330,N_35453);
or U44501 (N_44501,N_37458,N_38658);
and U44502 (N_44502,N_35342,N_36070);
nor U44503 (N_44503,N_36787,N_36160);
and U44504 (N_44504,N_38561,N_35564);
xor U44505 (N_44505,N_39940,N_39653);
and U44506 (N_44506,N_36151,N_37047);
xnor U44507 (N_44507,N_38897,N_38342);
and U44508 (N_44508,N_37772,N_38891);
nand U44509 (N_44509,N_38492,N_35484);
nor U44510 (N_44510,N_39862,N_37758);
and U44511 (N_44511,N_38185,N_36898);
nand U44512 (N_44512,N_36213,N_36390);
or U44513 (N_44513,N_38515,N_38367);
or U44514 (N_44514,N_39635,N_37971);
and U44515 (N_44515,N_36182,N_36860);
and U44516 (N_44516,N_38899,N_37070);
and U44517 (N_44517,N_38211,N_35459);
nand U44518 (N_44518,N_35930,N_38209);
and U44519 (N_44519,N_38309,N_35460);
and U44520 (N_44520,N_38400,N_38867);
nand U44521 (N_44521,N_37874,N_39963);
nor U44522 (N_44522,N_39796,N_37339);
nand U44523 (N_44523,N_35026,N_35687);
or U44524 (N_44524,N_39755,N_38795);
xnor U44525 (N_44525,N_38336,N_36355);
nand U44526 (N_44526,N_38256,N_37686);
or U44527 (N_44527,N_38563,N_36799);
nor U44528 (N_44528,N_39776,N_37127);
nand U44529 (N_44529,N_36133,N_38619);
xnor U44530 (N_44530,N_38544,N_35587);
nand U44531 (N_44531,N_38635,N_36546);
and U44532 (N_44532,N_39172,N_35519);
and U44533 (N_44533,N_35011,N_36309);
and U44534 (N_44534,N_36435,N_36723);
nand U44535 (N_44535,N_35842,N_36244);
nor U44536 (N_44536,N_38754,N_35085);
or U44537 (N_44537,N_38720,N_35659);
nand U44538 (N_44538,N_36393,N_36147);
nand U44539 (N_44539,N_36016,N_36211);
or U44540 (N_44540,N_39336,N_39457);
nor U44541 (N_44541,N_38096,N_35016);
and U44542 (N_44542,N_37735,N_38366);
or U44543 (N_44543,N_36998,N_38939);
nor U44544 (N_44544,N_38109,N_36737);
and U44545 (N_44545,N_39946,N_37644);
or U44546 (N_44546,N_36698,N_36546);
and U44547 (N_44547,N_36019,N_38193);
nor U44548 (N_44548,N_35125,N_39621);
or U44549 (N_44549,N_36324,N_39037);
nand U44550 (N_44550,N_38432,N_35031);
nor U44551 (N_44551,N_37673,N_35902);
or U44552 (N_44552,N_35264,N_37235);
or U44553 (N_44553,N_37923,N_39880);
xnor U44554 (N_44554,N_38998,N_37643);
nor U44555 (N_44555,N_39704,N_39490);
nor U44556 (N_44556,N_37442,N_35201);
or U44557 (N_44557,N_38078,N_36341);
xor U44558 (N_44558,N_36658,N_36397);
nand U44559 (N_44559,N_37595,N_39342);
xor U44560 (N_44560,N_35821,N_35594);
nand U44561 (N_44561,N_39148,N_39507);
and U44562 (N_44562,N_35122,N_38229);
nand U44563 (N_44563,N_36685,N_35613);
and U44564 (N_44564,N_38100,N_36870);
nand U44565 (N_44565,N_39025,N_39425);
or U44566 (N_44566,N_36050,N_39967);
nor U44567 (N_44567,N_38598,N_35831);
nand U44568 (N_44568,N_37198,N_39926);
or U44569 (N_44569,N_39374,N_37985);
nor U44570 (N_44570,N_38109,N_39766);
or U44571 (N_44571,N_35647,N_37044);
and U44572 (N_44572,N_38443,N_35482);
and U44573 (N_44573,N_39306,N_38094);
and U44574 (N_44574,N_37414,N_37320);
or U44575 (N_44575,N_37961,N_37953);
xnor U44576 (N_44576,N_35255,N_39590);
or U44577 (N_44577,N_35127,N_36716);
nand U44578 (N_44578,N_35409,N_37626);
nor U44579 (N_44579,N_39833,N_35704);
nand U44580 (N_44580,N_36385,N_37316);
and U44581 (N_44581,N_36612,N_36996);
and U44582 (N_44582,N_39297,N_37917);
nand U44583 (N_44583,N_36302,N_37448);
nand U44584 (N_44584,N_35638,N_39249);
nand U44585 (N_44585,N_39272,N_39053);
or U44586 (N_44586,N_36527,N_37533);
nand U44587 (N_44587,N_37296,N_37000);
nor U44588 (N_44588,N_36105,N_36589);
and U44589 (N_44589,N_39889,N_36025);
xor U44590 (N_44590,N_35552,N_38135);
xnor U44591 (N_44591,N_37509,N_37561);
or U44592 (N_44592,N_38849,N_36916);
or U44593 (N_44593,N_39813,N_37958);
nand U44594 (N_44594,N_35695,N_39111);
nand U44595 (N_44595,N_35110,N_39626);
and U44596 (N_44596,N_38469,N_35116);
xor U44597 (N_44597,N_36441,N_35798);
nor U44598 (N_44598,N_36622,N_39670);
nand U44599 (N_44599,N_35136,N_37459);
nor U44600 (N_44600,N_38157,N_38281);
nor U44601 (N_44601,N_38234,N_38958);
or U44602 (N_44602,N_35961,N_36164);
or U44603 (N_44603,N_38269,N_36566);
or U44604 (N_44604,N_36557,N_38162);
or U44605 (N_44605,N_36800,N_37167);
or U44606 (N_44606,N_39009,N_38296);
or U44607 (N_44607,N_36762,N_36965);
nand U44608 (N_44608,N_36806,N_36177);
nor U44609 (N_44609,N_35432,N_39135);
nand U44610 (N_44610,N_39601,N_37556);
and U44611 (N_44611,N_36812,N_37566);
nor U44612 (N_44612,N_39067,N_36018);
nor U44613 (N_44613,N_35657,N_38942);
nand U44614 (N_44614,N_39517,N_38694);
or U44615 (N_44615,N_37660,N_36466);
nor U44616 (N_44616,N_35324,N_39578);
and U44617 (N_44617,N_39377,N_35351);
nand U44618 (N_44618,N_37157,N_38565);
xnor U44619 (N_44619,N_37150,N_36926);
nand U44620 (N_44620,N_36844,N_39909);
nor U44621 (N_44621,N_37550,N_39604);
or U44622 (N_44622,N_37081,N_38520);
or U44623 (N_44623,N_35674,N_36972);
xor U44624 (N_44624,N_38616,N_38515);
nand U44625 (N_44625,N_38559,N_38435);
nor U44626 (N_44626,N_39014,N_38331);
nor U44627 (N_44627,N_38045,N_36246);
and U44628 (N_44628,N_39432,N_38511);
or U44629 (N_44629,N_38608,N_39637);
nand U44630 (N_44630,N_39828,N_39657);
and U44631 (N_44631,N_38587,N_35812);
nand U44632 (N_44632,N_36223,N_38273);
nand U44633 (N_44633,N_38263,N_35708);
or U44634 (N_44634,N_36491,N_38047);
nand U44635 (N_44635,N_35157,N_36583);
nor U44636 (N_44636,N_36939,N_39855);
or U44637 (N_44637,N_35662,N_37685);
or U44638 (N_44638,N_35368,N_36602);
nor U44639 (N_44639,N_37976,N_39091);
nand U44640 (N_44640,N_38136,N_35933);
nor U44641 (N_44641,N_36681,N_39540);
nor U44642 (N_44642,N_38150,N_38100);
nor U44643 (N_44643,N_35784,N_36753);
xor U44644 (N_44644,N_39878,N_37047);
nor U44645 (N_44645,N_37671,N_35284);
nor U44646 (N_44646,N_37811,N_35514);
nand U44647 (N_44647,N_36074,N_38807);
nand U44648 (N_44648,N_35683,N_35037);
nor U44649 (N_44649,N_35985,N_39431);
and U44650 (N_44650,N_35811,N_36832);
and U44651 (N_44651,N_35066,N_38826);
or U44652 (N_44652,N_35231,N_35717);
nor U44653 (N_44653,N_37618,N_36712);
nand U44654 (N_44654,N_37299,N_39432);
xnor U44655 (N_44655,N_38121,N_36501);
or U44656 (N_44656,N_38684,N_39538);
nand U44657 (N_44657,N_39440,N_36646);
nor U44658 (N_44658,N_39177,N_35671);
nor U44659 (N_44659,N_35290,N_36961);
xor U44660 (N_44660,N_38368,N_35215);
nor U44661 (N_44661,N_39897,N_36898);
nand U44662 (N_44662,N_37099,N_36969);
xor U44663 (N_44663,N_37017,N_36984);
nor U44664 (N_44664,N_37446,N_38962);
nor U44665 (N_44665,N_36898,N_37851);
nor U44666 (N_44666,N_36834,N_39990);
nand U44667 (N_44667,N_36835,N_39079);
or U44668 (N_44668,N_37050,N_38594);
and U44669 (N_44669,N_37348,N_35691);
and U44670 (N_44670,N_37080,N_36502);
and U44671 (N_44671,N_35608,N_38789);
nor U44672 (N_44672,N_35722,N_36650);
or U44673 (N_44673,N_37455,N_36771);
or U44674 (N_44674,N_38107,N_37181);
or U44675 (N_44675,N_35916,N_37090);
and U44676 (N_44676,N_39035,N_35481);
and U44677 (N_44677,N_36861,N_39310);
and U44678 (N_44678,N_37465,N_36428);
or U44679 (N_44679,N_39924,N_38311);
nor U44680 (N_44680,N_39455,N_35963);
and U44681 (N_44681,N_37604,N_38053);
or U44682 (N_44682,N_38584,N_38320);
xnor U44683 (N_44683,N_38688,N_36947);
or U44684 (N_44684,N_36736,N_37081);
or U44685 (N_44685,N_37451,N_39868);
or U44686 (N_44686,N_38656,N_39459);
nand U44687 (N_44687,N_35340,N_37713);
and U44688 (N_44688,N_38701,N_35032);
xnor U44689 (N_44689,N_36317,N_37400);
nand U44690 (N_44690,N_37001,N_37912);
xor U44691 (N_44691,N_36285,N_38214);
nand U44692 (N_44692,N_39407,N_36394);
nand U44693 (N_44693,N_39400,N_39246);
nand U44694 (N_44694,N_37695,N_35877);
xnor U44695 (N_44695,N_35931,N_38902);
and U44696 (N_44696,N_36263,N_38271);
and U44697 (N_44697,N_36192,N_37033);
nand U44698 (N_44698,N_39598,N_35665);
nor U44699 (N_44699,N_35505,N_35484);
and U44700 (N_44700,N_38605,N_38564);
nor U44701 (N_44701,N_35131,N_35947);
and U44702 (N_44702,N_37169,N_39301);
and U44703 (N_44703,N_35297,N_35912);
nor U44704 (N_44704,N_36732,N_35874);
xnor U44705 (N_44705,N_36660,N_36571);
and U44706 (N_44706,N_38355,N_38567);
or U44707 (N_44707,N_36734,N_36113);
nand U44708 (N_44708,N_38371,N_37080);
and U44709 (N_44709,N_37914,N_38896);
nor U44710 (N_44710,N_38453,N_38959);
or U44711 (N_44711,N_38974,N_36845);
or U44712 (N_44712,N_39567,N_39791);
nand U44713 (N_44713,N_38748,N_37298);
nor U44714 (N_44714,N_35631,N_39220);
nor U44715 (N_44715,N_39427,N_36774);
and U44716 (N_44716,N_38828,N_38616);
and U44717 (N_44717,N_35966,N_39587);
nor U44718 (N_44718,N_39778,N_37485);
or U44719 (N_44719,N_36600,N_38219);
or U44720 (N_44720,N_36775,N_35448);
xor U44721 (N_44721,N_38111,N_39565);
nor U44722 (N_44722,N_38209,N_38926);
nand U44723 (N_44723,N_37465,N_35298);
nand U44724 (N_44724,N_38765,N_37874);
or U44725 (N_44725,N_37226,N_37780);
or U44726 (N_44726,N_37634,N_39467);
or U44727 (N_44727,N_38477,N_35275);
and U44728 (N_44728,N_38520,N_35931);
or U44729 (N_44729,N_39807,N_39637);
nand U44730 (N_44730,N_39367,N_37265);
or U44731 (N_44731,N_38004,N_37621);
and U44732 (N_44732,N_35517,N_35828);
or U44733 (N_44733,N_39969,N_36313);
nor U44734 (N_44734,N_37845,N_38361);
nand U44735 (N_44735,N_35634,N_37468);
nand U44736 (N_44736,N_36588,N_39387);
nand U44737 (N_44737,N_36250,N_36192);
nand U44738 (N_44738,N_38725,N_38324);
or U44739 (N_44739,N_37603,N_38398);
and U44740 (N_44740,N_35668,N_35697);
xor U44741 (N_44741,N_37994,N_37105);
xnor U44742 (N_44742,N_35020,N_36500);
and U44743 (N_44743,N_35789,N_38987);
and U44744 (N_44744,N_37728,N_39656);
xnor U44745 (N_44745,N_37201,N_37407);
or U44746 (N_44746,N_36519,N_36023);
and U44747 (N_44747,N_36765,N_39866);
nand U44748 (N_44748,N_39664,N_37491);
nand U44749 (N_44749,N_38224,N_36941);
or U44750 (N_44750,N_38520,N_37311);
or U44751 (N_44751,N_35641,N_39563);
or U44752 (N_44752,N_36316,N_38555);
or U44753 (N_44753,N_36714,N_38503);
nor U44754 (N_44754,N_37235,N_38842);
nand U44755 (N_44755,N_37098,N_37379);
xnor U44756 (N_44756,N_39566,N_36595);
xnor U44757 (N_44757,N_38488,N_38173);
nor U44758 (N_44758,N_38827,N_36631);
xor U44759 (N_44759,N_37827,N_37246);
xor U44760 (N_44760,N_39752,N_37453);
and U44761 (N_44761,N_36253,N_37302);
nor U44762 (N_44762,N_38347,N_36359);
and U44763 (N_44763,N_38776,N_35764);
and U44764 (N_44764,N_36799,N_39955);
nor U44765 (N_44765,N_35021,N_38187);
or U44766 (N_44766,N_38266,N_36290);
and U44767 (N_44767,N_39409,N_35453);
nand U44768 (N_44768,N_39204,N_36288);
nand U44769 (N_44769,N_38567,N_36189);
nand U44770 (N_44770,N_35269,N_36058);
nand U44771 (N_44771,N_38739,N_35013);
nor U44772 (N_44772,N_39840,N_35031);
nor U44773 (N_44773,N_35379,N_37862);
nor U44774 (N_44774,N_38141,N_35328);
nand U44775 (N_44775,N_39620,N_39794);
and U44776 (N_44776,N_39558,N_37029);
nor U44777 (N_44777,N_39759,N_38291);
and U44778 (N_44778,N_36726,N_38555);
or U44779 (N_44779,N_36440,N_35655);
nor U44780 (N_44780,N_38785,N_36407);
xor U44781 (N_44781,N_39717,N_39662);
xor U44782 (N_44782,N_38296,N_37540);
nand U44783 (N_44783,N_36974,N_39749);
nand U44784 (N_44784,N_38254,N_36038);
nor U44785 (N_44785,N_35137,N_38348);
nor U44786 (N_44786,N_37771,N_37887);
and U44787 (N_44787,N_38295,N_39929);
nor U44788 (N_44788,N_37546,N_38820);
or U44789 (N_44789,N_37122,N_38567);
and U44790 (N_44790,N_35017,N_39589);
nand U44791 (N_44791,N_35654,N_36420);
or U44792 (N_44792,N_37260,N_38485);
nand U44793 (N_44793,N_38358,N_35201);
nand U44794 (N_44794,N_36505,N_37872);
or U44795 (N_44795,N_38780,N_35986);
nand U44796 (N_44796,N_35500,N_35513);
and U44797 (N_44797,N_39676,N_37638);
nor U44798 (N_44798,N_36122,N_37208);
nand U44799 (N_44799,N_37321,N_35429);
nor U44800 (N_44800,N_39433,N_36159);
or U44801 (N_44801,N_35387,N_35551);
or U44802 (N_44802,N_39384,N_39488);
nor U44803 (N_44803,N_36203,N_36071);
nand U44804 (N_44804,N_37846,N_36743);
or U44805 (N_44805,N_35542,N_38301);
nor U44806 (N_44806,N_36588,N_35029);
nand U44807 (N_44807,N_38482,N_39648);
nand U44808 (N_44808,N_36698,N_39707);
xnor U44809 (N_44809,N_35574,N_36521);
or U44810 (N_44810,N_35313,N_36080);
nor U44811 (N_44811,N_38515,N_36873);
nand U44812 (N_44812,N_35941,N_38279);
nor U44813 (N_44813,N_38342,N_38454);
and U44814 (N_44814,N_39977,N_37732);
or U44815 (N_44815,N_38057,N_35560);
nor U44816 (N_44816,N_38344,N_38304);
and U44817 (N_44817,N_39406,N_39462);
or U44818 (N_44818,N_36263,N_36223);
and U44819 (N_44819,N_36897,N_35121);
and U44820 (N_44820,N_35152,N_36751);
nand U44821 (N_44821,N_35312,N_38988);
and U44822 (N_44822,N_37476,N_35534);
nand U44823 (N_44823,N_36468,N_35761);
nand U44824 (N_44824,N_37502,N_38749);
or U44825 (N_44825,N_39491,N_37932);
nand U44826 (N_44826,N_39159,N_37502);
nor U44827 (N_44827,N_37981,N_38581);
nand U44828 (N_44828,N_35865,N_36185);
or U44829 (N_44829,N_38217,N_35883);
and U44830 (N_44830,N_39564,N_38860);
and U44831 (N_44831,N_35269,N_39541);
nor U44832 (N_44832,N_39090,N_37387);
or U44833 (N_44833,N_39148,N_37927);
nor U44834 (N_44834,N_37397,N_37717);
nor U44835 (N_44835,N_39564,N_39293);
nor U44836 (N_44836,N_37843,N_37630);
and U44837 (N_44837,N_37262,N_37737);
nor U44838 (N_44838,N_35639,N_39842);
or U44839 (N_44839,N_38227,N_38911);
nor U44840 (N_44840,N_38700,N_35935);
nor U44841 (N_44841,N_38374,N_37477);
and U44842 (N_44842,N_37628,N_38972);
or U44843 (N_44843,N_36171,N_38697);
and U44844 (N_44844,N_39120,N_36613);
xnor U44845 (N_44845,N_39680,N_35754);
and U44846 (N_44846,N_35662,N_35400);
nand U44847 (N_44847,N_35877,N_38741);
nand U44848 (N_44848,N_39956,N_38467);
nor U44849 (N_44849,N_36922,N_37032);
and U44850 (N_44850,N_36598,N_35806);
nor U44851 (N_44851,N_38298,N_39525);
nor U44852 (N_44852,N_35540,N_38375);
nand U44853 (N_44853,N_35681,N_35560);
and U44854 (N_44854,N_39237,N_35618);
or U44855 (N_44855,N_38274,N_38806);
nand U44856 (N_44856,N_39143,N_35299);
or U44857 (N_44857,N_39556,N_38548);
nor U44858 (N_44858,N_39793,N_36557);
nor U44859 (N_44859,N_38455,N_36486);
xor U44860 (N_44860,N_37587,N_37953);
nor U44861 (N_44861,N_36185,N_35350);
and U44862 (N_44862,N_38461,N_36723);
nand U44863 (N_44863,N_37807,N_37493);
or U44864 (N_44864,N_38637,N_37901);
xnor U44865 (N_44865,N_36759,N_35560);
and U44866 (N_44866,N_37017,N_36014);
or U44867 (N_44867,N_37068,N_39351);
and U44868 (N_44868,N_36710,N_39985);
xnor U44869 (N_44869,N_39148,N_37263);
and U44870 (N_44870,N_37825,N_38500);
nand U44871 (N_44871,N_38206,N_38577);
and U44872 (N_44872,N_38712,N_37517);
nor U44873 (N_44873,N_37584,N_37773);
and U44874 (N_44874,N_38054,N_35556);
or U44875 (N_44875,N_35191,N_38534);
or U44876 (N_44876,N_35013,N_35419);
nor U44877 (N_44877,N_38594,N_39026);
xor U44878 (N_44878,N_39525,N_39012);
or U44879 (N_44879,N_39098,N_35023);
nand U44880 (N_44880,N_36978,N_35661);
nand U44881 (N_44881,N_38231,N_38020);
and U44882 (N_44882,N_38811,N_36664);
and U44883 (N_44883,N_38325,N_38255);
nor U44884 (N_44884,N_36414,N_38004);
and U44885 (N_44885,N_36822,N_37057);
nor U44886 (N_44886,N_35225,N_39220);
nor U44887 (N_44887,N_36877,N_39256);
or U44888 (N_44888,N_38302,N_37668);
nor U44889 (N_44889,N_37938,N_37476);
nand U44890 (N_44890,N_38339,N_39458);
nor U44891 (N_44891,N_38712,N_35796);
and U44892 (N_44892,N_38977,N_37139);
xor U44893 (N_44893,N_36884,N_39456);
nor U44894 (N_44894,N_35270,N_38311);
or U44895 (N_44895,N_39730,N_37652);
xnor U44896 (N_44896,N_36037,N_36143);
nor U44897 (N_44897,N_35401,N_38356);
or U44898 (N_44898,N_37665,N_37363);
xor U44899 (N_44899,N_36414,N_39143);
xor U44900 (N_44900,N_36893,N_39254);
nor U44901 (N_44901,N_37950,N_38239);
xnor U44902 (N_44902,N_38075,N_37710);
or U44903 (N_44903,N_35211,N_36850);
nand U44904 (N_44904,N_35383,N_38694);
nor U44905 (N_44905,N_39876,N_38407);
nand U44906 (N_44906,N_35335,N_38713);
and U44907 (N_44907,N_38884,N_38362);
and U44908 (N_44908,N_39373,N_37920);
or U44909 (N_44909,N_39202,N_35394);
nor U44910 (N_44910,N_37937,N_37691);
and U44911 (N_44911,N_35153,N_39341);
nor U44912 (N_44912,N_36236,N_39138);
or U44913 (N_44913,N_38713,N_38139);
xnor U44914 (N_44914,N_39650,N_38307);
and U44915 (N_44915,N_36669,N_37752);
nor U44916 (N_44916,N_39360,N_39266);
nor U44917 (N_44917,N_38218,N_38041);
nor U44918 (N_44918,N_36268,N_39791);
nand U44919 (N_44919,N_36171,N_39224);
nand U44920 (N_44920,N_37240,N_36373);
or U44921 (N_44921,N_39426,N_36469);
nor U44922 (N_44922,N_36724,N_39057);
or U44923 (N_44923,N_35013,N_38871);
and U44924 (N_44924,N_39272,N_38359);
nand U44925 (N_44925,N_37103,N_38894);
nand U44926 (N_44926,N_36058,N_37539);
and U44927 (N_44927,N_38772,N_37467);
and U44928 (N_44928,N_38135,N_35637);
nand U44929 (N_44929,N_36426,N_39506);
and U44930 (N_44930,N_36897,N_39839);
nand U44931 (N_44931,N_35878,N_36957);
and U44932 (N_44932,N_35860,N_35764);
nor U44933 (N_44933,N_37448,N_36342);
nand U44934 (N_44934,N_39315,N_39907);
and U44935 (N_44935,N_39177,N_35514);
nand U44936 (N_44936,N_37996,N_39293);
nand U44937 (N_44937,N_36092,N_35211);
nand U44938 (N_44938,N_35523,N_36718);
or U44939 (N_44939,N_39463,N_37583);
and U44940 (N_44940,N_36379,N_39569);
and U44941 (N_44941,N_39032,N_35875);
or U44942 (N_44942,N_35177,N_37786);
nor U44943 (N_44943,N_39365,N_39701);
and U44944 (N_44944,N_36545,N_39827);
nand U44945 (N_44945,N_35561,N_39164);
nor U44946 (N_44946,N_38828,N_36144);
nand U44947 (N_44947,N_37025,N_37173);
xor U44948 (N_44948,N_38526,N_38696);
nand U44949 (N_44949,N_37927,N_39245);
or U44950 (N_44950,N_38280,N_35417);
nand U44951 (N_44951,N_38996,N_35967);
and U44952 (N_44952,N_36312,N_38831);
nand U44953 (N_44953,N_36281,N_39704);
nand U44954 (N_44954,N_37105,N_36105);
nor U44955 (N_44955,N_37320,N_37399);
nand U44956 (N_44956,N_38665,N_38853);
and U44957 (N_44957,N_38939,N_36059);
nand U44958 (N_44958,N_35307,N_38913);
xor U44959 (N_44959,N_36331,N_35749);
or U44960 (N_44960,N_36533,N_35080);
and U44961 (N_44961,N_39797,N_36447);
and U44962 (N_44962,N_38390,N_37175);
or U44963 (N_44963,N_35964,N_36606);
or U44964 (N_44964,N_39859,N_39498);
nor U44965 (N_44965,N_39428,N_36786);
xor U44966 (N_44966,N_37725,N_38077);
or U44967 (N_44967,N_35028,N_37845);
or U44968 (N_44968,N_37450,N_36839);
nand U44969 (N_44969,N_35819,N_36084);
or U44970 (N_44970,N_37005,N_38704);
and U44971 (N_44971,N_38564,N_35809);
nor U44972 (N_44972,N_37591,N_37296);
and U44973 (N_44973,N_36612,N_36095);
and U44974 (N_44974,N_37111,N_35231);
or U44975 (N_44975,N_39995,N_35180);
and U44976 (N_44976,N_37327,N_38737);
or U44977 (N_44977,N_37306,N_38725);
and U44978 (N_44978,N_36352,N_36410);
nand U44979 (N_44979,N_35485,N_36979);
and U44980 (N_44980,N_36498,N_36171);
nand U44981 (N_44981,N_38979,N_36467);
nor U44982 (N_44982,N_39179,N_35947);
nand U44983 (N_44983,N_37653,N_36209);
or U44984 (N_44984,N_39428,N_38789);
nand U44985 (N_44985,N_39729,N_39008);
nor U44986 (N_44986,N_37497,N_39493);
nand U44987 (N_44987,N_35193,N_36400);
or U44988 (N_44988,N_37033,N_38739);
nand U44989 (N_44989,N_39925,N_37696);
and U44990 (N_44990,N_38076,N_35231);
nand U44991 (N_44991,N_38481,N_38560);
xor U44992 (N_44992,N_36935,N_37904);
nand U44993 (N_44993,N_39078,N_38782);
or U44994 (N_44994,N_36805,N_35246);
or U44995 (N_44995,N_37799,N_38188);
or U44996 (N_44996,N_37709,N_38333);
and U44997 (N_44997,N_35168,N_37079);
nand U44998 (N_44998,N_38173,N_39833);
nor U44999 (N_44999,N_38691,N_37248);
nor U45000 (N_45000,N_44827,N_43211);
xnor U45001 (N_45001,N_43187,N_42518);
nand U45002 (N_45002,N_41171,N_41928);
nand U45003 (N_45003,N_44514,N_44067);
nor U45004 (N_45004,N_40766,N_41333);
or U45005 (N_45005,N_43286,N_41687);
or U45006 (N_45006,N_41257,N_42679);
and U45007 (N_45007,N_42204,N_41430);
xnor U45008 (N_45008,N_42510,N_44500);
or U45009 (N_45009,N_44178,N_44021);
nand U45010 (N_45010,N_40265,N_40723);
nor U45011 (N_45011,N_42630,N_40196);
nand U45012 (N_45012,N_40975,N_41410);
nand U45013 (N_45013,N_41168,N_43388);
or U45014 (N_45014,N_42911,N_41470);
or U45015 (N_45015,N_43750,N_42372);
and U45016 (N_45016,N_42476,N_43993);
nand U45017 (N_45017,N_43987,N_41938);
nor U45018 (N_45018,N_41269,N_44431);
or U45019 (N_45019,N_43975,N_42821);
nor U45020 (N_45020,N_43949,N_41455);
nand U45021 (N_45021,N_41622,N_40985);
nand U45022 (N_45022,N_44149,N_40057);
nand U45023 (N_45023,N_41434,N_40078);
nand U45024 (N_45024,N_43650,N_41179);
xor U45025 (N_45025,N_40001,N_44267);
nor U45026 (N_45026,N_40771,N_41981);
or U45027 (N_45027,N_41767,N_40520);
nor U45028 (N_45028,N_41173,N_40402);
nor U45029 (N_45029,N_44823,N_41140);
nand U45030 (N_45030,N_43494,N_41943);
or U45031 (N_45031,N_41777,N_40714);
and U45032 (N_45032,N_41639,N_42616);
and U45033 (N_45033,N_43027,N_40745);
and U45034 (N_45034,N_41485,N_42723);
and U45035 (N_45035,N_42035,N_43629);
or U45036 (N_45036,N_44009,N_44175);
nor U45037 (N_45037,N_41307,N_40240);
nand U45038 (N_45038,N_42099,N_42438);
or U45039 (N_45039,N_42364,N_40931);
and U45040 (N_45040,N_43342,N_42375);
and U45041 (N_45041,N_41715,N_43872);
or U45042 (N_45042,N_42383,N_40822);
nor U45043 (N_45043,N_44226,N_43435);
nand U45044 (N_45044,N_43285,N_43991);
xnor U45045 (N_45045,N_42084,N_42161);
and U45046 (N_45046,N_40942,N_41313);
nor U45047 (N_45047,N_42374,N_44727);
or U45048 (N_45048,N_41817,N_43045);
or U45049 (N_45049,N_41690,N_40691);
and U45050 (N_45050,N_44883,N_42982);
and U45051 (N_45051,N_42142,N_42920);
or U45052 (N_45052,N_40472,N_42443);
or U45053 (N_45053,N_41632,N_42685);
xor U45054 (N_45054,N_43674,N_41247);
and U45055 (N_45055,N_44454,N_42018);
nand U45056 (N_45056,N_43707,N_41031);
nor U45057 (N_45057,N_43527,N_41296);
xor U45058 (N_45058,N_44954,N_41862);
and U45059 (N_45059,N_43429,N_41824);
xnor U45060 (N_45060,N_42690,N_42980);
nor U45061 (N_45061,N_41655,N_41080);
xnor U45062 (N_45062,N_42988,N_40484);
or U45063 (N_45063,N_43295,N_41922);
or U45064 (N_45064,N_44768,N_42219);
or U45065 (N_45065,N_42494,N_42245);
nor U45066 (N_45066,N_41633,N_42160);
and U45067 (N_45067,N_44370,N_41570);
or U45068 (N_45068,N_43393,N_42893);
nor U45069 (N_45069,N_40033,N_43697);
nor U45070 (N_45070,N_43015,N_40067);
or U45071 (N_45071,N_44425,N_43655);
nor U45072 (N_45072,N_42754,N_40406);
nor U45073 (N_45073,N_43310,N_40419);
and U45074 (N_45074,N_44412,N_41323);
and U45075 (N_45075,N_40467,N_42267);
or U45076 (N_45076,N_43766,N_41787);
nor U45077 (N_45077,N_41857,N_40654);
nor U45078 (N_45078,N_42446,N_43708);
and U45079 (N_45079,N_43825,N_40254);
or U45080 (N_45080,N_43758,N_41162);
or U45081 (N_45081,N_41999,N_41825);
nand U45082 (N_45082,N_42167,N_44193);
xor U45083 (N_45083,N_44885,N_44169);
nor U45084 (N_45084,N_41615,N_41350);
nor U45085 (N_45085,N_40518,N_43212);
and U45086 (N_45086,N_41801,N_41720);
or U45087 (N_45087,N_44239,N_43856);
or U45088 (N_45088,N_40389,N_40159);
and U45089 (N_45089,N_42212,N_43831);
nand U45090 (N_45090,N_40512,N_42156);
or U45091 (N_45091,N_41714,N_41889);
nor U45092 (N_45092,N_41382,N_40628);
and U45093 (N_45093,N_41088,N_44018);
and U45094 (N_45094,N_44000,N_41920);
or U45095 (N_45095,N_44757,N_41065);
and U45096 (N_45096,N_42395,N_41166);
nor U45097 (N_45097,N_42825,N_44654);
nor U45098 (N_45098,N_40317,N_43622);
or U45099 (N_45099,N_41009,N_43118);
nor U45100 (N_45100,N_41285,N_43029);
or U45101 (N_45101,N_42089,N_42638);
nor U45102 (N_45102,N_40347,N_44908);
xor U45103 (N_45103,N_42491,N_43086);
nor U45104 (N_45104,N_41699,N_42803);
and U45105 (N_45105,N_41103,N_44300);
xor U45106 (N_45106,N_40874,N_42950);
and U45107 (N_45107,N_42465,N_41631);
nor U45108 (N_45108,N_43104,N_41159);
or U45109 (N_45109,N_44905,N_43402);
nor U45110 (N_45110,N_40411,N_40436);
nand U45111 (N_45111,N_41594,N_43502);
nand U45112 (N_45112,N_44420,N_41120);
nand U45113 (N_45113,N_41646,N_44333);
nor U45114 (N_45114,N_40720,N_43324);
nand U45115 (N_45115,N_41160,N_42523);
nor U45116 (N_45116,N_43190,N_42329);
and U45117 (N_45117,N_42484,N_42016);
nor U45118 (N_45118,N_44111,N_42037);
nor U45119 (N_45119,N_43314,N_44468);
nand U45120 (N_45120,N_43837,N_43325);
xnor U45121 (N_45121,N_43103,N_43366);
or U45122 (N_45122,N_44247,N_42056);
xor U45123 (N_45123,N_44354,N_41258);
and U45124 (N_45124,N_44352,N_41271);
nand U45125 (N_45125,N_44646,N_41573);
nand U45126 (N_45126,N_40938,N_41867);
or U45127 (N_45127,N_42781,N_40585);
and U45128 (N_45128,N_42753,N_43522);
nor U45129 (N_45129,N_40552,N_41925);
and U45130 (N_45130,N_43963,N_41517);
nand U45131 (N_45131,N_42336,N_42737);
or U45132 (N_45132,N_40601,N_43060);
and U45133 (N_45133,N_43642,N_42771);
or U45134 (N_45134,N_43634,N_42568);
or U45135 (N_45135,N_44177,N_43935);
nor U45136 (N_45136,N_44291,N_43733);
nor U45137 (N_45137,N_44887,N_43048);
and U45138 (N_45138,N_43292,N_42758);
xnor U45139 (N_45139,N_40266,N_43003);
or U45140 (N_45140,N_42976,N_43115);
or U45141 (N_45141,N_43698,N_43312);
nand U45142 (N_45142,N_42924,N_44898);
and U45143 (N_45143,N_43052,N_40217);
nand U45144 (N_45144,N_43226,N_41195);
xnor U45145 (N_45145,N_44019,N_40912);
or U45146 (N_45146,N_40903,N_42796);
nand U45147 (N_45147,N_40430,N_42457);
and U45148 (N_45148,N_44804,N_41339);
nand U45149 (N_45149,N_44976,N_42619);
nand U45150 (N_45150,N_41374,N_41521);
nor U45151 (N_45151,N_42557,N_44166);
or U45152 (N_45152,N_41396,N_44563);
nor U45153 (N_45153,N_42431,N_41189);
nor U45154 (N_45154,N_41984,N_42229);
nor U45155 (N_45155,N_43653,N_43789);
nand U45156 (N_45156,N_44606,N_43946);
or U45157 (N_45157,N_44229,N_44880);
and U45158 (N_45158,N_42517,N_44477);
and U45159 (N_45159,N_43817,N_43423);
nand U45160 (N_45160,N_44575,N_42461);
or U45161 (N_45161,N_44790,N_42519);
or U45162 (N_45162,N_41023,N_43084);
or U45163 (N_45163,N_43014,N_40987);
nor U45164 (N_45164,N_41582,N_42162);
nand U45165 (N_45165,N_44373,N_44847);
nor U45166 (N_45166,N_42861,N_41520);
nor U45167 (N_45167,N_43857,N_43185);
or U45168 (N_45168,N_41194,N_40207);
xor U45169 (N_45169,N_44488,N_40275);
nor U45170 (N_45170,N_42936,N_44508);
or U45171 (N_45171,N_40988,N_41856);
or U45172 (N_45172,N_43112,N_42618);
nor U45173 (N_45173,N_44743,N_41605);
nand U45174 (N_45174,N_42563,N_42330);
and U45175 (N_45175,N_44548,N_42290);
nand U45176 (N_45176,N_42571,N_44952);
or U45177 (N_45177,N_43517,N_44396);
or U45178 (N_45178,N_40305,N_40877);
and U45179 (N_45179,N_40362,N_42884);
or U45180 (N_45180,N_40417,N_40244);
and U45181 (N_45181,N_41513,N_42392);
nor U45182 (N_45182,N_41022,N_40536);
or U45183 (N_45183,N_41991,N_42774);
nand U45184 (N_45184,N_43034,N_40343);
nand U45185 (N_45185,N_43876,N_44301);
or U45186 (N_45186,N_40110,N_40360);
and U45187 (N_45187,N_41565,N_40172);
or U45188 (N_45188,N_40570,N_42964);
or U45189 (N_45189,N_44970,N_41716);
or U45190 (N_45190,N_43180,N_43705);
xnor U45191 (N_45191,N_44613,N_43834);
nand U45192 (N_45192,N_40867,N_41309);
xnor U45193 (N_45193,N_40846,N_40712);
nand U45194 (N_45194,N_40726,N_44503);
or U45195 (N_45195,N_40651,N_41230);
and U45196 (N_45196,N_40621,N_42974);
or U45197 (N_45197,N_41443,N_41536);
or U45198 (N_45198,N_41730,N_40584);
and U45199 (N_45199,N_41458,N_41502);
nor U45200 (N_45200,N_41368,N_42076);
and U45201 (N_45201,N_41365,N_40048);
or U45202 (N_45202,N_42214,N_44299);
and U45203 (N_45203,N_42011,N_44002);
and U45204 (N_45204,N_42263,N_42904);
xor U45205 (N_45205,N_40466,N_41979);
nor U45206 (N_45206,N_40205,N_43657);
nor U45207 (N_45207,N_44571,N_42732);
xor U45208 (N_45208,N_40073,N_44384);
nor U45209 (N_45209,N_40624,N_41937);
or U45210 (N_45210,N_42108,N_43070);
or U45211 (N_45211,N_42462,N_44184);
nor U45212 (N_45212,N_43780,N_41432);
and U45213 (N_45213,N_41074,N_41318);
nor U45214 (N_45214,N_41182,N_44723);
or U45215 (N_45215,N_44716,N_41289);
or U45216 (N_45216,N_44484,N_40587);
or U45217 (N_45217,N_42255,N_44469);
nand U45218 (N_45218,N_42891,N_41606);
or U45219 (N_45219,N_40225,N_41026);
and U45220 (N_45220,N_42086,N_42576);
nand U45221 (N_45221,N_42617,N_44141);
or U45222 (N_45222,N_41127,N_40192);
or U45223 (N_45223,N_44697,N_43056);
nor U45224 (N_45224,N_42736,N_41426);
and U45225 (N_45225,N_41897,N_43142);
or U45226 (N_45226,N_44553,N_41776);
nor U45227 (N_45227,N_44416,N_44751);
xor U45228 (N_45228,N_42473,N_40077);
nor U45229 (N_45229,N_44492,N_42733);
nor U45230 (N_45230,N_40390,N_43967);
xnor U45231 (N_45231,N_40120,N_42648);
nor U45232 (N_45232,N_43159,N_42237);
nand U45233 (N_45233,N_40463,N_41148);
nor U45234 (N_45234,N_44940,N_43004);
and U45235 (N_45235,N_42444,N_41243);
or U45236 (N_45236,N_44538,N_40134);
xor U45237 (N_45237,N_43897,N_44619);
and U45238 (N_45238,N_41390,N_41757);
and U45239 (N_45239,N_42034,N_41163);
or U45240 (N_45240,N_41844,N_42371);
or U45241 (N_45241,N_43980,N_40502);
or U45242 (N_45242,N_42173,N_42368);
or U45243 (N_45243,N_41841,N_40645);
nand U45244 (N_45244,N_40247,N_42554);
xor U45245 (N_45245,N_44734,N_44137);
nor U45246 (N_45246,N_42399,N_42468);
nand U45247 (N_45247,N_42001,N_42283);
nor U45248 (N_45248,N_43166,N_44878);
nand U45249 (N_45249,N_42671,N_40424);
and U45250 (N_45250,N_43518,N_41329);
nand U45251 (N_45251,N_43297,N_41858);
and U45252 (N_45252,N_40925,N_42532);
or U45253 (N_45253,N_43461,N_43986);
nand U45254 (N_45254,N_42958,N_44817);
and U45255 (N_45255,N_42642,N_44984);
or U45256 (N_45256,N_43638,N_43952);
xnor U45257 (N_45257,N_43068,N_42062);
nand U45258 (N_45258,N_42661,N_40015);
or U45259 (N_45259,N_41553,N_43270);
nor U45260 (N_45260,N_43951,N_42508);
nor U45261 (N_45261,N_40667,N_41064);
and U45262 (N_45262,N_42117,N_41854);
and U45263 (N_45263,N_41185,N_41244);
or U45264 (N_45264,N_43382,N_42624);
nand U45265 (N_45265,N_41558,N_43762);
nand U45266 (N_45266,N_40747,N_41516);
and U45267 (N_45267,N_43055,N_43581);
or U45268 (N_45268,N_42268,N_40250);
xor U45269 (N_45269,N_44609,N_40410);
or U45270 (N_45270,N_42952,N_41071);
nor U45271 (N_45271,N_42983,N_42080);
nand U45272 (N_45272,N_40005,N_43201);
nand U45273 (N_45273,N_44608,N_41771);
nor U45274 (N_45274,N_42451,N_40230);
and U45275 (N_45275,N_42136,N_41707);
or U45276 (N_45276,N_40344,N_40191);
and U45277 (N_45277,N_42900,N_44741);
and U45278 (N_45278,N_41005,N_41081);
xnor U45279 (N_45279,N_44766,N_41672);
nand U45280 (N_45280,N_40736,N_40095);
nor U45281 (N_45281,N_40642,N_41649);
or U45282 (N_45282,N_42720,N_44787);
nand U45283 (N_45283,N_41828,N_44685);
or U45284 (N_45284,N_43782,N_42751);
nor U45285 (N_45285,N_44956,N_40280);
and U45286 (N_45286,N_44277,N_40346);
or U45287 (N_45287,N_44753,N_40050);
or U45288 (N_45288,N_44459,N_43454);
and U45289 (N_45289,N_44088,N_40282);
nor U45290 (N_45290,N_41056,N_41997);
and U45291 (N_45291,N_40450,N_41813);
nor U45292 (N_45292,N_40418,N_44363);
nand U45293 (N_45293,N_41766,N_43647);
or U45294 (N_45294,N_43801,N_42186);
nand U45295 (N_45295,N_40944,N_42547);
xnor U45296 (N_45296,N_43498,N_43605);
nor U45297 (N_45297,N_40508,N_41033);
or U45298 (N_45298,N_44318,N_43443);
and U45299 (N_45299,N_44309,N_43533);
and U45300 (N_45300,N_44051,N_43909);
nand U45301 (N_45301,N_44680,N_43927);
or U45302 (N_45302,N_42742,N_43747);
nand U45303 (N_45303,N_41956,N_41221);
and U45304 (N_45304,N_40366,N_44865);
or U45305 (N_45305,N_42256,N_42073);
and U45306 (N_45306,N_43815,N_40501);
or U45307 (N_45307,N_44493,N_44465);
or U45308 (N_45308,N_43813,N_44520);
xnor U45309 (N_45309,N_42664,N_44513);
and U45310 (N_45310,N_40469,N_43209);
and U45311 (N_45311,N_40751,N_44607);
nor U45312 (N_45312,N_41336,N_42949);
and U45313 (N_45313,N_42063,N_42065);
nand U45314 (N_45314,N_43810,N_40089);
and U45315 (N_45315,N_40528,N_41412);
nand U45316 (N_45316,N_44549,N_43395);
nor U45317 (N_45317,N_41099,N_42581);
and U45318 (N_45318,N_41157,N_41609);
nor U45319 (N_45319,N_44181,N_44089);
nand U45320 (N_45320,N_43594,N_40034);
or U45321 (N_45321,N_44711,N_44460);
nand U45322 (N_45322,N_42349,N_40338);
and U45323 (N_45323,N_44470,N_41864);
or U45324 (N_45324,N_44863,N_41284);
or U45325 (N_45325,N_43922,N_43583);
xnor U45326 (N_45326,N_44602,N_44145);
and U45327 (N_45327,N_41543,N_42816);
nor U45328 (N_45328,N_42672,N_42441);
nor U45329 (N_45329,N_44758,N_41830);
nand U45330 (N_45330,N_42930,N_42354);
and U45331 (N_45331,N_42279,N_42487);
or U45332 (N_45332,N_42546,N_44934);
nand U45333 (N_45333,N_43841,N_41554);
and U45334 (N_45334,N_44410,N_40046);
or U45335 (N_45335,N_40190,N_41574);
nor U45336 (N_45336,N_42351,N_44877);
xnor U45337 (N_45337,N_42590,N_43722);
and U45338 (N_45338,N_43589,N_40929);
xor U45339 (N_45339,N_41484,N_42981);
nor U45340 (N_45340,N_43917,N_41262);
xnor U45341 (N_45341,N_44557,N_43346);
or U45342 (N_45342,N_40923,N_40594);
nor U45343 (N_45343,N_43095,N_41852);
and U45344 (N_45344,N_40401,N_41518);
and U45345 (N_45345,N_41164,N_42712);
nand U45346 (N_45346,N_42203,N_41394);
nand U45347 (N_45347,N_42639,N_41001);
xor U45348 (N_45348,N_43699,N_44891);
xnor U45349 (N_45349,N_44717,N_41196);
and U45350 (N_45350,N_41779,N_43303);
nand U45351 (N_45351,N_40861,N_40772);
nor U45352 (N_45352,N_43540,N_41397);
or U45353 (N_45353,N_44458,N_44864);
or U45354 (N_45354,N_44888,N_42848);
nand U45355 (N_45355,N_43066,N_41693);
or U45356 (N_45356,N_41488,N_43216);
nand U45357 (N_45357,N_41436,N_43000);
and U45358 (N_45358,N_42144,N_42217);
nand U45359 (N_45359,N_41256,N_43814);
nand U45360 (N_45360,N_41713,N_41017);
and U45361 (N_45361,N_41694,N_43221);
or U45362 (N_45362,N_43891,N_42944);
or U45363 (N_45363,N_44705,N_41599);
or U45364 (N_45364,N_40161,N_40836);
xnor U45365 (N_45365,N_43213,N_42340);
and U45366 (N_45366,N_44483,N_41040);
nor U45367 (N_45367,N_42418,N_40324);
nand U45368 (N_45368,N_40582,N_43901);
or U45369 (N_45369,N_43807,N_41132);
nand U45370 (N_45370,N_41569,N_43753);
xor U45371 (N_45371,N_40972,N_43374);
xor U45372 (N_45372,N_44429,N_44924);
or U45373 (N_45373,N_41172,N_42569);
or U45374 (N_45374,N_42646,N_41153);
nand U45375 (N_45375,N_41385,N_41832);
or U45376 (N_45376,N_41075,N_44190);
nand U45377 (N_45377,N_40635,N_41697);
nand U45378 (N_45378,N_42436,N_42947);
and U45379 (N_45379,N_43665,N_41363);
nand U45380 (N_45380,N_41449,N_40483);
nand U45381 (N_45381,N_44901,N_40248);
nor U45382 (N_45382,N_40882,N_40675);
nor U45383 (N_45383,N_41161,N_43693);
nand U45384 (N_45384,N_40128,N_40036);
and U45385 (N_45385,N_40039,N_41106);
and U45386 (N_45386,N_44104,N_42200);
and U45387 (N_45387,N_40328,N_40075);
nor U45388 (N_45388,N_43560,N_40810);
or U45389 (N_45389,N_41340,N_41263);
and U45390 (N_45390,N_44603,N_44312);
nor U45391 (N_45391,N_41060,N_40310);
or U45392 (N_45392,N_40540,N_42975);
or U45393 (N_45393,N_40604,N_41968);
and U45394 (N_45394,N_40560,N_41986);
xor U45395 (N_45395,N_40173,N_44675);
xnor U45396 (N_45396,N_43737,N_40127);
or U45397 (N_45397,N_40606,N_42497);
nor U45398 (N_45398,N_44574,N_43432);
xor U45399 (N_45399,N_44789,N_42898);
nand U45400 (N_45400,N_44385,N_43173);
nor U45401 (N_45401,N_42027,N_44875);
or U45402 (N_45402,N_40538,N_42138);
nand U45403 (N_45403,N_44985,N_44691);
or U45404 (N_45404,N_42660,N_44728);
or U45405 (N_45405,N_43976,N_43884);
nor U45406 (N_45406,N_42782,N_44873);
or U45407 (N_45407,N_43760,N_41966);
nand U45408 (N_45408,N_40638,N_40750);
and U45409 (N_45409,N_41010,N_42993);
and U45410 (N_45410,N_41403,N_44156);
nand U45411 (N_45411,N_43057,N_40672);
nand U45412 (N_45412,N_44497,N_43044);
or U45413 (N_45413,N_43727,N_41223);
nor U45414 (N_45414,N_42824,N_42480);
or U45415 (N_45415,N_43328,N_43352);
or U45416 (N_45416,N_43582,N_43408);
nand U45417 (N_45417,N_44610,N_44964);
and U45418 (N_45418,N_40984,N_42640);
nor U45419 (N_45419,N_41143,N_42230);
nor U45420 (N_45420,N_43883,N_44323);
nand U45421 (N_45421,N_42378,N_43691);
nand U45422 (N_45422,N_41028,N_40888);
or U45423 (N_45423,N_41461,N_42595);
and U45424 (N_45424,N_42676,N_42756);
nand U45425 (N_45425,N_41945,N_41109);
nor U45426 (N_45426,N_41840,N_43609);
or U45427 (N_45427,N_41621,N_41155);
xnor U45428 (N_45428,N_41015,N_41024);
xor U45429 (N_45429,N_42240,N_42453);
nand U45430 (N_45430,N_42054,N_41144);
nor U45431 (N_45431,N_44777,N_42622);
or U45432 (N_45432,N_43593,N_43337);
xor U45433 (N_45433,N_44369,N_44596);
nand U45434 (N_45434,N_44559,N_41052);
nor U45435 (N_45435,N_41535,N_44809);
nor U45436 (N_45436,N_41837,N_41698);
nor U45437 (N_45437,N_44818,N_40657);
nor U45438 (N_45438,N_43448,N_40676);
or U45439 (N_45439,N_44329,N_43827);
nor U45440 (N_45440,N_40576,N_40137);
xor U45441 (N_45441,N_44010,N_40849);
and U45442 (N_45442,N_44642,N_41197);
or U45443 (N_45443,N_42342,N_42668);
nand U45444 (N_45444,N_42310,N_40162);
nor U45445 (N_45445,N_44791,N_41653);
nand U45446 (N_45446,N_44573,N_41908);
and U45447 (N_45447,N_42629,N_42355);
nor U45448 (N_45448,N_40012,N_44890);
or U45449 (N_45449,N_42365,N_43063);
nor U45450 (N_45450,N_41217,N_44430);
xor U45451 (N_45451,N_41509,N_41280);
xnor U45452 (N_45452,N_41110,N_42812);
nor U45453 (N_45453,N_40889,N_43394);
nor U45454 (N_45454,N_43192,N_44733);
or U45455 (N_45455,N_40808,N_43203);
and U45456 (N_45456,N_41096,N_42560);
nand U45457 (N_45457,N_42085,N_40148);
nand U45458 (N_45458,N_42931,N_42303);
nor U45459 (N_45459,N_43422,N_41548);
and U45460 (N_45460,N_43610,N_43913);
xnor U45461 (N_45461,N_41077,N_43853);
nor U45462 (N_45462,N_42637,N_40364);
nor U45463 (N_45463,N_40835,N_40298);
and U45464 (N_45464,N_44266,N_42817);
nor U45465 (N_45465,N_40045,N_44496);
and U45466 (N_45466,N_43720,N_41718);
xnor U45467 (N_45467,N_41255,N_43050);
and U45468 (N_45468,N_40269,N_44411);
nand U45469 (N_45469,N_41067,N_40435);
or U45470 (N_45470,N_40996,N_44572);
xor U45471 (N_45471,N_42599,N_40742);
or U45472 (N_45472,N_42154,N_42585);
and U45473 (N_45473,N_42853,N_40449);
nand U45474 (N_45474,N_43033,N_43134);
nor U45475 (N_45475,N_41820,N_44035);
nor U45476 (N_45476,N_42338,N_40579);
xor U45477 (N_45477,N_40526,N_40897);
nand U45478 (N_45478,N_44029,N_44762);
nor U45479 (N_45479,N_40499,N_41082);
nor U45480 (N_45480,N_44550,N_42272);
nor U45481 (N_45481,N_41602,N_44135);
xnor U45482 (N_45482,N_43074,N_43444);
nand U45483 (N_45483,N_44906,N_43171);
nand U45484 (N_45484,N_44583,N_43711);
nor U45485 (N_45485,N_41932,N_42984);
nand U45486 (N_45486,N_42454,N_40107);
and U45487 (N_45487,N_44649,N_40633);
nand U45488 (N_45488,N_40837,N_41603);
nand U45489 (N_45489,N_44434,N_44714);
and U45490 (N_45490,N_40759,N_42973);
nor U45491 (N_45491,N_43974,N_41446);
and U45492 (N_45492,N_42564,N_40968);
nand U45493 (N_45493,N_40014,N_43848);
nor U45494 (N_45494,N_43918,N_41322);
nor U45495 (N_45495,N_41209,N_42247);
or U45496 (N_45496,N_42631,N_40541);
nand U45497 (N_45497,N_43955,N_44930);
or U45498 (N_45498,N_40256,N_44140);
and U45499 (N_45499,N_41346,N_44899);
nand U45500 (N_45500,N_44783,N_42201);
nand U45501 (N_45501,N_42029,N_42605);
or U45502 (N_45502,N_41706,N_43073);
xor U45503 (N_45503,N_41210,N_43777);
nand U45504 (N_45504,N_40363,N_44201);
or U45505 (N_45505,N_44249,N_44097);
or U45506 (N_45506,N_41654,N_44511);
and U45507 (N_45507,N_40037,N_42432);
nand U45508 (N_45508,N_44959,N_43802);
nor U45509 (N_45509,N_41732,N_43948);
nor U45510 (N_45510,N_40281,N_40227);
and U45511 (N_45511,N_44614,N_44661);
or U45512 (N_45512,N_40376,N_43521);
and U45513 (N_45513,N_41810,N_41624);
nor U45514 (N_45514,N_41772,N_40815);
xnor U45515 (N_45515,N_40811,N_42901);
nand U45516 (N_45516,N_43415,N_40199);
nand U45517 (N_45517,N_40590,N_41395);
nand U45518 (N_45518,N_44432,N_40748);
nand U45519 (N_45519,N_43679,N_43654);
and U45520 (N_45520,N_41473,N_43445);
or U45521 (N_45521,N_43828,N_44109);
nand U45522 (N_45522,N_44676,N_43754);
or U45523 (N_45523,N_42343,N_41768);
nor U45524 (N_45524,N_44545,N_43725);
xor U45525 (N_45525,N_41427,N_42641);
or U45526 (N_45526,N_40006,N_44016);
nor U45527 (N_45527,N_43531,N_43305);
xnor U45528 (N_45528,N_41689,N_43106);
and U45529 (N_45529,N_40229,N_41675);
or U45530 (N_45530,N_41523,N_42305);
or U45531 (N_45531,N_44355,N_40970);
and U45532 (N_45532,N_41051,N_42807);
or U45533 (N_45533,N_43411,N_40351);
and U45534 (N_45534,N_40238,N_43306);
and U45535 (N_45535,N_44413,N_42698);
nand U45536 (N_45536,N_41505,N_41617);
nor U45537 (N_45537,N_42579,N_41113);
or U45538 (N_45538,N_43500,N_44046);
nor U45539 (N_45539,N_42871,N_40821);
and U45540 (N_45540,N_41218,N_44050);
nand U45541 (N_45541,N_42189,N_42584);
or U45542 (N_45542,N_42926,N_40177);
and U45543 (N_45543,N_44012,N_42361);
or U45544 (N_45544,N_44589,N_42252);
nor U45545 (N_45545,N_42533,N_43123);
or U45546 (N_45546,N_40258,N_44911);
and U45547 (N_45547,N_40316,N_43623);
nand U45548 (N_45548,N_41447,N_42666);
and U45549 (N_45549,N_44895,N_44315);
nor U45550 (N_45550,N_42125,N_42942);
xnor U45551 (N_45551,N_42209,N_41250);
xor U45552 (N_45552,N_42914,N_40774);
nor U45553 (N_45553,N_43229,N_42066);
or U45554 (N_45554,N_44476,N_43736);
xnor U45555 (N_45555,N_41738,N_40044);
nor U45556 (N_45556,N_42257,N_40583);
nor U45557 (N_45557,N_40495,N_41585);
nor U45558 (N_45558,N_43250,N_44540);
nor U45559 (N_45559,N_43541,N_42677);
nor U45560 (N_45560,N_43178,N_43357);
nand U45561 (N_45561,N_44340,N_42360);
or U45562 (N_45562,N_41914,N_42667);
or U45563 (N_45563,N_40530,N_43836);
nand U45564 (N_45564,N_43889,N_41891);
nand U45565 (N_45565,N_42187,N_40522);
and U45566 (N_45566,N_40855,N_42105);
nor U45567 (N_45567,N_43706,N_40434);
or U45568 (N_45568,N_41883,N_41136);
xnor U45569 (N_45569,N_42297,N_43396);
and U45570 (N_45570,N_43863,N_40684);
and U45571 (N_45571,N_43726,N_44843);
or U45572 (N_45572,N_42079,N_43894);
nor U45573 (N_45573,N_42743,N_44130);
nand U45574 (N_45574,N_40525,N_44773);
nor U45575 (N_45575,N_44124,N_41095);
nand U45576 (N_45576,N_40476,N_42098);
and U45577 (N_45577,N_41278,N_41227);
and U45578 (N_45578,N_40547,N_40249);
and U45579 (N_45579,N_40578,N_40711);
nor U45580 (N_45580,N_44003,N_43473);
nand U45581 (N_45581,N_41090,N_44677);
nor U45582 (N_45582,N_40061,N_44975);
nor U45583 (N_45583,N_43480,N_43687);
nor U45584 (N_45584,N_41206,N_44760);
and U45585 (N_45585,N_43880,N_43266);
or U45586 (N_45586,N_43506,N_41831);
nor U45587 (N_45587,N_42434,N_44120);
nand U45588 (N_45588,N_41763,N_44052);
nor U45589 (N_45589,N_40490,N_44624);
nor U45590 (N_45590,N_40393,N_42058);
xor U45591 (N_45591,N_43005,N_42207);
nor U45592 (N_45592,N_44961,N_43253);
and U45593 (N_45593,N_43214,N_42868);
nand U45594 (N_45594,N_44802,N_41047);
or U45595 (N_45595,N_41324,N_43028);
or U45596 (N_45596,N_44701,N_44319);
nor U45597 (N_45597,N_42906,N_40831);
nand U45598 (N_45598,N_42347,N_41703);
xnor U45599 (N_45599,N_41851,N_42060);
and U45600 (N_45600,N_42225,N_41850);
and U45601 (N_45601,N_44879,N_41178);
nand U45602 (N_45602,N_40971,N_43102);
and U45603 (N_45603,N_44036,N_44403);
nand U45604 (N_45604,N_42932,N_41875);
xnor U45605 (N_45605,N_44541,N_44535);
and U45606 (N_45606,N_43511,N_43469);
nand U45607 (N_45607,N_40777,N_42918);
or U45608 (N_45608,N_42387,N_40480);
nor U45609 (N_45609,N_44629,N_42068);
nor U45610 (N_45610,N_40521,N_42358);
nand U45611 (N_45611,N_44065,N_40847);
nand U45612 (N_45612,N_41507,N_40063);
nand U45613 (N_45613,N_44837,N_42763);
nor U45614 (N_45614,N_41337,N_41202);
nor U45615 (N_45615,N_42919,N_42815);
or U45616 (N_45616,N_44982,N_43430);
nand U45617 (N_45617,N_40293,N_44147);
nor U45618 (N_45618,N_42994,N_42223);
nand U45619 (N_45619,N_40025,N_41728);
nor U45620 (N_45620,N_44116,N_42840);
nor U45621 (N_45621,N_44146,N_43893);
and U45622 (N_45622,N_43403,N_44811);
nor U45623 (N_45623,N_43367,N_41973);
nor U45624 (N_45624,N_44869,N_41960);
nor U45625 (N_45625,N_42860,N_43874);
and U45626 (N_45626,N_43569,N_40916);
and U45627 (N_45627,N_40438,N_40885);
nand U45628 (N_45628,N_43329,N_41399);
nand U45629 (N_45629,N_40274,N_41636);
and U45630 (N_45630,N_43959,N_44233);
and U45631 (N_45631,N_43464,N_40109);
and U45632 (N_45632,N_41982,N_44117);
and U45633 (N_45633,N_40122,N_41510);
xor U45634 (N_45634,N_44616,N_44128);
nand U45635 (N_45635,N_43718,N_43695);
or U45636 (N_45636,N_44807,N_44544);
nand U45637 (N_45637,N_43390,N_42206);
and U45638 (N_45638,N_43557,N_40092);
nor U45639 (N_45639,N_41036,N_44346);
nand U45640 (N_45640,N_41347,N_42987);
and U45641 (N_45641,N_41671,N_44779);
nand U45642 (N_45642,N_40209,N_41066);
xor U45643 (N_45643,N_41628,N_40455);
and U45644 (N_45644,N_40117,N_44382);
nand U45645 (N_45645,N_44360,N_44659);
and U45646 (N_45646,N_44217,N_44547);
and U45647 (N_45647,N_44265,N_43662);
or U45648 (N_45648,N_43684,N_41039);
or U45649 (N_45649,N_41955,N_44168);
nand U45650 (N_45650,N_44372,N_42966);
nand U45651 (N_45651,N_40296,N_40178);
nand U45652 (N_45652,N_43712,N_40135);
and U45653 (N_45653,N_42609,N_41796);
nand U45654 (N_45654,N_41135,N_42790);
nand U45655 (N_45655,N_41630,N_41808);
nand U45656 (N_45656,N_43839,N_44453);
xor U45657 (N_45657,N_40253,N_40103);
nor U45658 (N_45658,N_42332,N_44292);
and U45659 (N_45659,N_42178,N_42644);
xor U45660 (N_45660,N_41472,N_43341);
nand U45661 (N_45661,N_44253,N_44017);
nand U45662 (N_45662,N_44154,N_40622);
nor U45663 (N_45663,N_41465,N_43024);
or U45664 (N_45664,N_43645,N_42808);
xnor U45665 (N_45665,N_43288,N_43885);
nand U45666 (N_45666,N_43529,N_40279);
nand U45667 (N_45667,N_40631,N_40575);
nand U45668 (N_45668,N_42905,N_44077);
xnor U45669 (N_45669,N_44452,N_44251);
or U45670 (N_45670,N_40623,N_44143);
nor U45671 (N_45671,N_44594,N_41215);
nand U45672 (N_45672,N_43233,N_42916);
xor U45673 (N_45673,N_40817,N_44151);
nor U45674 (N_45674,N_41288,N_41044);
and U45675 (N_45675,N_41969,N_44829);
nand U45676 (N_45676,N_40749,N_40554);
and U45677 (N_45677,N_42695,N_44922);
nor U45678 (N_45678,N_43692,N_43345);
nor U45679 (N_45679,N_43321,N_44679);
nand U45680 (N_45680,N_40026,N_43590);
and U45681 (N_45681,N_41058,N_43438);
nor U45682 (N_45682,N_44592,N_43805);
and U45683 (N_45683,N_40548,N_41743);
or U45684 (N_45684,N_43206,N_40990);
nand U45685 (N_45685,N_41829,N_44107);
nand U45686 (N_45686,N_42047,N_43604);
nor U45687 (N_45687,N_42656,N_42198);
and U45688 (N_45688,N_41158,N_41134);
nand U45689 (N_45689,N_43965,N_42945);
nor U45690 (N_45690,N_40084,N_42493);
nand U45691 (N_45691,N_43619,N_44400);
or U45692 (N_45692,N_44365,N_40989);
or U45693 (N_45693,N_41377,N_43846);
and U45694 (N_45694,N_40394,N_40783);
and U45695 (N_45695,N_41559,N_40927);
nand U45696 (N_45696,N_42788,N_43031);
and U45697 (N_45697,N_41726,N_42543);
and U45698 (N_45698,N_42769,N_44706);
xor U45699 (N_45699,N_41249,N_42495);
nand U45700 (N_45700,N_41126,N_41093);
nand U45701 (N_45701,N_42837,N_41993);
nor U45702 (N_45702,N_44447,N_41165);
and U45703 (N_45703,N_40090,N_44296);
or U45704 (N_45704,N_42962,N_44311);
nor U45705 (N_45705,N_43961,N_40652);
xnor U45706 (N_45706,N_40333,N_43177);
nand U45707 (N_45707,N_43774,N_40756);
nand U45708 (N_45708,N_44059,N_41417);
nor U45709 (N_45709,N_44868,N_42516);
nor U45710 (N_45710,N_42692,N_44215);
and U45711 (N_45711,N_41793,N_43280);
nand U45712 (N_45712,N_44121,N_44349);
nand U45713 (N_45713,N_41881,N_43947);
and U45714 (N_45714,N_44442,N_40674);
nand U45715 (N_45715,N_43954,N_43937);
nand U45716 (N_45716,N_41468,N_44776);
nor U45717 (N_45717,N_40868,N_42353);
and U45718 (N_45718,N_43278,N_44945);
xnor U45719 (N_45719,N_42937,N_44440);
nand U45720 (N_45720,N_43702,N_40827);
or U45721 (N_45721,N_42165,N_41723);
xnor U45722 (N_45722,N_41742,N_40913);
nand U45723 (N_45723,N_44118,N_40709);
xnor U45724 (N_45724,N_40779,N_43356);
and U45725 (N_45725,N_40447,N_44338);
xor U45726 (N_45726,N_44546,N_43479);
xor U45727 (N_45727,N_43550,N_42243);
and U45728 (N_45728,N_43795,N_44580);
or U45729 (N_45729,N_40245,N_43580);
or U45730 (N_45730,N_44611,N_40863);
or U45731 (N_45731,N_44832,N_41025);
nor U45732 (N_45732,N_40195,N_40556);
nor U45733 (N_45733,N_41391,N_41686);
nor U45734 (N_45734,N_42362,N_40873);
nor U45735 (N_45735,N_44084,N_40679);
or U45736 (N_45736,N_44260,N_41059);
xnor U45737 (N_45737,N_42478,N_44637);
or U45738 (N_45738,N_40208,N_43175);
and U45739 (N_45739,N_40613,N_44562);
xor U45740 (N_45740,N_40257,N_44650);
or U45741 (N_45741,N_43493,N_40308);
nor U45742 (N_45742,N_42202,N_41006);
nor U45743 (N_45743,N_41627,N_42350);
or U45744 (N_45744,N_44798,N_41987);
nor U45745 (N_45745,N_40940,N_41827);
and U45746 (N_45746,N_43538,N_40669);
nor U45747 (N_45747,N_41648,N_40302);
or U45748 (N_45748,N_40066,N_41642);
and U45749 (N_45749,N_42104,N_42886);
nor U45750 (N_45750,N_43890,N_40838);
or U45751 (N_45751,N_43534,N_41939);
or U45752 (N_45752,N_44916,N_44893);
and U45753 (N_45753,N_41758,N_42725);
nand U45754 (N_45754,N_40787,N_43426);
nand U45755 (N_45755,N_41493,N_40079);
or U45756 (N_45756,N_44090,N_41949);
nor U45757 (N_45757,N_41384,N_41704);
nand U45758 (N_45758,N_43198,N_43658);
xor U45759 (N_45759,N_41236,N_40422);
nor U45760 (N_45760,N_41261,N_44836);
or U45761 (N_45761,N_41315,N_43713);
nand U45762 (N_45762,N_41692,N_44764);
nor U45763 (N_45763,N_43870,N_41188);
or U45764 (N_45764,N_43728,N_43009);
and U45765 (N_45765,N_42928,N_44977);
nor U45766 (N_45766,N_42752,N_41456);
nand U45767 (N_45767,N_44871,N_40222);
nand U45768 (N_45768,N_42525,N_43599);
nor U45769 (N_45769,N_43433,N_44722);
nor U45770 (N_45770,N_41885,N_41562);
xnor U45771 (N_45771,N_42039,N_40441);
nor U45772 (N_45772,N_41386,N_40610);
or U45773 (N_45773,N_41234,N_44913);
xnor U45774 (N_45774,N_43745,N_40524);
nand U45775 (N_45775,N_41740,N_44579);
nor U45776 (N_45776,N_43135,N_41119);
or U45777 (N_45777,N_44462,N_44034);
or U45778 (N_45778,N_43992,N_42735);
and U45779 (N_45779,N_42308,N_40958);
nor U45780 (N_45780,N_43824,N_40138);
nor U45781 (N_45781,N_44846,N_40796);
and U45782 (N_45782,N_42346,N_44939);
xor U45783 (N_45783,N_44784,N_41481);
and U45784 (N_45784,N_41054,N_42227);
nor U45785 (N_45785,N_43768,N_43792);
xnor U45786 (N_45786,N_42531,N_44819);
nand U45787 (N_45787,N_40342,N_40072);
and U45788 (N_45788,N_43405,N_42567);
or U45789 (N_45789,N_44856,N_42689);
or U45790 (N_45790,N_40881,N_41440);
or U45791 (N_45791,N_41102,N_44112);
nor U45792 (N_45792,N_41130,N_41169);
and U45793 (N_45793,N_41877,N_41531);
nand U45794 (N_45794,N_43808,N_42271);
xor U45795 (N_45795,N_41581,N_42957);
and U45796 (N_45796,N_40527,N_44748);
and U45797 (N_45797,N_40035,N_40442);
xnor U45798 (N_45798,N_43101,N_41133);
or U45799 (N_45799,N_43183,N_44030);
nor U45800 (N_45800,N_42304,N_43353);
nor U45801 (N_45801,N_44208,N_43997);
nor U45802 (N_45802,N_44317,N_43981);
nor U45803 (N_45803,N_43724,N_40687);
nor U45804 (N_45804,N_41823,N_41947);
or U45805 (N_45805,N_42922,N_43882);
nand U45806 (N_45806,N_41027,N_41604);
and U45807 (N_45807,N_42445,N_41868);
nand U45808 (N_45808,N_40202,N_41312);
and U45809 (N_45809,N_42071,N_44622);
nor U45810 (N_45810,N_41457,N_40517);
or U45811 (N_45811,N_42196,N_44221);
nand U45812 (N_45812,N_44020,N_41494);
xor U45813 (N_45813,N_42439,N_42273);
or U45814 (N_45814,N_44053,N_44058);
or U45815 (N_45815,N_44224,N_43365);
nor U45816 (N_45816,N_43656,N_43401);
and U45817 (N_45817,N_41367,N_42325);
and U45818 (N_45818,N_41474,N_40607);
nor U45819 (N_45819,N_41388,N_44289);
nor U45820 (N_45820,N_40311,N_44498);
xnor U45821 (N_45821,N_40567,N_44839);
and U45822 (N_45822,N_44228,N_43630);
nor U45823 (N_45823,N_41884,N_43261);
nor U45824 (N_45824,N_41297,N_40878);
nand U45825 (N_45825,N_41321,N_44245);
nand U45826 (N_45826,N_42009,N_42846);
and U45827 (N_45827,N_40697,N_40492);
nand U45828 (N_45828,N_43164,N_40616);
nand U45829 (N_45829,N_44910,N_44671);
nor U45830 (N_45830,N_43089,N_42721);
nor U45831 (N_45831,N_41674,N_44566);
or U45832 (N_45832,N_41673,N_41491);
and U45833 (N_45833,N_42366,N_43764);
nor U45834 (N_45834,N_40371,N_42634);
xor U45835 (N_45835,N_42499,N_42658);
and U45836 (N_45836,N_41944,N_41387);
nand U45837 (N_45837,N_43026,N_40784);
nor U45838 (N_45838,N_44343,N_41402);
or U45839 (N_45839,N_44564,N_40619);
xnor U45840 (N_45840,N_42074,N_41233);
xor U45841 (N_45841,N_40608,N_43349);
and U45842 (N_45842,N_41807,N_43677);
nand U45843 (N_45843,N_43300,N_42157);
nor U45844 (N_45844,N_42199,N_44989);
or U45845 (N_45845,N_43283,N_43694);
nand U45846 (N_45846,N_44657,N_44669);
and U45847 (N_45847,N_43640,N_44658);
or U45848 (N_45848,N_41291,N_44381);
nand U45849 (N_45849,N_44731,N_44192);
xnor U45850 (N_45850,N_40898,N_40288);
nor U45851 (N_45851,N_41319,N_41657);
or U45852 (N_45852,N_41664,N_42197);
or U45853 (N_45853,N_41916,N_43136);
and U45854 (N_45854,N_43021,N_42479);
and U45855 (N_45855,N_44045,N_43046);
and U45856 (N_45856,N_42285,N_44071);
and U45857 (N_45857,N_40529,N_44703);
xor U45858 (N_45858,N_40361,N_43895);
or U45859 (N_45859,N_43195,N_44040);
or U45860 (N_45860,N_43449,N_42472);
xor U45861 (N_45861,N_43282,N_41240);
or U45862 (N_45862,N_41555,N_41855);
nand U45863 (N_45863,N_43536,N_41086);
and U45864 (N_45864,N_40486,N_40982);
xor U45865 (N_45865,N_42548,N_40856);
nor U45866 (N_45866,N_42524,N_43983);
nor U45867 (N_45867,N_42158,N_42702);
nor U45868 (N_45868,N_42036,N_44761);
nand U45869 (N_45869,N_41590,N_40105);
nor U45870 (N_45870,N_43269,N_40315);
nand U45871 (N_45871,N_44951,N_43242);
and U45872 (N_45872,N_40895,N_42496);
or U45873 (N_45873,N_42805,N_40636);
nor U45874 (N_45874,N_40213,N_42578);
or U45875 (N_45875,N_42856,N_41198);
or U45876 (N_45876,N_41958,N_41659);
xnor U45877 (N_45877,N_42979,N_44744);
nor U45878 (N_45878,N_41724,N_40155);
nor U45879 (N_45879,N_42773,N_41866);
and U45880 (N_45880,N_40383,N_43043);
nor U45881 (N_45881,N_40510,N_42867);
xor U45882 (N_45882,N_42298,N_44219);
nor U45883 (N_45883,N_43888,N_44142);
and U45884 (N_45884,N_44889,N_44397);
nor U45885 (N_45885,N_43564,N_40917);
or U45886 (N_45886,N_44110,N_40778);
and U45887 (N_45887,N_43072,N_44222);
nand U45888 (N_45888,N_42101,N_43294);
and U45889 (N_45889,N_43476,N_44647);
xnor U45890 (N_45890,N_42764,N_41899);
nand U45891 (N_45891,N_44252,N_43597);
nor U45892 (N_45892,N_44339,N_44332);
and U45893 (N_45893,N_42334,N_43200);
xor U45894 (N_45894,N_40659,N_43994);
and U45895 (N_45895,N_43163,N_42768);
and U45896 (N_45896,N_40790,N_40555);
xnor U45897 (N_45897,N_44643,N_40118);
or U45898 (N_45898,N_40626,N_41383);
nand U45899 (N_45899,N_40010,N_44944);
nor U45900 (N_45900,N_43224,N_40785);
nand U45901 (N_45901,N_44955,N_40644);
nand U45902 (N_45902,N_42559,N_42382);
nor U45903 (N_45903,N_42669,N_40259);
and U45904 (N_45904,N_42706,N_41294);
nand U45905 (N_45905,N_44512,N_40233);
nor U45906 (N_45906,N_42386,N_41608);
nor U45907 (N_45907,N_40866,N_43899);
and U45908 (N_45908,N_41709,N_42313);
xor U45909 (N_45909,N_42107,N_43232);
xnor U45910 (N_45910,N_43600,N_44388);
or U45911 (N_45911,N_40145,N_42530);
or U45912 (N_45912,N_44958,N_42008);
nor U45913 (N_45913,N_43483,N_41308);
nor U45914 (N_45914,N_42582,N_40094);
nand U45915 (N_45915,N_42897,N_43819);
nor U45916 (N_45916,N_41781,N_44554);
and U45917 (N_45917,N_43785,N_40198);
nor U45918 (N_45918,N_44158,N_44163);
or U45919 (N_45919,N_44820,N_42522);
nor U45920 (N_45920,N_40219,N_40440);
nand U45921 (N_45921,N_41924,N_44287);
or U45922 (N_45922,N_40534,N_40763);
xnor U45923 (N_45923,N_40918,N_40731);
or U45924 (N_45924,N_43468,N_44516);
or U45925 (N_45925,N_40482,N_43490);
or U45926 (N_45926,N_41596,N_43381);
nor U45927 (N_45927,N_44328,N_41800);
xor U45928 (N_45928,N_40358,N_40108);
nand U45929 (N_45929,N_42356,N_42137);
nor U45930 (N_45930,N_40974,N_41967);
nor U45931 (N_45931,N_43263,N_42124);
nor U45932 (N_45932,N_44081,N_43752);
nand U45933 (N_45933,N_43119,N_41799);
nor U45934 (N_45934,N_42174,N_40979);
nand U45935 (N_45935,N_44375,N_40743);
nor U45936 (N_45936,N_40069,N_42862);
or U45937 (N_45937,N_43859,N_41888);
nor U45938 (N_45938,N_40149,N_44641);
or U45939 (N_45939,N_41727,N_42540);
nor U45940 (N_45940,N_41668,N_41839);
xnor U45941 (N_45941,N_41152,N_43377);
and U45942 (N_45942,N_43359,N_40869);
or U45943 (N_45943,N_41381,N_42727);
nand U45944 (N_45944,N_41349,N_40559);
and U45945 (N_45945,N_41873,N_42823);
nand U45946 (N_45946,N_43465,N_43956);
or U45947 (N_45947,N_41037,N_41544);
nor U45948 (N_45948,N_42526,N_42889);
or U45949 (N_45949,N_42429,N_42870);
xor U45950 (N_45950,N_44803,N_41863);
or U45951 (N_45951,N_42625,N_42100);
xnor U45952 (N_45952,N_40432,N_44894);
nor U45953 (N_45953,N_44276,N_43504);
xnor U45954 (N_45954,N_42112,N_42411);
nand U45955 (N_45955,N_44604,N_44037);
and U45956 (N_45956,N_40452,N_43105);
nand U45957 (N_45957,N_42427,N_44634);
nor U45958 (N_45958,N_40345,N_44129);
or U45959 (N_45959,N_42081,N_43734);
nand U45960 (N_45960,N_44845,N_40064);
nor U45961 (N_45961,N_44759,N_44200);
or U45962 (N_45962,N_43844,N_41380);
nand U45963 (N_45963,N_40761,N_42654);
nor U45964 (N_45964,N_44161,N_42917);
and U45965 (N_45965,N_40928,N_40655);
nor U45966 (N_45966,N_40773,N_41721);
nand U45967 (N_45967,N_44896,N_42843);
and U45968 (N_45968,N_43586,N_40268);
nor U45969 (N_45969,N_40549,N_42103);
nand U45970 (N_45970,N_41049,N_40936);
and U45971 (N_45971,N_44704,N_40906);
and U45972 (N_45972,N_41749,N_42025);
or U45973 (N_45973,N_42801,N_41332);
nand U45974 (N_45974,N_40278,N_41685);
xor U45975 (N_45975,N_44732,N_40937);
and U45976 (N_45976,N_42428,N_42789);
and U45977 (N_45977,N_44881,N_40719);
xor U45978 (N_45978,N_43627,N_42405);
and U45979 (N_45979,N_42022,N_41454);
and U45980 (N_45980,N_44080,N_42070);
nor U45981 (N_45981,N_41989,N_43495);
nand U45982 (N_45982,N_41935,N_42851);
nand U45983 (N_45983,N_41327,N_42147);
and U45984 (N_45984,N_43399,N_42593);
and U45985 (N_45985,N_41406,N_44518);
or U45986 (N_45986,N_42483,N_40334);
nor U45987 (N_45987,N_44786,N_44467);
nor U45988 (N_45988,N_40611,N_42614);
nor U45989 (N_45989,N_40098,N_43006);
nand U45990 (N_45990,N_41242,N_40312);
and U45991 (N_45991,N_40403,N_44395);
nor U45992 (N_45992,N_42007,N_42381);
nor U45993 (N_45993,N_42075,N_44038);
and U45994 (N_45994,N_43277,N_40646);
nor U45995 (N_45995,N_40121,N_44897);
or U45996 (N_45996,N_44555,N_44223);
or U45997 (N_45997,N_44792,N_43149);
nor U45998 (N_45998,N_43022,N_41783);
or U45999 (N_45999,N_44024,N_44682);
nor U46000 (N_46000,N_42111,N_44283);
or U46001 (N_46001,N_44485,N_44269);
nor U46002 (N_46002,N_40065,N_42699);
xor U46003 (N_46003,N_42492,N_43553);
nand U46004 (N_46004,N_42408,N_43896);
nand U46005 (N_46005,N_40727,N_43174);
xnor U46006 (N_46006,N_42146,N_42184);
xnor U46007 (N_46007,N_42110,N_43938);
and U46008 (N_46008,N_42220,N_41762);
nor U46009 (N_46009,N_44909,N_43532);
xnor U46010 (N_46010,N_43978,N_41007);
nand U46011 (N_46011,N_40123,N_43309);
nand U46012 (N_46012,N_40725,N_44294);
nor U46013 (N_46013,N_44517,N_41701);
nand U46014 (N_46014,N_44737,N_43196);
or U46015 (N_46015,N_43223,N_41343);
xor U46016 (N_46016,N_41115,N_41785);
and U46017 (N_46017,N_41201,N_40277);
or U46018 (N_46018,N_40532,N_44644);
nand U46019 (N_46019,N_40241,N_43338);
and U46020 (N_46020,N_40870,N_44957);
nor U46021 (N_46021,N_44139,N_42398);
nor U46022 (N_46022,N_41366,N_42367);
nor U46023 (N_46023,N_41826,N_40890);
xor U46024 (N_46024,N_42903,N_41849);
nand U46025 (N_46025,N_43011,N_42397);
nand U46026 (N_46026,N_43755,N_43962);
nand U46027 (N_46027,N_40707,N_44105);
and U46028 (N_46028,N_43775,N_42159);
nand U46029 (N_46029,N_41219,N_42948);
nor U46030 (N_46030,N_42419,N_40580);
or U46031 (N_46031,N_43575,N_43437);
and U46032 (N_46032,N_42985,N_41441);
nor U46033 (N_46033,N_41097,N_40042);
nor U46034 (N_46034,N_41498,N_41186);
nand U46035 (N_46035,N_41744,N_43133);
or U46036 (N_46036,N_43568,N_44551);
and U46037 (N_46037,N_41905,N_44288);
nor U46038 (N_46038,N_44082,N_43931);
or U46039 (N_46039,N_41711,N_40284);
and U46040 (N_46040,N_40729,N_44854);
and U46041 (N_46041,N_42515,N_41710);
or U46042 (N_46042,N_41917,N_44750);
and U46043 (N_46043,N_40313,N_42967);
xor U46044 (N_46044,N_41137,N_43923);
nor U46045 (N_46045,N_44973,N_42780);
nor U46046 (N_46046,N_42841,N_41122);
nand U46047 (N_46047,N_41078,N_42078);
nand U46048 (N_46048,N_41526,N_41869);
nand U46049 (N_46049,N_43716,N_44387);
and U46050 (N_46050,N_41677,N_40591);
or U46051 (N_46051,N_43649,N_44377);
nand U46052 (N_46052,N_43742,N_43615);
nor U46053 (N_46053,N_41466,N_44114);
and U46054 (N_46054,N_44255,N_42859);
or U46055 (N_46055,N_40919,N_40019);
and U46056 (N_46056,N_44719,N_42577);
and U46057 (N_46057,N_43945,N_40850);
and U46058 (N_46058,N_40085,N_40421);
and U46059 (N_46059,N_42067,N_43673);
nand U46060 (N_46060,N_41934,N_40291);
nand U46061 (N_46061,N_44093,N_44062);
nor U46062 (N_46062,N_41865,N_42574);
or U46063 (N_46063,N_40479,N_40454);
nor U46064 (N_46064,N_42048,N_43264);
or U46065 (N_46065,N_43117,N_44665);
nor U46066 (N_46066,N_41534,N_42224);
nand U46067 (N_46067,N_40041,N_41886);
nor U46068 (N_46068,N_43446,N_42299);
nand U46069 (N_46069,N_44534,N_44123);
or U46070 (N_46070,N_44907,N_44822);
nand U46071 (N_46071,N_44127,N_43546);
or U46072 (N_46072,N_42050,N_40031);
and U46073 (N_46073,N_41909,N_40349);
or U46074 (N_46074,N_40407,N_40519);
nor U46075 (N_46075,N_41539,N_43861);
nor U46076 (N_46076,N_40232,N_40027);
nand U46077 (N_46077,N_40325,N_41751);
nor U46078 (N_46078,N_42053,N_43208);
nor U46079 (N_46079,N_40924,N_40545);
or U46080 (N_46080,N_44884,N_41613);
nor U46081 (N_46081,N_43482,N_40614);
and U46082 (N_46082,N_41788,N_44188);
xor U46083 (N_46083,N_43069,N_40926);
xnor U46084 (N_46084,N_42226,N_43892);
xnor U46085 (N_46085,N_44923,N_44466);
nor U46086 (N_46086,N_41634,N_44521);
and U46087 (N_46087,N_42131,N_42437);
nor U46088 (N_46088,N_44305,N_40797);
and U46089 (N_46089,N_40694,N_44825);
nand U46090 (N_46090,N_42778,N_42026);
or U46091 (N_46091,N_41267,N_42328);
nor U46092 (N_46092,N_41971,N_40509);
nand U46093 (N_46093,N_42537,N_44904);
and U46094 (N_46094,N_41750,N_42270);
or U46095 (N_46095,N_41587,N_42838);
nor U46096 (N_46096,N_42762,N_44383);
nand U46097 (N_46097,N_41141,N_43501);
xor U46098 (N_46098,N_40693,N_43385);
nor U46099 (N_46099,N_40879,N_40488);
or U46100 (N_46100,N_42363,N_41550);
nand U46101 (N_46101,N_42040,N_43409);
nand U46102 (N_46102,N_40032,N_44995);
xnor U46103 (N_46103,N_43227,N_42738);
and U46104 (N_46104,N_41348,N_41421);
xnor U46105 (N_46105,N_44100,N_40543);
or U46106 (N_46106,N_43320,N_41138);
and U46107 (N_46107,N_43284,N_43018);
and U46108 (N_46108,N_43113,N_41116);
and U46109 (N_46109,N_43577,N_44993);
and U46110 (N_46110,N_40133,N_43441);
and U46111 (N_46111,N_44965,N_41842);
and U46112 (N_46112,N_44351,N_41614);
and U46113 (N_46113,N_43274,N_44234);
and U46114 (N_46114,N_44307,N_40911);
or U46115 (N_46115,N_44738,N_44927);
and U46116 (N_46116,N_41880,N_40008);
and U46117 (N_46117,N_42527,N_42061);
nor U46118 (N_46118,N_44974,N_44730);
or U46119 (N_46119,N_42592,N_42783);
xor U46120 (N_46120,N_43059,N_40553);
nand U46121 (N_46121,N_43966,N_43475);
nor U46122 (N_46122,N_41281,N_44073);
and U46123 (N_46123,N_41731,N_43410);
nand U46124 (N_46124,N_41463,N_44014);
and U46125 (N_46125,N_44695,N_41362);
nor U46126 (N_46126,N_41926,N_41287);
nand U46127 (N_46127,N_43413,N_40922);
and U46128 (N_46128,N_40262,N_41451);
or U46129 (N_46129,N_42102,N_41376);
or U46130 (N_46130,N_41264,N_43719);
nand U46131 (N_46131,N_41790,N_41068);
nor U46132 (N_46132,N_41479,N_42455);
and U46133 (N_46133,N_40056,N_44191);
nand U46134 (N_46134,N_42057,N_40059);
xnor U46135 (N_46135,N_42894,N_40744);
nor U46136 (N_46136,N_40365,N_40969);
xor U46137 (N_46137,N_40096,N_43833);
xnor U46138 (N_46138,N_42645,N_41442);
and U46139 (N_46139,N_44490,N_41252);
or U46140 (N_46140,N_42863,N_44876);
or U46141 (N_46141,N_40650,N_41876);
nor U46142 (N_46142,N_41092,N_40336);
and U46143 (N_46143,N_42127,N_40147);
nand U46144 (N_46144,N_43146,N_41414);
nor U46145 (N_46145,N_44259,N_43964);
nand U46146 (N_46146,N_44281,N_41439);
and U46147 (N_46147,N_42953,N_40602);
and U46148 (N_46148,N_43290,N_41149);
xnor U46149 (N_46149,N_44367,N_42095);
and U46150 (N_46150,N_40309,N_44203);
xor U46151 (N_46151,N_43865,N_40113);
nor U46152 (N_46152,N_40998,N_40183);
nor U46153 (N_46153,N_43572,N_43404);
or U46154 (N_46154,N_40605,N_42331);
nand U46155 (N_46155,N_42288,N_44054);
nand U46156 (N_46156,N_40632,N_44813);
nand U46157 (N_46157,N_44426,N_42293);
or U46158 (N_46158,N_44439,N_42873);
or U46159 (N_46159,N_43664,N_41556);
xor U46160 (N_46160,N_42475,N_41700);
nand U46161 (N_46161,N_42208,N_44990);
nand U46162 (N_46162,N_40537,N_42550);
nand U46163 (N_46163,N_44056,N_44049);
and U46164 (N_46164,N_42481,N_44912);
and U46165 (N_46165,N_44257,N_40609);
or U46166 (N_46166,N_41496,N_42426);
nand U46167 (N_46167,N_44745,N_44800);
nor U46168 (N_46168,N_40181,N_40563);
nor U46169 (N_46169,N_40353,N_40786);
nor U46170 (N_46170,N_42538,N_43873);
nand U46171 (N_46171,N_41253,N_41680);
nand U46172 (N_46172,N_41996,N_43344);
nor U46173 (N_46173,N_41688,N_43016);
nand U46174 (N_46174,N_41061,N_42500);
or U46175 (N_46175,N_41453,N_41833);
xnor U46176 (N_46176,N_42284,N_43351);
and U46177 (N_46177,N_41467,N_43614);
nand U46178 (N_46178,N_44670,N_44855);
or U46179 (N_46179,N_44126,N_40299);
nand U46180 (N_46180,N_41619,N_40243);
and U46181 (N_46181,N_43843,N_44625);
and U46182 (N_46182,N_44471,N_41974);
or U46183 (N_46183,N_42704,N_43757);
xor U46184 (N_46184,N_40550,N_42396);
or U46185 (N_46185,N_43879,N_41401);
and U46186 (N_46186,N_41225,N_42116);
xnor U46187 (N_46187,N_44172,N_40715);
nand U46188 (N_46188,N_44968,N_42403);
nand U46189 (N_46189,N_44552,N_44115);
nor U46190 (N_46190,N_40752,N_41741);
nor U46191 (N_46191,N_42015,N_40337);
and U46192 (N_46192,N_41124,N_40456);
or U46193 (N_46193,N_41460,N_42316);
nand U46194 (N_46194,N_42858,N_44063);
nor U46195 (N_46195,N_42710,N_41211);
nor U46196 (N_46196,N_43298,N_44341);
or U46197 (N_46197,N_42093,N_42261);
and U46198 (N_46198,N_41504,N_40197);
xor U46199 (N_46199,N_41797,N_43625);
or U46200 (N_46200,N_41915,N_43832);
nand U46201 (N_46201,N_40523,N_43111);
nand U46202 (N_46202,N_42719,N_42275);
and U46203 (N_46203,N_44026,N_40801);
or U46204 (N_46204,N_40546,N_41626);
xnor U46205 (N_46205,N_44216,N_44271);
and U46206 (N_46206,N_42278,N_42121);
xnor U46207 (N_46207,N_43555,N_43257);
or U46208 (N_46208,N_42134,N_40992);
and U46209 (N_46209,N_43602,N_41361);
and U46210 (N_46210,N_41199,N_40780);
nor U46211 (N_46211,N_42829,N_44407);
or U46212 (N_46212,N_44274,N_44359);
or U46213 (N_46213,N_42188,N_42806);
or U46214 (N_46214,N_42878,N_42874);
and U46215 (N_46215,N_44187,N_43666);
and U46216 (N_46216,N_43549,N_44008);
nor U46217 (N_46217,N_42377,N_44204);
nor U46218 (N_46218,N_43088,N_44240);
and U46219 (N_46219,N_43651,N_42417);
nor U46220 (N_46220,N_44627,N_43085);
nand U46221 (N_46221,N_40769,N_44102);
or U46222 (N_46222,N_42977,N_40504);
or U46223 (N_46223,N_43854,N_41667);
or U46224 (N_46224,N_42221,N_44821);
nand U46225 (N_46225,N_40179,N_41094);
xnor U46226 (N_46226,N_43851,N_44582);
or U46227 (N_46227,N_42151,N_44526);
nor U46228 (N_46228,N_44925,N_40625);
or U46229 (N_46229,N_40300,N_41212);
xnor U46230 (N_46230,N_40326,N_41584);
and U46231 (N_46231,N_41512,N_41580);
nor U46232 (N_46232,N_44948,N_41998);
nand U46233 (N_46233,N_42787,N_44455);
or U46234 (N_46234,N_43262,N_42090);
or U46235 (N_46235,N_42244,N_41293);
or U46236 (N_46236,N_43387,N_44683);
xor U46237 (N_46237,N_41745,N_44947);
nor U46238 (N_46238,N_44280,N_40887);
nor U46239 (N_46239,N_43919,N_42882);
or U46240 (N_46240,N_43704,N_40460);
and U46241 (N_46241,N_43421,N_41087);
nand U46242 (N_46242,N_44220,N_44648);
nor U46243 (N_46243,N_40569,N_41492);
nand U46244 (N_46244,N_44408,N_40915);
xnor U46245 (N_46245,N_40806,N_43740);
xnor U46246 (N_46246,N_44684,N_40706);
or U46247 (N_46247,N_44421,N_43322);
nor U46248 (N_46248,N_44450,N_40901);
xnor U46249 (N_46249,N_40058,N_42885);
xnor U46250 (N_46250,N_44816,N_44882);
xor U46251 (N_46251,N_42653,N_42447);
nor U46252 (N_46252,N_40721,N_42549);
or U46253 (N_46253,N_43220,N_40303);
or U46254 (N_46254,N_43165,N_41180);
and U46255 (N_46255,N_43773,N_44096);
and U46256 (N_46256,N_40960,N_41919);
nand U46257 (N_46257,N_41105,N_44724);
nand U46258 (N_46258,N_44963,N_42740);
and U46259 (N_46259,N_41691,N_43207);
nand U46260 (N_46260,N_41471,N_40933);
nor U46261 (N_46261,N_44330,N_43944);
nand U46262 (N_46262,N_41695,N_41375);
and U46263 (N_46263,N_44628,N_42318);
and U46264 (N_46264,N_43680,N_44584);
or U46265 (N_46265,N_42421,N_42175);
nor U46266 (N_46266,N_43121,N_43709);
nand U46267 (N_46267,N_44568,N_44033);
nor U46268 (N_46268,N_40690,N_40765);
and U46269 (N_46269,N_44079,N_42233);
nor U46270 (N_46270,N_44376,N_44165);
or U46271 (N_46271,N_40574,N_41251);
nor U46272 (N_46272,N_41392,N_40234);
nor U46273 (N_46273,N_43703,N_41229);
xor U46274 (N_46274,N_40593,N_40175);
nand U46275 (N_46275,N_42621,N_44886);
nand U46276 (N_46276,N_41013,N_40431);
nand U46277 (N_46277,N_41725,N_40813);
nand U46278 (N_46278,N_40981,N_44914);
or U46279 (N_46279,N_42819,N_41950);
xor U46280 (N_46280,N_42565,N_42169);
nor U46281 (N_46281,N_44164,N_42185);
nand U46282 (N_46282,N_42797,N_42746);
or U46283 (N_46283,N_41246,N_44103);
nand U46284 (N_46284,N_41503,N_43628);
or U46285 (N_46285,N_42164,N_42012);
or U46286 (N_46286,N_42014,N_40166);
nor U46287 (N_46287,N_43039,N_42246);
or U46288 (N_46288,N_42043,N_44707);
nor U46289 (N_46289,N_40273,N_43047);
or U46290 (N_46290,N_43484,N_42514);
or U46291 (N_46291,N_42655,N_44742);
or U46292 (N_46292,N_43820,N_42109);
xnor U46293 (N_46293,N_40399,N_43912);
xnor U46294 (N_46294,N_42561,N_41156);
or U46295 (N_46295,N_44656,N_43137);
or U46296 (N_46296,N_40021,N_44928);
nor U46297 (N_46297,N_44106,N_40475);
xnor U46298 (N_46298,N_44522,N_40807);
nand U46299 (N_46299,N_41753,N_44366);
and U46300 (N_46300,N_44258,N_43611);
nand U46301 (N_46301,N_40212,N_41929);
and U46302 (N_46302,N_43301,N_43414);
and U46303 (N_46303,N_43412,N_41754);
and U46304 (N_46304,N_43877,N_44337);
nand U46305 (N_46305,N_43255,N_43114);
xor U46306 (N_46306,N_44461,N_43019);
xnor U46307 (N_46307,N_44155,N_41566);
nor U46308 (N_46308,N_40615,N_40485);
nand U46309 (N_46309,N_44969,N_43023);
nor U46310 (N_46310,N_41957,N_44194);
nor U46311 (N_46311,N_40740,N_43457);
xor U46312 (N_46312,N_42341,N_41034);
xor U46313 (N_46313,N_41563,N_41030);
nand U46314 (N_46314,N_43781,N_40686);
and U46315 (N_46315,N_42876,N_43689);
and U46316 (N_46316,N_43926,N_40367);
or U46317 (N_46317,N_43688,N_42028);
or U46318 (N_46318,N_43829,N_43193);
nand U46319 (N_46319,N_41235,N_41379);
nor U46320 (N_46320,N_40872,N_43646);
nor U46321 (N_46321,N_41739,N_43339);
xnor U46322 (N_46322,N_40049,N_41623);
or U46323 (N_46323,N_40535,N_40789);
or U46324 (N_46324,N_44510,N_43246);
and U46325 (N_46325,N_42969,N_43143);
or U46326 (N_46326,N_43406,N_42369);
or U46327 (N_46327,N_42486,N_43928);
or U46328 (N_46328,N_40226,N_40194);
or U46329 (N_46329,N_42030,N_42665);
or U46330 (N_46330,N_42847,N_43098);
or U46331 (N_46331,N_42833,N_43767);
and U46332 (N_46332,N_41607,N_42005);
nor U46333 (N_46333,N_44399,N_42839);
nor U46334 (N_46334,N_42714,N_44331);
or U46335 (N_46335,N_42031,N_44709);
and U46336 (N_46336,N_44533,N_42678);
nor U46337 (N_46337,N_43617,N_42888);
or U46338 (N_46338,N_42291,N_40599);
or U46339 (N_46339,N_40106,N_41435);
xor U46340 (N_46340,N_40200,N_43109);
xor U46341 (N_46341,N_40062,N_42724);
nor U46342 (N_46342,N_43784,N_43254);
nand U46343 (N_46343,N_44527,N_42879);
nor U46344 (N_46344,N_44801,N_43478);
nand U46345 (N_46345,N_44074,N_42705);
nand U46346 (N_46346,N_40841,N_43953);
nor U46347 (N_46347,N_44919,N_40188);
or U46348 (N_46348,N_44264,N_41016);
nor U46349 (N_46349,N_41519,N_43507);
nand U46350 (N_46350,N_42359,N_43273);
and U46351 (N_46351,N_43081,N_44806);
or U46352 (N_46352,N_42896,N_40696);
nand U46353 (N_46353,N_43364,N_40639);
or U46354 (N_46354,N_40182,N_41811);
nor U46355 (N_46355,N_43881,N_43368);
and U46356 (N_46356,N_40865,N_41290);
xor U46357 (N_46357,N_43462,N_43249);
nand U46358 (N_46358,N_41870,N_43631);
nand U46359 (N_46359,N_40264,N_40130);
nor U46360 (N_46360,N_41542,N_43850);
xnor U46361 (N_46361,N_42253,N_41084);
nand U46362 (N_46362,N_41176,N_41423);
nor U46363 (N_46363,N_44171,N_42827);
nor U46364 (N_46364,N_44805,N_43578);
or U46365 (N_46365,N_40414,N_43452);
or U46366 (N_46366,N_43036,N_44921);
nor U46367 (N_46367,N_43238,N_43335);
and U46368 (N_46368,N_43902,N_41057);
nor U46369 (N_46369,N_41775,N_43145);
or U46370 (N_46370,N_42020,N_44364);
or U46371 (N_46371,N_42289,N_41644);
nor U46372 (N_46372,N_41370,N_44831);
or U46373 (N_46373,N_44651,N_43002);
nor U46374 (N_46374,N_44778,N_42951);
nand U46375 (N_46375,N_41330,N_42409);
nor U46376 (N_46376,N_43427,N_40444);
nor U46377 (N_46377,N_40640,N_42647);
nand U46378 (N_46378,N_41835,N_44091);
nand U46379 (N_46379,N_40080,N_43397);
nand U46380 (N_46380,N_42051,N_43373);
nor U46381 (N_46381,N_42177,N_42899);
nand U46382 (N_46382,N_40464,N_44039);
nor U46383 (N_46383,N_43215,N_40908);
nand U46384 (N_46384,N_44391,N_40218);
and U46385 (N_46385,N_41846,N_44231);
or U46386 (N_46386,N_42572,N_40795);
or U46387 (N_46387,N_44763,N_44176);
or U46388 (N_46388,N_40991,N_40458);
nor U46389 (N_46389,N_44499,N_40339);
or U46390 (N_46390,N_42997,N_40959);
or U46391 (N_46391,N_40453,N_41755);
and U46392 (N_46392,N_42939,N_43051);
nor U46393 (N_46393,N_42739,N_40251);
nor U46394 (N_46394,N_41764,N_41983);
nor U46395 (N_46395,N_42019,N_40682);
or U46396 (N_46396,N_44797,N_41962);
nor U46397 (N_46397,N_41142,N_41814);
nand U46398 (N_46398,N_43327,N_43343);
nand U46399 (N_46399,N_40900,N_43017);
xor U46400 (N_46400,N_40387,N_44828);
nor U46401 (N_46401,N_42254,N_44531);
or U46402 (N_46402,N_43287,N_42236);
or U46403 (N_46403,N_43739,N_43730);
and U46404 (N_46404,N_41647,N_40237);
or U46405 (N_46405,N_41002,N_43271);
xor U46406 (N_46406,N_42471,N_43307);
nand U46407 (N_46407,N_44320,N_41508);
nand U46408 (N_46408,N_41424,N_42611);
xnor U46409 (N_46409,N_44501,N_44491);
or U46410 (N_46410,N_44708,N_42002);
nor U46411 (N_46411,N_40101,N_42153);
and U46412 (N_46412,N_41438,N_41995);
nand U46413 (N_46413,N_42113,N_42832);
nor U46414 (N_46414,N_44688,N_41338);
nor U46415 (N_46415,N_42191,N_40506);
nand U46416 (N_46416,N_40986,N_40668);
nand U46417 (N_46417,N_42248,N_43570);
nor U46418 (N_46418,N_44966,N_44590);
or U46419 (N_46419,N_40818,N_42092);
nand U46420 (N_46420,N_43668,N_43369);
and U46421 (N_46421,N_41276,N_42845);
nand U46422 (N_46422,N_42306,N_43289);
nor U46423 (N_46423,N_40168,N_42315);
or U46424 (N_46424,N_44726,N_43574);
nor U46425 (N_46425,N_41560,N_42326);
nor U46426 (N_46426,N_40814,N_40286);
nor U46427 (N_46427,N_44371,N_44636);
nor U46428 (N_46428,N_44561,N_44402);
nor U46429 (N_46429,N_42234,N_42087);
nand U46430 (N_46430,N_42713,N_43867);
and U46431 (N_46431,N_43903,N_44393);
nor U46432 (N_46432,N_42179,N_43471);
nor U46433 (N_46433,N_40356,N_44183);
nor U46434 (N_46434,N_41612,N_41795);
and U46435 (N_46435,N_41717,N_42596);
nor U46436 (N_46436,N_40465,N_43181);
or U46437 (N_46437,N_44950,N_43761);
nand U46438 (N_46438,N_44066,N_44725);
and U46439 (N_46439,N_40301,N_43076);
nor U46440 (N_46440,N_42941,N_44630);
nor U46441 (N_46441,N_43686,N_42504);
and U46442 (N_46442,N_42895,N_40290);
or U46443 (N_46443,N_41975,N_41662);
nand U46444 (N_46444,N_43127,N_43240);
nor U46445 (N_46445,N_43663,N_43528);
nand U46446 (N_46446,N_41275,N_43508);
or U46447 (N_46447,N_40930,N_43116);
nand U46448 (N_46448,N_40493,N_40201);
nor U46449 (N_46449,N_43596,N_44525);
and U46450 (N_46450,N_42835,N_44929);
and U46451 (N_46451,N_42978,N_40187);
xor U46452 (N_46452,N_42608,N_40871);
nor U46453 (N_46453,N_43371,N_42684);
nand U46454 (N_46454,N_41041,N_42877);
nand U46455 (N_46455,N_42995,N_42875);
xor U46456 (N_46456,N_40221,N_42730);
or U46457 (N_46457,N_40804,N_43450);
and U46458 (N_46458,N_42176,N_43608);
nand U46459 (N_46459,N_41588,N_41226);
nand U46460 (N_46460,N_44057,N_43434);
nor U46461 (N_46461,N_43921,N_42681);
nor U46462 (N_46462,N_41954,N_43157);
or U46463 (N_46463,N_40803,N_40741);
xor U46464 (N_46464,N_42096,N_41859);
or U46465 (N_46465,N_44196,N_40851);
nor U46466 (N_46466,N_41635,N_40126);
and U46467 (N_46467,N_44386,N_40374);
and U46468 (N_46468,N_43779,N_42908);
or U46469 (N_46469,N_40185,N_40146);
or U46470 (N_46470,N_42192,N_44775);
or U46471 (N_46471,N_41098,N_40141);
xor U46472 (N_46472,N_43304,N_44419);
or U46473 (N_46473,N_41941,N_40184);
nor U46474 (N_46474,N_43251,N_43505);
nor U46475 (N_46475,N_43530,N_42320);
and U46476 (N_46476,N_41469,N_42766);
nor U46477 (N_46477,N_44015,N_43598);
or U46478 (N_46478,N_44986,N_43681);
or U46479 (N_46479,N_41988,N_40210);
and U46480 (N_46480,N_42970,N_41681);
xor U46481 (N_46481,N_40099,N_43260);
and U46482 (N_46482,N_43265,N_40666);
nor U46483 (N_46483,N_40588,N_42094);
nand U46484 (N_46484,N_43543,N_41568);
and U46485 (N_46485,N_42935,N_41769);
and U46486 (N_46486,N_44085,N_41004);
and U46487 (N_46487,N_41415,N_44482);
nand U46488 (N_46488,N_44297,N_40953);
nand U46489 (N_46489,N_42122,N_40053);
and U46490 (N_46490,N_40976,N_42804);
nand U46491 (N_46491,N_41511,N_41853);
or U46492 (N_46492,N_43756,N_42488);
nor U46493 (N_46493,N_43519,N_41806);
nand U46494 (N_46494,N_40564,N_43940);
or U46495 (N_46495,N_43510,N_41696);
nor U46496 (N_46496,N_43563,N_44626);
or U46497 (N_46497,N_42907,N_43272);
nand U46498 (N_46498,N_42566,N_40514);
nor U46499 (N_46499,N_40705,N_44414);
nor U46500 (N_46500,N_43460,N_43030);
and U46501 (N_46501,N_43091,N_40767);
nor U46502 (N_46502,N_43672,N_42458);
nand U46503 (N_46503,N_43652,N_44374);
nand U46504 (N_46504,N_44405,N_42711);
nor U46505 (N_46505,N_41483,N_40658);
nor U46506 (N_46506,N_44852,N_42091);
nand U46507 (N_46507,N_41561,N_42961);
nand U46508 (N_46508,N_43545,N_44560);
nor U46509 (N_46509,N_40905,N_44285);
or U46510 (N_46510,N_42149,N_41265);
nor U46511 (N_46511,N_42450,N_41354);
or U46512 (N_46512,N_40670,N_43503);
nand U46513 (N_46513,N_44378,N_44638);
nor U46514 (N_46514,N_43491,N_40070);
nor U46515 (N_46515,N_42379,N_44597);
nor U46516 (N_46516,N_40112,N_43244);
or U46517 (N_46517,N_42799,N_44075);
nor U46518 (N_46518,N_44949,N_41567);
or U46519 (N_46519,N_44999,N_43058);
xor U46520 (N_46520,N_42422,N_40020);
or U46521 (N_46521,N_40189,N_43499);
or U46522 (N_46522,N_43456,N_44932);
nor U46523 (N_46523,N_44043,N_42463);
nor U46524 (N_46524,N_40948,N_43520);
or U46525 (N_46525,N_40000,N_40966);
nand U46526 (N_46526,N_43556,N_43660);
and U46527 (N_46527,N_42794,N_41045);
and U46528 (N_46528,N_42887,N_44486);
nor U46529 (N_46529,N_41683,N_41317);
and U46530 (N_46530,N_44996,N_42238);
nor U46531 (N_46531,N_41872,N_42651);
and U46532 (N_46532,N_44427,N_42992);
or U46533 (N_46533,N_40144,N_42482);
nand U46534 (N_46534,N_43701,N_42755);
nor U46535 (N_46535,N_43915,N_41248);
and U46536 (N_46536,N_42956,N_40100);
nor U46537 (N_46537,N_42380,N_41048);
nand U46538 (N_46538,N_40136,N_42545);
or U46539 (N_46539,N_42800,N_43717);
and U46540 (N_46540,N_40016,N_43950);
or U46541 (N_46541,N_42542,N_43331);
nand U46542 (N_46542,N_43162,N_43007);
nor U46543 (N_46543,N_43363,N_41325);
or U46544 (N_46544,N_41546,N_41784);
nand U46545 (N_46545,N_40997,N_43147);
nor U46546 (N_46546,N_42553,N_40892);
xor U46547 (N_46547,N_44324,N_44211);
xnor U46548 (N_46548,N_41304,N_43806);
nor U46549 (N_46549,N_40272,N_41964);
nand U46550 (N_46550,N_42657,N_41444);
nand U46551 (N_46551,N_40776,N_43566);
nand U46552 (N_46552,N_41279,N_43302);
or U46553 (N_46553,N_42770,N_43700);
nand U46554 (N_46554,N_42989,N_41666);
or U46555 (N_46555,N_40573,N_43065);
nor U46556 (N_46556,N_44086,N_43973);
or U46557 (N_46557,N_40661,N_44356);
and U46558 (N_46558,N_42643,N_42384);
and U46559 (N_46559,N_42971,N_42077);
or U46560 (N_46560,N_42282,N_40713);
and U46561 (N_46561,N_42892,N_40557);
nor U46562 (N_46562,N_41564,N_43217);
and U46563 (N_46563,N_44133,N_40955);
xor U46564 (N_46564,N_43128,N_42152);
nor U46565 (N_46565,N_40060,N_41756);
nor U46566 (N_46566,N_41848,N_42416);
or U46567 (N_46567,N_42589,N_44023);
nor U46568 (N_46568,N_40980,N_44213);
and U46569 (N_46569,N_41464,N_42772);
nand U46570 (N_46570,N_44588,N_42394);
nand U46571 (N_46571,N_43141,N_44556);
nor U46572 (N_46572,N_42715,N_42986);
and U46573 (N_46573,N_42021,N_44180);
xnor U46574 (N_46574,N_44044,N_42575);
nand U46575 (N_46575,N_44900,N_42741);
nand U46576 (N_46576,N_40139,N_40457);
and U46577 (N_46577,N_43391,N_40662);
nor U46578 (N_46578,N_43451,N_43463);
and U46579 (N_46579,N_42141,N_43696);
nand U46580 (N_46580,N_44069,N_42686);
nor U46581 (N_46581,N_44225,N_41174);
nand U46582 (N_46582,N_40842,N_41224);
nand U46583 (N_46583,N_40663,N_43071);
nand U46584 (N_46584,N_40473,N_42281);
nor U46585 (N_46585,N_40692,N_40951);
or U46586 (N_46586,N_43900,N_43603);
and U46587 (N_46587,N_41303,N_43453);
nor U46588 (N_46588,N_42211,N_41552);
nand U46589 (N_46589,N_42536,N_44712);
or U46590 (N_46590,N_40321,N_40993);
nand U46591 (N_46591,N_43925,N_44310);
nand U46592 (N_46592,N_43497,N_40433);
or U46593 (N_46593,N_42317,N_41268);
or U46594 (N_46594,N_43799,N_40978);
and U46595 (N_46595,N_42784,N_42814);
xnor U46596 (N_46596,N_40701,N_40965);
xnor U46597 (N_46597,N_41283,N_40335);
or U46598 (N_46598,N_41678,N_42148);
or U46599 (N_46599,N_43738,N_40883);
or U46600 (N_46600,N_43911,N_44316);
or U46601 (N_46601,N_41951,N_41167);
or U46602 (N_46602,N_41540,N_43167);
nand U46603 (N_46603,N_42433,N_44720);
or U46604 (N_46604,N_41736,N_40494);
nor U46605 (N_46605,N_41773,N_41114);
or U46606 (N_46606,N_44199,N_44702);
xor U46607 (N_46607,N_42097,N_41940);
nand U46608 (N_46608,N_43245,N_40350);
and U46609 (N_46609,N_41921,N_44235);
nand U46610 (N_46610,N_44752,N_44782);
and U46611 (N_46611,N_42872,N_40341);
nor U46612 (N_46612,N_43790,N_44344);
or U46613 (N_46613,N_42385,N_44569);
nor U46614 (N_46614,N_40038,N_43156);
or U46615 (N_46615,N_41459,N_41735);
and U46616 (N_46616,N_44390,N_41794);
and U46617 (N_46617,N_44640,N_42470);
nor U46618 (N_46618,N_40487,N_43375);
nand U46619 (N_46619,N_42913,N_43231);
nor U46620 (N_46620,N_42696,N_44025);
nand U46621 (N_46621,N_42521,N_44027);
and U46622 (N_46622,N_40380,N_40884);
or U46623 (N_46623,N_42401,N_44686);
xnor U46624 (N_46624,N_40728,N_41618);
and U46625 (N_46625,N_41495,N_42759);
or U46626 (N_46626,N_43741,N_41670);
or U46627 (N_46627,N_44350,N_41369);
or U46628 (N_46628,N_42682,N_42163);
and U46629 (N_46629,N_43523,N_44841);
xor U46630 (N_46630,N_43370,N_41231);
xor U46631 (N_46631,N_41203,N_44988);
nand U46632 (N_46632,N_44667,N_40378);
nand U46633 (N_46633,N_43236,N_42302);
nand U46634 (N_46634,N_44754,N_40029);
or U46635 (N_46635,N_43138,N_43222);
or U46636 (N_46636,N_41489,N_42813);
or U46637 (N_46637,N_44001,N_42881);
or U46638 (N_46638,N_42506,N_41389);
nor U46639 (N_46639,N_42314,N_41593);
and U46640 (N_46640,N_41420,N_42335);
nor U46641 (N_46641,N_41342,N_44446);
and U46642 (N_46642,N_44254,N_44218);
nor U46643 (N_46643,N_40231,N_44838);
nand U46644 (N_46644,N_42489,N_44935);
nor U46645 (N_46645,N_42259,N_40571);
and U46646 (N_46646,N_42210,N_42615);
nand U46647 (N_46647,N_43419,N_43765);
or U46648 (N_46648,N_44746,N_41499);
nor U46649 (N_46649,N_43049,N_43749);
or U46650 (N_46650,N_44530,N_42370);
or U46651 (N_46651,N_44666,N_41525);
nand U46652 (N_46652,N_44631,N_44506);
nor U46653 (N_46653,N_42024,N_40853);
xnor U46654 (N_46654,N_42775,N_44844);
or U46655 (N_46655,N_42128,N_43539);
or U46656 (N_46656,N_42276,N_42600);
and U46657 (N_46657,N_41616,N_40236);
nor U46658 (N_46658,N_44595,N_44962);
or U46659 (N_46659,N_41679,N_42324);
and U46660 (N_46660,N_42135,N_40551);
and U46661 (N_46661,N_44417,N_42693);
or U46662 (N_46662,N_44131,N_41818);
nor U46663 (N_46663,N_41478,N_44445);
nor U46664 (N_46664,N_41985,N_43094);
xnor U46665 (N_46665,N_43682,N_41359);
or U46666 (N_46666,N_42059,N_41112);
nor U46667 (N_46667,N_40914,N_44261);
nor U46668 (N_46668,N_43330,N_41012);
or U46669 (N_46669,N_44772,N_44423);
and U46670 (N_46670,N_43010,N_44278);
nand U46671 (N_46671,N_41129,N_40285);
nor U46672 (N_46672,N_40382,N_41537);
nand U46673 (N_46673,N_43372,N_42120);
or U46674 (N_46674,N_40158,N_41431);
and U46675 (N_46675,N_40844,N_41191);
and U46676 (N_46676,N_41123,N_42205);
nor U46677 (N_46677,N_43097,N_43562);
nand U46678 (N_46678,N_42000,N_41207);
or U46679 (N_46679,N_42181,N_40637);
or U46680 (N_46680,N_41216,N_41904);
or U46681 (N_46681,N_40437,N_44198);
xnor U46682 (N_46682,N_44509,N_43822);
and U46683 (N_46683,N_40439,N_42583);
and U46684 (N_46684,N_43436,N_40111);
or U46685 (N_46685,N_40952,N_43513);
or U46686 (N_46686,N_44536,N_40396);
xnor U46687 (N_46687,N_42072,N_43778);
xor U46688 (N_46688,N_40983,N_43474);
nor U46689 (N_46689,N_42323,N_44543);
or U46690 (N_46690,N_44048,N_43204);
and U46691 (N_46691,N_41805,N_40577);
nor U46692 (N_46692,N_41802,N_41104);
xor U46693 (N_46693,N_44874,N_41450);
nand U46694 (N_46694,N_43988,N_44195);
and U46695 (N_46695,N_40950,N_41936);
and U46696 (N_46696,N_44437,N_43624);
nand U46697 (N_46697,N_40235,N_43078);
nor U46698 (N_46698,N_44699,N_40802);
or U46699 (N_46699,N_42934,N_40758);
or U46700 (N_46700,N_42512,N_40239);
nand U46701 (N_46701,N_40533,N_40381);
nor U46702 (N_46702,N_42505,N_43323);
or U46703 (N_46703,N_41021,N_43746);
nand U46704 (N_46704,N_44404,N_42598);
and U46705 (N_46705,N_42785,N_44793);
and U46706 (N_46706,N_41959,N_42235);
nor U46707 (N_46707,N_43035,N_42959);
nor U46708 (N_46708,N_42003,N_40051);
or U46709 (N_46709,N_41529,N_41295);
or U46710 (N_46710,N_43845,N_41437);
nor U46711 (N_46711,N_44739,N_43144);
and U46712 (N_46712,N_41400,N_42925);
nor U46713 (N_46713,N_44785,N_42777);
nand U46714 (N_46714,N_42296,N_43219);
and U46715 (N_46715,N_43678,N_43669);
nor U46716 (N_46716,N_43416,N_43186);
nor U46717 (N_46717,N_43258,N_42588);
nor U46718 (N_46718,N_41547,N_43830);
or U46719 (N_46719,N_40764,N_41100);
nor U46720 (N_46720,N_41089,N_40862);
and U46721 (N_46721,N_43093,N_41222);
xor U46722 (N_46722,N_44284,N_40391);
and U46723 (N_46723,N_41611,N_40737);
xnor U46724 (N_46724,N_43001,N_40426);
and U46725 (N_46725,N_41629,N_40040);
or U46726 (N_46726,N_43866,N_40733);
and U46727 (N_46727,N_41445,N_43906);
or U46728 (N_46728,N_41310,N_44593);
and U46729 (N_46729,N_42792,N_41895);
nand U46730 (N_46730,N_42749,N_41480);
nor U46731 (N_46731,N_41882,N_42049);
nor U46732 (N_46732,N_40630,N_42688);
or U46733 (N_46733,N_42921,N_44433);
and U46734 (N_46734,N_40017,N_44028);
nand U46735 (N_46735,N_43671,N_40496);
nand U46736 (N_46736,N_42933,N_40446);
xor U46737 (N_46737,N_43008,N_43110);
and U46738 (N_46738,N_43013,N_42415);
and U46739 (N_46739,N_41314,N_43916);
nor U46740 (N_46740,N_40375,N_43188);
nor U46741 (N_46741,N_42535,N_41232);
nor U46742 (N_46742,N_44994,N_44755);
nor U46743 (N_46743,N_43125,N_43907);
nor U46744 (N_46744,N_40372,N_42258);
and U46745 (N_46745,N_43267,N_40708);
and U46746 (N_46746,N_42623,N_41238);
nand U46747 (N_46747,N_43618,N_42830);
and U46748 (N_46748,N_41610,N_41861);
nor U46749 (N_46749,N_40242,N_44849);
nand U46750 (N_46750,N_43729,N_43898);
and U46751 (N_46751,N_42344,N_42083);
nand U46752 (N_46752,N_40875,N_42910);
nor U46753 (N_46753,N_43169,N_40400);
and U46754 (N_46754,N_42114,N_40329);
nand U46755 (N_46755,N_41272,N_41475);
nor U46756 (N_46756,N_40395,N_42193);
xor U46757 (N_46757,N_43431,N_43643);
or U46758 (N_46758,N_41404,N_44409);
nand U46759 (N_46759,N_42442,N_40429);
nand U46760 (N_46760,N_42606,N_43626);
xnor U46761 (N_46761,N_44565,N_40023);
or U46762 (N_46762,N_43407,N_44348);
and U46763 (N_46763,N_41408,N_40596);
nand U46764 (N_46764,N_41029,N_44174);
or U46765 (N_46765,N_42652,N_41948);
nor U46766 (N_46766,N_44401,N_42017);
nor U46767 (N_46767,N_40174,N_41487);
nor U46768 (N_46768,N_41042,N_41524);
nor U46769 (N_46769,N_43871,N_44834);
or U46770 (N_46770,N_42119,N_41302);
or U46771 (N_46771,N_43439,N_44690);
or U46772 (N_46772,N_43770,N_44747);
or U46773 (N_46773,N_44765,N_44424);
nor U46774 (N_46774,N_42166,N_42834);
or U46775 (N_46775,N_44302,N_42249);
nand U46776 (N_46776,N_44473,N_44304);
and U46777 (N_46777,N_41791,N_43197);
nand U46778 (N_46778,N_43122,N_40689);
xnor U46779 (N_46779,N_42155,N_41638);
and U46780 (N_46780,N_40677,N_43535);
nor U46781 (N_46781,N_42836,N_41416);
or U46782 (N_46782,N_40653,N_41306);
nand U46783 (N_46783,N_44047,N_43939);
and U46784 (N_46784,N_41816,N_42466);
or U46785 (N_46785,N_42927,N_43929);
and U46786 (N_46786,N_41506,N_43941);
xnor U46787 (N_46787,N_43979,N_44244);
or U46788 (N_46788,N_41737,N_42391);
nand U46789 (N_46789,N_40018,N_42309);
nand U46790 (N_46790,N_43386,N_40612);
nor U46791 (N_46791,N_43886,N_43130);
nand U46792 (N_46792,N_41011,N_43172);
nand U46793 (N_46793,N_44415,N_42448);
nor U46794 (N_46794,N_44119,N_41407);
nor U46795 (N_46795,N_40648,N_41965);
nor U46796 (N_46796,N_44489,N_41482);
nor U46797 (N_46797,N_42844,N_42126);
nor U46798 (N_46798,N_44850,N_44587);
and U46799 (N_46799,N_43887,N_40398);
or U46800 (N_46800,N_40114,N_44570);
or U46801 (N_46801,N_41154,N_40902);
nand U46802 (N_46802,N_42675,N_40459);
nand U46803 (N_46803,N_43633,N_43914);
or U46804 (N_46804,N_42555,N_42912);
nor U46805 (N_46805,N_43565,N_41911);
and U46806 (N_46806,N_43379,N_40932);
xnor U46807 (N_46807,N_40921,N_40964);
or U46808 (N_46808,N_43228,N_40055);
and U46809 (N_46809,N_41187,N_42464);
nand U46810 (N_46810,N_44558,N_44479);
xor U46811 (N_46811,N_42286,N_43054);
or U46812 (N_46812,N_43809,N_40086);
and U46813 (N_46813,N_42266,N_40833);
and U46814 (N_46814,N_40471,N_40899);
and U46815 (N_46815,N_44306,N_43383);
nand U46816 (N_46816,N_42456,N_43667);
xnor U46817 (N_46817,N_43333,N_42262);
or U46818 (N_46818,N_40798,N_44398);
nor U46819 (N_46819,N_40886,N_44268);
nor U46820 (N_46820,N_40656,N_43969);
xor U46821 (N_46821,N_42171,N_40097);
or U46822 (N_46822,N_40739,N_42425);
xor U46823 (N_46823,N_43525,N_43732);
or U46824 (N_46824,N_43243,N_42849);
nor U46825 (N_46825,N_42760,N_44347);
nand U46826 (N_46826,N_41008,N_43313);
nand U46827 (N_46827,N_40702,N_40531);
and U46828 (N_46828,N_42728,N_43588);
and U46829 (N_46829,N_42786,N_44721);
nor U46830 (N_46830,N_40408,N_43544);
nor U46831 (N_46831,N_43933,N_42082);
or U46832 (N_46832,N_43592,N_40753);
nand U46833 (N_46833,N_43786,N_42687);
nand U46834 (N_46834,N_43340,N_43075);
and U46835 (N_46835,N_40995,N_40409);
and U46836 (N_46836,N_42968,N_43384);
and U46837 (N_46837,N_40738,N_44248);
nor U46838 (N_46838,N_40935,N_42339);
and U46839 (N_46839,N_44740,N_40754);
nor U46840 (N_46840,N_40228,N_41351);
xor U46841 (N_46841,N_44428,N_41128);
or U46842 (N_46842,N_41497,N_40498);
nand U46843 (N_46843,N_43943,N_40204);
or U46844 (N_46844,N_43905,N_42477);
nand U46845 (N_46845,N_43488,N_44678);
and U46846 (N_46846,N_41301,N_42610);
nor U46847 (N_46847,N_42292,N_41239);
nand U46848 (N_46848,N_41320,N_41640);
nand U46849 (N_46849,N_44632,N_41770);
and U46850 (N_46850,N_41373,N_40003);
and U46851 (N_46851,N_41978,N_41658);
or U46852 (N_46852,N_44771,N_44830);
nor U46853 (N_46853,N_40143,N_42449);
nand U46854 (N_46854,N_41274,N_43077);
and U46855 (N_46855,N_41121,N_44006);
and U46856 (N_46856,N_42274,N_43120);
nand U46857 (N_46857,N_44620,N_44475);
and U46858 (N_46858,N_44842,N_40544);
and U46859 (N_46859,N_41760,N_41927);
nand U46860 (N_46860,N_43769,N_40762);
xnor U46861 (N_46861,N_40829,N_41907);
nand U46862 (N_46862,N_42406,N_41003);
nor U46863 (N_46863,N_40909,N_43400);
or U46864 (N_46864,N_44960,N_43567);
nor U46865 (N_46865,N_42580,N_43199);
or U46866 (N_46866,N_43576,N_44941);
xnor U46867 (N_46867,N_42541,N_44586);
nand U46868 (N_46868,N_43516,N_42902);
nand U46869 (N_46869,N_43205,N_40566);
and U46870 (N_46870,N_44238,N_41637);
or U46871 (N_46871,N_43053,N_41822);
nor U46872 (N_46872,N_42850,N_40081);
and U46873 (N_46873,N_44327,N_44451);
xor U46874 (N_46874,N_44639,N_43099);
nand U46875 (N_46875,N_41266,N_41845);
nand U46876 (N_46876,N_41729,N_43676);
and U46877 (N_46877,N_41125,N_40013);
xnor U46878 (N_46878,N_43772,N_44633);
and U46879 (N_46879,N_44537,N_41175);
nand U46880 (N_46880,N_41184,N_40420);
nand U46881 (N_46881,N_43467,N_43537);
nor U46882 (N_46882,N_42440,N_41541);
xor U46883 (N_46883,N_43160,N_44920);
xor U46884 (N_46884,N_43803,N_41298);
nand U46885 (N_46885,N_43612,N_42591);
nor U46886 (N_46886,N_41643,N_40734);
and U46887 (N_46887,N_42718,N_43061);
nor U46888 (N_46888,N_43920,N_43551);
nor U46889 (N_46889,N_43621,N_42795);
nand U46890 (N_46890,N_40627,N_44507);
nor U46891 (N_46891,N_40142,N_44443);
or U46892 (N_46892,N_41890,N_41335);
nand U46893 (N_46893,N_44072,N_42707);
nor U46894 (N_46894,N_41663,N_40009);
nor U46895 (N_46895,N_43798,N_43152);
or U46896 (N_46896,N_43970,N_40834);
nand U46897 (N_46897,N_41259,N_43930);
nand U46898 (N_46898,N_42779,N_40683);
or U46899 (N_46899,N_40203,N_44295);
xor U46900 (N_46900,N_43083,N_40562);
xor U46901 (N_46901,N_43972,N_44769);
nor U46902 (N_46902,N_43225,N_41183);
or U46903 (N_46903,N_40413,N_40323);
and U46904 (N_46904,N_44645,N_43032);
nand U46905 (N_46905,N_43275,N_40788);
and U46906 (N_46906,N_42701,N_41101);
or U46907 (N_46907,N_44815,N_40224);
nor U46908 (N_46908,N_44591,N_44250);
xnor U46909 (N_46909,N_44918,N_44279);
or U46910 (N_46910,N_42991,N_42802);
or U46911 (N_46911,N_42998,N_43878);
nand U46912 (N_46912,N_41371,N_44660);
nand U46913 (N_46913,N_44926,N_44011);
nand U46914 (N_46914,N_42562,N_44070);
and U46915 (N_46915,N_43168,N_42452);
nor U46916 (N_46916,N_40828,N_43418);
or U46917 (N_46917,N_43218,N_41476);
nand U46918 (N_46918,N_44157,N_44767);
nor U46919 (N_46919,N_40586,N_44502);
nand U46920 (N_46920,N_40368,N_42960);
nor U46921 (N_46921,N_44456,N_44946);
and U46922 (N_46922,N_40848,N_42708);
or U46923 (N_46923,N_40876,N_43148);
nor U46924 (N_46924,N_44689,N_41913);
and U46925 (N_46925,N_41018,N_44241);
and U46926 (N_46926,N_40304,N_42143);
xnor U46927 (N_46927,N_41641,N_44068);
nand U46928 (N_46928,N_40076,N_44700);
or U46929 (N_46929,N_42854,N_41946);
xor U46930 (N_46930,N_43319,N_43910);
nand U46931 (N_46931,N_44814,N_41625);
nor U46932 (N_46932,N_42038,N_41181);
nand U46933 (N_46933,N_40967,N_44243);
and U46934 (N_46934,N_41419,N_41073);
xnor U46935 (N_46935,N_41214,N_44858);
or U46936 (N_46936,N_40392,N_44206);
nor U46937 (N_46937,N_41992,N_40322);
nand U46938 (N_46938,N_43606,N_40513);
and U46939 (N_46939,N_44664,N_43202);
nand U46940 (N_46940,N_44060,N_44099);
and U46941 (N_46941,N_41972,N_44448);
nor U46942 (N_46942,N_42765,N_40620);
nor U46943 (N_46943,N_41241,N_41352);
and U46944 (N_46944,N_42552,N_44826);
nand U46945 (N_46945,N_44983,N_43509);
and U46946 (N_46946,N_41894,N_44242);
nand U46947 (N_46947,N_43020,N_44980);
or U46948 (N_46948,N_41035,N_44981);
nand U46949 (N_46949,N_42140,N_43350);
nor U46950 (N_46950,N_42046,N_43958);
nand U46951 (N_46951,N_44833,N_40357);
nor U46952 (N_46952,N_42044,N_40503);
and U46953 (N_46953,N_41583,N_41527);
or U46954 (N_46954,N_40618,N_43552);
or U46955 (N_46955,N_40685,N_40028);
nand U46956 (N_46956,N_43788,N_43299);
nor U46957 (N_46957,N_41786,N_42573);
and U46958 (N_46958,N_44256,N_40823);
xor U46959 (N_46959,N_42923,N_44808);
nor U46960 (N_46960,N_41530,N_43957);
xnor U46961 (N_46961,N_42586,N_43904);
nand U46962 (N_46962,N_42822,N_41411);
nor U46963 (N_46963,N_41759,N_40511);
or U46964 (N_46964,N_41722,N_41014);
or U46965 (N_46965,N_41600,N_43161);
nand U46966 (N_46966,N_44578,N_44150);
xor U46967 (N_46967,N_41076,N_42414);
nand U46968 (N_46968,N_41356,N_42680);
nor U46969 (N_46969,N_40091,N_43420);
or U46970 (N_46970,N_44481,N_43977);
xor U46971 (N_46971,N_40416,N_42228);
xnor U46972 (N_46972,N_44857,N_40252);
or U46973 (N_46973,N_41557,N_40140);
nor U46974 (N_46974,N_41069,N_40671);
nand U46975 (N_46975,N_41331,N_44605);
xnor U46976 (N_46976,N_41843,N_42055);
nor U46977 (N_46977,N_41656,N_44083);
or U46978 (N_46978,N_42242,N_43100);
or U46979 (N_46979,N_42459,N_40572);
or U46980 (N_46980,N_43794,N_42250);
or U46981 (N_46981,N_41334,N_40104);
xor U46982 (N_46982,N_43080,N_40180);
nor U46983 (N_46983,N_43477,N_41344);
nor U46984 (N_46984,N_41050,N_44308);
or U46985 (N_46985,N_40634,N_43189);
nor U46986 (N_46986,N_40680,N_40306);
or U46987 (N_46987,N_42745,N_43868);
and U46988 (N_46988,N_42915,N_43548);
nand U46989 (N_46989,N_40710,N_43632);
or U46990 (N_46990,N_40977,N_42880);
or U46991 (N_46991,N_44903,N_43040);
and U46992 (N_46992,N_40800,N_40973);
nand U46993 (N_46993,N_42424,N_43847);
xnor U46994 (N_46994,N_42269,N_42529);
nand U46995 (N_46995,N_40022,N_43685);
or U46996 (N_46996,N_43184,N_44230);
nand U46997 (N_46997,N_44943,N_41151);
or U46998 (N_46998,N_44457,N_41589);
nor U46999 (N_46999,N_40603,N_42534);
nand U47000 (N_47000,N_42955,N_40115);
or U47001 (N_47001,N_43318,N_42842);
or U47002 (N_47002,N_44064,N_44735);
and U47003 (N_47003,N_40589,N_40102);
or U47004 (N_47004,N_42650,N_40470);
or U47005 (N_47005,N_42999,N_40261);
and U47006 (N_47006,N_40768,N_40193);
xor U47007 (N_47007,N_40794,N_44693);
and U47008 (N_47008,N_43601,N_44005);
and U47009 (N_47009,N_43744,N_42006);
and U47010 (N_47010,N_41798,N_44353);
and U47011 (N_47011,N_43595,N_40999);
nor U47012 (N_47012,N_44357,N_40695);
nand U47013 (N_47013,N_43710,N_40370);
or U47014 (N_47014,N_42750,N_40083);
or U47015 (N_47015,N_44210,N_40373);
nor U47016 (N_47016,N_40474,N_44851);
nor U47017 (N_47017,N_40415,N_43811);
nor U47018 (N_47018,N_43025,N_41200);
or U47019 (N_47019,N_40386,N_40595);
nor U47020 (N_47020,N_40688,N_43132);
nand U47021 (N_47021,N_40840,N_43360);
nand U47022 (N_47022,N_41578,N_43607);
or U47023 (N_47023,N_41705,N_40153);
xnor U47024 (N_47024,N_44938,N_41748);
or U47025 (N_47025,N_41501,N_42659);
nand U47026 (N_47026,N_43472,N_44273);
or U47027 (N_47027,N_41918,N_42319);
and U47028 (N_47028,N_40830,N_42312);
nand U47029 (N_47029,N_42767,N_40893);
and U47030 (N_47030,N_41108,N_43924);
and U47031 (N_47031,N_41433,N_42023);
nor U47032 (N_47032,N_41708,N_41977);
and U47033 (N_47033,N_44615,N_40152);
and U47034 (N_47034,N_44655,N_40052);
nand U47035 (N_47035,N_43571,N_42232);
or U47036 (N_47036,N_42729,N_44031);
or U47037 (N_47037,N_43259,N_41213);
nor U47038 (N_47038,N_40678,N_44189);
nand U47039 (N_47039,N_41834,N_41204);
nor U47040 (N_47040,N_42709,N_41046);
and U47041 (N_47041,N_40283,N_41661);
xor U47042 (N_47042,N_42277,N_44581);
nor U47043 (N_47043,N_41933,N_43932);
nor U47044 (N_47044,N_40068,N_40864);
nor U47045 (N_47045,N_44275,N_44967);
nand U47046 (N_47046,N_42831,N_41838);
nand U47047 (N_47047,N_42809,N_42213);
nor U47048 (N_47048,N_42603,N_40379);
nor U47049 (N_47049,N_41874,N_40087);
nor U47050 (N_47050,N_40799,N_40167);
and U47051 (N_47051,N_41208,N_40845);
nor U47052 (N_47052,N_40340,N_44623);
nor U47053 (N_47053,N_43417,N_42570);
xor U47054 (N_47054,N_41145,N_40962);
and U47055 (N_47055,N_41538,N_43690);
nand U47056 (N_47056,N_40314,N_44715);
or U47057 (N_47057,N_43613,N_42307);
or U47058 (N_47058,N_40246,N_43158);
nand U47059 (N_47059,N_43748,N_40397);
or U47060 (N_47060,N_44618,N_43644);
and U47061 (N_47061,N_43818,N_41429);
and U47062 (N_47062,N_42963,N_41702);
and U47063 (N_47063,N_41665,N_44673);
nand U47064 (N_47064,N_41812,N_42757);
nor U47065 (N_47065,N_42376,N_44303);
or U47066 (N_47066,N_43348,N_42393);
and U47067 (N_47067,N_43759,N_40030);
or U47068 (N_47068,N_43585,N_40427);
or U47069 (N_47069,N_42683,N_44380);
nand U47070 (N_47070,N_40211,N_42490);
nor U47071 (N_47071,N_41070,N_40131);
or U47072 (N_47072,N_44505,N_41393);
nand U47073 (N_47073,N_42041,N_44710);
and U47074 (N_47074,N_41118,N_44321);
and U47075 (N_47075,N_40170,N_41131);
or U47076 (N_47076,N_44113,N_44635);
or U47077 (N_47077,N_40907,N_43731);
nor U47078 (N_47078,N_42612,N_42373);
nor U47079 (N_47079,N_44692,N_41792);
nand U47080 (N_47080,N_44861,N_44599);
nor U47081 (N_47081,N_40904,N_44061);
or U47082 (N_47082,N_41245,N_40332);
nand U47083 (N_47083,N_44840,N_44796);
nand U47084 (N_47084,N_44770,N_41780);
nor U47085 (N_47085,N_41528,N_43835);
nand U47086 (N_47086,N_44207,N_43108);
nor U47087 (N_47087,N_40597,N_44696);
xnor U47088 (N_47088,N_42194,N_41719);
or U47089 (N_47089,N_44101,N_40698);
or U47090 (N_47090,N_41292,N_41147);
nor U47091 (N_47091,N_41901,N_42129);
or U47092 (N_47092,N_44055,N_44173);
nor U47093 (N_47093,N_44270,N_43455);
and U47094 (N_47094,N_42321,N_40943);
or U47095 (N_47095,N_42601,N_43424);
xnor U47096 (N_47096,N_42133,N_41860);
or U47097 (N_47097,N_42857,N_43362);
and U47098 (N_47098,N_41591,N_40949);
xnor U47099 (N_47099,N_44668,N_40478);
or U47100 (N_47100,N_42938,N_41761);
xnor U47101 (N_47101,N_41821,N_42673);
nand U47102 (N_47102,N_41651,N_44799);
or U47103 (N_47103,N_44917,N_42132);
and U47104 (N_47104,N_40292,N_44436);
nor U47105 (N_47105,N_44612,N_43124);
and U47106 (N_47106,N_42602,N_44774);
nor U47107 (N_47107,N_40164,N_43392);
and U47108 (N_47108,N_41645,N_43376);
or U47109 (N_47109,N_41277,N_42311);
or U47110 (N_47110,N_42697,N_44167);
nor U47111 (N_47111,N_41898,N_43743);
nor U47112 (N_47112,N_44094,N_40852);
nor U47113 (N_47113,N_42627,N_42218);
nor U47114 (N_47114,N_40500,N_43155);
xor U47115 (N_47115,N_43855,N_43996);
nand U47116 (N_47116,N_41413,N_43150);
xnor U47117 (N_47117,N_40461,N_41765);
nand U47118 (N_47118,N_40295,N_41273);
and U47119 (N_47119,N_40894,N_41734);
and U47120 (N_47120,N_40860,N_42413);
or U47121 (N_47121,N_44756,N_40681);
and U47122 (N_47122,N_44335,N_44662);
or U47123 (N_47123,N_44246,N_40384);
or U47124 (N_47124,N_41072,N_43573);
nor U47125 (N_47125,N_44812,N_42865);
nor U47126 (N_47126,N_43486,N_41669);
nand U47127 (N_47127,N_44598,N_44148);
nand U47128 (N_47128,N_44998,N_41062);
and U47129 (N_47129,N_40507,N_42407);
and U47130 (N_47130,N_44444,N_40176);
nor U47131 (N_47131,N_42940,N_42866);
xnor U47132 (N_47132,N_44539,N_44480);
nor U47133 (N_47133,N_43934,N_43037);
and U47134 (N_47134,N_40223,N_43787);
nand U47135 (N_47135,N_41117,N_41579);
and U47136 (N_47136,N_44542,N_41299);
or U47137 (N_47137,N_40186,N_42033);
and U47138 (N_47138,N_40954,N_44933);
xnor U47139 (N_47139,N_41778,N_43714);
or U47140 (N_47140,N_43012,N_42420);
xnor U47141 (N_47141,N_42820,N_44153);
and U47142 (N_47142,N_43771,N_40405);
nand U47143 (N_47143,N_41428,N_42241);
and U47144 (N_47144,N_41355,N_40843);
nor U47145 (N_47145,N_44298,N_42731);
nand U47146 (N_47146,N_40722,N_42855);
and U47147 (N_47147,N_44290,N_41300);
or U47148 (N_47148,N_42402,N_44902);
or U47149 (N_47149,N_42633,N_41847);
nor U47150 (N_47150,N_43783,N_41592);
xnor U47151 (N_47151,N_43315,N_43293);
or U47152 (N_47152,N_44322,N_42587);
nand U47153 (N_47153,N_44672,N_40267);
and U47154 (N_47154,N_43191,N_43524);
nand U47155 (N_47155,N_41815,N_43326);
or U47156 (N_47156,N_41378,N_40717);
nor U47157 (N_47157,N_43281,N_43291);
nand U47158 (N_47158,N_43256,N_44232);
nor U47159 (N_47159,N_41892,N_44132);
or U47160 (N_47160,N_41789,N_41358);
or U47161 (N_47161,N_42348,N_41514);
and U47162 (N_47162,N_40896,N_42597);
xnor U47163 (N_47163,N_42635,N_43442);
xor U47164 (N_47164,N_44007,N_41326);
nand U47165 (N_47165,N_41341,N_41577);
and U47166 (N_47166,N_44144,N_43041);
and U47167 (N_47167,N_40641,N_40730);
and U47168 (N_47168,N_40124,N_42115);
xnor U47169 (N_47169,N_42145,N_40649);
or U47170 (N_47170,N_42747,N_44936);
nand U47171 (N_47171,N_43587,N_40348);
and U47172 (N_47172,N_43735,N_40781);
nor U47173 (N_47173,N_43591,N_43355);
and U47174 (N_47174,N_43675,N_42649);
nor U47175 (N_47175,N_42501,N_44134);
xnor U47176 (N_47176,N_43248,N_40809);
nand U47177 (N_47177,N_44472,N_40746);
nand U47178 (N_47178,N_43082,N_44532);
or U47179 (N_47179,N_44170,N_42322);
nor U47180 (N_47180,N_40941,N_44713);
or U47181 (N_47181,N_42670,N_41345);
and U47182 (N_47182,N_43378,N_43425);
nor U47183 (N_47183,N_42069,N_42828);
xor U47184 (N_47184,N_43821,N_41952);
nor U47185 (N_47185,N_40629,N_41360);
nand U47186 (N_47186,N_43440,N_44042);
nand U47187 (N_47187,N_40255,N_41190);
and U47188 (N_47188,N_44653,N_41660);
or U47189 (N_47189,N_44694,N_41364);
nor U47190 (N_47190,N_42662,N_40819);
and U47191 (N_47191,N_43481,N_44872);
and U47192 (N_47192,N_41500,N_43982);
or U47193 (N_47193,N_40718,N_44991);
nand U47194 (N_47194,N_41177,N_42943);
nor U47195 (N_47195,N_44185,N_41032);
nor U47196 (N_47196,N_41425,N_41942);
or U47197 (N_47197,N_40600,N_42852);
nand U47198 (N_47198,N_43458,N_40132);
or U47199 (N_47199,N_44214,N_43800);
or U47200 (N_47200,N_43334,N_42674);
or U47201 (N_47201,N_40947,N_41422);
and U47202 (N_47202,N_41963,N_40854);
nor U47203 (N_47203,N_42511,N_40825);
nor U47204 (N_47204,N_43554,N_43252);
and U47205 (N_47205,N_41900,N_44780);
or U47206 (N_47206,N_40116,N_42287);
or U47207 (N_47207,N_44078,N_40859);
or U47208 (N_47208,N_42264,N_44108);
and U47209 (N_47209,N_41572,N_44524);
nand U47210 (N_47210,N_40165,N_40491);
and U47211 (N_47211,N_44342,N_41486);
xor U47212 (N_47212,N_42620,N_40369);
nand U47213 (N_47213,N_42694,N_44179);
xor U47214 (N_47214,N_43816,N_41597);
and U47215 (N_47215,N_41912,N_44212);
nand U47216 (N_47216,N_40160,N_43751);
or U47217 (N_47217,N_43496,N_44463);
and U47218 (N_47218,N_40561,N_44449);
nor U47219 (N_47219,N_43354,N_42231);
or U47220 (N_47220,N_44892,N_40791);
or U47221 (N_47221,N_40647,N_42300);
nor U47222 (N_47222,N_42551,N_41085);
and U47223 (N_47223,N_44092,N_40735);
xor U47224 (N_47224,N_40891,N_44368);
xnor U47225 (N_47225,N_44122,N_40832);
xor U47226 (N_47226,N_43459,N_43140);
nand U47227 (N_47227,N_43347,N_44209);
nor U47228 (N_47228,N_40665,N_43336);
and U47229 (N_47229,N_40129,N_41533);
or U47230 (N_47230,N_44138,N_43995);
xor U47231 (N_47231,N_43179,N_40934);
nor U47232 (N_47232,N_43316,N_44848);
nor U47233 (N_47233,N_44729,N_40664);
nand U47234 (N_47234,N_41083,N_42182);
and U47235 (N_47235,N_40477,N_44004);
nor U47236 (N_47236,N_43670,N_42539);
nand U47237 (N_47237,N_44334,N_40125);
and U47238 (N_47238,N_42123,N_44159);
nor U47239 (N_47239,N_43908,N_43487);
nor U47240 (N_47240,N_40592,N_41684);
and U47241 (N_47241,N_41237,N_42294);
and U47242 (N_47242,N_43176,N_40151);
nor U47243 (N_47243,N_43247,N_41893);
nor U47244 (N_47244,N_41043,N_43234);
nor U47245 (N_47245,N_40581,N_43062);
xor U47246 (N_47246,N_44160,N_43276);
and U47247 (N_47247,N_43561,N_41398);
nand U47248 (N_47248,N_42042,N_40004);
nand U47249 (N_47249,N_41887,N_43989);
or U47250 (N_47250,N_40287,N_44835);
nor U47251 (N_47251,N_40839,N_44600);
nand U47252 (N_47252,N_44313,N_44435);
and U47253 (N_47253,N_43968,N_44389);
and U47254 (N_47254,N_41782,N_40704);
or U47255 (N_47255,N_43237,N_43999);
and U47256 (N_47256,N_41477,N_40220);
nor U47257 (N_47257,N_40319,N_40451);
nor U47258 (N_47258,N_40445,N_40961);
or U47259 (N_47259,N_43840,N_44866);
or U47260 (N_47260,N_40404,N_41311);
nand U47261 (N_47261,N_43637,N_41063);
and U47262 (N_47262,N_40359,N_40007);
xor U47263 (N_47263,N_43838,N_41551);
or U47264 (N_47264,N_42032,N_41328);
and U47265 (N_47265,N_41910,N_43332);
and U47266 (N_47266,N_44617,N_44336);
nor U47267 (N_47267,N_40215,N_44262);
nor U47268 (N_47268,N_42357,N_42485);
nand U47269 (N_47269,N_42703,N_41228);
nor U47270 (N_47270,N_41712,N_40565);
and U47271 (N_47271,N_44394,N_44263);
and U47272 (N_47272,N_42337,N_44915);
or U47273 (N_47273,N_42810,N_40294);
and U47274 (N_47274,N_41448,N_43984);
nand U47275 (N_47275,N_41220,N_43064);
or U47276 (N_47276,N_43092,N_40957);
nand U47277 (N_47277,N_41270,N_42170);
xnor U47278 (N_47278,N_44125,N_42864);
nor U47279 (N_47279,N_40331,N_43308);
or U47280 (N_47280,N_42423,N_42260);
or U47281 (N_47281,N_44795,N_40820);
and U47282 (N_47282,N_44942,N_44186);
nor U47283 (N_47283,N_40412,N_41903);
or U47284 (N_47284,N_44136,N_44358);
nand U47285 (N_47285,N_40826,N_43380);
or U47286 (N_47286,N_40002,N_44345);
nor U47287 (N_47287,N_44519,N_43182);
or U47288 (N_47288,N_40169,N_40539);
or U47289 (N_47289,N_44862,N_40327);
nor U47290 (N_47290,N_42632,N_44931);
xnor U47291 (N_47291,N_41079,N_43715);
nand U47292 (N_47292,N_43067,N_42388);
nor U47293 (N_47293,N_44718,N_43849);
or U47294 (N_47294,N_44293,N_44794);
xor U47295 (N_47295,N_42544,N_43526);
nand U47296 (N_47296,N_40805,N_44749);
and U47297 (N_47297,N_44197,N_40516);
nand U47298 (N_47298,N_43635,N_42172);
nand U47299 (N_47299,N_42513,N_42604);
and U47300 (N_47300,N_40824,N_43721);
and U47301 (N_47301,N_42507,N_42890);
and U47302 (N_47302,N_42010,N_41930);
xnor U47303 (N_47303,N_40307,N_41953);
or U47304 (N_47304,N_40088,N_42509);
nand U47305 (N_47305,N_44422,N_43268);
or U47306 (N_47306,N_41357,N_40956);
and U47307 (N_47307,N_40716,N_41896);
and U47308 (N_47308,N_42239,N_41931);
xor U47309 (N_47309,N_40355,N_44406);
nand U47310 (N_47310,N_41620,N_40505);
nand U47311 (N_47311,N_43661,N_41990);
xor U47312 (N_47312,N_40171,N_42520);
nor U47313 (N_47313,N_41139,N_41652);
xnor U47314 (N_47314,N_44325,N_42216);
and U47315 (N_47315,N_40793,N_42168);
or U47316 (N_47316,N_43683,N_41372);
nand U47317 (N_47317,N_44205,N_41774);
nand U47318 (N_47318,N_43842,N_42130);
or U47319 (N_47319,N_42626,N_41038);
nand U47320 (N_47320,N_44585,N_44162);
or U47321 (N_47321,N_42607,N_42929);
and U47322 (N_47322,N_44621,N_40673);
and U47323 (N_47323,N_41000,N_43659);
nor U47324 (N_47324,N_43547,N_43869);
and U47325 (N_47325,N_43558,N_43492);
nor U47326 (N_47326,N_42045,N_41586);
and U47327 (N_47327,N_43858,N_42636);
nor U47328 (N_47328,N_42811,N_40276);
or U47329 (N_47329,N_43428,N_43942);
nand U47330 (N_47330,N_43447,N_43311);
or U47331 (N_47331,N_42390,N_40385);
nor U47332 (N_47332,N_42106,N_44076);
nor U47333 (N_47333,N_44601,N_42748);
or U47334 (N_47334,N_43194,N_42195);
and U47335 (N_47335,N_42295,N_42333);
nand U47336 (N_47336,N_40770,N_42744);
nor U47337 (N_47337,N_42412,N_41598);
or U47338 (N_47338,N_42118,N_41752);
or U47339 (N_47339,N_40206,N_42183);
or U47340 (N_47340,N_43860,N_40939);
and U47341 (N_47341,N_41595,N_43579);
and U47342 (N_47342,N_41923,N_43960);
and U47343 (N_47343,N_43864,N_42474);
xnor U47344 (N_47344,N_40760,N_43154);
nor U47345 (N_47345,N_40119,N_42965);
nand U47346 (N_47346,N_40515,N_41286);
nor U47347 (N_47347,N_42528,N_40700);
nand U47348 (N_47348,N_41146,N_41650);
nand U47349 (N_47349,N_40074,N_41515);
nor U47350 (N_47350,N_41871,N_43852);
or U47351 (N_47351,N_40425,N_41305);
and U47352 (N_47352,N_41746,N_43485);
or U47353 (N_47353,N_40643,N_42327);
or U47354 (N_47354,N_44314,N_44326);
xor U47355 (N_47355,N_42410,N_41111);
or U47356 (N_47356,N_42726,N_41490);
or U47357 (N_47357,N_43317,N_44087);
or U47358 (N_47358,N_40910,N_40043);
nand U47359 (N_47359,N_41020,N_42716);
or U47360 (N_47360,N_44182,N_41545);
xnor U47361 (N_47361,N_44824,N_43470);
nor U47362 (N_47362,N_42180,N_42503);
and U47363 (N_47363,N_42251,N_41803);
nor U47364 (N_47364,N_44362,N_40568);
nand U47365 (N_47365,N_41316,N_44392);
nor U47366 (N_47366,N_42013,N_44652);
nor U47367 (N_47367,N_43723,N_44495);
xor U47368 (N_47368,N_40156,N_40775);
or U47369 (N_47369,N_43998,N_44674);
or U47370 (N_47370,N_42150,N_42430);
nand U47371 (N_47371,N_40320,N_44867);
nor U47372 (N_47372,N_40497,N_40260);
and U47373 (N_47373,N_43796,N_43466);
and U47374 (N_47374,N_43971,N_42088);
xor U47375 (N_47375,N_40755,N_42139);
or U47376 (N_47376,N_40468,N_40782);
xor U47377 (N_47377,N_40011,N_44286);
or U47378 (N_47378,N_44032,N_43239);
and U47379 (N_47379,N_42190,N_43129);
and U47380 (N_47380,N_41682,N_44474);
and U47381 (N_47381,N_40732,N_40617);
and U47382 (N_47382,N_43826,N_44987);
nor U47383 (N_47383,N_41462,N_42345);
nor U47384 (N_47384,N_44487,N_40558);
nor U47385 (N_47385,N_41576,N_43389);
nor U47386 (N_47386,N_43793,N_41836);
nor U47387 (N_47387,N_42734,N_42004);
xor U47388 (N_47388,N_42972,N_40443);
or U47389 (N_47389,N_44687,N_41819);
and U47390 (N_47390,N_43296,N_44464);
or U47391 (N_47391,N_40263,N_40994);
nor U47392 (N_47392,N_40724,N_43139);
nand U47393 (N_47393,N_41994,N_42064);
nand U47394 (N_47394,N_40054,N_43804);
and U47395 (N_47395,N_43096,N_40945);
and U47396 (N_47396,N_44227,N_44418);
or U47397 (N_47397,N_41980,N_41019);
nand U47398 (N_47398,N_44528,N_43776);
xnor U47399 (N_47399,N_42990,N_44992);
xor U47400 (N_47400,N_41053,N_41192);
nand U47401 (N_47401,N_40462,N_41409);
nand U47402 (N_47402,N_44504,N_44098);
nor U47403 (N_47403,N_41353,N_40271);
nand U47404 (N_47404,N_42467,N_43153);
or U47405 (N_47405,N_40157,N_43087);
nand U47406 (N_47406,N_44953,N_40858);
nand U47407 (N_47407,N_42691,N_43398);
or U47408 (N_47408,N_44095,N_40481);
nand U47409 (N_47409,N_43489,N_43131);
or U47410 (N_47410,N_40660,N_40920);
and U47411 (N_47411,N_41205,N_42946);
and U47412 (N_47412,N_44567,N_44282);
nand U47413 (N_47413,N_42469,N_43985);
nor U47414 (N_47414,N_43875,N_40946);
and U47415 (N_47415,N_42498,N_43514);
nor U47416 (N_47416,N_40216,N_43639);
and U47417 (N_47417,N_44859,N_40163);
nand U47418 (N_47418,N_40448,N_44860);
and U47419 (N_47419,N_40024,N_41170);
nand U47420 (N_47420,N_41976,N_43241);
nand U47421 (N_47421,N_42776,N_43584);
and U47422 (N_47422,N_43515,N_43616);
nand U47423 (N_47423,N_44810,N_44237);
and U47424 (N_47424,N_42793,N_43361);
and U47425 (N_47425,N_41260,N_44663);
nand U47426 (N_47426,N_44997,N_43107);
nand U47427 (N_47427,N_43279,N_42389);
xor U47428 (N_47428,N_40699,N_44978);
or U47429 (N_47429,N_41522,N_41878);
and U47430 (N_47430,N_43151,N_43823);
and U47431 (N_47431,N_42265,N_40857);
nand U47432 (N_47432,N_40297,N_41970);
nand U47433 (N_47433,N_42556,N_43990);
or U47434 (N_47434,N_40812,N_40289);
nand U47435 (N_47435,N_41254,N_40816);
nor U47436 (N_47436,N_40377,N_40214);
nor U47437 (N_47437,N_41405,N_40598);
nor U47438 (N_47438,N_43542,N_44041);
or U47439 (N_47439,N_43791,N_44438);
xor U47440 (N_47440,N_41961,N_41150);
or U47441 (N_47441,N_41747,N_43648);
nand U47442 (N_47442,N_43090,N_40428);
nand U47443 (N_47443,N_40703,N_42435);
nand U47444 (N_47444,N_40093,N_41282);
and U47445 (N_47445,N_42215,N_41804);
and U47446 (N_47446,N_42404,N_42663);
xnor U47447 (N_47447,N_40352,N_42460);
nand U47448 (N_47448,N_43862,N_41676);
and U47449 (N_47449,N_43641,N_44971);
or U47450 (N_47450,N_42761,N_42558);
xnor U47451 (N_47451,N_43620,N_42791);
nor U47452 (N_47452,N_40963,N_44379);
and U47453 (N_47453,N_44523,N_40150);
and U47454 (N_47454,N_41601,N_44576);
and U47455 (N_47455,N_41418,N_44494);
or U47456 (N_47456,N_41733,N_42301);
nand U47457 (N_47457,N_42909,N_40792);
or U47458 (N_47458,N_42883,N_42798);
nor U47459 (N_47459,N_44781,N_42352);
and U47460 (N_47460,N_42222,N_42722);
or U47461 (N_47461,N_40047,N_40757);
nand U47462 (N_47462,N_43797,N_43812);
nand U47463 (N_47463,N_42954,N_41091);
and U47464 (N_47464,N_40388,N_42996);
nor U47465 (N_47465,N_44698,N_44236);
nor U47466 (N_47466,N_43358,N_44272);
or U47467 (N_47467,N_43235,N_43079);
or U47468 (N_47468,N_40880,N_43763);
or U47469 (N_47469,N_44937,N_44361);
xor U47470 (N_47470,N_42700,N_44681);
nor U47471 (N_47471,N_41055,N_44478);
or U47472 (N_47472,N_42280,N_44022);
xnor U47473 (N_47473,N_41532,N_42826);
xor U47474 (N_47474,N_43559,N_43126);
nand U47475 (N_47475,N_43210,N_44202);
nor U47476 (N_47476,N_43230,N_41879);
nand U47477 (N_47477,N_44870,N_40354);
xor U47478 (N_47478,N_40082,N_41571);
or U47479 (N_47479,N_44736,N_41575);
and U47480 (N_47480,N_42052,N_40154);
xor U47481 (N_47481,N_40423,N_43170);
or U47482 (N_47482,N_40071,N_44013);
and U47483 (N_47483,N_43636,N_44577);
or U47484 (N_47484,N_41549,N_42717);
nand U47485 (N_47485,N_41193,N_41107);
nand U47486 (N_47486,N_41452,N_40489);
nand U47487 (N_47487,N_44788,N_40330);
and U47488 (N_47488,N_42628,N_44972);
nand U47489 (N_47489,N_42613,N_40318);
or U47490 (N_47490,N_44853,N_41906);
nor U47491 (N_47491,N_43512,N_42400);
or U47492 (N_47492,N_41902,N_43936);
xnor U47493 (N_47493,N_42869,N_44441);
and U47494 (N_47494,N_44515,N_42502);
or U47495 (N_47495,N_40542,N_44979);
nor U47496 (N_47496,N_43042,N_41809);
or U47497 (N_47497,N_44529,N_43038);
nor U47498 (N_47498,N_40270,N_42818);
or U47499 (N_47499,N_44152,N_42594);
nor U47500 (N_47500,N_43081,N_41406);
or U47501 (N_47501,N_40067,N_40551);
nand U47502 (N_47502,N_41181,N_41425);
and U47503 (N_47503,N_42220,N_44419);
nand U47504 (N_47504,N_42788,N_44612);
and U47505 (N_47505,N_41874,N_41655);
or U47506 (N_47506,N_42278,N_40735);
nand U47507 (N_47507,N_42140,N_44567);
nor U47508 (N_47508,N_41045,N_42498);
nand U47509 (N_47509,N_41137,N_41675);
nor U47510 (N_47510,N_43035,N_40614);
nand U47511 (N_47511,N_41372,N_43346);
xnor U47512 (N_47512,N_42430,N_40589);
and U47513 (N_47513,N_44810,N_44942);
and U47514 (N_47514,N_41394,N_44508);
nand U47515 (N_47515,N_43072,N_42452);
and U47516 (N_47516,N_43749,N_43551);
nand U47517 (N_47517,N_40443,N_43598);
or U47518 (N_47518,N_41435,N_44099);
or U47519 (N_47519,N_44872,N_40394);
and U47520 (N_47520,N_44963,N_43189);
nor U47521 (N_47521,N_44099,N_44663);
nor U47522 (N_47522,N_41492,N_42073);
nor U47523 (N_47523,N_41192,N_42582);
nand U47524 (N_47524,N_42817,N_41453);
nor U47525 (N_47525,N_43052,N_42281);
xnor U47526 (N_47526,N_42131,N_41000);
or U47527 (N_47527,N_43394,N_41839);
nand U47528 (N_47528,N_41631,N_40127);
xnor U47529 (N_47529,N_44441,N_42881);
or U47530 (N_47530,N_43392,N_42908);
nor U47531 (N_47531,N_40403,N_42870);
xor U47532 (N_47532,N_41969,N_42672);
or U47533 (N_47533,N_41193,N_41190);
nand U47534 (N_47534,N_44682,N_43680);
and U47535 (N_47535,N_40808,N_40427);
nor U47536 (N_47536,N_41867,N_42641);
xor U47537 (N_47537,N_41808,N_43233);
nand U47538 (N_47538,N_43178,N_42193);
nor U47539 (N_47539,N_41271,N_40112);
or U47540 (N_47540,N_43680,N_41584);
nand U47541 (N_47541,N_44513,N_40849);
xor U47542 (N_47542,N_41892,N_44363);
nand U47543 (N_47543,N_44427,N_42193);
nor U47544 (N_47544,N_41512,N_42441);
xnor U47545 (N_47545,N_42526,N_43733);
nand U47546 (N_47546,N_40254,N_44767);
and U47547 (N_47547,N_43936,N_44293);
nand U47548 (N_47548,N_43203,N_44356);
xor U47549 (N_47549,N_40184,N_40907);
nand U47550 (N_47550,N_42821,N_43635);
nand U47551 (N_47551,N_43769,N_44418);
or U47552 (N_47552,N_40992,N_41412);
xor U47553 (N_47553,N_41741,N_41084);
nor U47554 (N_47554,N_42538,N_43833);
nand U47555 (N_47555,N_40674,N_41833);
and U47556 (N_47556,N_43503,N_43733);
or U47557 (N_47557,N_41188,N_43473);
and U47558 (N_47558,N_43885,N_40996);
or U47559 (N_47559,N_41416,N_43757);
and U47560 (N_47560,N_44791,N_43078);
and U47561 (N_47561,N_43478,N_43869);
nand U47562 (N_47562,N_41016,N_44118);
nor U47563 (N_47563,N_43968,N_43563);
nand U47564 (N_47564,N_44408,N_43149);
nand U47565 (N_47565,N_42403,N_40593);
nand U47566 (N_47566,N_42483,N_40920);
nor U47567 (N_47567,N_44565,N_41534);
and U47568 (N_47568,N_41664,N_43387);
nor U47569 (N_47569,N_44255,N_40809);
xor U47570 (N_47570,N_40678,N_43743);
nor U47571 (N_47571,N_40295,N_42369);
nand U47572 (N_47572,N_44740,N_41090);
xor U47573 (N_47573,N_44831,N_44200);
or U47574 (N_47574,N_42390,N_42715);
or U47575 (N_47575,N_42213,N_41426);
nand U47576 (N_47576,N_42456,N_44030);
nand U47577 (N_47577,N_43431,N_43179);
xnor U47578 (N_47578,N_42254,N_44074);
nand U47579 (N_47579,N_43929,N_42475);
and U47580 (N_47580,N_40978,N_43618);
xor U47581 (N_47581,N_44253,N_40663);
xor U47582 (N_47582,N_44402,N_44977);
or U47583 (N_47583,N_44167,N_44090);
nand U47584 (N_47584,N_40170,N_40110);
nand U47585 (N_47585,N_41810,N_43491);
nand U47586 (N_47586,N_41813,N_43520);
and U47587 (N_47587,N_42650,N_41314);
nand U47588 (N_47588,N_44360,N_44246);
and U47589 (N_47589,N_44260,N_41754);
and U47590 (N_47590,N_40385,N_43879);
xnor U47591 (N_47591,N_41429,N_40726);
or U47592 (N_47592,N_43456,N_42685);
nor U47593 (N_47593,N_40918,N_40455);
nand U47594 (N_47594,N_44822,N_40173);
nand U47595 (N_47595,N_41211,N_41176);
xor U47596 (N_47596,N_40984,N_41190);
or U47597 (N_47597,N_44731,N_41059);
nand U47598 (N_47598,N_44232,N_43515);
or U47599 (N_47599,N_40871,N_42888);
or U47600 (N_47600,N_44344,N_41157);
and U47601 (N_47601,N_44211,N_40397);
nor U47602 (N_47602,N_40627,N_43661);
nand U47603 (N_47603,N_43861,N_43882);
and U47604 (N_47604,N_43596,N_40790);
or U47605 (N_47605,N_40748,N_44769);
or U47606 (N_47606,N_41416,N_41629);
and U47607 (N_47607,N_43323,N_43884);
or U47608 (N_47608,N_41240,N_42382);
or U47609 (N_47609,N_42319,N_40565);
nor U47610 (N_47610,N_43869,N_40135);
or U47611 (N_47611,N_43302,N_43061);
or U47612 (N_47612,N_42435,N_42892);
nand U47613 (N_47613,N_43996,N_44554);
nand U47614 (N_47614,N_40390,N_43420);
and U47615 (N_47615,N_41201,N_44118);
nand U47616 (N_47616,N_41884,N_44449);
or U47617 (N_47617,N_42105,N_43281);
and U47618 (N_47618,N_40484,N_43106);
or U47619 (N_47619,N_41644,N_41067);
nor U47620 (N_47620,N_42749,N_42615);
nand U47621 (N_47621,N_43638,N_43788);
and U47622 (N_47622,N_43249,N_40803);
nand U47623 (N_47623,N_42629,N_41755);
xnor U47624 (N_47624,N_44079,N_42681);
or U47625 (N_47625,N_42165,N_44109);
and U47626 (N_47626,N_43423,N_40820);
nor U47627 (N_47627,N_43461,N_44544);
and U47628 (N_47628,N_42713,N_41844);
nand U47629 (N_47629,N_43077,N_43670);
and U47630 (N_47630,N_40059,N_44728);
nand U47631 (N_47631,N_41447,N_43219);
or U47632 (N_47632,N_43263,N_41423);
and U47633 (N_47633,N_43268,N_40112);
nor U47634 (N_47634,N_42800,N_40766);
or U47635 (N_47635,N_40926,N_43723);
or U47636 (N_47636,N_43948,N_42661);
xor U47637 (N_47637,N_44371,N_43719);
and U47638 (N_47638,N_43056,N_40379);
or U47639 (N_47639,N_40559,N_42070);
nand U47640 (N_47640,N_43224,N_42775);
nand U47641 (N_47641,N_40963,N_42926);
and U47642 (N_47642,N_44799,N_44195);
xor U47643 (N_47643,N_41297,N_43430);
and U47644 (N_47644,N_44556,N_43728);
and U47645 (N_47645,N_40154,N_40714);
or U47646 (N_47646,N_43325,N_43106);
nor U47647 (N_47647,N_42513,N_43533);
xnor U47648 (N_47648,N_44173,N_40202);
or U47649 (N_47649,N_41446,N_41984);
nor U47650 (N_47650,N_44517,N_44353);
xnor U47651 (N_47651,N_41647,N_43528);
and U47652 (N_47652,N_41342,N_44570);
and U47653 (N_47653,N_42005,N_44618);
or U47654 (N_47654,N_41665,N_42312);
and U47655 (N_47655,N_40858,N_43815);
nand U47656 (N_47656,N_43409,N_41318);
and U47657 (N_47657,N_44048,N_40504);
xor U47658 (N_47658,N_42088,N_42502);
and U47659 (N_47659,N_42874,N_43744);
and U47660 (N_47660,N_41266,N_41192);
nand U47661 (N_47661,N_41154,N_41248);
nand U47662 (N_47662,N_41987,N_40215);
nand U47663 (N_47663,N_42816,N_40132);
or U47664 (N_47664,N_40598,N_40488);
and U47665 (N_47665,N_41104,N_41992);
nor U47666 (N_47666,N_41232,N_44017);
or U47667 (N_47667,N_44806,N_44145);
and U47668 (N_47668,N_44539,N_42010);
xnor U47669 (N_47669,N_40817,N_41411);
or U47670 (N_47670,N_42294,N_40461);
and U47671 (N_47671,N_44207,N_42667);
nor U47672 (N_47672,N_43646,N_41420);
or U47673 (N_47673,N_42247,N_43547);
nand U47674 (N_47674,N_43049,N_43690);
or U47675 (N_47675,N_44420,N_43374);
and U47676 (N_47676,N_44786,N_43372);
xnor U47677 (N_47677,N_40793,N_40759);
xnor U47678 (N_47678,N_40331,N_43505);
or U47679 (N_47679,N_40423,N_44534);
or U47680 (N_47680,N_42625,N_42676);
nor U47681 (N_47681,N_41281,N_40936);
nor U47682 (N_47682,N_41368,N_41645);
nor U47683 (N_47683,N_43455,N_40641);
nor U47684 (N_47684,N_41421,N_43945);
nor U47685 (N_47685,N_40514,N_42192);
nor U47686 (N_47686,N_44805,N_44087);
xor U47687 (N_47687,N_42933,N_41586);
xnor U47688 (N_47688,N_42362,N_44275);
xor U47689 (N_47689,N_40648,N_43920);
and U47690 (N_47690,N_42481,N_42249);
nor U47691 (N_47691,N_42592,N_44914);
and U47692 (N_47692,N_42698,N_44583);
nand U47693 (N_47693,N_42533,N_43963);
nand U47694 (N_47694,N_42489,N_41991);
nor U47695 (N_47695,N_41751,N_43241);
or U47696 (N_47696,N_41124,N_43891);
or U47697 (N_47697,N_44839,N_40593);
or U47698 (N_47698,N_44356,N_44792);
nand U47699 (N_47699,N_44641,N_41126);
or U47700 (N_47700,N_44633,N_40228);
nand U47701 (N_47701,N_43954,N_43162);
nand U47702 (N_47702,N_41437,N_42963);
nor U47703 (N_47703,N_42752,N_42486);
nor U47704 (N_47704,N_44535,N_41805);
nor U47705 (N_47705,N_43940,N_43394);
or U47706 (N_47706,N_42994,N_44831);
nand U47707 (N_47707,N_43669,N_44553);
and U47708 (N_47708,N_43867,N_40094);
xnor U47709 (N_47709,N_44067,N_44058);
and U47710 (N_47710,N_41986,N_40082);
nor U47711 (N_47711,N_40036,N_43270);
nand U47712 (N_47712,N_43482,N_41429);
nor U47713 (N_47713,N_42825,N_41697);
nand U47714 (N_47714,N_43068,N_42396);
nor U47715 (N_47715,N_41585,N_43172);
nor U47716 (N_47716,N_43712,N_42544);
and U47717 (N_47717,N_44613,N_41091);
nor U47718 (N_47718,N_44214,N_44984);
nor U47719 (N_47719,N_41872,N_44894);
xnor U47720 (N_47720,N_40886,N_43694);
or U47721 (N_47721,N_41730,N_41017);
xnor U47722 (N_47722,N_42396,N_40432);
and U47723 (N_47723,N_41553,N_42653);
and U47724 (N_47724,N_42779,N_41183);
or U47725 (N_47725,N_43993,N_44228);
and U47726 (N_47726,N_44376,N_42682);
nor U47727 (N_47727,N_44716,N_41622);
nor U47728 (N_47728,N_44434,N_41774);
and U47729 (N_47729,N_40988,N_43197);
nand U47730 (N_47730,N_44865,N_42213);
and U47731 (N_47731,N_42320,N_44685);
nor U47732 (N_47732,N_43102,N_41367);
or U47733 (N_47733,N_43549,N_42506);
nand U47734 (N_47734,N_43350,N_43031);
nand U47735 (N_47735,N_41418,N_44346);
xor U47736 (N_47736,N_40001,N_41262);
or U47737 (N_47737,N_41123,N_42981);
or U47738 (N_47738,N_41486,N_42235);
nor U47739 (N_47739,N_40570,N_42094);
and U47740 (N_47740,N_40522,N_44779);
nor U47741 (N_47741,N_43194,N_41453);
nor U47742 (N_47742,N_41423,N_44955);
xor U47743 (N_47743,N_40363,N_42270);
nand U47744 (N_47744,N_42852,N_42871);
and U47745 (N_47745,N_42435,N_41653);
or U47746 (N_47746,N_43398,N_42254);
xor U47747 (N_47747,N_44506,N_40062);
or U47748 (N_47748,N_44031,N_41371);
nand U47749 (N_47749,N_42731,N_43420);
nor U47750 (N_47750,N_41377,N_40072);
nor U47751 (N_47751,N_42745,N_40472);
and U47752 (N_47752,N_42621,N_43547);
and U47753 (N_47753,N_42117,N_41701);
and U47754 (N_47754,N_44417,N_44905);
nand U47755 (N_47755,N_42127,N_40305);
nand U47756 (N_47756,N_41757,N_41247);
nor U47757 (N_47757,N_40299,N_42014);
nand U47758 (N_47758,N_43814,N_42825);
and U47759 (N_47759,N_44750,N_40614);
or U47760 (N_47760,N_40646,N_44634);
or U47761 (N_47761,N_44576,N_43407);
and U47762 (N_47762,N_44582,N_43617);
and U47763 (N_47763,N_42551,N_41613);
nor U47764 (N_47764,N_41273,N_40189);
or U47765 (N_47765,N_42206,N_41311);
or U47766 (N_47766,N_43169,N_42166);
nor U47767 (N_47767,N_44867,N_43418);
nor U47768 (N_47768,N_40081,N_44909);
nand U47769 (N_47769,N_43041,N_43911);
nand U47770 (N_47770,N_44977,N_44665);
and U47771 (N_47771,N_43507,N_42317);
nor U47772 (N_47772,N_40566,N_41509);
and U47773 (N_47773,N_41343,N_40822);
and U47774 (N_47774,N_42783,N_41363);
or U47775 (N_47775,N_44229,N_44896);
nor U47776 (N_47776,N_41638,N_41959);
nor U47777 (N_47777,N_44523,N_44896);
or U47778 (N_47778,N_42121,N_44179);
and U47779 (N_47779,N_40993,N_44607);
nand U47780 (N_47780,N_42266,N_40881);
nor U47781 (N_47781,N_42828,N_43472);
nor U47782 (N_47782,N_41723,N_43718);
nand U47783 (N_47783,N_40557,N_43248);
nor U47784 (N_47784,N_42395,N_42062);
nor U47785 (N_47785,N_44005,N_44427);
or U47786 (N_47786,N_43391,N_41444);
xor U47787 (N_47787,N_44295,N_44825);
nor U47788 (N_47788,N_44410,N_40295);
or U47789 (N_47789,N_41191,N_44885);
nor U47790 (N_47790,N_44437,N_44536);
and U47791 (N_47791,N_40857,N_40409);
nand U47792 (N_47792,N_40324,N_41286);
nor U47793 (N_47793,N_41108,N_44542);
nand U47794 (N_47794,N_43311,N_41352);
or U47795 (N_47795,N_42334,N_44974);
nor U47796 (N_47796,N_41842,N_42538);
nand U47797 (N_47797,N_44632,N_41933);
nand U47798 (N_47798,N_41881,N_41810);
or U47799 (N_47799,N_40579,N_41061);
or U47800 (N_47800,N_43285,N_43625);
or U47801 (N_47801,N_42177,N_41866);
xor U47802 (N_47802,N_40619,N_40699);
and U47803 (N_47803,N_41215,N_43862);
or U47804 (N_47804,N_40562,N_43793);
or U47805 (N_47805,N_41901,N_43832);
nor U47806 (N_47806,N_42291,N_44991);
nor U47807 (N_47807,N_43258,N_43168);
and U47808 (N_47808,N_44837,N_42691);
and U47809 (N_47809,N_43571,N_40337);
nand U47810 (N_47810,N_41339,N_42538);
or U47811 (N_47811,N_43537,N_42212);
and U47812 (N_47812,N_42608,N_40074);
and U47813 (N_47813,N_42534,N_43420);
nand U47814 (N_47814,N_44875,N_43640);
nand U47815 (N_47815,N_40636,N_44977);
nor U47816 (N_47816,N_41537,N_43712);
nor U47817 (N_47817,N_43599,N_40574);
or U47818 (N_47818,N_41915,N_44520);
and U47819 (N_47819,N_42183,N_44756);
nor U47820 (N_47820,N_42473,N_41912);
and U47821 (N_47821,N_42291,N_42829);
and U47822 (N_47822,N_44595,N_42703);
or U47823 (N_47823,N_44062,N_41125);
or U47824 (N_47824,N_42259,N_43418);
nor U47825 (N_47825,N_42093,N_42309);
or U47826 (N_47826,N_40636,N_44483);
nor U47827 (N_47827,N_44582,N_42568);
xor U47828 (N_47828,N_44493,N_44468);
and U47829 (N_47829,N_40320,N_43324);
nor U47830 (N_47830,N_43559,N_41598);
or U47831 (N_47831,N_41914,N_43081);
or U47832 (N_47832,N_40803,N_42379);
and U47833 (N_47833,N_41851,N_40385);
nand U47834 (N_47834,N_43402,N_43558);
or U47835 (N_47835,N_44169,N_41681);
xnor U47836 (N_47836,N_42603,N_40397);
or U47837 (N_47837,N_41793,N_43410);
and U47838 (N_47838,N_43447,N_44203);
and U47839 (N_47839,N_43246,N_42806);
nor U47840 (N_47840,N_44407,N_44600);
or U47841 (N_47841,N_41368,N_43323);
nor U47842 (N_47842,N_44965,N_44581);
and U47843 (N_47843,N_44341,N_44748);
and U47844 (N_47844,N_40134,N_44272);
or U47845 (N_47845,N_40127,N_40623);
nor U47846 (N_47846,N_40859,N_43603);
nand U47847 (N_47847,N_43809,N_41926);
or U47848 (N_47848,N_44416,N_40957);
nor U47849 (N_47849,N_44361,N_42120);
nand U47850 (N_47850,N_44871,N_42538);
nor U47851 (N_47851,N_44975,N_41993);
and U47852 (N_47852,N_44716,N_43166);
xnor U47853 (N_47853,N_44853,N_40326);
and U47854 (N_47854,N_40050,N_40404);
and U47855 (N_47855,N_44003,N_41637);
nor U47856 (N_47856,N_42921,N_41213);
nor U47857 (N_47857,N_40442,N_41241);
and U47858 (N_47858,N_42998,N_41319);
and U47859 (N_47859,N_40317,N_42058);
and U47860 (N_47860,N_43135,N_41671);
xor U47861 (N_47861,N_41255,N_44898);
or U47862 (N_47862,N_43164,N_43617);
or U47863 (N_47863,N_41112,N_42928);
or U47864 (N_47864,N_41630,N_43491);
xnor U47865 (N_47865,N_44724,N_41475);
nand U47866 (N_47866,N_41931,N_43612);
nor U47867 (N_47867,N_42410,N_41529);
or U47868 (N_47868,N_42864,N_41089);
nand U47869 (N_47869,N_44015,N_43943);
nor U47870 (N_47870,N_44396,N_42357);
and U47871 (N_47871,N_43897,N_42286);
or U47872 (N_47872,N_42791,N_40759);
nand U47873 (N_47873,N_44948,N_43496);
xnor U47874 (N_47874,N_41039,N_42192);
xor U47875 (N_47875,N_41073,N_41887);
and U47876 (N_47876,N_41274,N_40338);
or U47877 (N_47877,N_41602,N_43043);
nor U47878 (N_47878,N_41416,N_41880);
nand U47879 (N_47879,N_41953,N_40834);
xnor U47880 (N_47880,N_44055,N_43530);
nor U47881 (N_47881,N_40313,N_41669);
and U47882 (N_47882,N_41713,N_40804);
and U47883 (N_47883,N_44785,N_44523);
xnor U47884 (N_47884,N_40905,N_43840);
nand U47885 (N_47885,N_43639,N_42556);
xnor U47886 (N_47886,N_41329,N_44391);
and U47887 (N_47887,N_41714,N_41299);
or U47888 (N_47888,N_41055,N_41412);
and U47889 (N_47889,N_40685,N_43481);
nor U47890 (N_47890,N_43221,N_40123);
and U47891 (N_47891,N_40809,N_43027);
or U47892 (N_47892,N_44581,N_40990);
nand U47893 (N_47893,N_42595,N_44803);
and U47894 (N_47894,N_43952,N_43253);
or U47895 (N_47895,N_42682,N_40003);
xnor U47896 (N_47896,N_41612,N_44961);
or U47897 (N_47897,N_40947,N_42720);
and U47898 (N_47898,N_43801,N_41998);
or U47899 (N_47899,N_41471,N_44122);
nand U47900 (N_47900,N_40056,N_40877);
or U47901 (N_47901,N_44708,N_44786);
or U47902 (N_47902,N_44803,N_40563);
and U47903 (N_47903,N_41171,N_42694);
or U47904 (N_47904,N_40158,N_41601);
nor U47905 (N_47905,N_43381,N_44365);
and U47906 (N_47906,N_40955,N_40621);
or U47907 (N_47907,N_42919,N_42453);
or U47908 (N_47908,N_44512,N_41056);
nor U47909 (N_47909,N_41421,N_40170);
nor U47910 (N_47910,N_44024,N_40851);
nand U47911 (N_47911,N_42261,N_41032);
and U47912 (N_47912,N_44272,N_43553);
nand U47913 (N_47913,N_41637,N_40810);
nand U47914 (N_47914,N_41335,N_44461);
nand U47915 (N_47915,N_41908,N_43893);
or U47916 (N_47916,N_40603,N_40440);
or U47917 (N_47917,N_40637,N_42751);
xnor U47918 (N_47918,N_44622,N_43169);
xor U47919 (N_47919,N_44348,N_40771);
or U47920 (N_47920,N_41773,N_44636);
or U47921 (N_47921,N_43917,N_44008);
nand U47922 (N_47922,N_41685,N_40888);
nor U47923 (N_47923,N_42329,N_44634);
nor U47924 (N_47924,N_40380,N_44056);
and U47925 (N_47925,N_41143,N_41629);
nand U47926 (N_47926,N_42547,N_43469);
or U47927 (N_47927,N_41039,N_41971);
or U47928 (N_47928,N_40861,N_42109);
or U47929 (N_47929,N_43754,N_41084);
nor U47930 (N_47930,N_44863,N_42343);
nand U47931 (N_47931,N_40937,N_41402);
or U47932 (N_47932,N_41145,N_41500);
xnor U47933 (N_47933,N_40567,N_42780);
nor U47934 (N_47934,N_41829,N_43430);
and U47935 (N_47935,N_41804,N_42368);
or U47936 (N_47936,N_40554,N_43815);
and U47937 (N_47937,N_42059,N_43661);
nand U47938 (N_47938,N_43249,N_41907);
nor U47939 (N_47939,N_42351,N_40724);
xnor U47940 (N_47940,N_44361,N_42718);
and U47941 (N_47941,N_44819,N_41295);
nand U47942 (N_47942,N_41049,N_43995);
nand U47943 (N_47943,N_40596,N_40266);
nand U47944 (N_47944,N_42192,N_40107);
nand U47945 (N_47945,N_44680,N_41526);
or U47946 (N_47946,N_41973,N_43092);
and U47947 (N_47947,N_42874,N_42691);
nor U47948 (N_47948,N_40758,N_43442);
nor U47949 (N_47949,N_40361,N_44611);
and U47950 (N_47950,N_41795,N_41990);
xnor U47951 (N_47951,N_43008,N_44577);
and U47952 (N_47952,N_40399,N_44245);
or U47953 (N_47953,N_42567,N_43221);
or U47954 (N_47954,N_42791,N_40859);
or U47955 (N_47955,N_41689,N_40811);
and U47956 (N_47956,N_42240,N_41928);
nand U47957 (N_47957,N_41246,N_42144);
nand U47958 (N_47958,N_44833,N_40154);
or U47959 (N_47959,N_44822,N_42500);
nand U47960 (N_47960,N_40144,N_42347);
and U47961 (N_47961,N_42104,N_40864);
nand U47962 (N_47962,N_42433,N_41367);
nor U47963 (N_47963,N_41490,N_44533);
nor U47964 (N_47964,N_43124,N_41869);
or U47965 (N_47965,N_41655,N_43536);
nand U47966 (N_47966,N_41549,N_43082);
and U47967 (N_47967,N_44414,N_42032);
nor U47968 (N_47968,N_44061,N_43925);
nor U47969 (N_47969,N_42175,N_44887);
and U47970 (N_47970,N_42240,N_42192);
nand U47971 (N_47971,N_43401,N_44604);
nor U47972 (N_47972,N_40916,N_40234);
xor U47973 (N_47973,N_41749,N_44346);
nand U47974 (N_47974,N_41681,N_41321);
nand U47975 (N_47975,N_42348,N_43124);
nand U47976 (N_47976,N_41047,N_41988);
or U47977 (N_47977,N_44705,N_42823);
nand U47978 (N_47978,N_40204,N_44798);
xor U47979 (N_47979,N_43574,N_40098);
or U47980 (N_47980,N_42722,N_41450);
xor U47981 (N_47981,N_41694,N_44878);
nand U47982 (N_47982,N_43656,N_40452);
nor U47983 (N_47983,N_40833,N_40381);
xor U47984 (N_47984,N_42165,N_40498);
xnor U47985 (N_47985,N_43055,N_41750);
nor U47986 (N_47986,N_42228,N_43891);
and U47987 (N_47987,N_44639,N_43784);
or U47988 (N_47988,N_42608,N_40545);
or U47989 (N_47989,N_44077,N_42974);
or U47990 (N_47990,N_44434,N_43668);
or U47991 (N_47991,N_40930,N_41076);
and U47992 (N_47992,N_40747,N_40802);
or U47993 (N_47993,N_43748,N_44370);
or U47994 (N_47994,N_42868,N_40818);
nand U47995 (N_47995,N_43183,N_43669);
nor U47996 (N_47996,N_42364,N_41998);
or U47997 (N_47997,N_42402,N_42777);
xnor U47998 (N_47998,N_41692,N_43908);
nand U47999 (N_47999,N_44035,N_40637);
or U48000 (N_48000,N_44250,N_40682);
and U48001 (N_48001,N_42937,N_43376);
or U48002 (N_48002,N_43524,N_40451);
or U48003 (N_48003,N_44907,N_43480);
or U48004 (N_48004,N_43641,N_44751);
or U48005 (N_48005,N_41118,N_42215);
and U48006 (N_48006,N_44458,N_44623);
nor U48007 (N_48007,N_42086,N_44022);
and U48008 (N_48008,N_40891,N_40281);
xnor U48009 (N_48009,N_43634,N_42446);
nand U48010 (N_48010,N_43818,N_42468);
xor U48011 (N_48011,N_43016,N_43560);
nor U48012 (N_48012,N_42708,N_44870);
or U48013 (N_48013,N_44555,N_40415);
or U48014 (N_48014,N_43685,N_44608);
nor U48015 (N_48015,N_40625,N_41739);
nand U48016 (N_48016,N_43843,N_40226);
nand U48017 (N_48017,N_41231,N_43106);
and U48018 (N_48018,N_40323,N_41892);
and U48019 (N_48019,N_43520,N_40897);
and U48020 (N_48020,N_43486,N_44447);
and U48021 (N_48021,N_41875,N_44234);
and U48022 (N_48022,N_44053,N_44130);
or U48023 (N_48023,N_44093,N_41668);
xnor U48024 (N_48024,N_40846,N_44313);
nor U48025 (N_48025,N_42758,N_40271);
or U48026 (N_48026,N_43375,N_41405);
nand U48027 (N_48027,N_40078,N_41789);
or U48028 (N_48028,N_44502,N_40519);
nor U48029 (N_48029,N_41345,N_41450);
or U48030 (N_48030,N_42945,N_40536);
and U48031 (N_48031,N_43836,N_42692);
xor U48032 (N_48032,N_40874,N_41431);
and U48033 (N_48033,N_42552,N_42319);
or U48034 (N_48034,N_44510,N_43718);
and U48035 (N_48035,N_43946,N_43865);
nor U48036 (N_48036,N_41131,N_44244);
xor U48037 (N_48037,N_44713,N_42784);
nand U48038 (N_48038,N_42530,N_43656);
or U48039 (N_48039,N_40442,N_44920);
or U48040 (N_48040,N_44619,N_41934);
and U48041 (N_48041,N_43227,N_40016);
nor U48042 (N_48042,N_41553,N_42549);
xnor U48043 (N_48043,N_41428,N_42069);
nor U48044 (N_48044,N_44585,N_41593);
and U48045 (N_48045,N_44435,N_44857);
xor U48046 (N_48046,N_42012,N_42194);
and U48047 (N_48047,N_42167,N_42518);
nand U48048 (N_48048,N_42519,N_44963);
or U48049 (N_48049,N_43401,N_43610);
and U48050 (N_48050,N_41227,N_41081);
nand U48051 (N_48051,N_40060,N_42783);
and U48052 (N_48052,N_43819,N_40085);
xor U48053 (N_48053,N_43236,N_40083);
nor U48054 (N_48054,N_43269,N_44754);
nand U48055 (N_48055,N_42942,N_44975);
or U48056 (N_48056,N_44487,N_44733);
nor U48057 (N_48057,N_42188,N_42613);
and U48058 (N_48058,N_41345,N_41575);
nand U48059 (N_48059,N_40084,N_42751);
nand U48060 (N_48060,N_43107,N_42692);
nand U48061 (N_48061,N_42170,N_44575);
nor U48062 (N_48062,N_43926,N_42586);
nand U48063 (N_48063,N_43075,N_42860);
nand U48064 (N_48064,N_42226,N_42479);
or U48065 (N_48065,N_40592,N_42866);
and U48066 (N_48066,N_43552,N_44849);
nand U48067 (N_48067,N_41851,N_43468);
or U48068 (N_48068,N_41580,N_40320);
nor U48069 (N_48069,N_44472,N_40554);
nand U48070 (N_48070,N_42858,N_41747);
or U48071 (N_48071,N_40637,N_41043);
and U48072 (N_48072,N_43631,N_40879);
nand U48073 (N_48073,N_40974,N_43091);
nor U48074 (N_48074,N_44221,N_42622);
nand U48075 (N_48075,N_44861,N_42873);
nor U48076 (N_48076,N_44332,N_42515);
or U48077 (N_48077,N_43888,N_42909);
or U48078 (N_48078,N_42761,N_41639);
nor U48079 (N_48079,N_42012,N_44625);
nor U48080 (N_48080,N_44302,N_40662);
nor U48081 (N_48081,N_43765,N_42029);
nand U48082 (N_48082,N_42049,N_42435);
nor U48083 (N_48083,N_43888,N_41883);
nor U48084 (N_48084,N_42428,N_44224);
or U48085 (N_48085,N_40881,N_44094);
nand U48086 (N_48086,N_41405,N_41077);
nor U48087 (N_48087,N_43457,N_42850);
nor U48088 (N_48088,N_42586,N_42840);
nor U48089 (N_48089,N_43073,N_40013);
nor U48090 (N_48090,N_42630,N_43254);
and U48091 (N_48091,N_44772,N_41211);
or U48092 (N_48092,N_41192,N_42608);
xnor U48093 (N_48093,N_41422,N_42186);
nand U48094 (N_48094,N_43637,N_42623);
xnor U48095 (N_48095,N_44286,N_42053);
and U48096 (N_48096,N_44154,N_40028);
nand U48097 (N_48097,N_42344,N_40489);
and U48098 (N_48098,N_40737,N_40519);
or U48099 (N_48099,N_42628,N_44655);
and U48100 (N_48100,N_42297,N_41919);
or U48101 (N_48101,N_40336,N_44554);
nor U48102 (N_48102,N_41862,N_42927);
nand U48103 (N_48103,N_40075,N_40151);
nand U48104 (N_48104,N_41291,N_40519);
and U48105 (N_48105,N_41633,N_42865);
nand U48106 (N_48106,N_43005,N_40311);
nor U48107 (N_48107,N_43240,N_40160);
nand U48108 (N_48108,N_44306,N_42631);
or U48109 (N_48109,N_42086,N_43138);
nand U48110 (N_48110,N_43519,N_44163);
or U48111 (N_48111,N_41546,N_43444);
xor U48112 (N_48112,N_41443,N_40094);
nand U48113 (N_48113,N_44163,N_42988);
nor U48114 (N_48114,N_40075,N_43710);
nor U48115 (N_48115,N_42521,N_40266);
xor U48116 (N_48116,N_41056,N_42507);
nand U48117 (N_48117,N_44108,N_41908);
and U48118 (N_48118,N_40935,N_42437);
and U48119 (N_48119,N_42256,N_44843);
nor U48120 (N_48120,N_42988,N_42039);
and U48121 (N_48121,N_42138,N_42981);
or U48122 (N_48122,N_42872,N_44312);
nor U48123 (N_48123,N_43424,N_43775);
nand U48124 (N_48124,N_44752,N_40432);
nor U48125 (N_48125,N_42570,N_40049);
nand U48126 (N_48126,N_42738,N_40126);
or U48127 (N_48127,N_44723,N_40063);
xor U48128 (N_48128,N_41233,N_42567);
nor U48129 (N_48129,N_40650,N_43047);
and U48130 (N_48130,N_44387,N_42159);
or U48131 (N_48131,N_42060,N_41663);
nand U48132 (N_48132,N_40529,N_44768);
and U48133 (N_48133,N_43824,N_41843);
or U48134 (N_48134,N_41130,N_42021);
nor U48135 (N_48135,N_42103,N_44013);
or U48136 (N_48136,N_40573,N_40779);
and U48137 (N_48137,N_42596,N_42983);
nand U48138 (N_48138,N_44241,N_41813);
nand U48139 (N_48139,N_41482,N_41514);
and U48140 (N_48140,N_40162,N_44867);
or U48141 (N_48141,N_40890,N_42659);
xor U48142 (N_48142,N_43090,N_40246);
or U48143 (N_48143,N_41972,N_41716);
or U48144 (N_48144,N_40722,N_41579);
or U48145 (N_48145,N_44216,N_44089);
or U48146 (N_48146,N_40730,N_42809);
xnor U48147 (N_48147,N_40770,N_40565);
nand U48148 (N_48148,N_44968,N_40500);
and U48149 (N_48149,N_41607,N_44500);
or U48150 (N_48150,N_41052,N_44414);
nor U48151 (N_48151,N_41599,N_41862);
nand U48152 (N_48152,N_40503,N_40125);
nor U48153 (N_48153,N_42770,N_43300);
and U48154 (N_48154,N_41090,N_40505);
or U48155 (N_48155,N_42261,N_41962);
and U48156 (N_48156,N_44172,N_43994);
or U48157 (N_48157,N_44635,N_40907);
xor U48158 (N_48158,N_41539,N_42287);
xnor U48159 (N_48159,N_42211,N_42816);
nor U48160 (N_48160,N_40755,N_41142);
or U48161 (N_48161,N_40007,N_43812);
nor U48162 (N_48162,N_43203,N_40350);
and U48163 (N_48163,N_40157,N_43224);
xnor U48164 (N_48164,N_43891,N_40061);
nor U48165 (N_48165,N_40887,N_44244);
or U48166 (N_48166,N_41910,N_41402);
nand U48167 (N_48167,N_43777,N_43646);
nand U48168 (N_48168,N_42311,N_43678);
and U48169 (N_48169,N_43877,N_44318);
nand U48170 (N_48170,N_44000,N_44439);
and U48171 (N_48171,N_42330,N_44186);
nand U48172 (N_48172,N_44153,N_40244);
nor U48173 (N_48173,N_43882,N_44520);
and U48174 (N_48174,N_40559,N_42281);
nor U48175 (N_48175,N_43723,N_44930);
or U48176 (N_48176,N_40038,N_41726);
or U48177 (N_48177,N_42894,N_42497);
nand U48178 (N_48178,N_44461,N_43621);
or U48179 (N_48179,N_42455,N_42710);
nand U48180 (N_48180,N_43821,N_44685);
or U48181 (N_48181,N_44343,N_43604);
and U48182 (N_48182,N_44818,N_41711);
nor U48183 (N_48183,N_40363,N_43244);
nand U48184 (N_48184,N_44420,N_40811);
nor U48185 (N_48185,N_43751,N_42373);
nor U48186 (N_48186,N_43569,N_44780);
nor U48187 (N_48187,N_40602,N_43482);
or U48188 (N_48188,N_43704,N_41317);
nand U48189 (N_48189,N_42165,N_40733);
nand U48190 (N_48190,N_44755,N_43769);
nor U48191 (N_48191,N_42251,N_43715);
nand U48192 (N_48192,N_42777,N_43447);
nor U48193 (N_48193,N_40177,N_44830);
nor U48194 (N_48194,N_44825,N_42972);
and U48195 (N_48195,N_42380,N_44383);
nor U48196 (N_48196,N_42406,N_40151);
xor U48197 (N_48197,N_40560,N_42035);
nand U48198 (N_48198,N_40008,N_41422);
nand U48199 (N_48199,N_41465,N_43746);
nand U48200 (N_48200,N_40478,N_43280);
nor U48201 (N_48201,N_43511,N_43353);
or U48202 (N_48202,N_42598,N_43680);
nand U48203 (N_48203,N_43151,N_43274);
and U48204 (N_48204,N_42128,N_42471);
nor U48205 (N_48205,N_42065,N_44069);
and U48206 (N_48206,N_44807,N_42342);
nand U48207 (N_48207,N_42921,N_40345);
nor U48208 (N_48208,N_41890,N_44146);
nor U48209 (N_48209,N_41536,N_42161);
or U48210 (N_48210,N_43183,N_41071);
nand U48211 (N_48211,N_43986,N_41755);
and U48212 (N_48212,N_40500,N_41493);
nor U48213 (N_48213,N_40685,N_43007);
and U48214 (N_48214,N_40695,N_44150);
xor U48215 (N_48215,N_40572,N_43861);
nor U48216 (N_48216,N_43572,N_44354);
nor U48217 (N_48217,N_44732,N_43160);
nor U48218 (N_48218,N_41011,N_41004);
or U48219 (N_48219,N_42649,N_44432);
nand U48220 (N_48220,N_41928,N_44680);
nor U48221 (N_48221,N_41493,N_42159);
nor U48222 (N_48222,N_42475,N_42926);
or U48223 (N_48223,N_42554,N_44458);
or U48224 (N_48224,N_41844,N_42616);
nand U48225 (N_48225,N_41592,N_41104);
nand U48226 (N_48226,N_40415,N_41003);
nand U48227 (N_48227,N_42066,N_43575);
nor U48228 (N_48228,N_41891,N_40816);
nand U48229 (N_48229,N_40053,N_40650);
nor U48230 (N_48230,N_42454,N_43638);
nor U48231 (N_48231,N_42642,N_40594);
nand U48232 (N_48232,N_41219,N_42253);
nor U48233 (N_48233,N_43645,N_42086);
nand U48234 (N_48234,N_43326,N_43415);
or U48235 (N_48235,N_44195,N_42781);
nand U48236 (N_48236,N_41104,N_41771);
nor U48237 (N_48237,N_43574,N_41719);
nand U48238 (N_48238,N_40298,N_44025);
and U48239 (N_48239,N_43847,N_42293);
or U48240 (N_48240,N_43836,N_40237);
and U48241 (N_48241,N_41740,N_41530);
xor U48242 (N_48242,N_44092,N_41948);
and U48243 (N_48243,N_43878,N_43910);
nand U48244 (N_48244,N_42624,N_41914);
nand U48245 (N_48245,N_40383,N_41903);
nand U48246 (N_48246,N_41979,N_40285);
and U48247 (N_48247,N_42072,N_41477);
xnor U48248 (N_48248,N_41633,N_40461);
and U48249 (N_48249,N_43568,N_43873);
and U48250 (N_48250,N_41622,N_40733);
nand U48251 (N_48251,N_40519,N_44356);
nand U48252 (N_48252,N_44987,N_42411);
and U48253 (N_48253,N_42151,N_41586);
nand U48254 (N_48254,N_44308,N_40201);
and U48255 (N_48255,N_41581,N_40770);
or U48256 (N_48256,N_42914,N_44075);
nor U48257 (N_48257,N_40941,N_42055);
nand U48258 (N_48258,N_41420,N_44502);
nand U48259 (N_48259,N_43448,N_41362);
nor U48260 (N_48260,N_41441,N_43653);
xor U48261 (N_48261,N_40963,N_43232);
nor U48262 (N_48262,N_41775,N_41514);
and U48263 (N_48263,N_41925,N_43191);
and U48264 (N_48264,N_43769,N_42680);
nor U48265 (N_48265,N_44263,N_41876);
nand U48266 (N_48266,N_40333,N_44579);
nand U48267 (N_48267,N_40159,N_41961);
and U48268 (N_48268,N_42599,N_42274);
nor U48269 (N_48269,N_44677,N_44396);
nor U48270 (N_48270,N_40343,N_43338);
nand U48271 (N_48271,N_42231,N_43718);
nand U48272 (N_48272,N_42481,N_43310);
nand U48273 (N_48273,N_40534,N_42082);
or U48274 (N_48274,N_43479,N_41402);
and U48275 (N_48275,N_40120,N_40696);
nor U48276 (N_48276,N_44174,N_40301);
nor U48277 (N_48277,N_40779,N_42341);
nand U48278 (N_48278,N_40029,N_41666);
nand U48279 (N_48279,N_40496,N_42152);
or U48280 (N_48280,N_40253,N_40229);
nand U48281 (N_48281,N_44775,N_40307);
nor U48282 (N_48282,N_42183,N_43303);
nor U48283 (N_48283,N_43498,N_42607);
nor U48284 (N_48284,N_41361,N_41247);
xnor U48285 (N_48285,N_42175,N_41234);
nand U48286 (N_48286,N_41146,N_41332);
xor U48287 (N_48287,N_41635,N_43757);
or U48288 (N_48288,N_41522,N_42377);
and U48289 (N_48289,N_44416,N_41513);
nand U48290 (N_48290,N_43874,N_41328);
nor U48291 (N_48291,N_40619,N_43803);
and U48292 (N_48292,N_41610,N_41608);
or U48293 (N_48293,N_41622,N_43982);
xnor U48294 (N_48294,N_42896,N_41965);
xnor U48295 (N_48295,N_41831,N_43032);
or U48296 (N_48296,N_40454,N_44416);
or U48297 (N_48297,N_44541,N_40037);
nand U48298 (N_48298,N_40091,N_44106);
nand U48299 (N_48299,N_42959,N_41342);
nand U48300 (N_48300,N_42738,N_40807);
nor U48301 (N_48301,N_41533,N_40279);
and U48302 (N_48302,N_40320,N_43275);
nor U48303 (N_48303,N_42008,N_42649);
and U48304 (N_48304,N_40857,N_44511);
or U48305 (N_48305,N_43388,N_42934);
xnor U48306 (N_48306,N_43606,N_44565);
nor U48307 (N_48307,N_42438,N_42698);
nor U48308 (N_48308,N_40129,N_41854);
nand U48309 (N_48309,N_40002,N_44471);
nor U48310 (N_48310,N_41262,N_42949);
and U48311 (N_48311,N_40823,N_42200);
and U48312 (N_48312,N_42092,N_41074);
nand U48313 (N_48313,N_41206,N_44338);
nand U48314 (N_48314,N_42664,N_41797);
nand U48315 (N_48315,N_41305,N_44415);
and U48316 (N_48316,N_42451,N_40192);
nand U48317 (N_48317,N_44124,N_44770);
and U48318 (N_48318,N_43574,N_42955);
or U48319 (N_48319,N_43713,N_41612);
and U48320 (N_48320,N_40311,N_43329);
xnor U48321 (N_48321,N_43955,N_43666);
and U48322 (N_48322,N_40487,N_44156);
or U48323 (N_48323,N_41520,N_41178);
xor U48324 (N_48324,N_43167,N_41955);
xnor U48325 (N_48325,N_44903,N_41351);
and U48326 (N_48326,N_43699,N_44409);
nor U48327 (N_48327,N_42181,N_41927);
nor U48328 (N_48328,N_41964,N_41938);
and U48329 (N_48329,N_42075,N_44557);
or U48330 (N_48330,N_44501,N_43461);
nor U48331 (N_48331,N_43260,N_41534);
and U48332 (N_48332,N_44124,N_44298);
nand U48333 (N_48333,N_42259,N_40893);
nor U48334 (N_48334,N_40167,N_42485);
and U48335 (N_48335,N_43340,N_44929);
nor U48336 (N_48336,N_42306,N_41488);
nand U48337 (N_48337,N_40490,N_40103);
nand U48338 (N_48338,N_43268,N_44490);
nand U48339 (N_48339,N_43251,N_44833);
nor U48340 (N_48340,N_44671,N_41325);
or U48341 (N_48341,N_44114,N_43583);
nand U48342 (N_48342,N_41020,N_44231);
nor U48343 (N_48343,N_40563,N_40810);
nand U48344 (N_48344,N_43473,N_40330);
and U48345 (N_48345,N_40285,N_40442);
and U48346 (N_48346,N_40188,N_44019);
nor U48347 (N_48347,N_41843,N_42895);
nor U48348 (N_48348,N_41780,N_43128);
or U48349 (N_48349,N_40228,N_44536);
nor U48350 (N_48350,N_43586,N_42421);
nor U48351 (N_48351,N_42665,N_40667);
nor U48352 (N_48352,N_40518,N_44502);
and U48353 (N_48353,N_43541,N_43874);
nor U48354 (N_48354,N_43020,N_44167);
nor U48355 (N_48355,N_44435,N_43795);
nand U48356 (N_48356,N_44242,N_43862);
and U48357 (N_48357,N_44685,N_43980);
and U48358 (N_48358,N_43668,N_41837);
nor U48359 (N_48359,N_44910,N_41235);
nor U48360 (N_48360,N_41915,N_44053);
nor U48361 (N_48361,N_40950,N_43583);
nor U48362 (N_48362,N_42957,N_44583);
nand U48363 (N_48363,N_40331,N_41405);
nor U48364 (N_48364,N_41526,N_44373);
nor U48365 (N_48365,N_44738,N_42967);
nor U48366 (N_48366,N_43990,N_43539);
nor U48367 (N_48367,N_43485,N_40307);
nand U48368 (N_48368,N_42791,N_40391);
nand U48369 (N_48369,N_43928,N_44191);
nor U48370 (N_48370,N_43865,N_44498);
nor U48371 (N_48371,N_42787,N_44017);
nand U48372 (N_48372,N_41880,N_43800);
and U48373 (N_48373,N_42658,N_44002);
nor U48374 (N_48374,N_40237,N_42266);
xor U48375 (N_48375,N_42625,N_44027);
nor U48376 (N_48376,N_42975,N_42829);
and U48377 (N_48377,N_44690,N_42638);
nor U48378 (N_48378,N_40760,N_42481);
xor U48379 (N_48379,N_44242,N_41661);
and U48380 (N_48380,N_42281,N_43409);
nor U48381 (N_48381,N_40470,N_44530);
nand U48382 (N_48382,N_41378,N_40343);
xor U48383 (N_48383,N_41825,N_41456);
nand U48384 (N_48384,N_44960,N_42075);
xor U48385 (N_48385,N_41595,N_42787);
or U48386 (N_48386,N_44395,N_44452);
or U48387 (N_48387,N_40823,N_44972);
and U48388 (N_48388,N_41685,N_44336);
and U48389 (N_48389,N_43739,N_44819);
nand U48390 (N_48390,N_40026,N_43253);
nor U48391 (N_48391,N_41251,N_44610);
and U48392 (N_48392,N_43998,N_42776);
and U48393 (N_48393,N_40486,N_43614);
and U48394 (N_48394,N_40165,N_41623);
xnor U48395 (N_48395,N_44496,N_42394);
or U48396 (N_48396,N_40441,N_44610);
or U48397 (N_48397,N_44572,N_44988);
nand U48398 (N_48398,N_41219,N_41912);
xnor U48399 (N_48399,N_40221,N_41165);
or U48400 (N_48400,N_42158,N_44567);
and U48401 (N_48401,N_40965,N_40848);
nor U48402 (N_48402,N_41770,N_43511);
nand U48403 (N_48403,N_44250,N_44451);
or U48404 (N_48404,N_41781,N_40728);
or U48405 (N_48405,N_43462,N_42477);
or U48406 (N_48406,N_44577,N_41675);
xor U48407 (N_48407,N_40149,N_41345);
and U48408 (N_48408,N_42468,N_40991);
and U48409 (N_48409,N_40362,N_42758);
nand U48410 (N_48410,N_43959,N_41339);
nor U48411 (N_48411,N_40198,N_43398);
nand U48412 (N_48412,N_43793,N_40439);
or U48413 (N_48413,N_43136,N_41606);
xnor U48414 (N_48414,N_42642,N_42307);
and U48415 (N_48415,N_40074,N_44628);
nor U48416 (N_48416,N_44474,N_41876);
nor U48417 (N_48417,N_42380,N_42446);
nor U48418 (N_48418,N_41487,N_43351);
and U48419 (N_48419,N_44693,N_44140);
and U48420 (N_48420,N_43397,N_41090);
or U48421 (N_48421,N_42789,N_40188);
or U48422 (N_48422,N_41309,N_42895);
and U48423 (N_48423,N_41119,N_43781);
xor U48424 (N_48424,N_44346,N_43638);
or U48425 (N_48425,N_40568,N_42860);
and U48426 (N_48426,N_42147,N_41421);
nand U48427 (N_48427,N_41428,N_43112);
and U48428 (N_48428,N_44797,N_42790);
nor U48429 (N_48429,N_43935,N_42227);
nand U48430 (N_48430,N_44685,N_41122);
and U48431 (N_48431,N_42967,N_43619);
xor U48432 (N_48432,N_42811,N_43351);
xor U48433 (N_48433,N_44580,N_43080);
nor U48434 (N_48434,N_40563,N_42893);
or U48435 (N_48435,N_41346,N_41538);
nand U48436 (N_48436,N_42189,N_44357);
nor U48437 (N_48437,N_41588,N_44899);
nor U48438 (N_48438,N_40881,N_41594);
xnor U48439 (N_48439,N_42802,N_41614);
and U48440 (N_48440,N_44737,N_43106);
nand U48441 (N_48441,N_41651,N_44002);
nand U48442 (N_48442,N_43400,N_42154);
nor U48443 (N_48443,N_42905,N_40596);
or U48444 (N_48444,N_40652,N_41219);
nor U48445 (N_48445,N_43459,N_44598);
and U48446 (N_48446,N_44819,N_40163);
or U48447 (N_48447,N_44708,N_40649);
nor U48448 (N_48448,N_40201,N_42744);
or U48449 (N_48449,N_40543,N_43376);
and U48450 (N_48450,N_41042,N_44220);
nand U48451 (N_48451,N_41488,N_44477);
nor U48452 (N_48452,N_43020,N_43966);
nor U48453 (N_48453,N_42046,N_43485);
and U48454 (N_48454,N_42385,N_43241);
nand U48455 (N_48455,N_44976,N_43183);
nand U48456 (N_48456,N_40253,N_41299);
xnor U48457 (N_48457,N_40926,N_44864);
nand U48458 (N_48458,N_43841,N_43965);
and U48459 (N_48459,N_42731,N_43526);
nand U48460 (N_48460,N_41359,N_43442);
and U48461 (N_48461,N_40947,N_42002);
nand U48462 (N_48462,N_40532,N_43898);
xnor U48463 (N_48463,N_40920,N_40883);
nand U48464 (N_48464,N_43448,N_41257);
nand U48465 (N_48465,N_42481,N_42928);
nand U48466 (N_48466,N_41622,N_40804);
nand U48467 (N_48467,N_43197,N_41106);
and U48468 (N_48468,N_42646,N_40619);
and U48469 (N_48469,N_43589,N_42172);
and U48470 (N_48470,N_43223,N_42757);
and U48471 (N_48471,N_41099,N_43267);
or U48472 (N_48472,N_40272,N_41693);
nand U48473 (N_48473,N_43893,N_44119);
xor U48474 (N_48474,N_42405,N_44782);
or U48475 (N_48475,N_42546,N_43206);
nand U48476 (N_48476,N_40527,N_41379);
nand U48477 (N_48477,N_43439,N_42024);
nor U48478 (N_48478,N_40131,N_44995);
nor U48479 (N_48479,N_44238,N_40712);
nand U48480 (N_48480,N_41401,N_40871);
nor U48481 (N_48481,N_40361,N_41756);
and U48482 (N_48482,N_44966,N_40864);
and U48483 (N_48483,N_43137,N_43572);
and U48484 (N_48484,N_41206,N_44109);
or U48485 (N_48485,N_42233,N_41253);
or U48486 (N_48486,N_42779,N_44713);
or U48487 (N_48487,N_43044,N_40644);
or U48488 (N_48488,N_42572,N_42685);
nand U48489 (N_48489,N_42427,N_41381);
and U48490 (N_48490,N_40681,N_42282);
nand U48491 (N_48491,N_41383,N_41125);
nor U48492 (N_48492,N_43956,N_40265);
or U48493 (N_48493,N_44623,N_43507);
and U48494 (N_48494,N_42138,N_40851);
and U48495 (N_48495,N_42711,N_43149);
xor U48496 (N_48496,N_44967,N_43445);
or U48497 (N_48497,N_40169,N_44101);
nor U48498 (N_48498,N_41237,N_44792);
nor U48499 (N_48499,N_40329,N_44491);
or U48500 (N_48500,N_44654,N_40798);
nand U48501 (N_48501,N_44668,N_42373);
xor U48502 (N_48502,N_42873,N_44779);
nor U48503 (N_48503,N_41552,N_44182);
nor U48504 (N_48504,N_44001,N_43915);
and U48505 (N_48505,N_40953,N_40796);
nand U48506 (N_48506,N_40469,N_42327);
and U48507 (N_48507,N_40668,N_40190);
or U48508 (N_48508,N_41765,N_44979);
and U48509 (N_48509,N_41155,N_42604);
nor U48510 (N_48510,N_44577,N_42154);
nor U48511 (N_48511,N_41035,N_41867);
and U48512 (N_48512,N_41996,N_43127);
nor U48513 (N_48513,N_42241,N_41400);
nor U48514 (N_48514,N_42243,N_42858);
nor U48515 (N_48515,N_44829,N_43732);
and U48516 (N_48516,N_43010,N_42146);
nand U48517 (N_48517,N_40326,N_42466);
or U48518 (N_48518,N_43631,N_43266);
and U48519 (N_48519,N_40418,N_41411);
nor U48520 (N_48520,N_41544,N_42450);
nor U48521 (N_48521,N_44204,N_44621);
and U48522 (N_48522,N_43903,N_41263);
xnor U48523 (N_48523,N_41426,N_43317);
xnor U48524 (N_48524,N_42669,N_42080);
nor U48525 (N_48525,N_40523,N_42273);
and U48526 (N_48526,N_42662,N_44135);
xor U48527 (N_48527,N_43575,N_40813);
or U48528 (N_48528,N_42867,N_43257);
xnor U48529 (N_48529,N_44988,N_40820);
and U48530 (N_48530,N_44180,N_42215);
nor U48531 (N_48531,N_44973,N_44433);
or U48532 (N_48532,N_40656,N_41255);
and U48533 (N_48533,N_43874,N_43128);
nand U48534 (N_48534,N_41710,N_43336);
nor U48535 (N_48535,N_41752,N_43523);
and U48536 (N_48536,N_42576,N_41104);
or U48537 (N_48537,N_42230,N_43748);
nor U48538 (N_48538,N_41320,N_44659);
or U48539 (N_48539,N_40986,N_44752);
nand U48540 (N_48540,N_44330,N_40694);
nand U48541 (N_48541,N_42048,N_40079);
nand U48542 (N_48542,N_41318,N_42847);
nor U48543 (N_48543,N_40354,N_44562);
nor U48544 (N_48544,N_43209,N_42245);
nor U48545 (N_48545,N_42710,N_40121);
and U48546 (N_48546,N_41981,N_44590);
nor U48547 (N_48547,N_43039,N_43330);
nor U48548 (N_48548,N_41973,N_40259);
and U48549 (N_48549,N_42083,N_43531);
or U48550 (N_48550,N_41628,N_44955);
or U48551 (N_48551,N_43072,N_42644);
or U48552 (N_48552,N_44281,N_42472);
nand U48553 (N_48553,N_41549,N_44758);
nand U48554 (N_48554,N_41993,N_42303);
and U48555 (N_48555,N_44381,N_44419);
or U48556 (N_48556,N_44639,N_42304);
nand U48557 (N_48557,N_44155,N_43328);
nor U48558 (N_48558,N_42760,N_43690);
nor U48559 (N_48559,N_43348,N_40146);
and U48560 (N_48560,N_41995,N_41028);
and U48561 (N_48561,N_44395,N_42931);
xor U48562 (N_48562,N_40764,N_42340);
xnor U48563 (N_48563,N_44566,N_42351);
nor U48564 (N_48564,N_43138,N_43069);
and U48565 (N_48565,N_41947,N_44479);
and U48566 (N_48566,N_44267,N_44983);
and U48567 (N_48567,N_40221,N_43977);
or U48568 (N_48568,N_43731,N_44121);
nand U48569 (N_48569,N_44102,N_43732);
and U48570 (N_48570,N_40852,N_43847);
nand U48571 (N_48571,N_44473,N_44114);
or U48572 (N_48572,N_44830,N_44988);
nor U48573 (N_48573,N_44534,N_44991);
or U48574 (N_48574,N_41437,N_41972);
or U48575 (N_48575,N_43541,N_41597);
nand U48576 (N_48576,N_41351,N_44980);
and U48577 (N_48577,N_42750,N_42585);
xnor U48578 (N_48578,N_44523,N_43800);
and U48579 (N_48579,N_44716,N_41425);
xor U48580 (N_48580,N_44611,N_42268);
nor U48581 (N_48581,N_43216,N_42260);
and U48582 (N_48582,N_40951,N_41492);
nand U48583 (N_48583,N_44085,N_44775);
nor U48584 (N_48584,N_44146,N_41386);
or U48585 (N_48585,N_40564,N_42548);
nand U48586 (N_48586,N_40278,N_40976);
and U48587 (N_48587,N_44980,N_43741);
nor U48588 (N_48588,N_42172,N_43862);
nor U48589 (N_48589,N_40121,N_42461);
nand U48590 (N_48590,N_44303,N_43258);
or U48591 (N_48591,N_41691,N_40478);
nand U48592 (N_48592,N_44244,N_41603);
and U48593 (N_48593,N_43854,N_43564);
or U48594 (N_48594,N_43222,N_43819);
nor U48595 (N_48595,N_43239,N_43432);
or U48596 (N_48596,N_43448,N_42047);
or U48597 (N_48597,N_42553,N_42384);
nor U48598 (N_48598,N_42470,N_43903);
nor U48599 (N_48599,N_44310,N_41608);
and U48600 (N_48600,N_41306,N_42315);
and U48601 (N_48601,N_41736,N_40028);
nand U48602 (N_48602,N_41171,N_44391);
xor U48603 (N_48603,N_43133,N_43009);
nor U48604 (N_48604,N_40264,N_43509);
nand U48605 (N_48605,N_44742,N_40837);
or U48606 (N_48606,N_41760,N_44163);
or U48607 (N_48607,N_41528,N_43559);
nor U48608 (N_48608,N_40639,N_44009);
and U48609 (N_48609,N_40950,N_42879);
and U48610 (N_48610,N_43498,N_44373);
nand U48611 (N_48611,N_44710,N_41253);
nand U48612 (N_48612,N_43534,N_42878);
nor U48613 (N_48613,N_43336,N_43294);
nor U48614 (N_48614,N_44729,N_40607);
nand U48615 (N_48615,N_40055,N_44112);
nand U48616 (N_48616,N_40816,N_43770);
nand U48617 (N_48617,N_44322,N_40210);
or U48618 (N_48618,N_40958,N_41404);
nand U48619 (N_48619,N_41330,N_44151);
and U48620 (N_48620,N_42125,N_40593);
or U48621 (N_48621,N_40878,N_42657);
xnor U48622 (N_48622,N_43318,N_43290);
and U48623 (N_48623,N_41494,N_43118);
nand U48624 (N_48624,N_41198,N_42018);
and U48625 (N_48625,N_40386,N_43165);
nand U48626 (N_48626,N_42645,N_44323);
or U48627 (N_48627,N_41171,N_40197);
or U48628 (N_48628,N_44442,N_40396);
nor U48629 (N_48629,N_44503,N_44889);
nand U48630 (N_48630,N_40710,N_44972);
nor U48631 (N_48631,N_43822,N_41169);
or U48632 (N_48632,N_43153,N_41353);
nand U48633 (N_48633,N_41532,N_44987);
nor U48634 (N_48634,N_42876,N_42964);
xor U48635 (N_48635,N_42544,N_40546);
or U48636 (N_48636,N_41468,N_44712);
or U48637 (N_48637,N_41848,N_40304);
nand U48638 (N_48638,N_43726,N_44693);
nand U48639 (N_48639,N_40136,N_44602);
nand U48640 (N_48640,N_44131,N_42735);
nand U48641 (N_48641,N_44027,N_40446);
nor U48642 (N_48642,N_44234,N_43659);
or U48643 (N_48643,N_42804,N_44163);
nor U48644 (N_48644,N_42377,N_44358);
nor U48645 (N_48645,N_42774,N_44556);
and U48646 (N_48646,N_42277,N_43355);
nor U48647 (N_48647,N_42841,N_44168);
nor U48648 (N_48648,N_43872,N_41343);
nand U48649 (N_48649,N_42258,N_44300);
and U48650 (N_48650,N_41988,N_40696);
nand U48651 (N_48651,N_42801,N_44457);
and U48652 (N_48652,N_41750,N_44594);
nor U48653 (N_48653,N_43075,N_43306);
or U48654 (N_48654,N_44646,N_43072);
nor U48655 (N_48655,N_41812,N_41746);
or U48656 (N_48656,N_43114,N_41258);
nand U48657 (N_48657,N_42012,N_43681);
nor U48658 (N_48658,N_40143,N_41366);
nand U48659 (N_48659,N_40280,N_44200);
nor U48660 (N_48660,N_41493,N_42407);
nor U48661 (N_48661,N_42057,N_43166);
nand U48662 (N_48662,N_40829,N_44538);
xnor U48663 (N_48663,N_40460,N_42426);
nor U48664 (N_48664,N_42197,N_42291);
nor U48665 (N_48665,N_42060,N_40964);
nor U48666 (N_48666,N_41496,N_43289);
or U48667 (N_48667,N_42610,N_44308);
or U48668 (N_48668,N_43479,N_44352);
or U48669 (N_48669,N_43282,N_41624);
and U48670 (N_48670,N_43985,N_42090);
nand U48671 (N_48671,N_43242,N_42117);
nor U48672 (N_48672,N_40036,N_44060);
nand U48673 (N_48673,N_42168,N_44684);
xnor U48674 (N_48674,N_43585,N_43811);
and U48675 (N_48675,N_40436,N_40194);
nor U48676 (N_48676,N_43044,N_42828);
xor U48677 (N_48677,N_43763,N_43180);
nand U48678 (N_48678,N_41227,N_43240);
nand U48679 (N_48679,N_41337,N_42987);
nand U48680 (N_48680,N_41921,N_43647);
nand U48681 (N_48681,N_40218,N_43106);
and U48682 (N_48682,N_43177,N_40186);
or U48683 (N_48683,N_44583,N_41313);
or U48684 (N_48684,N_43931,N_44012);
or U48685 (N_48685,N_43005,N_41249);
nand U48686 (N_48686,N_43240,N_41845);
and U48687 (N_48687,N_41096,N_42817);
or U48688 (N_48688,N_40168,N_41183);
nand U48689 (N_48689,N_40044,N_43269);
nor U48690 (N_48690,N_40776,N_42858);
nor U48691 (N_48691,N_43053,N_44945);
nand U48692 (N_48692,N_40490,N_41753);
and U48693 (N_48693,N_40869,N_41855);
nor U48694 (N_48694,N_40745,N_41095);
nand U48695 (N_48695,N_43920,N_44072);
nor U48696 (N_48696,N_42149,N_44937);
nor U48697 (N_48697,N_44829,N_42507);
xnor U48698 (N_48698,N_44307,N_40792);
or U48699 (N_48699,N_44419,N_44052);
nand U48700 (N_48700,N_43832,N_43247);
and U48701 (N_48701,N_40600,N_44276);
nor U48702 (N_48702,N_44155,N_40939);
and U48703 (N_48703,N_42217,N_44608);
nand U48704 (N_48704,N_40505,N_40830);
and U48705 (N_48705,N_43179,N_44048);
nor U48706 (N_48706,N_41276,N_41571);
and U48707 (N_48707,N_43607,N_42144);
or U48708 (N_48708,N_42939,N_42537);
and U48709 (N_48709,N_40240,N_44657);
xnor U48710 (N_48710,N_43802,N_43382);
and U48711 (N_48711,N_42983,N_40382);
or U48712 (N_48712,N_42497,N_40530);
nand U48713 (N_48713,N_42186,N_43051);
nor U48714 (N_48714,N_42038,N_41526);
xnor U48715 (N_48715,N_40010,N_43106);
nand U48716 (N_48716,N_43681,N_42379);
or U48717 (N_48717,N_41896,N_43808);
nor U48718 (N_48718,N_40158,N_42899);
nor U48719 (N_48719,N_43641,N_40053);
nor U48720 (N_48720,N_42994,N_43268);
and U48721 (N_48721,N_42586,N_40434);
nand U48722 (N_48722,N_43069,N_42088);
nor U48723 (N_48723,N_40397,N_44744);
or U48724 (N_48724,N_44488,N_41418);
nor U48725 (N_48725,N_42927,N_40756);
and U48726 (N_48726,N_43348,N_43231);
xor U48727 (N_48727,N_43964,N_42759);
nor U48728 (N_48728,N_41496,N_43627);
nor U48729 (N_48729,N_44590,N_43295);
nor U48730 (N_48730,N_41657,N_40992);
or U48731 (N_48731,N_42904,N_42797);
and U48732 (N_48732,N_43153,N_40572);
xnor U48733 (N_48733,N_42609,N_42817);
and U48734 (N_48734,N_43616,N_40591);
or U48735 (N_48735,N_41196,N_42230);
and U48736 (N_48736,N_44926,N_44748);
or U48737 (N_48737,N_40542,N_40828);
nand U48738 (N_48738,N_41470,N_43338);
and U48739 (N_48739,N_43185,N_41737);
or U48740 (N_48740,N_41883,N_43031);
xnor U48741 (N_48741,N_41178,N_44857);
xnor U48742 (N_48742,N_40678,N_41766);
xor U48743 (N_48743,N_40942,N_42635);
and U48744 (N_48744,N_42156,N_43569);
or U48745 (N_48745,N_42629,N_42366);
nand U48746 (N_48746,N_42144,N_40792);
and U48747 (N_48747,N_44913,N_41044);
nor U48748 (N_48748,N_44313,N_41544);
and U48749 (N_48749,N_43362,N_43971);
or U48750 (N_48750,N_43023,N_41636);
or U48751 (N_48751,N_44003,N_42731);
nor U48752 (N_48752,N_41773,N_43842);
or U48753 (N_48753,N_44123,N_41807);
xnor U48754 (N_48754,N_43625,N_40517);
or U48755 (N_48755,N_40938,N_43695);
nand U48756 (N_48756,N_44985,N_41039);
nand U48757 (N_48757,N_40603,N_43260);
xnor U48758 (N_48758,N_44605,N_44024);
or U48759 (N_48759,N_44288,N_42137);
and U48760 (N_48760,N_41746,N_44139);
and U48761 (N_48761,N_44802,N_40898);
nor U48762 (N_48762,N_43857,N_41562);
nand U48763 (N_48763,N_42925,N_44584);
and U48764 (N_48764,N_40789,N_43215);
and U48765 (N_48765,N_43744,N_43024);
or U48766 (N_48766,N_44411,N_41546);
nor U48767 (N_48767,N_43449,N_44043);
nand U48768 (N_48768,N_41514,N_44941);
or U48769 (N_48769,N_41215,N_44460);
or U48770 (N_48770,N_40287,N_44521);
and U48771 (N_48771,N_40967,N_42298);
xnor U48772 (N_48772,N_44158,N_41506);
nor U48773 (N_48773,N_41658,N_44517);
or U48774 (N_48774,N_41757,N_41455);
nand U48775 (N_48775,N_44780,N_41346);
nand U48776 (N_48776,N_40390,N_40648);
or U48777 (N_48777,N_44591,N_43516);
or U48778 (N_48778,N_42223,N_44501);
nand U48779 (N_48779,N_42636,N_41174);
nor U48780 (N_48780,N_42301,N_43625);
and U48781 (N_48781,N_42020,N_44757);
or U48782 (N_48782,N_41326,N_41138);
or U48783 (N_48783,N_40465,N_40292);
nor U48784 (N_48784,N_42031,N_41203);
and U48785 (N_48785,N_42021,N_41746);
nor U48786 (N_48786,N_41246,N_44496);
nand U48787 (N_48787,N_41041,N_40525);
and U48788 (N_48788,N_44262,N_44815);
nand U48789 (N_48789,N_42982,N_44954);
nor U48790 (N_48790,N_41863,N_43421);
nor U48791 (N_48791,N_40672,N_41811);
and U48792 (N_48792,N_40764,N_40405);
nor U48793 (N_48793,N_40812,N_41198);
or U48794 (N_48794,N_42788,N_42032);
nand U48795 (N_48795,N_40493,N_44515);
or U48796 (N_48796,N_44524,N_41353);
nor U48797 (N_48797,N_40900,N_40439);
nand U48798 (N_48798,N_44733,N_41258);
nand U48799 (N_48799,N_40874,N_44941);
and U48800 (N_48800,N_44297,N_40164);
or U48801 (N_48801,N_42167,N_40689);
and U48802 (N_48802,N_41839,N_42210);
nor U48803 (N_48803,N_41206,N_42300);
xor U48804 (N_48804,N_43938,N_42185);
nor U48805 (N_48805,N_41711,N_43786);
and U48806 (N_48806,N_42878,N_43805);
nand U48807 (N_48807,N_42808,N_42326);
and U48808 (N_48808,N_40753,N_42800);
xnor U48809 (N_48809,N_40509,N_41886);
and U48810 (N_48810,N_44690,N_43693);
xnor U48811 (N_48811,N_40284,N_44216);
or U48812 (N_48812,N_43923,N_44408);
and U48813 (N_48813,N_41754,N_43558);
or U48814 (N_48814,N_40535,N_40035);
or U48815 (N_48815,N_43595,N_40792);
xnor U48816 (N_48816,N_44060,N_42138);
and U48817 (N_48817,N_43478,N_44694);
or U48818 (N_48818,N_43939,N_41930);
or U48819 (N_48819,N_41659,N_43943);
and U48820 (N_48820,N_41813,N_40427);
nand U48821 (N_48821,N_40305,N_42241);
and U48822 (N_48822,N_44842,N_43748);
xnor U48823 (N_48823,N_43666,N_40279);
and U48824 (N_48824,N_43332,N_43161);
xnor U48825 (N_48825,N_44486,N_40314);
nand U48826 (N_48826,N_43182,N_42938);
nand U48827 (N_48827,N_42255,N_41306);
nand U48828 (N_48828,N_42494,N_43720);
xnor U48829 (N_48829,N_40599,N_42403);
and U48830 (N_48830,N_44024,N_44198);
nand U48831 (N_48831,N_42408,N_42050);
nor U48832 (N_48832,N_42060,N_40720);
nor U48833 (N_48833,N_44765,N_42303);
and U48834 (N_48834,N_44979,N_41437);
or U48835 (N_48835,N_41098,N_44420);
or U48836 (N_48836,N_43254,N_42208);
and U48837 (N_48837,N_43560,N_40862);
and U48838 (N_48838,N_44421,N_41569);
and U48839 (N_48839,N_40871,N_40611);
nand U48840 (N_48840,N_41706,N_42400);
or U48841 (N_48841,N_44984,N_40090);
nor U48842 (N_48842,N_40095,N_43270);
or U48843 (N_48843,N_40648,N_44957);
or U48844 (N_48844,N_44162,N_43005);
nand U48845 (N_48845,N_42189,N_41412);
nand U48846 (N_48846,N_40454,N_43483);
or U48847 (N_48847,N_44164,N_41099);
and U48848 (N_48848,N_41439,N_43542);
and U48849 (N_48849,N_44669,N_42674);
nor U48850 (N_48850,N_42808,N_43269);
nand U48851 (N_48851,N_43184,N_41194);
or U48852 (N_48852,N_43333,N_42342);
or U48853 (N_48853,N_41892,N_43732);
and U48854 (N_48854,N_40955,N_42960);
nand U48855 (N_48855,N_43736,N_44847);
or U48856 (N_48856,N_42489,N_44267);
xor U48857 (N_48857,N_41566,N_41977);
xor U48858 (N_48858,N_40362,N_44491);
nor U48859 (N_48859,N_41791,N_40995);
xor U48860 (N_48860,N_44594,N_41551);
or U48861 (N_48861,N_43510,N_41779);
and U48862 (N_48862,N_42766,N_41269);
nor U48863 (N_48863,N_41011,N_41052);
and U48864 (N_48864,N_41027,N_43774);
or U48865 (N_48865,N_40136,N_42622);
or U48866 (N_48866,N_43295,N_42615);
nand U48867 (N_48867,N_42844,N_44621);
and U48868 (N_48868,N_41637,N_44390);
nor U48869 (N_48869,N_40935,N_42808);
nor U48870 (N_48870,N_44195,N_40848);
nor U48871 (N_48871,N_43308,N_41231);
nand U48872 (N_48872,N_41548,N_43658);
xnor U48873 (N_48873,N_43022,N_41314);
and U48874 (N_48874,N_40821,N_41847);
or U48875 (N_48875,N_43939,N_42705);
nand U48876 (N_48876,N_40800,N_40123);
xnor U48877 (N_48877,N_40959,N_40898);
or U48878 (N_48878,N_40595,N_41236);
and U48879 (N_48879,N_43877,N_43514);
nand U48880 (N_48880,N_40634,N_44298);
and U48881 (N_48881,N_43892,N_40595);
nand U48882 (N_48882,N_43250,N_43486);
or U48883 (N_48883,N_43540,N_44651);
and U48884 (N_48884,N_43184,N_42821);
nand U48885 (N_48885,N_40425,N_43257);
nand U48886 (N_48886,N_40704,N_42826);
nand U48887 (N_48887,N_44478,N_44903);
and U48888 (N_48888,N_40628,N_42859);
nor U48889 (N_48889,N_41448,N_43637);
or U48890 (N_48890,N_44861,N_40363);
and U48891 (N_48891,N_41425,N_40957);
or U48892 (N_48892,N_42465,N_41961);
nor U48893 (N_48893,N_42425,N_44367);
and U48894 (N_48894,N_44755,N_44715);
nand U48895 (N_48895,N_42741,N_42960);
nand U48896 (N_48896,N_43558,N_43524);
nand U48897 (N_48897,N_42463,N_43428);
nand U48898 (N_48898,N_41351,N_42552);
nand U48899 (N_48899,N_41865,N_40913);
and U48900 (N_48900,N_43178,N_41805);
nand U48901 (N_48901,N_42050,N_44364);
or U48902 (N_48902,N_40281,N_44096);
and U48903 (N_48903,N_43702,N_40823);
or U48904 (N_48904,N_40908,N_42301);
and U48905 (N_48905,N_40901,N_42118);
nor U48906 (N_48906,N_40217,N_44324);
or U48907 (N_48907,N_40525,N_42159);
or U48908 (N_48908,N_42814,N_44187);
nand U48909 (N_48909,N_43655,N_40879);
nor U48910 (N_48910,N_44543,N_43331);
or U48911 (N_48911,N_40697,N_41421);
or U48912 (N_48912,N_44331,N_41184);
nor U48913 (N_48913,N_44163,N_42458);
and U48914 (N_48914,N_41655,N_40186);
or U48915 (N_48915,N_40612,N_43827);
nand U48916 (N_48916,N_44119,N_40005);
nor U48917 (N_48917,N_40825,N_43642);
nor U48918 (N_48918,N_41167,N_41879);
nand U48919 (N_48919,N_40265,N_40655);
nor U48920 (N_48920,N_43006,N_41287);
and U48921 (N_48921,N_43035,N_42080);
nor U48922 (N_48922,N_42049,N_40695);
xnor U48923 (N_48923,N_44868,N_43284);
nor U48924 (N_48924,N_43929,N_41624);
nand U48925 (N_48925,N_42339,N_43082);
or U48926 (N_48926,N_43108,N_40795);
or U48927 (N_48927,N_41878,N_42160);
or U48928 (N_48928,N_40616,N_41966);
nand U48929 (N_48929,N_44829,N_43720);
and U48930 (N_48930,N_43928,N_40396);
nor U48931 (N_48931,N_40690,N_42028);
or U48932 (N_48932,N_42713,N_41702);
and U48933 (N_48933,N_41056,N_42526);
nand U48934 (N_48934,N_44329,N_40988);
nand U48935 (N_48935,N_42059,N_44746);
nor U48936 (N_48936,N_41112,N_40928);
nand U48937 (N_48937,N_42599,N_44427);
and U48938 (N_48938,N_44480,N_42149);
nand U48939 (N_48939,N_40753,N_42677);
nor U48940 (N_48940,N_44177,N_43383);
nand U48941 (N_48941,N_44823,N_42560);
nor U48942 (N_48942,N_42998,N_41867);
or U48943 (N_48943,N_40715,N_44439);
nor U48944 (N_48944,N_42436,N_40526);
and U48945 (N_48945,N_44298,N_40922);
nor U48946 (N_48946,N_41239,N_43405);
nor U48947 (N_48947,N_41624,N_44038);
and U48948 (N_48948,N_40213,N_40393);
nand U48949 (N_48949,N_41610,N_44293);
xnor U48950 (N_48950,N_44412,N_44090);
nor U48951 (N_48951,N_41473,N_42944);
nand U48952 (N_48952,N_44661,N_41055);
and U48953 (N_48953,N_43002,N_40462);
nand U48954 (N_48954,N_43755,N_42067);
xnor U48955 (N_48955,N_40641,N_41414);
nand U48956 (N_48956,N_41008,N_43265);
nand U48957 (N_48957,N_40146,N_43524);
nor U48958 (N_48958,N_44482,N_42078);
nand U48959 (N_48959,N_42171,N_41518);
and U48960 (N_48960,N_41785,N_40381);
or U48961 (N_48961,N_44585,N_43369);
and U48962 (N_48962,N_42613,N_43862);
nand U48963 (N_48963,N_42440,N_40918);
or U48964 (N_48964,N_40825,N_44145);
nand U48965 (N_48965,N_43825,N_40919);
nand U48966 (N_48966,N_43765,N_44121);
or U48967 (N_48967,N_44354,N_42874);
nand U48968 (N_48968,N_42411,N_40898);
nand U48969 (N_48969,N_41804,N_42453);
nand U48970 (N_48970,N_43207,N_42543);
and U48971 (N_48971,N_42830,N_41861);
or U48972 (N_48972,N_40093,N_43583);
nand U48973 (N_48973,N_41308,N_40994);
or U48974 (N_48974,N_44456,N_44352);
nand U48975 (N_48975,N_44193,N_44860);
and U48976 (N_48976,N_44163,N_43253);
nor U48977 (N_48977,N_40719,N_40431);
nor U48978 (N_48978,N_42496,N_41379);
and U48979 (N_48979,N_40107,N_40782);
or U48980 (N_48980,N_41205,N_44598);
nand U48981 (N_48981,N_41553,N_43817);
nand U48982 (N_48982,N_40216,N_44153);
xnor U48983 (N_48983,N_42949,N_41225);
and U48984 (N_48984,N_44942,N_42438);
nor U48985 (N_48985,N_41487,N_40584);
or U48986 (N_48986,N_40891,N_42983);
nor U48987 (N_48987,N_44278,N_41956);
nand U48988 (N_48988,N_42794,N_44775);
nand U48989 (N_48989,N_42317,N_40506);
nand U48990 (N_48990,N_43445,N_42646);
nand U48991 (N_48991,N_42787,N_43520);
nor U48992 (N_48992,N_41627,N_42755);
nor U48993 (N_48993,N_41050,N_41730);
or U48994 (N_48994,N_44797,N_42715);
nor U48995 (N_48995,N_43562,N_43337);
xnor U48996 (N_48996,N_40906,N_41943);
and U48997 (N_48997,N_44249,N_43041);
and U48998 (N_48998,N_44752,N_41027);
and U48999 (N_48999,N_41732,N_40400);
or U49000 (N_49000,N_42159,N_44068);
nand U49001 (N_49001,N_43246,N_43015);
nor U49002 (N_49002,N_40000,N_44312);
nor U49003 (N_49003,N_40104,N_40111);
nor U49004 (N_49004,N_42870,N_43373);
and U49005 (N_49005,N_41423,N_42142);
nor U49006 (N_49006,N_44980,N_42518);
nor U49007 (N_49007,N_41227,N_43668);
and U49008 (N_49008,N_40727,N_40784);
nand U49009 (N_49009,N_44693,N_40404);
and U49010 (N_49010,N_41001,N_43340);
or U49011 (N_49011,N_43357,N_43444);
and U49012 (N_49012,N_41231,N_40125);
or U49013 (N_49013,N_41031,N_44351);
nor U49014 (N_49014,N_44628,N_41426);
nand U49015 (N_49015,N_44959,N_44627);
or U49016 (N_49016,N_41146,N_41852);
nor U49017 (N_49017,N_41645,N_42976);
or U49018 (N_49018,N_40578,N_44918);
xnor U49019 (N_49019,N_43660,N_42685);
and U49020 (N_49020,N_43455,N_44786);
nor U49021 (N_49021,N_42950,N_40662);
or U49022 (N_49022,N_41649,N_42530);
nor U49023 (N_49023,N_40087,N_43706);
nand U49024 (N_49024,N_44512,N_44654);
and U49025 (N_49025,N_40732,N_43449);
nor U49026 (N_49026,N_42551,N_43322);
or U49027 (N_49027,N_40558,N_41419);
nand U49028 (N_49028,N_41338,N_41482);
and U49029 (N_49029,N_41103,N_40734);
or U49030 (N_49030,N_40017,N_42964);
or U49031 (N_49031,N_42430,N_44055);
or U49032 (N_49032,N_44609,N_42339);
and U49033 (N_49033,N_43263,N_42671);
nor U49034 (N_49034,N_43553,N_43236);
nor U49035 (N_49035,N_40096,N_40023);
nand U49036 (N_49036,N_42986,N_44624);
and U49037 (N_49037,N_41515,N_40501);
nor U49038 (N_49038,N_44068,N_41640);
and U49039 (N_49039,N_44975,N_41568);
nor U49040 (N_49040,N_40453,N_44478);
nand U49041 (N_49041,N_42754,N_41832);
xor U49042 (N_49042,N_43430,N_40627);
nand U49043 (N_49043,N_40412,N_41513);
nand U49044 (N_49044,N_42897,N_44395);
nor U49045 (N_49045,N_43668,N_44980);
and U49046 (N_49046,N_40075,N_44441);
nor U49047 (N_49047,N_40824,N_42488);
or U49048 (N_49048,N_43904,N_40464);
nor U49049 (N_49049,N_43754,N_40115);
and U49050 (N_49050,N_41844,N_40982);
nand U49051 (N_49051,N_40147,N_44682);
or U49052 (N_49052,N_43223,N_42617);
xor U49053 (N_49053,N_42541,N_44103);
nand U49054 (N_49054,N_41121,N_41649);
or U49055 (N_49055,N_41726,N_41217);
or U49056 (N_49056,N_42579,N_44705);
and U49057 (N_49057,N_40798,N_43148);
nor U49058 (N_49058,N_43401,N_40109);
nand U49059 (N_49059,N_43736,N_41939);
and U49060 (N_49060,N_43433,N_43469);
nand U49061 (N_49061,N_40958,N_44959);
nor U49062 (N_49062,N_42856,N_44215);
xnor U49063 (N_49063,N_42660,N_41391);
nand U49064 (N_49064,N_44905,N_43890);
xor U49065 (N_49065,N_42120,N_42524);
nand U49066 (N_49066,N_44557,N_44765);
and U49067 (N_49067,N_40797,N_44064);
xnor U49068 (N_49068,N_43866,N_40516);
xor U49069 (N_49069,N_40837,N_40023);
xor U49070 (N_49070,N_41080,N_42529);
nor U49071 (N_49071,N_43167,N_44708);
xnor U49072 (N_49072,N_44466,N_42061);
and U49073 (N_49073,N_43895,N_41583);
or U49074 (N_49074,N_40769,N_42296);
or U49075 (N_49075,N_41588,N_42229);
xor U49076 (N_49076,N_42791,N_42209);
nand U49077 (N_49077,N_43141,N_42007);
nor U49078 (N_49078,N_44727,N_43188);
nand U49079 (N_49079,N_42583,N_44572);
nor U49080 (N_49080,N_40590,N_42335);
or U49081 (N_49081,N_44883,N_41954);
and U49082 (N_49082,N_41865,N_41417);
nand U49083 (N_49083,N_42206,N_43967);
nand U49084 (N_49084,N_40301,N_43302);
nor U49085 (N_49085,N_42750,N_40329);
nor U49086 (N_49086,N_40370,N_41884);
or U49087 (N_49087,N_43939,N_40606);
xnor U49088 (N_49088,N_41256,N_43976);
xor U49089 (N_49089,N_43096,N_40559);
or U49090 (N_49090,N_42283,N_44048);
or U49091 (N_49091,N_42859,N_44566);
nand U49092 (N_49092,N_43855,N_42747);
and U49093 (N_49093,N_44281,N_43171);
nand U49094 (N_49094,N_43242,N_43249);
nor U49095 (N_49095,N_42160,N_42817);
or U49096 (N_49096,N_41912,N_42914);
and U49097 (N_49097,N_43159,N_42213);
or U49098 (N_49098,N_41291,N_41582);
or U49099 (N_49099,N_43988,N_41209);
and U49100 (N_49100,N_41020,N_40980);
nand U49101 (N_49101,N_42060,N_43043);
xnor U49102 (N_49102,N_43059,N_44476);
or U49103 (N_49103,N_43849,N_40670);
and U49104 (N_49104,N_43960,N_41944);
nand U49105 (N_49105,N_44613,N_40156);
xnor U49106 (N_49106,N_42713,N_41287);
nand U49107 (N_49107,N_43703,N_42690);
nor U49108 (N_49108,N_42326,N_40139);
nor U49109 (N_49109,N_41033,N_43848);
or U49110 (N_49110,N_42054,N_43837);
or U49111 (N_49111,N_42734,N_42887);
or U49112 (N_49112,N_43561,N_40136);
and U49113 (N_49113,N_42525,N_42727);
nor U49114 (N_49114,N_44046,N_40647);
and U49115 (N_49115,N_43333,N_42244);
xor U49116 (N_49116,N_40165,N_40161);
nor U49117 (N_49117,N_43674,N_40443);
nor U49118 (N_49118,N_42835,N_41545);
and U49119 (N_49119,N_42212,N_44163);
xor U49120 (N_49120,N_42754,N_41152);
xor U49121 (N_49121,N_44893,N_44542);
and U49122 (N_49122,N_43085,N_40332);
or U49123 (N_49123,N_42924,N_42336);
nor U49124 (N_49124,N_42212,N_43601);
nor U49125 (N_49125,N_44834,N_44530);
nand U49126 (N_49126,N_42864,N_43749);
nand U49127 (N_49127,N_41534,N_41980);
or U49128 (N_49128,N_40461,N_41592);
or U49129 (N_49129,N_44816,N_44516);
and U49130 (N_49130,N_41155,N_40057);
and U49131 (N_49131,N_42347,N_44839);
and U49132 (N_49132,N_42658,N_43960);
and U49133 (N_49133,N_42757,N_43230);
nor U49134 (N_49134,N_43843,N_41346);
and U49135 (N_49135,N_42817,N_41299);
nand U49136 (N_49136,N_40291,N_40683);
nand U49137 (N_49137,N_42506,N_44530);
and U49138 (N_49138,N_42050,N_43794);
or U49139 (N_49139,N_44310,N_41724);
or U49140 (N_49140,N_44816,N_42701);
nor U49141 (N_49141,N_43876,N_43825);
and U49142 (N_49142,N_42393,N_40999);
and U49143 (N_49143,N_43270,N_42092);
nor U49144 (N_49144,N_43805,N_40541);
and U49145 (N_49145,N_44684,N_42843);
or U49146 (N_49146,N_40752,N_43642);
nor U49147 (N_49147,N_43966,N_44798);
xnor U49148 (N_49148,N_42687,N_44812);
and U49149 (N_49149,N_40720,N_44717);
nor U49150 (N_49150,N_42972,N_42481);
and U49151 (N_49151,N_44528,N_40831);
nor U49152 (N_49152,N_43187,N_44711);
nand U49153 (N_49153,N_42269,N_44799);
nor U49154 (N_49154,N_41061,N_42172);
nand U49155 (N_49155,N_40014,N_43884);
xnor U49156 (N_49156,N_42465,N_43869);
nor U49157 (N_49157,N_42069,N_40894);
or U49158 (N_49158,N_42040,N_44128);
and U49159 (N_49159,N_43916,N_44312);
and U49160 (N_49160,N_41676,N_42706);
nand U49161 (N_49161,N_42513,N_44714);
xor U49162 (N_49162,N_41679,N_40061);
and U49163 (N_49163,N_40749,N_40776);
and U49164 (N_49164,N_40711,N_41802);
and U49165 (N_49165,N_42563,N_40743);
nand U49166 (N_49166,N_43978,N_43462);
nand U49167 (N_49167,N_44012,N_41843);
or U49168 (N_49168,N_42184,N_44151);
and U49169 (N_49169,N_43546,N_40143);
nor U49170 (N_49170,N_43059,N_40588);
nor U49171 (N_49171,N_44673,N_44136);
nand U49172 (N_49172,N_41455,N_41909);
or U49173 (N_49173,N_41549,N_43733);
and U49174 (N_49174,N_41636,N_44102);
nor U49175 (N_49175,N_43907,N_43386);
or U49176 (N_49176,N_44743,N_42723);
and U49177 (N_49177,N_42050,N_44444);
xor U49178 (N_49178,N_43602,N_43329);
xor U49179 (N_49179,N_43255,N_41382);
nor U49180 (N_49180,N_43743,N_40218);
and U49181 (N_49181,N_41477,N_42998);
or U49182 (N_49182,N_40102,N_40252);
nand U49183 (N_49183,N_40767,N_42600);
and U49184 (N_49184,N_42283,N_43392);
nor U49185 (N_49185,N_40204,N_41716);
nor U49186 (N_49186,N_42990,N_42720);
and U49187 (N_49187,N_42732,N_41625);
or U49188 (N_49188,N_40351,N_44159);
or U49189 (N_49189,N_42434,N_44733);
nor U49190 (N_49190,N_40148,N_41080);
nand U49191 (N_49191,N_42729,N_43376);
xnor U49192 (N_49192,N_40670,N_44116);
or U49193 (N_49193,N_43402,N_43712);
and U49194 (N_49194,N_43491,N_42320);
and U49195 (N_49195,N_41268,N_44235);
or U49196 (N_49196,N_44061,N_42845);
or U49197 (N_49197,N_44111,N_40459);
or U49198 (N_49198,N_42769,N_44373);
nand U49199 (N_49199,N_43785,N_43102);
or U49200 (N_49200,N_40608,N_43709);
nand U49201 (N_49201,N_41624,N_42812);
or U49202 (N_49202,N_41326,N_43676);
nor U49203 (N_49203,N_41869,N_41251);
and U49204 (N_49204,N_40864,N_42437);
or U49205 (N_49205,N_42154,N_42861);
or U49206 (N_49206,N_43690,N_42784);
nand U49207 (N_49207,N_44887,N_41569);
or U49208 (N_49208,N_41040,N_44881);
and U49209 (N_49209,N_41848,N_44482);
nand U49210 (N_49210,N_43439,N_41835);
and U49211 (N_49211,N_44805,N_43462);
nand U49212 (N_49212,N_41430,N_42432);
nand U49213 (N_49213,N_42710,N_44333);
and U49214 (N_49214,N_43889,N_42012);
or U49215 (N_49215,N_43384,N_43139);
or U49216 (N_49216,N_44237,N_43044);
nor U49217 (N_49217,N_44421,N_42036);
nand U49218 (N_49218,N_41583,N_42726);
nor U49219 (N_49219,N_44635,N_43381);
and U49220 (N_49220,N_40197,N_41910);
or U49221 (N_49221,N_42423,N_40742);
nand U49222 (N_49222,N_43417,N_44351);
nor U49223 (N_49223,N_44693,N_43520);
nor U49224 (N_49224,N_44104,N_41133);
nor U49225 (N_49225,N_43371,N_42038);
xnor U49226 (N_49226,N_40520,N_41911);
xnor U49227 (N_49227,N_41151,N_44549);
and U49228 (N_49228,N_44950,N_41950);
nand U49229 (N_49229,N_40271,N_40915);
and U49230 (N_49230,N_40277,N_43753);
and U49231 (N_49231,N_44920,N_42539);
nor U49232 (N_49232,N_41470,N_43894);
nor U49233 (N_49233,N_43394,N_44434);
and U49234 (N_49234,N_44816,N_44992);
and U49235 (N_49235,N_44175,N_40924);
and U49236 (N_49236,N_41945,N_44909);
nor U49237 (N_49237,N_43845,N_40108);
or U49238 (N_49238,N_41382,N_42744);
and U49239 (N_49239,N_41786,N_44737);
xor U49240 (N_49240,N_42671,N_42013);
nor U49241 (N_49241,N_40897,N_44419);
nor U49242 (N_49242,N_43317,N_40638);
nor U49243 (N_49243,N_42468,N_41508);
nand U49244 (N_49244,N_43662,N_43695);
nor U49245 (N_49245,N_43307,N_41129);
and U49246 (N_49246,N_41284,N_41398);
or U49247 (N_49247,N_40008,N_42735);
xnor U49248 (N_49248,N_41909,N_43057);
or U49249 (N_49249,N_41385,N_44777);
or U49250 (N_49250,N_40892,N_44574);
nor U49251 (N_49251,N_42683,N_44489);
or U49252 (N_49252,N_41669,N_43642);
nand U49253 (N_49253,N_40792,N_41504);
and U49254 (N_49254,N_44281,N_44197);
or U49255 (N_49255,N_42243,N_43605);
or U49256 (N_49256,N_42069,N_42094);
or U49257 (N_49257,N_40609,N_40403);
or U49258 (N_49258,N_44699,N_40814);
nor U49259 (N_49259,N_40920,N_44357);
nor U49260 (N_49260,N_42794,N_43130);
and U49261 (N_49261,N_41551,N_43963);
or U49262 (N_49262,N_40883,N_40696);
nor U49263 (N_49263,N_40536,N_40716);
and U49264 (N_49264,N_40017,N_41523);
or U49265 (N_49265,N_40616,N_41376);
xnor U49266 (N_49266,N_42106,N_44901);
or U49267 (N_49267,N_43667,N_44847);
nor U49268 (N_49268,N_40242,N_44998);
and U49269 (N_49269,N_42381,N_41204);
or U49270 (N_49270,N_43880,N_41302);
or U49271 (N_49271,N_41841,N_43929);
nor U49272 (N_49272,N_41661,N_42940);
or U49273 (N_49273,N_40058,N_42900);
nor U49274 (N_49274,N_42238,N_41207);
nor U49275 (N_49275,N_40009,N_40349);
and U49276 (N_49276,N_44639,N_41091);
nor U49277 (N_49277,N_41929,N_41446);
nand U49278 (N_49278,N_42481,N_40739);
nand U49279 (N_49279,N_41888,N_41578);
and U49280 (N_49280,N_40997,N_43223);
nand U49281 (N_49281,N_41239,N_41344);
and U49282 (N_49282,N_44651,N_43597);
nor U49283 (N_49283,N_40082,N_42223);
or U49284 (N_49284,N_44707,N_43406);
nor U49285 (N_49285,N_42301,N_40605);
and U49286 (N_49286,N_44015,N_42680);
nand U49287 (N_49287,N_42096,N_42202);
nand U49288 (N_49288,N_42800,N_43226);
nand U49289 (N_49289,N_40414,N_44693);
or U49290 (N_49290,N_42241,N_44145);
nand U49291 (N_49291,N_43236,N_42572);
nand U49292 (N_49292,N_42073,N_43461);
and U49293 (N_49293,N_43829,N_42888);
or U49294 (N_49294,N_43896,N_43702);
nand U49295 (N_49295,N_41052,N_43764);
xnor U49296 (N_49296,N_40438,N_41833);
or U49297 (N_49297,N_43921,N_43529);
and U49298 (N_49298,N_44097,N_44950);
and U49299 (N_49299,N_42963,N_41418);
nand U49300 (N_49300,N_41747,N_40047);
and U49301 (N_49301,N_41125,N_43145);
and U49302 (N_49302,N_43369,N_40617);
or U49303 (N_49303,N_42997,N_44712);
and U49304 (N_49304,N_43085,N_41289);
xnor U49305 (N_49305,N_40525,N_44839);
nor U49306 (N_49306,N_41062,N_44782);
or U49307 (N_49307,N_42596,N_41523);
and U49308 (N_49308,N_40050,N_44278);
and U49309 (N_49309,N_42951,N_43096);
nand U49310 (N_49310,N_44180,N_40302);
nor U49311 (N_49311,N_42847,N_43675);
or U49312 (N_49312,N_44528,N_40646);
nand U49313 (N_49313,N_44727,N_43864);
nor U49314 (N_49314,N_42609,N_44849);
and U49315 (N_49315,N_42873,N_40945);
or U49316 (N_49316,N_41759,N_40875);
and U49317 (N_49317,N_44857,N_42061);
or U49318 (N_49318,N_42407,N_42109);
nand U49319 (N_49319,N_40929,N_40949);
and U49320 (N_49320,N_44971,N_42276);
or U49321 (N_49321,N_42008,N_40542);
nand U49322 (N_49322,N_40549,N_41298);
or U49323 (N_49323,N_40463,N_41885);
nand U49324 (N_49324,N_41067,N_42585);
and U49325 (N_49325,N_43826,N_43389);
nor U49326 (N_49326,N_44406,N_42622);
xnor U49327 (N_49327,N_41150,N_43785);
and U49328 (N_49328,N_40376,N_43680);
or U49329 (N_49329,N_42800,N_41675);
nand U49330 (N_49330,N_40486,N_40152);
xor U49331 (N_49331,N_44602,N_43093);
nor U49332 (N_49332,N_40932,N_41417);
nand U49333 (N_49333,N_44655,N_41065);
and U49334 (N_49334,N_40897,N_42815);
and U49335 (N_49335,N_42596,N_41064);
and U49336 (N_49336,N_43801,N_40672);
and U49337 (N_49337,N_41967,N_42099);
or U49338 (N_49338,N_41771,N_42408);
nor U49339 (N_49339,N_42168,N_40094);
xnor U49340 (N_49340,N_44945,N_42655);
nor U49341 (N_49341,N_40287,N_42015);
nor U49342 (N_49342,N_40893,N_40305);
nand U49343 (N_49343,N_40305,N_41175);
nand U49344 (N_49344,N_42345,N_42981);
and U49345 (N_49345,N_40066,N_44932);
nor U49346 (N_49346,N_43880,N_41042);
nor U49347 (N_49347,N_43826,N_41637);
xnor U49348 (N_49348,N_40835,N_44831);
nor U49349 (N_49349,N_41827,N_40829);
and U49350 (N_49350,N_40567,N_40274);
and U49351 (N_49351,N_41742,N_44672);
xnor U49352 (N_49352,N_41423,N_42951);
nand U49353 (N_49353,N_44018,N_42937);
xor U49354 (N_49354,N_44020,N_44467);
nor U49355 (N_49355,N_44749,N_40002);
xnor U49356 (N_49356,N_43833,N_40158);
nor U49357 (N_49357,N_40514,N_41480);
nand U49358 (N_49358,N_43275,N_44614);
xnor U49359 (N_49359,N_41470,N_41091);
nor U49360 (N_49360,N_41591,N_41351);
nand U49361 (N_49361,N_40207,N_40397);
nor U49362 (N_49362,N_44169,N_42700);
nor U49363 (N_49363,N_44647,N_42440);
nand U49364 (N_49364,N_40389,N_44243);
and U49365 (N_49365,N_43203,N_43535);
nand U49366 (N_49366,N_41733,N_41602);
and U49367 (N_49367,N_40695,N_42224);
xor U49368 (N_49368,N_43074,N_43648);
xnor U49369 (N_49369,N_41376,N_42046);
xnor U49370 (N_49370,N_44613,N_41473);
nand U49371 (N_49371,N_43842,N_42797);
and U49372 (N_49372,N_42722,N_43155);
nand U49373 (N_49373,N_43977,N_40790);
and U49374 (N_49374,N_43023,N_40882);
nand U49375 (N_49375,N_43003,N_44009);
nand U49376 (N_49376,N_44695,N_43458);
xor U49377 (N_49377,N_42999,N_43916);
or U49378 (N_49378,N_41153,N_44291);
and U49379 (N_49379,N_43466,N_40064);
and U49380 (N_49380,N_42989,N_42980);
nand U49381 (N_49381,N_42292,N_43095);
nand U49382 (N_49382,N_41546,N_42999);
or U49383 (N_49383,N_42704,N_43369);
and U49384 (N_49384,N_44390,N_40031);
or U49385 (N_49385,N_43220,N_43639);
xor U49386 (N_49386,N_43096,N_43569);
nor U49387 (N_49387,N_41086,N_43485);
or U49388 (N_49388,N_41049,N_43479);
and U49389 (N_49389,N_40412,N_41920);
or U49390 (N_49390,N_44123,N_43675);
and U49391 (N_49391,N_42804,N_44678);
or U49392 (N_49392,N_41293,N_40200);
nand U49393 (N_49393,N_43196,N_42971);
and U49394 (N_49394,N_40934,N_42756);
nor U49395 (N_49395,N_44063,N_43507);
or U49396 (N_49396,N_41522,N_43781);
and U49397 (N_49397,N_44057,N_44485);
or U49398 (N_49398,N_44407,N_43621);
and U49399 (N_49399,N_42179,N_43939);
and U49400 (N_49400,N_44483,N_41782);
or U49401 (N_49401,N_44535,N_42736);
and U49402 (N_49402,N_43808,N_42231);
and U49403 (N_49403,N_44383,N_44602);
xnor U49404 (N_49404,N_41697,N_41078);
nand U49405 (N_49405,N_40974,N_40952);
nand U49406 (N_49406,N_41839,N_41259);
nand U49407 (N_49407,N_43692,N_40418);
or U49408 (N_49408,N_41898,N_43863);
nor U49409 (N_49409,N_40195,N_44525);
xnor U49410 (N_49410,N_41849,N_40589);
nor U49411 (N_49411,N_41614,N_43820);
xor U49412 (N_49412,N_44895,N_40674);
and U49413 (N_49413,N_42880,N_41816);
nor U49414 (N_49414,N_42742,N_44624);
and U49415 (N_49415,N_41312,N_43197);
nor U49416 (N_49416,N_41706,N_42493);
nand U49417 (N_49417,N_42477,N_43766);
nor U49418 (N_49418,N_40477,N_43562);
nor U49419 (N_49419,N_44460,N_41115);
or U49420 (N_49420,N_44329,N_42358);
nor U49421 (N_49421,N_41694,N_41800);
nand U49422 (N_49422,N_40008,N_43617);
nor U49423 (N_49423,N_41012,N_43893);
and U49424 (N_49424,N_42421,N_44979);
nor U49425 (N_49425,N_43740,N_44772);
nor U49426 (N_49426,N_41290,N_41128);
nor U49427 (N_49427,N_44967,N_40006);
or U49428 (N_49428,N_41179,N_43251);
nor U49429 (N_49429,N_42773,N_42342);
nor U49430 (N_49430,N_42962,N_43583);
nand U49431 (N_49431,N_43386,N_43810);
nor U49432 (N_49432,N_40691,N_44429);
nand U49433 (N_49433,N_42030,N_43495);
nand U49434 (N_49434,N_42967,N_43983);
nand U49435 (N_49435,N_43924,N_42570);
and U49436 (N_49436,N_41709,N_42031);
nand U49437 (N_49437,N_41588,N_42179);
nor U49438 (N_49438,N_40912,N_42630);
xor U49439 (N_49439,N_41816,N_42780);
and U49440 (N_49440,N_41623,N_40519);
nand U49441 (N_49441,N_42457,N_44031);
nor U49442 (N_49442,N_42873,N_41514);
nand U49443 (N_49443,N_43461,N_43108);
nor U49444 (N_49444,N_43253,N_42729);
nand U49445 (N_49445,N_40983,N_44061);
nor U49446 (N_49446,N_41277,N_43189);
nand U49447 (N_49447,N_44192,N_41122);
nor U49448 (N_49448,N_44858,N_44344);
nand U49449 (N_49449,N_42336,N_42686);
and U49450 (N_49450,N_40135,N_43982);
or U49451 (N_49451,N_44769,N_41044);
nor U49452 (N_49452,N_44342,N_44903);
and U49453 (N_49453,N_42487,N_43611);
or U49454 (N_49454,N_43850,N_43436);
and U49455 (N_49455,N_44811,N_41723);
nor U49456 (N_49456,N_44665,N_44510);
or U49457 (N_49457,N_40862,N_44304);
nor U49458 (N_49458,N_44322,N_42775);
nand U49459 (N_49459,N_42874,N_44185);
nor U49460 (N_49460,N_42952,N_42744);
nor U49461 (N_49461,N_44179,N_43281);
or U49462 (N_49462,N_42739,N_40446);
xor U49463 (N_49463,N_41622,N_44470);
nor U49464 (N_49464,N_43872,N_44469);
nor U49465 (N_49465,N_40739,N_42693);
and U49466 (N_49466,N_42531,N_44564);
nand U49467 (N_49467,N_40860,N_43648);
nor U49468 (N_49468,N_42577,N_43881);
and U49469 (N_49469,N_42877,N_43069);
or U49470 (N_49470,N_42690,N_44761);
and U49471 (N_49471,N_43793,N_42323);
or U49472 (N_49472,N_40648,N_43775);
or U49473 (N_49473,N_44801,N_44200);
nand U49474 (N_49474,N_43298,N_43942);
nor U49475 (N_49475,N_44771,N_42104);
nand U49476 (N_49476,N_42235,N_40427);
and U49477 (N_49477,N_44103,N_43737);
or U49478 (N_49478,N_41544,N_43024);
and U49479 (N_49479,N_41384,N_41463);
nand U49480 (N_49480,N_43830,N_41213);
nor U49481 (N_49481,N_44392,N_40499);
nor U49482 (N_49482,N_42563,N_41767);
and U49483 (N_49483,N_42965,N_44224);
nor U49484 (N_49484,N_41296,N_41499);
nand U49485 (N_49485,N_43127,N_44116);
and U49486 (N_49486,N_43969,N_43498);
and U49487 (N_49487,N_41788,N_42874);
and U49488 (N_49488,N_41724,N_40115);
nor U49489 (N_49489,N_41353,N_43847);
or U49490 (N_49490,N_41781,N_44814);
or U49491 (N_49491,N_43456,N_41096);
and U49492 (N_49492,N_40405,N_44819);
nor U49493 (N_49493,N_40088,N_42076);
or U49494 (N_49494,N_40870,N_44649);
and U49495 (N_49495,N_43336,N_42177);
nor U49496 (N_49496,N_43006,N_43346);
or U49497 (N_49497,N_41785,N_41663);
nor U49498 (N_49498,N_44278,N_43314);
nand U49499 (N_49499,N_43550,N_44638);
xor U49500 (N_49500,N_44344,N_40472);
nor U49501 (N_49501,N_44751,N_43906);
nor U49502 (N_49502,N_43118,N_44698);
nor U49503 (N_49503,N_41747,N_41248);
and U49504 (N_49504,N_41882,N_42916);
or U49505 (N_49505,N_43634,N_41810);
and U49506 (N_49506,N_43161,N_41570);
nor U49507 (N_49507,N_43601,N_44254);
nand U49508 (N_49508,N_44386,N_42243);
nor U49509 (N_49509,N_41960,N_43204);
and U49510 (N_49510,N_40166,N_40404);
or U49511 (N_49511,N_43998,N_40172);
nand U49512 (N_49512,N_40213,N_43333);
and U49513 (N_49513,N_42507,N_42312);
or U49514 (N_49514,N_43888,N_40677);
nand U49515 (N_49515,N_40543,N_44958);
nand U49516 (N_49516,N_41175,N_43080);
xor U49517 (N_49517,N_43847,N_43903);
or U49518 (N_49518,N_44361,N_41300);
nor U49519 (N_49519,N_40899,N_42897);
nand U49520 (N_49520,N_44274,N_44352);
nor U49521 (N_49521,N_43729,N_43528);
or U49522 (N_49522,N_42877,N_40353);
and U49523 (N_49523,N_40701,N_41343);
xnor U49524 (N_49524,N_40484,N_40212);
nor U49525 (N_49525,N_40348,N_43003);
nand U49526 (N_49526,N_41317,N_41414);
and U49527 (N_49527,N_44263,N_42865);
xnor U49528 (N_49528,N_40326,N_42372);
and U49529 (N_49529,N_40870,N_44133);
nand U49530 (N_49530,N_44452,N_40276);
or U49531 (N_49531,N_44423,N_43387);
nor U49532 (N_49532,N_41283,N_40615);
and U49533 (N_49533,N_42689,N_42949);
and U49534 (N_49534,N_42530,N_43969);
nor U49535 (N_49535,N_40508,N_41686);
xor U49536 (N_49536,N_42375,N_41937);
and U49537 (N_49537,N_43974,N_43388);
nor U49538 (N_49538,N_44885,N_43095);
nor U49539 (N_49539,N_43385,N_42268);
and U49540 (N_49540,N_43198,N_43397);
xnor U49541 (N_49541,N_41284,N_44770);
nor U49542 (N_49542,N_44284,N_40148);
nand U49543 (N_49543,N_44460,N_42166);
nand U49544 (N_49544,N_41671,N_44697);
nand U49545 (N_49545,N_40396,N_41179);
or U49546 (N_49546,N_42470,N_40504);
and U49547 (N_49547,N_42375,N_40519);
xor U49548 (N_49548,N_42806,N_42479);
or U49549 (N_49549,N_42703,N_41282);
xor U49550 (N_49550,N_43432,N_40827);
or U49551 (N_49551,N_41093,N_42864);
and U49552 (N_49552,N_40661,N_41276);
and U49553 (N_49553,N_44131,N_41107);
xnor U49554 (N_49554,N_42078,N_43783);
or U49555 (N_49555,N_43771,N_44085);
or U49556 (N_49556,N_44072,N_41568);
and U49557 (N_49557,N_40635,N_44622);
or U49558 (N_49558,N_44051,N_40222);
nand U49559 (N_49559,N_40040,N_43985);
or U49560 (N_49560,N_42418,N_40454);
or U49561 (N_49561,N_44704,N_42384);
nor U49562 (N_49562,N_42792,N_40039);
or U49563 (N_49563,N_42743,N_43893);
nand U49564 (N_49564,N_40434,N_42655);
nand U49565 (N_49565,N_42897,N_44406);
or U49566 (N_49566,N_40276,N_44033);
and U49567 (N_49567,N_41428,N_41457);
and U49568 (N_49568,N_43749,N_42385);
and U49569 (N_49569,N_44095,N_42779);
xor U49570 (N_49570,N_40982,N_43392);
xnor U49571 (N_49571,N_42659,N_41299);
nor U49572 (N_49572,N_40038,N_44434);
nor U49573 (N_49573,N_40065,N_44907);
or U49574 (N_49574,N_44596,N_41434);
nor U49575 (N_49575,N_42222,N_40426);
and U49576 (N_49576,N_43822,N_42335);
xor U49577 (N_49577,N_41243,N_41581);
nor U49578 (N_49578,N_44149,N_42999);
nor U49579 (N_49579,N_40919,N_40561);
nor U49580 (N_49580,N_42163,N_41076);
xnor U49581 (N_49581,N_44130,N_43306);
or U49582 (N_49582,N_43399,N_42724);
or U49583 (N_49583,N_43987,N_44075);
or U49584 (N_49584,N_43637,N_43204);
nand U49585 (N_49585,N_44879,N_40977);
or U49586 (N_49586,N_40785,N_42783);
nor U49587 (N_49587,N_44115,N_41481);
or U49588 (N_49588,N_43422,N_42944);
and U49589 (N_49589,N_40692,N_42234);
nor U49590 (N_49590,N_42107,N_40527);
nand U49591 (N_49591,N_44911,N_41477);
nor U49592 (N_49592,N_40556,N_43845);
and U49593 (N_49593,N_42726,N_40449);
and U49594 (N_49594,N_41716,N_44486);
nand U49595 (N_49595,N_41419,N_44993);
or U49596 (N_49596,N_44365,N_43235);
nor U49597 (N_49597,N_40664,N_44574);
and U49598 (N_49598,N_44191,N_44817);
nand U49599 (N_49599,N_44220,N_40366);
nor U49600 (N_49600,N_40837,N_41801);
xnor U49601 (N_49601,N_42367,N_41394);
nand U49602 (N_49602,N_40478,N_42139);
nor U49603 (N_49603,N_44140,N_43054);
nand U49604 (N_49604,N_40609,N_43084);
and U49605 (N_49605,N_40279,N_44564);
nand U49606 (N_49606,N_42691,N_41758);
nand U49607 (N_49607,N_40346,N_40820);
and U49608 (N_49608,N_42199,N_40750);
xnor U49609 (N_49609,N_43286,N_44867);
and U49610 (N_49610,N_43068,N_40252);
nor U49611 (N_49611,N_44034,N_42657);
nand U49612 (N_49612,N_41683,N_42965);
or U49613 (N_49613,N_40025,N_44923);
xor U49614 (N_49614,N_44642,N_41978);
nand U49615 (N_49615,N_40979,N_43178);
nand U49616 (N_49616,N_41837,N_42170);
and U49617 (N_49617,N_40376,N_42304);
and U49618 (N_49618,N_44359,N_44220);
nand U49619 (N_49619,N_43971,N_43349);
nor U49620 (N_49620,N_40502,N_42325);
nor U49621 (N_49621,N_41461,N_41794);
nand U49622 (N_49622,N_43571,N_44980);
nand U49623 (N_49623,N_42210,N_41565);
nand U49624 (N_49624,N_40275,N_40867);
and U49625 (N_49625,N_40206,N_40797);
nor U49626 (N_49626,N_43122,N_40354);
nand U49627 (N_49627,N_41469,N_42253);
or U49628 (N_49628,N_41780,N_41403);
and U49629 (N_49629,N_40499,N_42993);
nand U49630 (N_49630,N_42134,N_42841);
nand U49631 (N_49631,N_40640,N_42680);
xnor U49632 (N_49632,N_42830,N_42666);
nand U49633 (N_49633,N_43702,N_40017);
nor U49634 (N_49634,N_40338,N_41946);
nor U49635 (N_49635,N_43692,N_44670);
nor U49636 (N_49636,N_42548,N_41401);
nor U49637 (N_49637,N_42420,N_44895);
and U49638 (N_49638,N_40807,N_44477);
and U49639 (N_49639,N_43372,N_42490);
nand U49640 (N_49640,N_42576,N_41824);
and U49641 (N_49641,N_44200,N_41674);
xor U49642 (N_49642,N_42061,N_40663);
or U49643 (N_49643,N_44057,N_44859);
nand U49644 (N_49644,N_44838,N_41543);
or U49645 (N_49645,N_41323,N_40661);
nor U49646 (N_49646,N_41637,N_41062);
nor U49647 (N_49647,N_41819,N_41510);
and U49648 (N_49648,N_44829,N_42935);
xnor U49649 (N_49649,N_41462,N_41568);
or U49650 (N_49650,N_40208,N_44447);
and U49651 (N_49651,N_41408,N_41525);
or U49652 (N_49652,N_43808,N_44163);
and U49653 (N_49653,N_41125,N_40206);
nand U49654 (N_49654,N_43983,N_41965);
or U49655 (N_49655,N_43373,N_42317);
xor U49656 (N_49656,N_40185,N_44056);
or U49657 (N_49657,N_41339,N_41116);
or U49658 (N_49658,N_41531,N_44476);
or U49659 (N_49659,N_40719,N_41081);
nand U49660 (N_49660,N_44482,N_41476);
nor U49661 (N_49661,N_42417,N_42251);
nand U49662 (N_49662,N_42999,N_44269);
or U49663 (N_49663,N_42274,N_40011);
nand U49664 (N_49664,N_42151,N_41691);
nor U49665 (N_49665,N_44758,N_44917);
or U49666 (N_49666,N_43440,N_41181);
nor U49667 (N_49667,N_43371,N_40520);
or U49668 (N_49668,N_41085,N_43120);
nor U49669 (N_49669,N_43523,N_42097);
and U49670 (N_49670,N_42349,N_42842);
or U49671 (N_49671,N_44997,N_41615);
and U49672 (N_49672,N_42158,N_42895);
xor U49673 (N_49673,N_42661,N_43371);
or U49674 (N_49674,N_40982,N_41752);
and U49675 (N_49675,N_43743,N_44747);
nand U49676 (N_49676,N_40114,N_41819);
nand U49677 (N_49677,N_43167,N_43260);
nor U49678 (N_49678,N_43013,N_44465);
and U49679 (N_49679,N_44637,N_44346);
and U49680 (N_49680,N_42931,N_41907);
nor U49681 (N_49681,N_43072,N_44912);
and U49682 (N_49682,N_44591,N_40753);
nor U49683 (N_49683,N_43001,N_40753);
or U49684 (N_49684,N_43060,N_43525);
or U49685 (N_49685,N_40610,N_41871);
nand U49686 (N_49686,N_43476,N_43801);
xor U49687 (N_49687,N_41846,N_40496);
nand U49688 (N_49688,N_41558,N_42200);
nor U49689 (N_49689,N_40671,N_44114);
and U49690 (N_49690,N_40634,N_41559);
nor U49691 (N_49691,N_42395,N_43595);
nand U49692 (N_49692,N_40516,N_42659);
and U49693 (N_49693,N_43718,N_44646);
or U49694 (N_49694,N_43798,N_42327);
and U49695 (N_49695,N_44522,N_43031);
nor U49696 (N_49696,N_44404,N_43070);
xor U49697 (N_49697,N_43873,N_43254);
nor U49698 (N_49698,N_43648,N_40531);
nand U49699 (N_49699,N_41507,N_40196);
nor U49700 (N_49700,N_42923,N_42951);
xor U49701 (N_49701,N_42613,N_42385);
xnor U49702 (N_49702,N_41079,N_42814);
nand U49703 (N_49703,N_41226,N_40869);
and U49704 (N_49704,N_40385,N_44018);
nor U49705 (N_49705,N_42690,N_40497);
and U49706 (N_49706,N_44403,N_43356);
and U49707 (N_49707,N_42308,N_41275);
and U49708 (N_49708,N_44512,N_41072);
or U49709 (N_49709,N_40136,N_42384);
and U49710 (N_49710,N_44273,N_40072);
or U49711 (N_49711,N_42832,N_42905);
and U49712 (N_49712,N_42057,N_43886);
or U49713 (N_49713,N_43085,N_42142);
nor U49714 (N_49714,N_43063,N_40311);
or U49715 (N_49715,N_44731,N_44532);
and U49716 (N_49716,N_42005,N_42083);
nor U49717 (N_49717,N_41249,N_40532);
or U49718 (N_49718,N_42498,N_42529);
xnor U49719 (N_49719,N_44783,N_41059);
or U49720 (N_49720,N_42865,N_43024);
and U49721 (N_49721,N_43084,N_43435);
nand U49722 (N_49722,N_44603,N_41049);
and U49723 (N_49723,N_43368,N_40688);
nand U49724 (N_49724,N_40495,N_44459);
nand U49725 (N_49725,N_40286,N_43102);
or U49726 (N_49726,N_43395,N_41435);
and U49727 (N_49727,N_44344,N_41193);
xnor U49728 (N_49728,N_44735,N_43049);
and U49729 (N_49729,N_40193,N_42744);
nor U49730 (N_49730,N_41523,N_41859);
nor U49731 (N_49731,N_40443,N_40804);
nor U49732 (N_49732,N_42211,N_43962);
nand U49733 (N_49733,N_44295,N_41547);
nand U49734 (N_49734,N_41365,N_44658);
nor U49735 (N_49735,N_42848,N_40917);
or U49736 (N_49736,N_43685,N_41631);
nor U49737 (N_49737,N_44619,N_41936);
or U49738 (N_49738,N_43300,N_41213);
nor U49739 (N_49739,N_40704,N_44527);
nor U49740 (N_49740,N_41405,N_40193);
nor U49741 (N_49741,N_42858,N_42945);
nand U49742 (N_49742,N_40957,N_44464);
nand U49743 (N_49743,N_41844,N_43034);
or U49744 (N_49744,N_42164,N_41163);
nand U49745 (N_49745,N_43801,N_44317);
and U49746 (N_49746,N_40987,N_44048);
and U49747 (N_49747,N_42057,N_43971);
or U49748 (N_49748,N_43411,N_42412);
or U49749 (N_49749,N_43096,N_43941);
and U49750 (N_49750,N_42217,N_40598);
nor U49751 (N_49751,N_44646,N_44444);
nor U49752 (N_49752,N_41037,N_44331);
nand U49753 (N_49753,N_43822,N_40306);
nor U49754 (N_49754,N_41950,N_40477);
nand U49755 (N_49755,N_40164,N_41080);
nor U49756 (N_49756,N_43658,N_42894);
or U49757 (N_49757,N_42536,N_43427);
nand U49758 (N_49758,N_40786,N_41551);
or U49759 (N_49759,N_40621,N_43220);
nand U49760 (N_49760,N_41399,N_42448);
or U49761 (N_49761,N_41648,N_41925);
nor U49762 (N_49762,N_41808,N_40102);
nor U49763 (N_49763,N_40013,N_40128);
nand U49764 (N_49764,N_44778,N_42402);
xnor U49765 (N_49765,N_40792,N_44965);
nand U49766 (N_49766,N_44726,N_41459);
or U49767 (N_49767,N_42226,N_44641);
and U49768 (N_49768,N_42958,N_43817);
and U49769 (N_49769,N_43264,N_40803);
nand U49770 (N_49770,N_41733,N_40549);
and U49771 (N_49771,N_43313,N_44064);
nand U49772 (N_49772,N_43697,N_42698);
xor U49773 (N_49773,N_41565,N_44226);
nor U49774 (N_49774,N_43681,N_41206);
or U49775 (N_49775,N_44728,N_40860);
or U49776 (N_49776,N_40605,N_43213);
nor U49777 (N_49777,N_42853,N_44415);
nor U49778 (N_49778,N_40989,N_43735);
nor U49779 (N_49779,N_44073,N_40504);
xor U49780 (N_49780,N_43502,N_43210);
xnor U49781 (N_49781,N_43829,N_42996);
or U49782 (N_49782,N_40051,N_42367);
nand U49783 (N_49783,N_43877,N_43087);
or U49784 (N_49784,N_42184,N_44108);
nand U49785 (N_49785,N_40416,N_40279);
or U49786 (N_49786,N_41495,N_41006);
nor U49787 (N_49787,N_41000,N_41196);
xor U49788 (N_49788,N_41955,N_44988);
and U49789 (N_49789,N_43876,N_40665);
and U49790 (N_49790,N_43827,N_43201);
or U49791 (N_49791,N_44884,N_42218);
and U49792 (N_49792,N_40483,N_40289);
nor U49793 (N_49793,N_41891,N_44004);
or U49794 (N_49794,N_44337,N_44116);
xnor U49795 (N_49795,N_42480,N_44730);
or U49796 (N_49796,N_43766,N_41175);
nor U49797 (N_49797,N_42077,N_42304);
nand U49798 (N_49798,N_40725,N_44166);
and U49799 (N_49799,N_41143,N_42090);
or U49800 (N_49800,N_40006,N_40809);
nor U49801 (N_49801,N_43633,N_43980);
nor U49802 (N_49802,N_44064,N_42564);
nand U49803 (N_49803,N_44012,N_43919);
and U49804 (N_49804,N_42784,N_42936);
nor U49805 (N_49805,N_44740,N_42511);
or U49806 (N_49806,N_40531,N_44659);
nand U49807 (N_49807,N_40444,N_43817);
and U49808 (N_49808,N_41298,N_41643);
and U49809 (N_49809,N_44790,N_40523);
and U49810 (N_49810,N_43309,N_40350);
or U49811 (N_49811,N_40577,N_41181);
nand U49812 (N_49812,N_40790,N_43252);
nand U49813 (N_49813,N_40677,N_41306);
nand U49814 (N_49814,N_44744,N_43893);
or U49815 (N_49815,N_43195,N_42759);
and U49816 (N_49816,N_44728,N_40311);
nand U49817 (N_49817,N_42984,N_44255);
nor U49818 (N_49818,N_40615,N_41510);
nand U49819 (N_49819,N_42675,N_44025);
xnor U49820 (N_49820,N_44755,N_40811);
xor U49821 (N_49821,N_41679,N_42325);
or U49822 (N_49822,N_44618,N_44577);
nand U49823 (N_49823,N_44353,N_43723);
nand U49824 (N_49824,N_40599,N_40381);
or U49825 (N_49825,N_40608,N_40852);
nand U49826 (N_49826,N_42067,N_44254);
or U49827 (N_49827,N_42991,N_43308);
or U49828 (N_49828,N_40571,N_40814);
nand U49829 (N_49829,N_43703,N_40415);
nand U49830 (N_49830,N_44989,N_40145);
or U49831 (N_49831,N_42019,N_41407);
nor U49832 (N_49832,N_43678,N_40886);
and U49833 (N_49833,N_42894,N_40222);
and U49834 (N_49834,N_42424,N_44344);
or U49835 (N_49835,N_42441,N_43142);
nand U49836 (N_49836,N_43197,N_42127);
nand U49837 (N_49837,N_43782,N_44618);
nor U49838 (N_49838,N_40570,N_44531);
and U49839 (N_49839,N_41981,N_44936);
or U49840 (N_49840,N_43795,N_42876);
and U49841 (N_49841,N_41865,N_42232);
or U49842 (N_49842,N_44614,N_44670);
nor U49843 (N_49843,N_42665,N_44563);
nor U49844 (N_49844,N_44556,N_42850);
and U49845 (N_49845,N_41050,N_42798);
nor U49846 (N_49846,N_42377,N_43905);
nor U49847 (N_49847,N_43663,N_43553);
and U49848 (N_49848,N_44519,N_43832);
or U49849 (N_49849,N_40395,N_41010);
or U49850 (N_49850,N_41210,N_43344);
and U49851 (N_49851,N_43861,N_43347);
nand U49852 (N_49852,N_44087,N_41597);
nand U49853 (N_49853,N_43973,N_42889);
and U49854 (N_49854,N_43847,N_42580);
nand U49855 (N_49855,N_41173,N_40002);
and U49856 (N_49856,N_41463,N_43044);
nor U49857 (N_49857,N_41905,N_40300);
nand U49858 (N_49858,N_41650,N_42745);
nand U49859 (N_49859,N_41115,N_43611);
or U49860 (N_49860,N_44834,N_43812);
and U49861 (N_49861,N_40803,N_40870);
and U49862 (N_49862,N_41159,N_44266);
and U49863 (N_49863,N_40789,N_42501);
and U49864 (N_49864,N_43439,N_42257);
nor U49865 (N_49865,N_42826,N_44478);
or U49866 (N_49866,N_44901,N_41224);
or U49867 (N_49867,N_42536,N_44797);
nor U49868 (N_49868,N_42682,N_42773);
and U49869 (N_49869,N_43294,N_42488);
and U49870 (N_49870,N_43246,N_43225);
and U49871 (N_49871,N_43524,N_43514);
nor U49872 (N_49872,N_41031,N_43392);
or U49873 (N_49873,N_42235,N_41961);
nand U49874 (N_49874,N_43109,N_43744);
and U49875 (N_49875,N_41337,N_41604);
nand U49876 (N_49876,N_42700,N_44347);
nor U49877 (N_49877,N_40478,N_42369);
nor U49878 (N_49878,N_42466,N_43156);
nor U49879 (N_49879,N_43605,N_44545);
nor U49880 (N_49880,N_44742,N_42984);
xnor U49881 (N_49881,N_41605,N_40447);
or U49882 (N_49882,N_42876,N_43373);
nor U49883 (N_49883,N_40653,N_44574);
nor U49884 (N_49884,N_40649,N_43878);
or U49885 (N_49885,N_41064,N_44821);
xor U49886 (N_49886,N_44571,N_41357);
nor U49887 (N_49887,N_43880,N_43036);
nor U49888 (N_49888,N_40632,N_42447);
nand U49889 (N_49889,N_43681,N_41739);
or U49890 (N_49890,N_43678,N_41031);
and U49891 (N_49891,N_44823,N_40200);
or U49892 (N_49892,N_42304,N_42061);
nand U49893 (N_49893,N_44615,N_42190);
nand U49894 (N_49894,N_43677,N_44066);
nor U49895 (N_49895,N_43151,N_41511);
xor U49896 (N_49896,N_42163,N_41995);
nand U49897 (N_49897,N_42880,N_40234);
and U49898 (N_49898,N_41446,N_42361);
nor U49899 (N_49899,N_44057,N_43673);
nor U49900 (N_49900,N_42193,N_44705);
and U49901 (N_49901,N_42590,N_43280);
or U49902 (N_49902,N_44590,N_41242);
nor U49903 (N_49903,N_40122,N_42839);
or U49904 (N_49904,N_44335,N_43724);
xnor U49905 (N_49905,N_44742,N_44142);
nor U49906 (N_49906,N_41274,N_40426);
or U49907 (N_49907,N_44492,N_43779);
nand U49908 (N_49908,N_41724,N_42099);
or U49909 (N_49909,N_42796,N_42715);
nand U49910 (N_49910,N_44649,N_42245);
nor U49911 (N_49911,N_44929,N_44771);
or U49912 (N_49912,N_40605,N_41247);
nand U49913 (N_49913,N_41308,N_44437);
or U49914 (N_49914,N_42987,N_44322);
nand U49915 (N_49915,N_43199,N_40007);
nand U49916 (N_49916,N_41589,N_40411);
and U49917 (N_49917,N_40235,N_44273);
and U49918 (N_49918,N_43643,N_41984);
and U49919 (N_49919,N_43860,N_40591);
and U49920 (N_49920,N_41303,N_44404);
nand U49921 (N_49921,N_43110,N_43875);
or U49922 (N_49922,N_44160,N_40932);
or U49923 (N_49923,N_44312,N_44188);
nand U49924 (N_49924,N_40788,N_42851);
nor U49925 (N_49925,N_42247,N_42557);
and U49926 (N_49926,N_41583,N_40630);
or U49927 (N_49927,N_43172,N_44250);
or U49928 (N_49928,N_44500,N_44569);
and U49929 (N_49929,N_42054,N_42548);
or U49930 (N_49930,N_42583,N_44813);
xnor U49931 (N_49931,N_43140,N_40896);
or U49932 (N_49932,N_42766,N_41865);
nand U49933 (N_49933,N_44869,N_43520);
or U49934 (N_49934,N_41289,N_42925);
nor U49935 (N_49935,N_42317,N_44075);
nand U49936 (N_49936,N_43248,N_41301);
nand U49937 (N_49937,N_40676,N_43972);
or U49938 (N_49938,N_43755,N_41632);
or U49939 (N_49939,N_42388,N_43727);
and U49940 (N_49940,N_40333,N_40055);
xor U49941 (N_49941,N_42301,N_43877);
nor U49942 (N_49942,N_41313,N_41314);
nor U49943 (N_49943,N_42047,N_40229);
or U49944 (N_49944,N_42331,N_40533);
nand U49945 (N_49945,N_40233,N_44969);
and U49946 (N_49946,N_44529,N_40113);
nor U49947 (N_49947,N_41009,N_41316);
and U49948 (N_49948,N_41537,N_43259);
and U49949 (N_49949,N_41431,N_40728);
nand U49950 (N_49950,N_42965,N_40528);
nor U49951 (N_49951,N_44527,N_44135);
nand U49952 (N_49952,N_40064,N_41144);
or U49953 (N_49953,N_43365,N_41215);
and U49954 (N_49954,N_44836,N_41576);
nand U49955 (N_49955,N_40423,N_43467);
nor U49956 (N_49956,N_43700,N_42829);
or U49957 (N_49957,N_42249,N_41091);
xor U49958 (N_49958,N_41355,N_41212);
nor U49959 (N_49959,N_40099,N_42890);
nor U49960 (N_49960,N_40718,N_42854);
and U49961 (N_49961,N_40480,N_44519);
and U49962 (N_49962,N_44345,N_42238);
nand U49963 (N_49963,N_40879,N_41432);
nor U49964 (N_49964,N_40189,N_42140);
xnor U49965 (N_49965,N_44970,N_44734);
nand U49966 (N_49966,N_41012,N_40887);
nor U49967 (N_49967,N_42772,N_41792);
nand U49968 (N_49968,N_43585,N_43581);
nor U49969 (N_49969,N_41238,N_40155);
nand U49970 (N_49970,N_41331,N_44702);
nand U49971 (N_49971,N_41415,N_40895);
or U49972 (N_49972,N_44350,N_42124);
or U49973 (N_49973,N_43787,N_40167);
and U49974 (N_49974,N_43191,N_44083);
nor U49975 (N_49975,N_44626,N_44027);
nand U49976 (N_49976,N_42187,N_40358);
nor U49977 (N_49977,N_44056,N_44232);
xnor U49978 (N_49978,N_40967,N_40637);
or U49979 (N_49979,N_44338,N_44937);
nor U49980 (N_49980,N_42996,N_41245);
or U49981 (N_49981,N_41439,N_41290);
or U49982 (N_49982,N_41786,N_42747);
or U49983 (N_49983,N_43897,N_40790);
or U49984 (N_49984,N_43184,N_44651);
nor U49985 (N_49985,N_41387,N_44845);
nand U49986 (N_49986,N_41385,N_41549);
nor U49987 (N_49987,N_42591,N_41590);
nand U49988 (N_49988,N_44463,N_44852);
or U49989 (N_49989,N_43449,N_42014);
xor U49990 (N_49990,N_44947,N_44617);
nor U49991 (N_49991,N_41427,N_43740);
and U49992 (N_49992,N_40386,N_43089);
nor U49993 (N_49993,N_40328,N_44589);
or U49994 (N_49994,N_42487,N_43815);
or U49995 (N_49995,N_42054,N_44390);
and U49996 (N_49996,N_41391,N_41650);
and U49997 (N_49997,N_42804,N_40498);
xnor U49998 (N_49998,N_41108,N_44987);
and U49999 (N_49999,N_43030,N_43047);
and UO_0 (O_0,N_47092,N_46289);
nor UO_1 (O_1,N_48426,N_46707);
nor UO_2 (O_2,N_49683,N_47093);
or UO_3 (O_3,N_47099,N_48890);
or UO_4 (O_4,N_46900,N_49777);
nand UO_5 (O_5,N_47055,N_49858);
nand UO_6 (O_6,N_46672,N_47188);
nand UO_7 (O_7,N_46710,N_47841);
or UO_8 (O_8,N_48462,N_49091);
nor UO_9 (O_9,N_45611,N_45795);
nor UO_10 (O_10,N_45086,N_46074);
or UO_11 (O_11,N_46040,N_46475);
and UO_12 (O_12,N_49714,N_49972);
and UO_13 (O_13,N_47699,N_48522);
and UO_14 (O_14,N_46474,N_45155);
nand UO_15 (O_15,N_46940,N_45183);
and UO_16 (O_16,N_48040,N_45461);
or UO_17 (O_17,N_47508,N_49307);
nor UO_18 (O_18,N_46658,N_48549);
nand UO_19 (O_19,N_47962,N_46220);
nor UO_20 (O_20,N_49973,N_47660);
nor UO_21 (O_21,N_45434,N_46336);
nor UO_22 (O_22,N_47686,N_48799);
or UO_23 (O_23,N_45585,N_45015);
or UO_24 (O_24,N_48452,N_47587);
nor UO_25 (O_25,N_45697,N_48018);
nor UO_26 (O_26,N_49521,N_49348);
nor UO_27 (O_27,N_49891,N_49810);
xor UO_28 (O_28,N_47189,N_47240);
and UO_29 (O_29,N_47907,N_49320);
and UO_30 (O_30,N_47580,N_45624);
nor UO_31 (O_31,N_46813,N_49577);
and UO_32 (O_32,N_46833,N_46134);
xnor UO_33 (O_33,N_46688,N_49042);
nor UO_34 (O_34,N_46614,N_46534);
nor UO_35 (O_35,N_49076,N_45390);
and UO_36 (O_36,N_46723,N_45582);
nor UO_37 (O_37,N_48245,N_46440);
nor UO_38 (O_38,N_46817,N_46633);
and UO_39 (O_39,N_46943,N_47884);
or UO_40 (O_40,N_47017,N_47346);
or UO_41 (O_41,N_49877,N_45309);
and UO_42 (O_42,N_45347,N_47060);
nor UO_43 (O_43,N_49574,N_47338);
or UO_44 (O_44,N_48223,N_45030);
nand UO_45 (O_45,N_45707,N_48399);
nand UO_46 (O_46,N_49483,N_45272);
nor UO_47 (O_47,N_45836,N_46741);
and UO_48 (O_48,N_49189,N_47140);
and UO_49 (O_49,N_47859,N_49466);
and UO_50 (O_50,N_46554,N_45603);
or UO_51 (O_51,N_48185,N_46061);
or UO_52 (O_52,N_48049,N_48374);
and UO_53 (O_53,N_47864,N_45524);
and UO_54 (O_54,N_49619,N_45923);
nand UO_55 (O_55,N_45291,N_49132);
or UO_56 (O_56,N_48918,N_49075);
nand UO_57 (O_57,N_46635,N_49729);
and UO_58 (O_58,N_46523,N_45289);
or UO_59 (O_59,N_46133,N_48866);
and UO_60 (O_60,N_47023,N_49799);
nor UO_61 (O_61,N_47305,N_46222);
nor UO_62 (O_62,N_48017,N_48105);
or UO_63 (O_63,N_45467,N_46893);
or UO_64 (O_64,N_48054,N_49908);
nor UO_65 (O_65,N_46231,N_49916);
nand UO_66 (O_66,N_46985,N_46766);
nand UO_67 (O_67,N_48818,N_45798);
xor UO_68 (O_68,N_45148,N_46693);
or UO_69 (O_69,N_46454,N_49816);
or UO_70 (O_70,N_46153,N_48016);
or UO_71 (O_71,N_45997,N_47571);
xor UO_72 (O_72,N_48046,N_45075);
nor UO_73 (O_73,N_47169,N_45587);
nand UO_74 (O_74,N_45371,N_48839);
nand UO_75 (O_75,N_47177,N_47697);
nand UO_76 (O_76,N_45479,N_48526);
and UO_77 (O_77,N_46564,N_46364);
and UO_78 (O_78,N_45592,N_45646);
xor UO_79 (O_79,N_49443,N_49438);
nand UO_80 (O_80,N_45310,N_46448);
nor UO_81 (O_81,N_48699,N_47341);
nand UO_82 (O_82,N_45964,N_45385);
nor UO_83 (O_83,N_47952,N_49603);
nor UO_84 (O_84,N_49399,N_46405);
nand UO_85 (O_85,N_45073,N_48989);
nand UO_86 (O_86,N_46768,N_47637);
xnor UO_87 (O_87,N_46158,N_47021);
nor UO_88 (O_88,N_46851,N_47829);
or UO_89 (O_89,N_47225,N_47701);
or UO_90 (O_90,N_46856,N_49802);
or UO_91 (O_91,N_46292,N_46677);
nor UO_92 (O_92,N_46749,N_46241);
nand UO_93 (O_93,N_49665,N_46545);
nor UO_94 (O_94,N_48630,N_49808);
or UO_95 (O_95,N_46065,N_45223);
nor UO_96 (O_96,N_47524,N_45166);
and UO_97 (O_97,N_45049,N_47256);
nand UO_98 (O_98,N_45410,N_45335);
or UO_99 (O_99,N_45729,N_45100);
nor UO_100 (O_100,N_45138,N_47591);
and UO_101 (O_101,N_46675,N_48525);
or UO_102 (O_102,N_46835,N_45508);
nor UO_103 (O_103,N_48030,N_48910);
or UO_104 (O_104,N_47726,N_45115);
nor UO_105 (O_105,N_49990,N_49261);
or UO_106 (O_106,N_45366,N_45175);
or UO_107 (O_107,N_49650,N_48567);
xnor UO_108 (O_108,N_49966,N_49145);
or UO_109 (O_109,N_45786,N_45572);
and UO_110 (O_110,N_48550,N_47249);
nor UO_111 (O_111,N_45614,N_48832);
nand UO_112 (O_112,N_49664,N_45243);
and UO_113 (O_113,N_46301,N_47437);
or UO_114 (O_114,N_46462,N_47152);
nor UO_115 (O_115,N_49372,N_46145);
or UO_116 (O_116,N_47570,N_47011);
nand UO_117 (O_117,N_47657,N_46172);
and UO_118 (O_118,N_45452,N_45355);
and UO_119 (O_119,N_49149,N_47815);
and UO_120 (O_120,N_47037,N_49028);
nand UO_121 (O_121,N_49449,N_46910);
or UO_122 (O_122,N_47654,N_46684);
or UO_123 (O_123,N_49484,N_46589);
nor UO_124 (O_124,N_45986,N_48651);
xnor UO_125 (O_125,N_47538,N_48347);
and UO_126 (O_126,N_47431,N_46109);
nor UO_127 (O_127,N_49964,N_48093);
or UO_128 (O_128,N_45456,N_49516);
nand UO_129 (O_129,N_47960,N_49981);
or UO_130 (O_130,N_46908,N_48156);
nor UO_131 (O_131,N_46959,N_47958);
nor UO_132 (O_132,N_46681,N_49989);
nor UO_133 (O_133,N_45544,N_47927);
nor UO_134 (O_134,N_45333,N_46206);
nor UO_135 (O_135,N_46007,N_47110);
nor UO_136 (O_136,N_49366,N_47557);
nand UO_137 (O_137,N_48358,N_49188);
xor UO_138 (O_138,N_49159,N_45717);
and UO_139 (O_139,N_49226,N_47880);
nor UO_140 (O_140,N_48899,N_45915);
xor UO_141 (O_141,N_47360,N_48132);
and UO_142 (O_142,N_46769,N_49783);
or UO_143 (O_143,N_49104,N_45616);
xor UO_144 (O_144,N_47752,N_48411);
and UO_145 (O_145,N_46154,N_49613);
xor UO_146 (O_146,N_47123,N_49138);
nor UO_147 (O_147,N_48702,N_46692);
nor UO_148 (O_148,N_45612,N_49067);
nand UO_149 (O_149,N_48831,N_49626);
or UO_150 (O_150,N_48743,N_48577);
xor UO_151 (O_151,N_45302,N_45742);
or UO_152 (O_152,N_47273,N_47247);
and UO_153 (O_153,N_49288,N_45424);
nor UO_154 (O_154,N_47222,N_47635);
nor UO_155 (O_155,N_48515,N_46088);
nor UO_156 (O_156,N_45562,N_48341);
nand UO_157 (O_157,N_46955,N_45249);
nor UO_158 (O_158,N_49486,N_46214);
xnor UO_159 (O_159,N_48469,N_45312);
nor UO_160 (O_160,N_45083,N_46712);
xnor UO_161 (O_161,N_45160,N_47412);
and UO_162 (O_162,N_46213,N_48642);
nand UO_163 (O_163,N_49924,N_45525);
and UO_164 (O_164,N_47615,N_46471);
xnor UO_165 (O_165,N_49183,N_47742);
xnor UO_166 (O_166,N_47393,N_48034);
or UO_167 (O_167,N_49755,N_47838);
or UO_168 (O_168,N_46411,N_47084);
or UO_169 (O_169,N_49277,N_49295);
xnor UO_170 (O_170,N_49734,N_46035);
xor UO_171 (O_171,N_47381,N_49184);
nand UO_172 (O_172,N_49287,N_45801);
nor UO_173 (O_173,N_48151,N_46574);
or UO_174 (O_174,N_49493,N_49682);
nand UO_175 (O_175,N_49697,N_49616);
or UO_176 (O_176,N_48619,N_47766);
and UO_177 (O_177,N_49835,N_46782);
and UO_178 (O_178,N_47835,N_45045);
nor UO_179 (O_179,N_48383,N_49914);
and UO_180 (O_180,N_49929,N_48148);
or UO_181 (O_181,N_47767,N_46901);
xnor UO_182 (O_182,N_47708,N_48301);
and UO_183 (O_183,N_49994,N_47039);
and UO_184 (O_184,N_45214,N_47854);
and UO_185 (O_185,N_48896,N_49244);
xor UO_186 (O_186,N_45698,N_47146);
xor UO_187 (O_187,N_49046,N_48086);
and UO_188 (O_188,N_46227,N_45809);
nor UO_189 (O_189,N_49100,N_49312);
nand UO_190 (O_190,N_46530,N_49782);
and UO_191 (O_191,N_45730,N_49940);
nand UO_192 (O_192,N_45430,N_49114);
nand UO_193 (O_193,N_48451,N_47245);
and UO_194 (O_194,N_49815,N_48145);
or UO_195 (O_195,N_47083,N_48995);
or UO_196 (O_196,N_49901,N_45949);
or UO_197 (O_197,N_47403,N_48837);
nand UO_198 (O_198,N_47432,N_48260);
and UO_199 (O_199,N_46425,N_45884);
and UO_200 (O_200,N_47241,N_45770);
or UO_201 (O_201,N_49880,N_47034);
or UO_202 (O_202,N_47300,N_46797);
or UO_203 (O_203,N_49719,N_48594);
nor UO_204 (O_204,N_46042,N_45263);
and UO_205 (O_205,N_46143,N_45095);
or UO_206 (O_206,N_45899,N_46353);
xor UO_207 (O_207,N_46493,N_49241);
nor UO_208 (O_208,N_47905,N_49367);
or UO_209 (O_209,N_49198,N_46935);
and UO_210 (O_210,N_46915,N_46198);
or UO_211 (O_211,N_46647,N_45131);
or UO_212 (O_212,N_47542,N_46458);
and UO_213 (O_213,N_48931,N_46611);
xnor UO_214 (O_214,N_47170,N_45292);
nand UO_215 (O_215,N_48098,N_48179);
and UO_216 (O_216,N_45259,N_47940);
and UO_217 (O_217,N_46089,N_48107);
nor UO_218 (O_218,N_48415,N_48945);
nor UO_219 (O_219,N_47866,N_48486);
or UO_220 (O_220,N_49131,N_48723);
nor UO_221 (O_221,N_47218,N_47168);
or UO_222 (O_222,N_49462,N_46827);
nand UO_223 (O_223,N_46731,N_49576);
and UO_224 (O_224,N_48888,N_47285);
xor UO_225 (O_225,N_45182,N_46778);
or UO_226 (O_226,N_47574,N_49881);
nand UO_227 (O_227,N_47978,N_48494);
or UO_228 (O_228,N_47743,N_49999);
nand UO_229 (O_229,N_45920,N_46247);
or UO_230 (O_230,N_46550,N_49242);
nor UO_231 (O_231,N_49886,N_49101);
nand UO_232 (O_232,N_48907,N_46793);
or UO_233 (O_233,N_48344,N_49544);
and UO_234 (O_234,N_49831,N_49398);
nor UO_235 (O_235,N_49548,N_46632);
or UO_236 (O_236,N_47024,N_47228);
and UO_237 (O_237,N_46097,N_47374);
or UO_238 (O_238,N_47428,N_49645);
and UO_239 (O_239,N_46698,N_47390);
or UO_240 (O_240,N_47577,N_49748);
nor UO_241 (O_241,N_46274,N_48122);
nand UO_242 (O_242,N_46587,N_47843);
or UO_243 (O_243,N_47821,N_46481);
and UO_244 (O_244,N_48072,N_45265);
or UO_245 (O_245,N_49873,N_45577);
and UO_246 (O_246,N_49098,N_48733);
and UO_247 (O_247,N_45752,N_48765);
and UO_248 (O_248,N_49174,N_47179);
xor UO_249 (O_249,N_47925,N_47278);
nand UO_250 (O_250,N_48271,N_47072);
nand UO_251 (O_251,N_49432,N_46019);
and UO_252 (O_252,N_46976,N_46515);
nor UO_253 (O_253,N_47204,N_46713);
nor UO_254 (O_254,N_49454,N_47471);
nand UO_255 (O_255,N_48956,N_49502);
nor UO_256 (O_256,N_47913,N_48708);
or UO_257 (O_257,N_47857,N_48756);
and UO_258 (O_258,N_47299,N_48787);
nand UO_259 (O_259,N_48328,N_48474);
and UO_260 (O_260,N_49803,N_45590);
nand UO_261 (O_261,N_46037,N_48089);
and UO_262 (O_262,N_48511,N_48395);
nor UO_263 (O_263,N_47281,N_49379);
and UO_264 (O_264,N_46244,N_45609);
and UO_265 (O_265,N_48563,N_47178);
nand UO_266 (O_266,N_45613,N_47100);
nor UO_267 (O_267,N_46776,N_48304);
nand UO_268 (O_268,N_47347,N_45256);
and UO_269 (O_269,N_46914,N_46001);
nor UO_270 (O_270,N_45651,N_47109);
and UO_271 (O_271,N_49843,N_48169);
nor UO_272 (O_272,N_47718,N_49048);
nor UO_273 (O_273,N_46862,N_46946);
nand UO_274 (O_274,N_49027,N_48114);
nand UO_275 (O_275,N_45196,N_48934);
nand UO_276 (O_276,N_49662,N_47561);
nor UO_277 (O_277,N_48479,N_45981);
or UO_278 (O_278,N_48429,N_46280);
nor UO_279 (O_279,N_47194,N_46730);
and UO_280 (O_280,N_49476,N_49250);
and UO_281 (O_281,N_48102,N_46294);
and UO_282 (O_282,N_47845,N_46881);
or UO_283 (O_283,N_45888,N_46127);
or UO_284 (O_284,N_49837,N_48460);
nor UO_285 (O_285,N_47087,N_48578);
nor UO_286 (O_286,N_46287,N_45762);
or UO_287 (O_287,N_48144,N_46014);
nor UO_288 (O_288,N_45031,N_49272);
and UO_289 (O_289,N_46234,N_48942);
and UO_290 (O_290,N_48750,N_49670);
nand UO_291 (O_291,N_48561,N_48661);
and UO_292 (O_292,N_49125,N_49086);
and UO_293 (O_293,N_48311,N_46815);
and UO_294 (O_294,N_49479,N_47141);
or UO_295 (O_295,N_47250,N_46447);
nand UO_296 (O_296,N_49518,N_49463);
or UO_297 (O_297,N_47401,N_47205);
nand UO_298 (O_298,N_46956,N_45515);
and UO_299 (O_299,N_45995,N_47186);
nand UO_300 (O_300,N_49833,N_48854);
nand UO_301 (O_301,N_48143,N_49325);
and UO_302 (O_302,N_49988,N_46099);
or UO_303 (O_303,N_45689,N_47460);
or UO_304 (O_304,N_49968,N_47722);
and UO_305 (O_305,N_45172,N_45617);
nor UO_306 (O_306,N_46066,N_46062);
or UO_307 (O_307,N_47762,N_49531);
or UO_308 (O_308,N_49495,N_48700);
and UO_309 (O_309,N_49378,N_47400);
and UO_310 (O_310,N_47662,N_45566);
xor UO_311 (O_311,N_45431,N_49246);
or UO_312 (O_312,N_46580,N_47568);
or UO_313 (O_313,N_45376,N_49381);
or UO_314 (O_314,N_48720,N_48597);
nand UO_315 (O_315,N_47203,N_48565);
and UO_316 (O_316,N_49275,N_47549);
nor UO_317 (O_317,N_47071,N_49137);
nand UO_318 (O_318,N_45297,N_49085);
or UO_319 (O_319,N_49439,N_48969);
or UO_320 (O_320,N_49687,N_47214);
and UO_321 (O_321,N_49955,N_48305);
nand UO_322 (O_322,N_45691,N_48496);
nand UO_323 (O_323,N_47944,N_47018);
and UO_324 (O_324,N_49934,N_49072);
and UO_325 (O_325,N_49666,N_48189);
or UO_326 (O_326,N_47379,N_47727);
nand UO_327 (O_327,N_48187,N_49889);
or UO_328 (O_328,N_45020,N_47288);
or UO_329 (O_329,N_47387,N_49927);
and UO_330 (O_330,N_47610,N_46535);
nor UO_331 (O_331,N_45134,N_45639);
nor UO_332 (O_332,N_48716,N_49844);
and UO_333 (O_333,N_49862,N_48346);
or UO_334 (O_334,N_48976,N_45618);
or UO_335 (O_335,N_45268,N_48729);
and UO_336 (O_336,N_46786,N_49663);
or UO_337 (O_337,N_47490,N_48300);
nand UO_338 (O_338,N_45489,N_48695);
nand UO_339 (O_339,N_49821,N_48530);
nor UO_340 (O_340,N_45758,N_48119);
and UO_341 (O_341,N_46013,N_48901);
or UO_342 (O_342,N_49062,N_48617);
xor UO_343 (O_343,N_46996,N_48192);
and UO_344 (O_344,N_47807,N_49382);
or UO_345 (O_345,N_46697,N_45350);
xnor UO_346 (O_346,N_48435,N_48568);
nand UO_347 (O_347,N_45386,N_49515);
nor UO_348 (O_348,N_47450,N_45914);
nand UO_349 (O_349,N_45829,N_46537);
and UO_350 (O_350,N_47030,N_47182);
nand UO_351 (O_351,N_47923,N_49195);
or UO_352 (O_352,N_45975,N_49407);
nor UO_353 (O_353,N_49834,N_48076);
nor UO_354 (O_354,N_48096,N_46196);
nand UO_355 (O_355,N_45427,N_46250);
nor UO_356 (O_356,N_47676,N_48769);
or UO_357 (O_357,N_49087,N_49411);
nor UO_358 (O_358,N_48365,N_46842);
or UO_359 (O_359,N_48330,N_48937);
and UO_360 (O_360,N_49676,N_46740);
and UO_361 (O_361,N_48442,N_45293);
nand UO_362 (O_362,N_49809,N_45513);
xor UO_363 (O_363,N_47628,N_46478);
nor UO_364 (O_364,N_49280,N_48984);
and UO_365 (O_365,N_46655,N_45307);
or UO_366 (O_366,N_48570,N_46029);
nor UO_367 (O_367,N_49509,N_45046);
nor UO_368 (O_368,N_45442,N_46906);
xnor UO_369 (O_369,N_48283,N_45586);
and UO_370 (O_370,N_47778,N_47348);
or UO_371 (O_371,N_48372,N_45678);
xor UO_372 (O_372,N_48378,N_48274);
nor UO_373 (O_373,N_49582,N_49725);
and UO_374 (O_374,N_47029,N_48183);
nor UO_375 (O_375,N_47794,N_49453);
nand UO_376 (O_376,N_49170,N_48580);
nand UO_377 (O_377,N_48176,N_45823);
nand UO_378 (O_378,N_46466,N_46983);
or UO_379 (O_379,N_49201,N_46569);
nand UO_380 (O_380,N_47190,N_46063);
or UO_381 (O_381,N_47114,N_45145);
nor UO_382 (O_382,N_48241,N_49309);
nor UO_383 (O_383,N_46563,N_45969);
nor UO_384 (O_384,N_45666,N_45731);
nand UO_385 (O_385,N_45535,N_46331);
nor UO_386 (O_386,N_46790,N_46657);
nor UO_387 (O_387,N_45526,N_48803);
and UO_388 (O_388,N_45890,N_45184);
and UO_389 (O_389,N_47519,N_49129);
nand UO_390 (O_390,N_49464,N_45325);
nor UO_391 (O_391,N_48256,N_49147);
nor UO_392 (O_392,N_49614,N_45542);
nand UO_393 (O_393,N_47493,N_49945);
xor UO_394 (O_394,N_45018,N_47066);
nand UO_395 (O_395,N_47010,N_45408);
and UO_396 (O_396,N_45925,N_46395);
xor UO_397 (O_397,N_45242,N_48585);
nor UO_398 (O_398,N_49305,N_49984);
xor UO_399 (O_399,N_45853,N_47881);
or UO_400 (O_400,N_47995,N_46075);
or UO_401 (O_401,N_47137,N_45488);
nor UO_402 (O_402,N_48645,N_49173);
xnor UO_403 (O_403,N_46455,N_48622);
nor UO_404 (O_404,N_46004,N_48006);
nand UO_405 (O_405,N_45527,N_49043);
xnor UO_406 (O_406,N_46439,N_47830);
nand UO_407 (O_407,N_45747,N_47627);
nor UO_408 (O_408,N_45168,N_47407);
nor UO_409 (O_409,N_47098,N_48504);
nor UO_410 (O_410,N_46207,N_49900);
and UO_411 (O_411,N_45276,N_46918);
nor UO_412 (O_412,N_48202,N_48336);
nand UO_413 (O_413,N_45159,N_45240);
and UO_414 (O_414,N_49735,N_48432);
nor UO_415 (O_415,N_49960,N_47625);
nor UO_416 (O_416,N_49055,N_49290);
and UO_417 (O_417,N_48427,N_47440);
xor UO_418 (O_418,N_46041,N_48009);
xnor UO_419 (O_419,N_49866,N_47920);
nand UO_420 (O_420,N_49607,N_48846);
or UO_421 (O_421,N_47918,N_47414);
nand UO_422 (O_422,N_47648,N_47038);
and UO_423 (O_423,N_46806,N_46516);
xnor UO_424 (O_424,N_49501,N_47311);
nor UO_425 (O_425,N_45339,N_47477);
nor UO_426 (O_426,N_49329,N_49526);
or UO_427 (O_427,N_47721,N_46205);
nand UO_428 (O_428,N_46416,N_48895);
or UO_429 (O_429,N_48412,N_48444);
or UO_430 (O_430,N_46663,N_49135);
nand UO_431 (O_431,N_48652,N_45475);
or UO_432 (O_432,N_49296,N_45912);
and UO_433 (O_433,N_46795,N_46579);
and UO_434 (O_434,N_47646,N_46131);
and UO_435 (O_435,N_47789,N_47891);
and UO_436 (O_436,N_45939,N_48506);
and UO_437 (O_437,N_48685,N_47784);
or UO_438 (O_438,N_46077,N_46626);
xnor UO_439 (O_439,N_48862,N_49639);
and UO_440 (O_440,N_49690,N_46964);
nor UO_441 (O_441,N_45320,N_47623);
xnor UO_442 (O_442,N_45207,N_48903);
nor UO_443 (O_443,N_46577,N_47313);
nor UO_444 (O_444,N_46122,N_47380);
xor UO_445 (O_445,N_46272,N_46796);
and UO_446 (O_446,N_48491,N_48424);
nor UO_447 (O_447,N_48215,N_49073);
nand UO_448 (O_448,N_48828,N_49232);
nor UO_449 (O_449,N_49757,N_47659);
or UO_450 (O_450,N_48291,N_47861);
nor UO_451 (O_451,N_48884,N_49434);
nor UO_452 (O_452,N_46708,N_45827);
nand UO_453 (O_453,N_48882,N_46139);
nor UO_454 (O_454,N_46819,N_47424);
nand UO_455 (O_455,N_45474,N_49389);
nor UO_456 (O_456,N_46188,N_49818);
or UO_457 (O_457,N_48200,N_49094);
nand UO_458 (O_458,N_45094,N_48588);
nand UO_459 (O_459,N_45980,N_47397);
nand UO_460 (O_460,N_45640,N_46746);
nand UO_461 (O_461,N_49304,N_46832);
or UO_462 (O_462,N_48255,N_48704);
or UO_463 (O_463,N_46662,N_47201);
nand UO_464 (O_464,N_46000,N_49693);
nand UO_465 (O_465,N_47343,N_46430);
nor UO_466 (O_466,N_46499,N_47198);
and UO_467 (O_467,N_46674,N_48680);
and UO_468 (O_468,N_47227,N_45540);
xor UO_469 (O_469,N_49743,N_49217);
nand UO_470 (O_470,N_49878,N_45945);
and UO_471 (O_471,N_47602,N_45460);
nor UO_472 (O_472,N_47936,N_49139);
nand UO_473 (O_473,N_46892,N_46977);
or UO_474 (O_474,N_48898,N_46111);
nand UO_475 (O_475,N_47924,N_45803);
and UO_476 (O_476,N_48238,N_46086);
xor UO_477 (O_477,N_48941,N_46816);
or UO_478 (O_478,N_49252,N_47297);
nand UO_479 (O_479,N_45720,N_45652);
nor UO_480 (O_480,N_45622,N_47293);
nor UO_481 (O_481,N_48725,N_49642);
and UO_482 (O_482,N_45314,N_46733);
nor UO_483 (O_483,N_45568,N_46903);
and UO_484 (O_484,N_49884,N_49146);
nand UO_485 (O_485,N_47284,N_49970);
or UO_486 (O_486,N_49907,N_46619);
xor UO_487 (O_487,N_47257,N_45529);
or UO_488 (O_488,N_49513,N_47675);
or UO_489 (O_489,N_45687,N_46069);
xor UO_490 (O_490,N_48891,N_45271);
nand UO_491 (O_491,N_47790,N_46483);
nand UO_492 (O_492,N_46546,N_47756);
nor UO_493 (O_493,N_45204,N_49196);
nor UO_494 (O_494,N_48992,N_47695);
or UO_495 (O_495,N_45667,N_49632);
or UO_496 (O_496,N_48463,N_47565);
nor UO_497 (O_497,N_45677,N_47875);
nor UO_498 (O_498,N_47406,N_45534);
nor UO_499 (O_499,N_46627,N_47454);
and UO_500 (O_500,N_48686,N_46605);
nor UO_501 (O_501,N_49596,N_45751);
and UO_502 (O_502,N_47753,N_47349);
nand UO_503 (O_503,N_45202,N_49016);
and UO_504 (O_504,N_46699,N_48674);
xor UO_505 (O_505,N_47455,N_45907);
nor UO_506 (O_506,N_47351,N_49359);
and UO_507 (O_507,N_48035,N_46664);
and UO_508 (O_508,N_45007,N_49216);
nor UO_509 (O_509,N_45322,N_49455);
nand UO_510 (O_510,N_49396,N_45607);
nor UO_511 (O_511,N_46020,N_45088);
nand UO_512 (O_512,N_47933,N_45569);
or UO_513 (O_513,N_47199,N_49008);
and UO_514 (O_514,N_45069,N_48523);
or UO_515 (O_515,N_48108,N_47714);
xor UO_516 (O_516,N_45288,N_45212);
and UO_517 (O_517,N_46195,N_47078);
or UO_518 (O_518,N_48163,N_48873);
nor UO_519 (O_519,N_49847,N_48671);
or UO_520 (O_520,N_46607,N_46055);
nor UO_521 (O_521,N_47617,N_47116);
nand UO_522 (O_522,N_49897,N_45298);
or UO_523 (O_523,N_46686,N_45942);
nand UO_524 (O_524,N_47649,N_48340);
nand UO_525 (O_525,N_47441,N_46048);
nand UO_526 (O_526,N_49801,N_48084);
and UO_527 (O_527,N_46347,N_48562);
nand UO_528 (O_528,N_46103,N_48312);
nand UO_529 (O_529,N_47765,N_47286);
and UO_530 (O_530,N_45739,N_45631);
nor UO_531 (O_531,N_46053,N_45749);
xnor UO_532 (O_532,N_48414,N_48536);
nor UO_533 (O_533,N_48448,N_47128);
nor UO_534 (O_534,N_46264,N_47971);
nand UO_535 (O_535,N_46146,N_47622);
nand UO_536 (O_536,N_48778,N_46486);
nand UO_537 (O_537,N_47283,N_48961);
nand UO_538 (O_538,N_48827,N_47504);
nor UO_539 (O_539,N_48109,N_48705);
nand UO_540 (O_540,N_47748,N_48690);
nand UO_541 (O_541,N_47946,N_45664);
or UO_542 (O_542,N_48277,N_48558);
nor UO_543 (O_543,N_47014,N_48904);
xor UO_544 (O_544,N_46329,N_49942);
and UO_545 (O_545,N_47149,N_48919);
xor UO_546 (O_546,N_47153,N_45137);
and UO_547 (O_547,N_46370,N_47801);
nor UO_548 (O_548,N_49123,N_49025);
nand UO_549 (O_549,N_49733,N_45104);
nor UO_550 (O_550,N_48653,N_45399);
or UO_551 (O_551,N_48861,N_46362);
nand UO_552 (O_552,N_45559,N_47535);
nand UO_553 (O_553,N_49221,N_45701);
nand UO_554 (O_554,N_48973,N_47174);
xnor UO_555 (O_555,N_47655,N_48154);
xnor UO_556 (O_556,N_46271,N_45336);
or UO_557 (O_557,N_48618,N_45725);
or UO_558 (O_558,N_45567,N_47248);
xnor UO_559 (O_559,N_45663,N_48269);
nor UO_560 (O_560,N_45685,N_47027);
nand UO_561 (O_561,N_45736,N_49959);
nand UO_562 (O_562,N_49776,N_46868);
xor UO_563 (O_563,N_45187,N_47849);
nand UO_564 (O_564,N_48316,N_47626);
and UO_565 (O_565,N_45278,N_49040);
and UO_566 (O_566,N_47665,N_46745);
xor UO_567 (O_567,N_45052,N_49499);
or UO_568 (O_568,N_46552,N_47238);
nand UO_569 (O_569,N_48650,N_46937);
nor UO_570 (O_570,N_49158,N_49871);
xnor UO_571 (O_571,N_46254,N_45373);
and UO_572 (O_572,N_48129,N_48218);
nand UO_573 (O_573,N_48422,N_45850);
nor UO_574 (O_574,N_46360,N_47295);
or UO_575 (O_575,N_45197,N_49951);
or UO_576 (O_576,N_46757,N_48943);
nor UO_577 (O_577,N_47558,N_49391);
and UO_578 (O_578,N_48540,N_46283);
and UO_579 (O_579,N_45668,N_48106);
or UO_580 (O_580,N_47945,N_45846);
and UO_581 (O_581,N_48795,N_45043);
nand UO_582 (O_582,N_47272,N_45181);
or UO_583 (O_583,N_45423,N_47365);
nor UO_584 (O_584,N_47994,N_46238);
nand UO_585 (O_585,N_46240,N_45469);
nand UO_586 (O_586,N_45791,N_45573);
or UO_587 (O_587,N_48669,N_45711);
nor UO_588 (O_588,N_46369,N_45224);
and UO_589 (O_589,N_46352,N_45228);
nand UO_590 (O_590,N_47498,N_48259);
nor UO_591 (O_591,N_46303,N_47077);
and UO_592 (O_592,N_46700,N_47405);
nor UO_593 (O_593,N_46379,N_47470);
and UO_594 (O_594,N_46812,N_47419);
nor UO_595 (O_595,N_46163,N_47512);
xor UO_596 (O_596,N_46896,N_48998);
nand UO_597 (O_597,N_48505,N_49532);
nand UO_598 (O_598,N_45188,N_46293);
nor UO_599 (O_599,N_47922,N_46006);
and UO_600 (O_600,N_48968,N_48867);
nand UO_601 (O_601,N_47266,N_47310);
nor UO_602 (O_602,N_48793,N_45062);
and UO_603 (O_603,N_45955,N_47867);
nor UO_604 (O_604,N_46583,N_45723);
or UO_605 (O_605,N_46027,N_49107);
nor UO_606 (O_606,N_47687,N_48471);
nor UO_607 (O_607,N_45695,N_49322);
xnor UO_608 (O_608,N_49565,N_48607);
nor UO_609 (O_609,N_47062,N_45713);
and UO_610 (O_610,N_47267,N_47427);
nand UO_611 (O_611,N_45634,N_49556);
and UO_612 (O_612,N_47871,N_49279);
or UO_613 (O_613,N_46934,N_48220);
nor UO_614 (O_614,N_49161,N_45236);
or UO_615 (O_615,N_45476,N_49563);
nor UO_616 (O_616,N_47409,N_47669);
and UO_617 (O_617,N_46920,N_49144);
nor UO_618 (O_618,N_46810,N_49826);
or UO_619 (O_619,N_46050,N_49219);
and UO_620 (O_620,N_49022,N_47475);
or UO_621 (O_621,N_48656,N_46210);
and UO_622 (O_622,N_49321,N_49249);
nor UO_623 (O_623,N_45655,N_48041);
and UO_624 (O_624,N_45035,N_48800);
nor UO_625 (O_625,N_45235,N_49268);
nor UO_626 (O_626,N_48579,N_45260);
or UO_627 (O_627,N_49681,N_45113);
nand UO_628 (O_628,N_49442,N_49292);
nor UO_629 (O_629,N_46124,N_47763);
or UO_630 (O_630,N_45943,N_49197);
nand UO_631 (O_631,N_47410,N_47262);
or UO_632 (O_632,N_45541,N_45454);
and UO_633 (O_633,N_45550,N_46999);
and UO_634 (O_634,N_48728,N_45311);
and UO_635 (O_635,N_48191,N_49018);
or UO_636 (O_636,N_48150,N_49247);
nor UO_637 (O_637,N_45818,N_48052);
nand UO_638 (O_638,N_46268,N_48772);
and UO_639 (O_639,N_47582,N_46358);
and UO_640 (O_640,N_47877,N_45505);
and UO_641 (O_641,N_47673,N_45163);
and UO_642 (O_642,N_49842,N_45543);
nand UO_643 (O_643,N_46427,N_48332);
nor UO_644 (O_644,N_46223,N_45564);
nor UO_645 (O_645,N_45102,N_49954);
nand UO_646 (O_646,N_47423,N_49203);
nor UO_647 (O_647,N_46504,N_46636);
and UO_648 (O_648,N_47548,N_47882);
nor UO_649 (O_649,N_47425,N_45316);
and UO_650 (O_650,N_47159,N_47876);
and UO_651 (O_651,N_49696,N_49202);
xor UO_652 (O_652,N_48235,N_45773);
nor UO_653 (O_653,N_45305,N_47231);
and UO_654 (O_654,N_45509,N_48446);
nand UO_655 (O_655,N_45238,N_47820);
and UO_656 (O_656,N_48139,N_47860);
nand UO_657 (O_657,N_45067,N_46511);
xor UO_658 (O_658,N_46084,N_47773);
or UO_659 (O_659,N_46199,N_47355);
nor UO_660 (O_660,N_45784,N_45738);
nand UO_661 (O_661,N_47651,N_47304);
nor UO_662 (O_662,N_47497,N_46137);
nand UO_663 (O_663,N_46413,N_48718);
or UO_664 (O_664,N_48289,N_46297);
and UO_665 (O_665,N_45185,N_45416);
nor UO_666 (O_666,N_47890,N_47808);
or UO_667 (O_667,N_48282,N_47725);
and UO_668 (O_668,N_48730,N_49660);
xor UO_669 (O_669,N_48965,N_46646);
or UO_670 (O_670,N_48755,N_49053);
or UO_671 (O_671,N_46773,N_45744);
xor UO_672 (O_672,N_45436,N_47122);
nor UO_673 (O_673,N_48514,N_48015);
nand UO_674 (O_674,N_49302,N_49600);
and UO_675 (O_675,N_49383,N_49500);
xor UO_676 (O_676,N_48309,N_45963);
nor UO_677 (O_677,N_49636,N_45860);
nand UO_678 (O_678,N_49165,N_49263);
and UO_679 (O_679,N_47326,N_49931);
xor UO_680 (O_680,N_48302,N_47048);
nand UO_681 (O_681,N_45841,N_45061);
nand UO_682 (O_682,N_48027,N_48796);
and UO_683 (O_683,N_48662,N_48337);
xnor UO_684 (O_684,N_49525,N_45578);
nand UO_685 (O_685,N_47354,N_49409);
and UO_686 (O_686,N_46253,N_48394);
nor UO_687 (O_687,N_47301,N_45472);
or UO_688 (O_688,N_48036,N_47126);
or UO_689 (O_689,N_46125,N_49498);
xnor UO_690 (O_690,N_49224,N_48643);
or UO_691 (O_691,N_45295,N_48880);
or UO_692 (O_692,N_46818,N_45909);
nor UO_693 (O_693,N_45139,N_49278);
nand UO_694 (O_694,N_46882,N_47208);
or UO_695 (O_695,N_48342,N_47526);
nand UO_696 (O_696,N_45497,N_46459);
nand UO_697 (O_697,N_48364,N_46245);
nor UO_698 (O_698,N_48508,N_47395);
nand UO_699 (O_699,N_48930,N_48465);
or UO_700 (O_700,N_45001,N_46406);
and UO_701 (O_701,N_47435,N_48935);
and UO_702 (O_702,N_47371,N_45555);
or UO_703 (O_703,N_45112,N_47171);
xor UO_704 (O_704,N_49694,N_46219);
nand UO_705 (O_705,N_46175,N_49172);
nand UO_706 (O_706,N_48236,N_46852);
and UO_707 (O_707,N_45107,N_49938);
and UO_708 (O_708,N_47361,N_46620);
and UO_709 (O_709,N_47661,N_47690);
nand UO_710 (O_710,N_49774,N_46368);
nand UO_711 (O_711,N_47948,N_48925);
nor UO_712 (O_712,N_45483,N_48079);
nand UO_713 (O_713,N_49005,N_45003);
nor UO_714 (O_714,N_46808,N_48039);
and UO_715 (O_715,N_47902,N_48205);
and UO_716 (O_716,N_46047,N_47992);
nand UO_717 (O_717,N_47466,N_49851);
or UO_718 (O_718,N_45946,N_46855);
nor UO_719 (O_719,N_49408,N_49155);
and UO_720 (O_720,N_48559,N_45961);
and UO_721 (O_721,N_48834,N_46610);
nor UO_722 (O_722,N_48641,N_46437);
nand UO_723 (O_723,N_49431,N_46644);
nand UO_724 (O_724,N_49127,N_48061);
nand UO_725 (O_725,N_48073,N_46415);
and UO_726 (O_726,N_47731,N_46434);
or UO_727 (O_727,N_47547,N_47691);
and UO_728 (O_728,N_49394,N_45806);
and UO_729 (O_729,N_48470,N_49424);
or UO_730 (O_730,N_45372,N_47465);
nor UO_731 (O_731,N_47608,N_48263);
nand UO_732 (O_732,N_45447,N_46276);
xor UO_733 (O_733,N_49731,N_46031);
or UO_734 (O_734,N_49669,N_49634);
nor UO_735 (O_735,N_47677,N_48319);
xor UO_736 (O_736,N_45519,N_47230);
or UO_737 (O_737,N_47827,N_45781);
nor UO_738 (O_738,N_49110,N_46721);
nor UO_739 (O_739,N_49883,N_47434);
xor UO_740 (O_740,N_48953,N_45771);
nor UO_741 (O_741,N_45896,N_48621);
nand UO_742 (O_742,N_45748,N_48055);
nor UO_743 (O_743,N_48761,N_48459);
xnor UO_744 (O_744,N_49404,N_48315);
or UO_745 (O_745,N_47996,N_45852);
xnor UO_746 (O_746,N_45438,N_45296);
nand UO_747 (O_747,N_48626,N_45610);
nand UO_748 (O_748,N_49793,N_46735);
and UO_749 (O_749,N_46104,N_46969);
and UO_750 (O_750,N_46948,N_48829);
nand UO_751 (O_751,N_45231,N_49092);
xnor UO_752 (O_752,N_48631,N_48639);
nor UO_753 (O_753,N_46777,N_45504);
or UO_754 (O_754,N_46665,N_49905);
xnor UO_755 (O_755,N_48008,N_49163);
nor UO_756 (O_756,N_47388,N_48044);
or UO_757 (O_757,N_46321,N_46344);
or UO_758 (O_758,N_48753,N_48975);
or UO_759 (O_759,N_48221,N_45724);
nor UO_760 (O_760,N_45022,N_47917);
or UO_761 (O_761,N_47730,N_48198);
and UO_762 (O_762,N_45768,N_49976);
nand UO_763 (O_763,N_48352,N_48028);
or UO_764 (O_764,N_48467,N_46136);
nand UO_765 (O_765,N_45282,N_47439);
and UO_766 (O_766,N_49356,N_49962);
nor UO_767 (O_767,N_45118,N_48967);
nand UO_768 (O_768,N_49069,N_47715);
nor UO_769 (O_769,N_48264,N_46702);
or UO_770 (O_770,N_47485,N_47474);
or UO_771 (O_771,N_48845,N_49156);
xor UO_772 (O_772,N_46886,N_47206);
or UO_773 (O_773,N_48476,N_47612);
nand UO_774 (O_774,N_45737,N_48001);
nor UO_775 (O_775,N_45574,N_49162);
and UO_776 (O_776,N_49311,N_45261);
xor UO_777 (O_777,N_47327,N_49338);
or UO_778 (O_778,N_46661,N_48575);
or UO_779 (O_779,N_48384,N_46034);
nor UO_780 (O_780,N_45971,N_46711);
or UO_781 (O_781,N_49640,N_48848);
and UO_782 (O_782,N_47133,N_45952);
xor UO_783 (O_783,N_46376,N_49742);
nor UO_784 (O_784,N_47003,N_45632);
nand UO_785 (O_785,N_48637,N_48234);
nor UO_786 (O_786,N_48092,N_46970);
or UO_787 (O_787,N_47102,N_49572);
or UO_788 (O_788,N_45209,N_45468);
and UO_789 (O_789,N_48094,N_47375);
nor UO_790 (O_790,N_46239,N_47167);
nand UO_791 (O_791,N_48182,N_48920);
nor UO_792 (O_792,N_47148,N_47051);
nor UO_793 (O_793,N_47544,N_48177);
nand UO_794 (O_794,N_45121,N_49708);
or UO_795 (O_795,N_46978,N_46414);
or UO_796 (O_796,N_45033,N_45560);
and UO_797 (O_797,N_45580,N_45140);
nand UO_798 (O_798,N_46101,N_48966);
nand UO_799 (O_799,N_46193,N_48548);
and UO_800 (O_800,N_46221,N_45480);
nand UO_801 (O_801,N_45084,N_49281);
and UO_802 (O_802,N_47585,N_48894);
or UO_803 (O_803,N_49651,N_49345);
and UO_804 (O_804,N_46363,N_45321);
or UO_805 (O_805,N_47545,N_45647);
nand UO_806 (O_806,N_48461,N_48533);
nand UO_807 (O_807,N_48553,N_45871);
or UO_808 (O_808,N_45974,N_45435);
or UO_809 (O_809,N_48776,N_46215);
and UO_810 (O_810,N_48911,N_47516);
or UO_811 (O_811,N_46926,N_47350);
or UO_812 (O_812,N_48947,N_49054);
nand UO_813 (O_813,N_49986,N_47223);
or UO_814 (O_814,N_47892,N_47941);
nor UO_815 (O_815,N_45805,N_49026);
nor UO_816 (O_816,N_46553,N_46168);
and UO_817 (O_817,N_45344,N_46243);
nor UO_818 (O_818,N_45763,N_46668);
nand UO_819 (O_819,N_48402,N_46469);
or UO_820 (O_820,N_47942,N_48991);
nand UO_821 (O_821,N_45537,N_49204);
nand UO_822 (O_822,N_48490,N_47274);
or UO_823 (O_823,N_46570,N_48811);
or UO_824 (O_824,N_47068,N_48120);
and UO_825 (O_825,N_47531,N_46834);
nand UO_826 (O_826,N_49066,N_46667);
and UO_827 (O_827,N_46155,N_46057);
nand UO_828 (O_828,N_45873,N_47443);
and UO_829 (O_829,N_49001,N_48868);
and UO_830 (O_830,N_45226,N_45150);
nor UO_831 (O_831,N_47950,N_47173);
nor UO_832 (O_832,N_48872,N_49504);
nor UO_833 (O_833,N_48797,N_48038);
nand UO_834 (O_834,N_45128,N_46157);
nor UO_835 (O_835,N_49798,N_45523);
nand UO_836 (O_836,N_46850,N_48926);
nand UO_837 (O_837,N_49346,N_47729);
nor UO_838 (O_838,N_45071,N_48000);
xor UO_839 (O_839,N_45799,N_45532);
or UO_840 (O_840,N_49331,N_48393);
nor UO_841 (O_841,N_45477,N_49788);
nor UO_842 (O_842,N_45485,N_45448);
nand UO_843 (O_843,N_48466,N_48031);
or UO_844 (O_844,N_49117,N_49441);
nor UO_845 (O_845,N_46100,N_46994);
and UO_846 (O_846,N_45716,N_47207);
and UO_847 (O_847,N_47142,N_49507);
or UO_848 (O_848,N_48529,N_45164);
or UO_849 (O_849,N_48306,N_49351);
nor UO_850 (O_850,N_46847,N_49928);
nor UO_851 (O_851,N_47467,N_46373);
and UO_852 (O_852,N_45596,N_48972);
or UO_853 (O_853,N_48859,N_49538);
xor UO_854 (O_854,N_49444,N_48707);
nand UO_855 (O_855,N_49341,N_45777);
nand UO_856 (O_856,N_49925,N_45028);
and UO_857 (O_857,N_49448,N_46539);
nor UO_858 (O_858,N_47378,N_47679);
nand UO_859 (O_859,N_47987,N_45976);
or UO_860 (O_860,N_47529,N_47914);
nor UO_861 (O_861,N_49235,N_45859);
and UO_862 (O_862,N_45746,N_49060);
or UO_863 (O_863,N_47085,N_45126);
nor UO_864 (O_864,N_49688,N_48963);
xnor UO_865 (O_865,N_45388,N_45085);
nand UO_866 (O_866,N_48881,N_49786);
or UO_867 (O_867,N_47345,N_46555);
nor UO_868 (O_868,N_46407,N_48404);
or UO_869 (O_869,N_48408,N_49385);
xor UO_870 (O_870,N_46839,N_45017);
nor UO_871 (O_871,N_46021,N_49384);
or UO_872 (O_872,N_45709,N_48870);
nand UO_873 (O_873,N_45750,N_46849);
nand UO_874 (O_874,N_47251,N_45405);
nor UO_875 (O_875,N_47685,N_48174);
nor UO_876 (O_876,N_46717,N_47586);
nand UO_877 (O_877,N_49849,N_48286);
and UO_878 (O_878,N_48824,N_47101);
nand UO_879 (O_879,N_45332,N_45384);
xnor UO_880 (O_880,N_46083,N_45047);
nor UO_881 (O_881,N_48988,N_47255);
and UO_882 (O_882,N_46325,N_46108);
xnor UO_883 (O_883,N_45802,N_49912);
or UO_884 (O_884,N_49059,N_46957);
and UO_885 (O_885,N_46148,N_47964);
nor UO_886 (O_886,N_49206,N_49376);
and UO_887 (O_887,N_49691,N_48922);
nand UO_888 (O_888,N_46003,N_48292);
and UO_889 (O_889,N_45218,N_46939);
nor UO_890 (O_890,N_45757,N_45533);
or UO_891 (O_891,N_45552,N_47736);
nor UO_892 (O_892,N_46609,N_47546);
or UO_893 (O_893,N_46183,N_45064);
and UO_894 (O_894,N_48477,N_45225);
nand UO_895 (O_895,N_47812,N_47983);
and UO_896 (O_896,N_45835,N_46822);
and UO_897 (O_897,N_48214,N_47252);
xor UO_898 (O_898,N_48021,N_45200);
and UO_899 (O_899,N_45794,N_46278);
nor UO_900 (O_900,N_46525,N_46252);
and UO_901 (O_901,N_46911,N_49610);
nor UO_902 (O_902,N_45947,N_48711);
and UO_903 (O_903,N_46005,N_45146);
xor UO_904 (O_904,N_46257,N_48133);
nor UO_905 (O_905,N_48014,N_45637);
nor UO_906 (O_906,N_49922,N_48022);
or UO_907 (O_907,N_45324,N_49037);
nand UO_908 (O_908,N_46694,N_47620);
or UO_909 (O_909,N_47553,N_48293);
nor UO_910 (O_910,N_47020,N_49140);
nand UO_911 (O_911,N_46774,N_47989);
or UO_912 (O_912,N_48308,N_47031);
nand UO_913 (O_913,N_47595,N_48363);
and UO_914 (O_914,N_46138,N_49002);
or UO_915 (O_915,N_48168,N_46428);
or UO_916 (O_916,N_48503,N_46631);
nor UO_917 (O_917,N_49867,N_47576);
xor UO_918 (O_918,N_49344,N_48654);
nor UO_919 (O_919,N_49894,N_47127);
xnor UO_920 (O_920,N_47160,N_48667);
nand UO_921 (O_921,N_48267,N_46002);
nor UO_922 (O_922,N_47492,N_49306);
nand UO_923 (O_923,N_47195,N_45960);
nor UO_924 (O_924,N_49692,N_47478);
nand UO_925 (O_925,N_46426,N_46317);
and UO_926 (O_926,N_45576,N_45522);
and UO_927 (O_927,N_49143,N_45420);
or UO_928 (O_928,N_47344,N_46338);
nor UO_929 (O_929,N_47575,N_48361);
or UO_930 (O_930,N_47013,N_45558);
nor UO_931 (O_931,N_47334,N_49763);
or UO_932 (O_932,N_46039,N_47486);
xor UO_933 (O_933,N_47684,N_47555);
nand UO_934 (O_934,N_46600,N_45317);
or UO_935 (O_935,N_49365,N_48698);
nor UO_936 (O_936,N_47511,N_48745);
xor UO_937 (O_937,N_47834,N_49419);
or UO_938 (O_938,N_48280,N_48217);
and UO_939 (O_939,N_45455,N_45674);
or UO_940 (O_940,N_46443,N_45602);
or UO_941 (O_941,N_46606,N_49589);
or UO_942 (O_942,N_47420,N_47581);
xnor UO_943 (O_943,N_48788,N_49418);
and UO_944 (O_944,N_49349,N_47798);
or UO_945 (O_945,N_45645,N_45834);
and UO_946 (O_946,N_48771,N_45938);
nor UO_947 (O_947,N_46931,N_47314);
and UO_948 (O_948,N_48497,N_46805);
or UO_949 (O_949,N_49324,N_48510);
and UO_950 (O_950,N_49336,N_45715);
and UO_951 (O_951,N_45034,N_47564);
nand UO_952 (O_952,N_48592,N_48297);
nor UO_953 (O_953,N_47540,N_48171);
xnor UO_954 (O_954,N_45516,N_45521);
nand UO_955 (O_955,N_48481,N_47445);
xnor UO_956 (O_956,N_45832,N_45755);
nor UO_957 (O_957,N_47046,N_49253);
nor UO_958 (O_958,N_46059,N_49327);
nor UO_959 (O_959,N_47398,N_45864);
nor UO_960 (O_960,N_49580,N_45136);
or UO_961 (O_961,N_45929,N_48980);
and UO_962 (O_962,N_45988,N_46263);
nor UO_963 (O_963,N_47746,N_47253);
nand UO_964 (O_964,N_46342,N_45267);
nand UO_965 (O_965,N_48003,N_46705);
nand UO_966 (O_966,N_46080,N_45005);
nor UO_967 (O_967,N_45154,N_48949);
xor UO_968 (O_968,N_48043,N_46764);
nor UO_969 (O_969,N_46547,N_46696);
or UO_970 (O_970,N_48789,N_47541);
nand UO_971 (O_971,N_45065,N_46298);
nor UO_972 (O_972,N_47572,N_48240);
or UO_973 (O_973,N_49364,N_45703);
nand UO_974 (O_974,N_45229,N_49630);
nand UO_975 (O_975,N_45091,N_46785);
and UO_976 (O_976,N_48193,N_45370);
or UO_977 (O_977,N_49936,N_45693);
and UO_978 (O_978,N_48137,N_45009);
and UO_979 (O_979,N_47926,N_49033);
or UO_980 (O_980,N_45308,N_49079);
xnor UO_981 (O_981,N_49481,N_47342);
nor UO_982 (O_982,N_49350,N_49848);
or UO_983 (O_983,N_48636,N_47916);
and UO_984 (O_984,N_48914,N_48369);
and UO_985 (O_985,N_47970,N_49430);
nand UO_986 (O_986,N_48272,N_46510);
xnor UO_987 (O_987,N_49181,N_49904);
or UO_988 (O_988,N_49554,N_47322);
nor UO_989 (O_989,N_49604,N_46540);
and UO_990 (O_990,N_49111,N_47588);
or UO_991 (O_991,N_47738,N_46404);
and UO_992 (O_992,N_46169,N_47449);
nor UO_993 (O_993,N_49417,N_48757);
nand UO_994 (O_994,N_45141,N_45077);
xor UO_995 (O_995,N_49004,N_48296);
xor UO_996 (O_996,N_46477,N_49435);
and UO_997 (O_997,N_49014,N_46235);
and UO_998 (O_998,N_48457,N_49795);
nor UO_999 (O_999,N_45970,N_49315);
nor UO_1000 (O_1000,N_46473,N_45649);
and UO_1001 (O_1001,N_47758,N_47386);
or UO_1002 (O_1002,N_49609,N_47075);
nor UO_1003 (O_1003,N_47263,N_47781);
or UO_1004 (O_1004,N_45165,N_47733);
and UO_1005 (O_1005,N_47692,N_48409);
and UO_1006 (O_1006,N_47638,N_49393);
or UO_1007 (O_1007,N_47680,N_47154);
nor UO_1008 (O_1008,N_45735,N_46194);
nand UO_1009 (O_1009,N_47176,N_47672);
and UO_1010 (O_1010,N_49926,N_47049);
or UO_1011 (O_1011,N_48519,N_48840);
nand UO_1012 (O_1012,N_48254,N_47500);
nand UO_1013 (O_1013,N_46738,N_46046);
or UO_1014 (O_1014,N_48142,N_45341);
xor UO_1015 (O_1015,N_49071,N_48858);
nand UO_1016 (O_1016,N_45233,N_48543);
nor UO_1017 (O_1017,N_47329,N_46873);
nand UO_1018 (O_1018,N_49510,N_47720);
or UO_1019 (O_1019,N_49857,N_49944);
and UO_1020 (O_1020,N_49126,N_45323);
nor UO_1021 (O_1021,N_47782,N_46296);
nand UO_1022 (O_1022,N_45418,N_48646);
nor UO_1023 (O_1023,N_48222,N_48013);
xnor UO_1024 (O_1024,N_45721,N_49401);
nand UO_1025 (O_1025,N_48951,N_49643);
and UO_1026 (O_1026,N_45565,N_45173);
nand UO_1027 (O_1027,N_48770,N_49963);
nand UO_1028 (O_1028,N_46256,N_48266);
nand UO_1029 (O_1029,N_49737,N_49677);
nor UO_1030 (O_1030,N_48545,N_46394);
and UO_1031 (O_1031,N_46506,N_47332);
nand UO_1032 (O_1032,N_45548,N_47217);
and UO_1033 (O_1033,N_48835,N_49185);
xnor UO_1034 (O_1034,N_45753,N_45252);
and UO_1035 (O_1035,N_48939,N_49567);
or UO_1036 (O_1036,N_48774,N_49746);
xor UO_1037 (O_1037,N_47220,N_46928);
nor UO_1038 (O_1038,N_47858,N_45286);
or UO_1039 (O_1039,N_47276,N_48900);
nor UO_1040 (O_1040,N_46431,N_46544);
and UO_1041 (O_1041,N_46442,N_49034);
nor UO_1042 (O_1042,N_49537,N_47972);
or UO_1043 (O_1043,N_46685,N_48045);
nand UO_1044 (O_1044,N_47934,N_46267);
or UO_1045 (O_1045,N_48583,N_46854);
xnor UO_1046 (O_1046,N_46310,N_48211);
and UO_1047 (O_1047,N_45108,N_47442);
and UO_1048 (O_1048,N_46549,N_49520);
nor UO_1049 (O_1049,N_49257,N_48668);
nand UO_1050 (O_1050,N_46938,N_48541);
xor UO_1051 (O_1051,N_45174,N_45626);
nor UO_1052 (O_1052,N_45605,N_49298);
and UO_1053 (O_1053,N_45012,N_47979);
xnor UO_1054 (O_1054,N_48051,N_47394);
and UO_1055 (O_1055,N_49433,N_46590);
nor UO_1056 (O_1056,N_48628,N_46557);
nand UO_1057 (O_1057,N_49234,N_48874);
nor UO_1058 (O_1058,N_45547,N_49210);
xnor UO_1059 (O_1059,N_46690,N_45038);
nand UO_1060 (O_1060,N_47458,N_49840);
or UO_1061 (O_1061,N_47671,N_49712);
nor UO_1062 (O_1062,N_47799,N_49868);
nor UO_1063 (O_1063,N_47840,N_48059);
or UO_1064 (O_1064,N_46952,N_45845);
nor UO_1065 (O_1065,N_46780,N_49919);
nand UO_1066 (O_1066,N_47863,N_49222);
nor UO_1067 (O_1067,N_49566,N_46679);
or UO_1068 (O_1068,N_46361,N_46909);
or UO_1069 (O_1069,N_47596,N_49941);
nand UO_1070 (O_1070,N_46340,N_48418);
nand UO_1071 (O_1071,N_47494,N_46436);
or UO_1072 (O_1072,N_47912,N_48186);
or UO_1073 (O_1073,N_46598,N_47532);
or UO_1074 (O_1074,N_47872,N_46595);
nand UO_1075 (O_1075,N_48517,N_48527);
xor UO_1076 (O_1076,N_49212,N_48954);
and UO_1077 (O_1077,N_48847,N_48262);
nor UO_1078 (O_1078,N_48781,N_48212);
nor UO_1079 (O_1079,N_49050,N_49797);
nor UO_1080 (O_1080,N_49120,N_47740);
and UO_1081 (O_1081,N_45520,N_48468);
and UO_1082 (O_1082,N_45239,N_45093);
nor UO_1083 (O_1083,N_48433,N_45919);
nor UO_1084 (O_1084,N_48285,N_49063);
nor UO_1085 (O_1085,N_46261,N_46836);
nor UO_1086 (O_1086,N_48946,N_49529);
or UO_1087 (O_1087,N_45063,N_49180);
and UO_1088 (O_1088,N_48644,N_46803);
and UO_1089 (O_1089,N_47724,N_47775);
or UO_1090 (O_1090,N_48440,N_45989);
or UO_1091 (O_1091,N_47408,N_47389);
and UO_1092 (O_1092,N_48638,N_48323);
xnor UO_1093 (O_1093,N_49678,N_46290);
or UO_1094 (O_1094,N_49134,N_45208);
or UO_1095 (O_1095,N_48130,N_49074);
nor UO_1096 (O_1096,N_45158,N_48964);
nand UO_1097 (O_1097,N_49122,N_47739);
nand UO_1098 (O_1098,N_45124,N_45380);
xor UO_1099 (O_1099,N_48860,N_45648);
nand UO_1100 (O_1100,N_49471,N_47124);
nand UO_1101 (O_1101,N_48688,N_49828);
and UO_1102 (O_1102,N_48478,N_47421);
and UO_1103 (O_1103,N_46073,N_45453);
or UO_1104 (O_1104,N_45152,N_48819);
or UO_1105 (O_1105,N_49105,N_46656);
xnor UO_1106 (O_1106,N_48375,N_46582);
nand UO_1107 (O_1107,N_47399,N_49330);
nor UO_1108 (O_1108,N_49133,N_47593);
nor UO_1109 (O_1109,N_45167,N_48348);
nor UO_1110 (O_1110,N_49505,N_48706);
or UO_1111 (O_1111,N_49768,N_45998);
nor UO_1112 (O_1112,N_47606,N_48806);
or UO_1113 (O_1113,N_46008,N_47851);
nand UO_1114 (O_1114,N_46623,N_49388);
and UO_1115 (O_1115,N_45222,N_46880);
and UO_1116 (O_1116,N_48833,N_49254);
or UO_1117 (O_1117,N_49655,N_48225);
or UO_1118 (O_1118,N_48250,N_47331);
and UO_1119 (O_1119,N_46993,N_48841);
or UO_1120 (O_1120,N_48842,N_46857);
or UO_1121 (O_1121,N_46599,N_47594);
nand UO_1122 (O_1122,N_45319,N_46226);
or UO_1123 (O_1123,N_45982,N_45215);
and UO_1124 (O_1124,N_49061,N_46912);
nand UO_1125 (O_1125,N_47396,N_49593);
nor UO_1126 (O_1126,N_47583,N_49767);
nand UO_1127 (O_1127,N_46566,N_49652);
nand UO_1128 (O_1128,N_48320,N_49011);
or UO_1129 (O_1129,N_45694,N_49657);
nand UO_1130 (O_1130,N_46259,N_45633);
nor UO_1131 (O_1131,N_46865,N_48996);
and UO_1132 (O_1132,N_45996,N_47870);
nor UO_1133 (O_1133,N_45866,N_45728);
or UO_1134 (O_1134,N_49624,N_45849);
xor UO_1135 (O_1135,N_48090,N_48161);
nor UO_1136 (O_1136,N_46174,N_45922);
and UO_1137 (O_1137,N_49689,N_49465);
or UO_1138 (O_1138,N_48095,N_46085);
and UO_1139 (O_1139,N_46232,N_46965);
or UO_1140 (O_1140,N_46660,N_45902);
or UO_1141 (O_1141,N_45506,N_48170);
nor UO_1142 (O_1142,N_47459,N_46743);
nor UO_1143 (O_1143,N_45406,N_45401);
nand UO_1144 (O_1144,N_48391,N_46591);
nor UO_1145 (O_1145,N_49715,N_46492);
or UO_1146 (O_1146,N_48625,N_49360);
or UO_1147 (O_1147,N_46998,N_45459);
nand UO_1148 (O_1148,N_45466,N_49540);
xor UO_1149 (O_1149,N_48735,N_45170);
nand UO_1150 (O_1150,N_45869,N_47064);
or UO_1151 (O_1151,N_49412,N_47991);
nor UO_1152 (O_1152,N_48715,N_49511);
or UO_1153 (O_1153,N_47162,N_46095);
nand UO_1154 (O_1154,N_47734,N_47613);
nand UO_1155 (O_1155,N_47308,N_46637);
nor UO_1156 (O_1156,N_46666,N_45338);
nand UO_1157 (O_1157,N_45891,N_46102);
and UO_1158 (O_1158,N_46517,N_49452);
and UO_1159 (O_1159,N_48754,N_47507);
nand UO_1160 (O_1160,N_45510,N_47333);
nand UO_1161 (O_1161,N_46130,N_48970);
and UO_1162 (O_1162,N_46033,N_46596);
or UO_1163 (O_1163,N_49024,N_45362);
nand UO_1164 (O_1164,N_45002,N_48537);
xor UO_1165 (O_1165,N_49112,N_48566);
nor UO_1166 (O_1166,N_45783,N_46932);
nor UO_1167 (O_1167,N_45439,N_49947);
or UO_1168 (O_1168,N_46752,N_45389);
nor UO_1169 (O_1169,N_46845,N_45412);
and UO_1170 (O_1170,N_45650,N_49578);
and UO_1171 (O_1171,N_48851,N_48546);
nor UO_1172 (O_1172,N_48664,N_45660);
or UO_1173 (O_1173,N_49870,N_49559);
or UO_1174 (O_1174,N_45491,N_46863);
and UO_1175 (O_1175,N_46453,N_47104);
nor UO_1176 (O_1176,N_46305,N_48609);
nor UO_1177 (O_1177,N_45042,N_47647);
nand UO_1178 (O_1178,N_45881,N_46351);
nand UO_1179 (O_1179,N_48552,N_48153);
and UO_1180 (O_1180,N_48231,N_47862);
nor UO_1181 (O_1181,N_49096,N_45636);
and UO_1182 (O_1182,N_46771,N_47562);
and UO_1183 (O_1183,N_47847,N_48889);
and UO_1184 (O_1184,N_48048,N_49539);
nor UO_1185 (O_1185,N_47844,N_46185);
or UO_1186 (O_1186,N_46883,N_45669);
nor UO_1187 (O_1187,N_48237,N_49673);
or UO_1188 (O_1188,N_49380,N_48197);
or UO_1189 (O_1189,N_46792,N_49459);
nand UO_1190 (O_1190,N_47839,N_49888);
nand UO_1191 (O_1191,N_46639,N_46971);
or UO_1192 (O_1192,N_49933,N_47197);
or UO_1193 (O_1193,N_49007,N_48809);
nand UO_1194 (O_1194,N_49524,N_47956);
nand UO_1195 (O_1195,N_49387,N_47236);
nor UO_1196 (O_1196,N_46421,N_48524);
or UO_1197 (O_1197,N_48902,N_49508);
or UO_1198 (O_1198,N_47113,N_49225);
nor UO_1199 (O_1199,N_48366,N_45304);
xnor UO_1200 (O_1200,N_49756,N_46984);
and UO_1201 (O_1201,N_47009,N_45690);
nor UO_1202 (O_1202,N_45630,N_45462);
or UO_1203 (O_1203,N_47433,N_47473);
nor UO_1204 (O_1204,N_48892,N_49512);
nand UO_1205 (O_1205,N_46417,N_48441);
or UO_1206 (O_1206,N_47036,N_47786);
nand UO_1207 (O_1207,N_48157,N_46218);
and UO_1208 (O_1208,N_46485,N_47103);
nand UO_1209 (O_1209,N_45911,N_47515);
nor UO_1210 (O_1210,N_46837,N_47209);
nor UO_1211 (O_1211,N_45097,N_49766);
nor UO_1212 (O_1212,N_49570,N_47070);
and UO_1213 (O_1213,N_46734,N_48389);
or UO_1214 (O_1214,N_46187,N_49902);
or UO_1215 (O_1215,N_49446,N_47073);
or UO_1216 (O_1216,N_47129,N_49882);
or UO_1217 (O_1217,N_46314,N_45563);
and UO_1218 (O_1218,N_46536,N_48982);
and UO_1219 (O_1219,N_49239,N_46659);
nor UO_1220 (O_1220,N_45843,N_48485);
nand UO_1221 (O_1221,N_49547,N_49906);
xnor UO_1222 (O_1222,N_46967,N_46332);
and UO_1223 (O_1223,N_47640,N_48081);
or UO_1224 (O_1224,N_47155,N_47134);
and UO_1225 (O_1225,N_46804,N_49332);
nand UO_1226 (O_1226,N_46638,N_45255);
or UO_1227 (O_1227,N_48830,N_48502);
and UO_1228 (O_1228,N_47219,N_48317);
nand UO_1229 (O_1229,N_46217,N_45381);
nor UO_1230 (O_1230,N_46328,N_49804);
and UO_1231 (O_1231,N_49237,N_45792);
and UO_1232 (O_1232,N_46568,N_46457);
or UO_1233 (O_1233,N_48499,N_48140);
nand UO_1234 (O_1234,N_46275,N_47528);
or UO_1235 (O_1235,N_46341,N_45898);
or UO_1236 (O_1236,N_45700,N_46951);
and UO_1237 (O_1237,N_47705,N_49490);
nand UO_1238 (O_1238,N_49865,N_47280);
or UO_1239 (O_1239,N_45014,N_48683);
or UO_1240 (O_1240,N_49334,N_45706);
xor UO_1241 (O_1241,N_47819,N_49373);
or UO_1242 (O_1242,N_47264,N_49363);
nand UO_1243 (O_1243,N_47416,N_49357);
xnor UO_1244 (O_1244,N_49819,N_48232);
nand UO_1245 (O_1245,N_47377,N_49467);
and UO_1246 (O_1246,N_49314,N_47609);
xor UO_1247 (O_1247,N_47105,N_49598);
or UO_1248 (O_1248,N_48380,N_47193);
nand UO_1249 (O_1249,N_49724,N_47879);
xor UO_1250 (O_1250,N_47759,N_48593);
xor UO_1251 (O_1251,N_45502,N_47496);
xnor UO_1252 (O_1252,N_45396,N_46871);
nor UO_1253 (O_1253,N_47004,N_45941);
nor UO_1254 (O_1254,N_45861,N_48213);
nor UO_1255 (O_1255,N_47683,N_49711);
nand UO_1256 (O_1256,N_46753,N_47809);
nor UO_1257 (O_1257,N_46958,N_47771);
or UO_1258 (O_1258,N_48278,N_49790);
nor UO_1259 (O_1259,N_45839,N_48345);
or UO_1260 (O_1260,N_46772,N_49308);
nor UO_1261 (O_1261,N_47832,N_46162);
nand UO_1262 (O_1262,N_46082,N_47138);
nand UO_1263 (O_1263,N_47242,N_48697);
nand UO_1264 (O_1264,N_47598,N_49265);
xor UO_1265 (O_1265,N_45876,N_46831);
nor UO_1266 (O_1266,N_48265,N_48838);
nand UO_1267 (O_1267,N_49517,N_46560);
and UO_1268 (O_1268,N_47261,N_46190);
nand UO_1269 (O_1269,N_49977,N_47796);
nor UO_1270 (O_1270,N_45854,N_46843);
nand UO_1271 (O_1271,N_49347,N_49282);
and UO_1272 (O_1272,N_47664,N_46840);
xnor UO_1273 (O_1273,N_47244,N_46801);
nand UO_1274 (O_1274,N_48696,N_45591);
and UO_1275 (O_1275,N_47259,N_45331);
nand UO_1276 (O_1276,N_47975,N_47041);
nor UO_1277 (O_1277,N_46754,N_46023);
or UO_1278 (O_1278,N_46781,N_49220);
nor UO_1279 (O_1279,N_45353,N_49545);
nand UO_1280 (O_1280,N_45144,N_47040);
nand UO_1281 (O_1281,N_49553,N_47793);
and UO_1282 (O_1282,N_45797,N_45300);
or UO_1283 (O_1283,N_46787,N_45279);
nand UO_1284 (O_1284,N_49923,N_49301);
and UO_1285 (O_1285,N_49166,N_46356);
and UO_1286 (O_1286,N_47614,N_47294);
nor UO_1287 (O_1287,N_45889,N_49667);
nor UO_1288 (O_1288,N_46116,N_46233);
or UO_1289 (O_1289,N_48307,N_48605);
or UO_1290 (O_1290,N_48528,N_45821);
xor UO_1291 (O_1291,N_48538,N_49557);
nor UO_1292 (O_1292,N_47822,N_47631);
nor UO_1293 (O_1293,N_45761,N_47968);
xor UO_1294 (O_1294,N_47131,N_46119);
nor UO_1295 (O_1295,N_48713,N_46601);
and UO_1296 (O_1296,N_48165,N_48206);
and UO_1297 (O_1297,N_45581,N_48324);
or UO_1298 (O_1298,N_48826,N_48373);
nor UO_1299 (O_1299,N_48836,N_45360);
and UO_1300 (O_1300,N_49289,N_46299);
or UO_1301 (O_1301,N_48760,N_45865);
nor UO_1302 (O_1302,N_48986,N_45778);
or UO_1303 (O_1303,N_45354,N_48802);
nor UO_1304 (O_1304,N_47921,N_48447);
nand UO_1305 (O_1305,N_47112,N_49601);
nor UO_1306 (O_1306,N_49637,N_49915);
and UO_1307 (O_1307,N_45484,N_48632);
nand UO_1308 (O_1308,N_48203,N_48333);
or UO_1309 (O_1309,N_47518,N_48376);
nand UO_1310 (O_1310,N_49468,N_47797);
and UO_1311 (O_1311,N_49228,N_45556);
or UO_1312 (O_1312,N_45813,N_47883);
xnor UO_1313 (O_1313,N_47452,N_45247);
xor UO_1314 (O_1314,N_48909,N_49017);
nand UO_1315 (O_1315,N_45673,N_45414);
and UO_1316 (O_1316,N_45856,N_46565);
or UO_1317 (O_1317,N_49506,N_45363);
and UO_1318 (O_1318,N_49403,N_49648);
nand UO_1319 (O_1319,N_49825,N_48917);
or UO_1320 (O_1320,N_46986,N_45868);
and UO_1321 (O_1321,N_46070,N_46482);
xnor UO_1322 (O_1322,N_45874,N_45000);
or UO_1323 (O_1323,N_46897,N_48682);
or UO_1324 (O_1324,N_48944,N_45019);
nor UO_1325 (O_1325,N_48790,N_48663);
nand UO_1326 (O_1326,N_48062,N_47117);
xor UO_1327 (O_1327,N_47761,N_46824);
and UO_1328 (O_1328,N_48400,N_46496);
or UO_1329 (O_1329,N_48766,N_47296);
nand UO_1330 (O_1330,N_45189,N_47707);
and UO_1331 (O_1331,N_45089,N_45284);
or UO_1332 (O_1332,N_47984,N_48396);
and UO_1333 (O_1333,N_48569,N_46744);
xor UO_1334 (O_1334,N_48019,N_47130);
nand UO_1335 (O_1335,N_48434,N_47269);
nand UO_1336 (O_1336,N_47237,N_49794);
and UO_1337 (O_1337,N_47780,N_48815);
and UO_1338 (O_1338,N_45984,N_49473);
and UO_1339 (O_1339,N_49082,N_47323);
or UO_1340 (O_1340,N_49397,N_48581);
nand UO_1341 (O_1341,N_48979,N_46309);
nor UO_1342 (O_1342,N_45726,N_48064);
nor UO_1343 (O_1343,N_47997,N_48056);
or UO_1344 (O_1344,N_45110,N_48940);
nand UO_1345 (O_1345,N_48741,N_48678);
nand UO_1346 (O_1346,N_46472,N_47063);
and UO_1347 (O_1347,N_49390,N_48734);
and UO_1348 (O_1348,N_47569,N_48500);
nand UO_1349 (O_1349,N_46015,N_46345);
nor UO_1350 (O_1350,N_49200,N_46704);
xnor UO_1351 (O_1351,N_49375,N_46399);
nor UO_1352 (O_1352,N_45036,N_46410);
and UO_1353 (O_1353,N_45194,N_48253);
or UO_1354 (O_1354,N_45916,N_45826);
or UO_1355 (O_1355,N_45940,N_46202);
nand UO_1356 (O_1356,N_47047,N_49093);
nor UO_1357 (O_1357,N_49890,N_48005);
or UO_1358 (O_1358,N_46548,N_48817);
and UO_1359 (O_1359,N_47764,N_47505);
nand UO_1360 (O_1360,N_46683,N_47258);
or UO_1361 (O_1361,N_49732,N_48763);
nor UO_1362 (O_1362,N_46567,N_45306);
and UO_1363 (O_1363,N_45692,N_49323);
or UO_1364 (O_1364,N_46500,N_46494);
nand UO_1365 (O_1365,N_46468,N_48419);
or UO_1366 (O_1366,N_45551,N_47464);
nand UO_1367 (O_1367,N_49789,N_47802);
nand UO_1368 (O_1368,N_49775,N_46480);
and UO_1369 (O_1369,N_45671,N_45553);
and UO_1370 (O_1370,N_46211,N_45105);
nand UO_1371 (O_1371,N_47510,N_48258);
nor UO_1372 (O_1372,N_46879,N_47320);
nand UO_1373 (O_1373,N_46502,N_48228);
nand UO_1374 (O_1374,N_45594,N_46389);
nor UO_1375 (O_1375,N_45294,N_48343);
nor UO_1376 (O_1376,N_47076,N_46575);
or UO_1377 (O_1377,N_45248,N_47487);
and UO_1378 (O_1378,N_46974,N_48379);
and UO_1379 (O_1379,N_48673,N_45400);
nand UO_1380 (O_1380,N_49142,N_46334);
and UO_1381 (O_1381,N_48655,N_46173);
nor UO_1382 (O_1382,N_48821,N_48572);
nand UO_1383 (O_1383,N_49751,N_47590);
nor UO_1384 (O_1384,N_48960,N_48748);
or UO_1385 (O_1385,N_49099,N_45351);
nand UO_1386 (O_1386,N_48912,N_46501);
nand UO_1387 (O_1387,N_49425,N_48099);
nand UO_1388 (O_1388,N_46538,N_49267);
nand UO_1389 (O_1389,N_47362,N_47957);
nor UO_1390 (O_1390,N_49611,N_48242);
and UO_1391 (O_1391,N_46076,N_48149);
and UO_1392 (O_1392,N_47653,N_45011);
nor UO_1393 (O_1393,N_45766,N_46204);
and UO_1394 (O_1394,N_45368,N_49319);
nor UO_1395 (O_1395,N_47319,N_45040);
xnor UO_1396 (O_1396,N_46242,N_49039);
xor UO_1397 (O_1397,N_47479,N_45530);
xor UO_1398 (O_1398,N_46923,N_45894);
xnor UO_1399 (O_1399,N_49458,N_45027);
and UO_1400 (O_1400,N_48879,N_45710);
or UO_1401 (O_1401,N_45157,N_49010);
nor UO_1402 (O_1402,N_45081,N_48740);
nand UO_1403 (O_1403,N_48146,N_49745);
nand UO_1404 (O_1404,N_46755,N_47422);
nand UO_1405 (O_1405,N_45575,N_48539);
nand UO_1406 (O_1406,N_47383,N_45833);
nor UO_1407 (O_1407,N_46673,N_46763);
nor UO_1408 (O_1408,N_45359,N_46121);
nand UO_1409 (O_1409,N_49470,N_47364);
and UO_1410 (O_1410,N_48416,N_49012);
nand UO_1411 (O_1411,N_46807,N_46182);
and UO_1412 (O_1412,N_48012,N_49186);
or UO_1413 (O_1413,N_48906,N_46112);
or UO_1414 (O_1414,N_49077,N_46423);
nand UO_1415 (O_1415,N_49488,N_45059);
nor UO_1416 (O_1416,N_49038,N_47533);
nor UO_1417 (O_1417,N_47850,N_45600);
and UO_1418 (O_1418,N_48810,N_47713);
nand UO_1419 (O_1419,N_49784,N_45375);
xnor UO_1420 (O_1420,N_48825,N_46980);
nand UO_1421 (O_1421,N_45847,N_46775);
nor UO_1422 (O_1422,N_47363,N_46114);
xnor UO_1423 (O_1423,N_45774,N_48853);
or UO_1424 (O_1424,N_47951,N_45855);
nor UO_1425 (O_1425,N_49949,N_49584);
nor UO_1426 (O_1426,N_49415,N_47483);
or UO_1427 (O_1427,N_45044,N_48121);
or UO_1428 (O_1428,N_48353,N_49070);
nor UO_1429 (O_1429,N_48110,N_48633);
nor UO_1430 (O_1430,N_45629,N_47976);
nand UO_1431 (O_1431,N_45910,N_47814);
xor UO_1432 (O_1432,N_49041,N_45672);
nand UO_1433 (O_1433,N_47865,N_47894);
nand UO_1434 (O_1434,N_47963,N_48814);
nand UO_1435 (O_1435,N_49800,N_49921);
and UO_1436 (O_1436,N_48011,N_46947);
xnor UO_1437 (O_1437,N_48657,N_46315);
nor UO_1438 (O_1438,N_46071,N_46044);
and UO_1439 (O_1439,N_47804,N_46966);
nand UO_1440 (O_1440,N_49920,N_47919);
xnor UO_1441 (O_1441,N_48923,N_45450);
and UO_1442 (O_1442,N_45862,N_49130);
or UO_1443 (O_1443,N_47373,N_49869);
or UO_1444 (O_1444,N_46126,N_47682);
and UO_1445 (O_1445,N_47552,N_48464);
or UO_1446 (O_1446,N_49352,N_45983);
or UO_1447 (O_1447,N_48115,N_49656);
nand UO_1448 (O_1448,N_48691,N_49861);
and UO_1449 (O_1449,N_48257,N_49588);
and UO_1450 (O_1450,N_48070,N_45776);
nor UO_1451 (O_1451,N_45451,N_47067);
or UO_1452 (O_1452,N_47666,N_48112);
or UO_1453 (O_1453,N_45473,N_46859);
nor UO_1454 (O_1454,N_46630,N_46343);
nor UO_1455 (O_1455,N_49276,N_48679);
xnor UO_1456 (O_1456,N_48327,N_48640);
nand UO_1457 (O_1457,N_48883,N_49191);
and UO_1458 (O_1458,N_46973,N_45050);
and UO_1459 (O_1459,N_46715,N_46161);
nand UO_1460 (O_1460,N_49672,N_47050);
and UO_1461 (O_1461,N_45931,N_46495);
nor UO_1462 (O_1462,N_47472,N_47592);
or UO_1463 (O_1463,N_45772,N_46446);
nor UO_1464 (O_1464,N_48807,N_49903);
nor UO_1465 (O_1465,N_46578,N_46374);
or UO_1466 (O_1466,N_48249,N_49832);
and UO_1467 (O_1467,N_48590,N_47463);
nand UO_1468 (O_1468,N_46716,N_45409);
and UO_1469 (O_1469,N_47368,N_49264);
nor UO_1470 (O_1470,N_46281,N_48489);
or UO_1471 (O_1471,N_47706,N_46386);
nor UO_1472 (O_1472,N_46024,N_46526);
or UO_1473 (O_1473,N_45262,N_46200);
or UO_1474 (O_1474,N_47750,N_46645);
or UO_1475 (O_1475,N_47887,N_48602);
or UO_1476 (O_1476,N_48574,N_45584);
and UO_1477 (O_1477,N_49723,N_45217);
nor UO_1478 (O_1478,N_46400,N_46490);
or UO_1479 (O_1479,N_46230,N_45815);
nor UO_1480 (O_1480,N_46602,N_46981);
or UO_1481 (O_1481,N_49176,N_46049);
nor UO_1482 (O_1482,N_46450,N_47097);
xor UO_1483 (O_1483,N_46895,N_49003);
nor UO_1484 (O_1484,N_45867,N_45213);
or UO_1485 (O_1485,N_45732,N_46179);
nand UO_1486 (O_1486,N_49478,N_48893);
and UO_1487 (O_1487,N_45283,N_45994);
or UO_1488 (O_1488,N_46017,N_47823);
nor UO_1489 (O_1489,N_45244,N_45392);
and UO_1490 (O_1490,N_49855,N_49617);
or UO_1491 (O_1491,N_47965,N_46106);
nor UO_1492 (O_1492,N_47069,N_48518);
nand UO_1493 (O_1493,N_48855,N_49492);
nor UO_1494 (O_1494,N_49661,N_49293);
or UO_1495 (O_1495,N_48813,N_49227);
nand UO_1496 (O_1496,N_45977,N_48162);
nand UO_1497 (O_1497,N_45070,N_48204);
or UO_1498 (O_1498,N_45702,N_47579);
or UO_1499 (O_1499,N_45441,N_46498);
nand UO_1500 (O_1500,N_46422,N_49423);
or UO_1501 (O_1501,N_46068,N_47404);
nor UO_1502 (O_1502,N_46641,N_48390);
or UO_1503 (O_1503,N_49807,N_47893);
and UO_1504 (O_1504,N_47755,N_48623);
or UO_1505 (O_1505,N_49622,N_47316);
nor UO_1506 (O_1506,N_46917,N_46258);
nor UO_1507 (O_1507,N_48762,N_49102);
nand UO_1508 (O_1508,N_46489,N_45993);
xor UO_1509 (O_1509,N_48955,N_49946);
xnor UO_1510 (O_1510,N_47856,N_47151);
or UO_1511 (O_1511,N_45281,N_49702);
nor UO_1512 (O_1512,N_48050,N_48270);
and UO_1513 (O_1513,N_49852,N_45026);
or UO_1514 (O_1514,N_45039,N_46887);
nor UO_1515 (O_1515,N_46167,N_48207);
xor UO_1516 (O_1516,N_49587,N_47514);
xnor UO_1517 (O_1517,N_45893,N_47370);
nor UO_1518 (O_1518,N_47658,N_46078);
and UO_1519 (O_1519,N_47776,N_46424);
nor UO_1520 (O_1520,N_46514,N_46260);
or UO_1521 (O_1521,N_48024,N_46176);
nor UO_1522 (O_1522,N_47641,N_45978);
and UO_1523 (O_1523,N_48160,N_48712);
xnor UO_1524 (O_1524,N_48010,N_48977);
or UO_1525 (O_1525,N_48629,N_47161);
nor UO_1526 (O_1526,N_47988,N_45358);
and UO_1527 (O_1527,N_49342,N_47828);
nand UO_1528 (O_1528,N_47429,N_46279);
nor UO_1529 (O_1529,N_47986,N_45950);
xnor UO_1530 (O_1530,N_46401,N_49854);
and UO_1531 (O_1531,N_45880,N_46603);
or UO_1532 (O_1532,N_49113,N_45642);
or UO_1533 (O_1533,N_46110,N_48226);
or UO_1534 (O_1534,N_46018,N_45092);
nand UO_1535 (O_1535,N_49796,N_45793);
xor UO_1536 (O_1536,N_45090,N_48273);
nand UO_1537 (O_1537,N_47909,N_47943);
or UO_1538 (O_1538,N_49879,N_47749);
or UO_1539 (O_1539,N_48498,N_48058);
nand UO_1540 (O_1540,N_45277,N_49822);
and UO_1541 (O_1541,N_48721,N_48736);
or UO_1542 (O_1542,N_49760,N_48227);
and UO_1543 (O_1543,N_46921,N_47215);
or UO_1544 (O_1544,N_45496,N_48438);
or UO_1545 (O_1545,N_46320,N_48584);
nor UO_1546 (O_1546,N_48103,N_45101);
and UO_1547 (O_1547,N_46255,N_49957);
nand UO_1548 (O_1548,N_45055,N_45122);
and UO_1549 (O_1549,N_47451,N_49658);
nor UO_1550 (O_1550,N_49047,N_45619);
nand UO_1551 (O_1551,N_46051,N_47937);
or UO_1552 (O_1552,N_45733,N_48351);
or UO_1553 (O_1553,N_45162,N_45948);
and UO_1554 (O_1554,N_47694,N_48437);
or UO_1555 (O_1555,N_48275,N_49169);
or UO_1556 (O_1556,N_45417,N_46491);
and UO_1557 (O_1557,N_49413,N_48687);
xnor UO_1558 (O_1558,N_48908,N_47693);
or UO_1559 (O_1559,N_49813,N_46941);
or UO_1560 (O_1560,N_48425,N_46593);
xnor UO_1561 (O_1561,N_46383,N_48600);
or UO_1562 (O_1562,N_47702,N_45478);
nand UO_1563 (O_1563,N_47115,N_46732);
xnor UO_1564 (O_1564,N_49983,N_46372);
or UO_1565 (O_1565,N_48582,N_46117);
and UO_1566 (O_1566,N_46586,N_47757);
and UO_1567 (O_1567,N_48492,N_48509);
or UO_1568 (O_1568,N_45932,N_47456);
nand UO_1569 (O_1569,N_48385,N_49675);
and UO_1570 (O_1570,N_48614,N_46339);
nor UO_1571 (O_1571,N_49823,N_46724);
nand UO_1572 (O_1572,N_49284,N_48786);
or UO_1573 (O_1573,N_45905,N_45048);
and UO_1574 (O_1574,N_46487,N_46113);
or UO_1575 (O_1575,N_48123,N_48612);
nor UO_1576 (O_1576,N_45882,N_49674);
or UO_1577 (O_1577,N_46616,N_48684);
nor UO_1578 (O_1578,N_48359,N_48246);
nor UO_1579 (O_1579,N_48196,N_46687);
nor UO_1580 (O_1580,N_48849,N_45514);
nor UO_1581 (O_1581,N_48785,N_48852);
or UO_1582 (O_1582,N_45722,N_47366);
and UO_1583 (O_1583,N_48180,N_48950);
nand UO_1584 (O_1584,N_46060,N_47852);
or UO_1585 (O_1585,N_49581,N_47915);
nor UO_1586 (O_1586,N_46949,N_48857);
nand UO_1587 (O_1587,N_48598,N_46357);
xor UO_1588 (O_1588,N_46933,N_49758);
nor UO_1589 (O_1589,N_46092,N_47298);
and UO_1590 (O_1590,N_48071,N_48060);
nor UO_1591 (O_1591,N_47357,N_49971);
nand UO_1592 (O_1592,N_48381,N_46676);
or UO_1593 (O_1593,N_47180,N_48556);
or UO_1594 (O_1594,N_48224,N_47723);
nor UO_1595 (O_1595,N_48665,N_45571);
or UO_1596 (O_1596,N_45877,N_47745);
xnor UO_1597 (O_1597,N_48025,N_47232);
nor UO_1598 (O_1598,N_47032,N_47788);
and UO_1599 (O_1599,N_46079,N_48281);
and UO_1600 (O_1600,N_49370,N_46067);
nand UO_1601 (O_1601,N_47846,N_49106);
or UO_1602 (O_1602,N_47417,N_45087);
and UO_1603 (O_1603,N_46032,N_48020);
and UO_1604 (O_1604,N_49874,N_46728);
or UO_1605 (O_1605,N_48535,N_46573);
or UO_1606 (O_1606,N_48974,N_47328);
nand UO_1607 (O_1607,N_47033,N_49633);
nand UO_1608 (O_1608,N_48284,N_49684);
or UO_1609 (O_1609,N_46784,N_47183);
nand UO_1610 (O_1610,N_46987,N_45892);
nand UO_1611 (O_1611,N_46420,N_46968);
or UO_1612 (O_1612,N_47202,N_47754);
xnor UO_1613 (O_1613,N_48420,N_45068);
or UO_1614 (O_1614,N_48127,N_48078);
nor UO_1615 (O_1615,N_48331,N_48928);
xor UO_1616 (O_1616,N_45142,N_46624);
and UO_1617 (O_1617,N_47457,N_49541);
nor UO_1618 (O_1618,N_49791,N_46925);
and UO_1619 (O_1619,N_49771,N_49961);
or UO_1620 (O_1620,N_49958,N_48472);
nor UO_1621 (O_1621,N_49514,N_45037);
nand UO_1622 (O_1622,N_47772,N_46899);
nand UO_1623 (O_1623,N_46330,N_45334);
nor UO_1624 (O_1624,N_48053,N_49558);
nor UO_1625 (O_1625,N_48501,N_46972);
nand UO_1626 (O_1626,N_45211,N_47953);
or UO_1627 (O_1627,N_48660,N_46380);
or UO_1628 (O_1628,N_48401,N_46470);
or UO_1629 (O_1629,N_48749,N_49248);
or UO_1630 (O_1630,N_46091,N_48201);
and UO_1631 (O_1631,N_46642,N_47165);
and UO_1632 (O_1632,N_47448,N_47530);
nor UO_1633 (O_1633,N_47045,N_46888);
or UO_1634 (O_1634,N_48595,N_48586);
and UO_1635 (O_1635,N_45076,N_49597);
or UO_1636 (O_1636,N_45290,N_47282);
nand UO_1637 (O_1637,N_47760,N_46950);
nor UO_1638 (O_1638,N_49207,N_46282);
nand UO_1639 (O_1639,N_48243,N_45116);
and UO_1640 (O_1640,N_48877,N_48087);
and UO_1641 (O_1641,N_49726,N_49629);
nand UO_1642 (O_1642,N_46316,N_45273);
and UO_1643 (O_1643,N_49550,N_46844);
and UO_1644 (O_1644,N_47527,N_49899);
xnor UO_1645 (O_1645,N_46864,N_48326);
and UO_1646 (O_1646,N_46201,N_49229);
or UO_1647 (O_1647,N_45129,N_45130);
and UO_1648 (O_1648,N_48913,N_46585);
xor UO_1649 (O_1649,N_46273,N_48990);
and UO_1650 (O_1650,N_46052,N_45471);
or UO_1651 (O_1651,N_46192,N_47949);
or UO_1652 (O_1652,N_46907,N_45176);
and UO_1653 (O_1653,N_45464,N_49496);
nand UO_1654 (O_1654,N_48077,N_46988);
xnor UO_1655 (O_1655,N_45595,N_45901);
or UO_1656 (O_1656,N_49535,N_47150);
nor UO_1657 (O_1657,N_46979,N_48726);
nand UO_1658 (O_1658,N_47059,N_49967);
or UO_1659 (O_1659,N_47560,N_49953);
nor UO_1660 (O_1660,N_48417,N_46142);
nor UO_1661 (O_1661,N_47254,N_46799);
nor UO_1662 (O_1662,N_47826,N_47042);
nor UO_1663 (O_1663,N_49343,N_48475);
nand UO_1664 (O_1664,N_45013,N_47321);
nand UO_1665 (O_1665,N_46265,N_49410);
or UO_1666 (O_1666,N_49021,N_45879);
or UO_1667 (O_1667,N_48775,N_48329);
nor UO_1668 (O_1668,N_46324,N_49779);
nand UO_1669 (O_1669,N_49187,N_47650);
and UO_1670 (O_1670,N_45432,N_49979);
and UO_1671 (O_1671,N_45539,N_49316);
or UO_1672 (O_1672,N_47589,N_47340);
nand UO_1673 (O_1673,N_49551,N_49056);
and UO_1674 (O_1674,N_48777,N_47501);
or UO_1675 (O_1675,N_45518,N_47289);
or UO_1676 (O_1676,N_46012,N_45494);
nand UO_1677 (O_1677,N_48719,N_49846);
or UO_1678 (O_1678,N_47022,N_48310);
nor UO_1679 (O_1679,N_48488,N_46036);
or UO_1680 (O_1680,N_47889,N_45804);
nor UO_1681 (O_1681,N_46543,N_45760);
nor UO_1682 (O_1682,N_48573,N_46512);
nor UO_1683 (O_1683,N_49262,N_47853);
or UO_1684 (O_1684,N_45810,N_45153);
nand UO_1685 (O_1685,N_48128,N_46991);
or UO_1686 (O_1686,N_47095,N_49440);
xnor UO_1687 (O_1687,N_47816,N_46147);
nand UO_1688 (O_1688,N_47330,N_46521);
nor UO_1689 (O_1689,N_45025,N_45053);
nor UO_1690 (O_1690,N_47939,N_48322);
nand UO_1691 (O_1691,N_49780,N_47157);
nand UO_1692 (O_1692,N_47106,N_45658);
nand UO_1693 (O_1693,N_49969,N_48647);
and UO_1694 (O_1694,N_45990,N_47903);
and UO_1695 (O_1695,N_46556,N_48350);
and UO_1696 (O_1696,N_45029,N_46212);
or UO_1697 (O_1697,N_46181,N_49215);
nand UO_1698 (O_1698,N_47356,N_48747);
nand UO_1699 (O_1699,N_47482,N_49103);
xor UO_1700 (O_1700,N_48355,N_46922);
and UO_1701 (O_1701,N_48244,N_49753);
and UO_1702 (O_1702,N_49910,N_49575);
and UO_1703 (O_1703,N_48413,N_45109);
and UO_1704 (O_1704,N_49709,N_49177);
nor UO_1705 (O_1705,N_46518,N_45659);
and UO_1706 (O_1706,N_46890,N_45117);
nand UO_1707 (O_1707,N_48978,N_46311);
and UO_1708 (O_1708,N_45402,N_46141);
and UO_1709 (O_1709,N_46826,N_46465);
or UO_1710 (O_1710,N_48173,N_49885);
nand UO_1711 (O_1711,N_45147,N_49592);
and UO_1712 (O_1712,N_48155,N_47352);
and UO_1713 (O_1713,N_49231,N_46156);
or UO_1714 (O_1714,N_46307,N_48587);
and UO_1715 (O_1715,N_47094,N_46629);
nor UO_1716 (O_1716,N_47239,N_45428);
and UO_1717 (O_1717,N_47520,N_47074);
and UO_1718 (O_1718,N_49477,N_47488);
or UO_1719 (O_1719,N_48948,N_46894);
nand UO_1720 (O_1720,N_49447,N_48649);
nand UO_1721 (O_1721,N_48816,N_47536);
nor UO_1722 (O_1722,N_45719,N_47667);
nor UO_1723 (O_1723,N_46869,N_45951);
and UO_1724 (O_1724,N_47044,N_47054);
or UO_1725 (O_1725,N_46393,N_47633);
and UO_1726 (O_1726,N_49615,N_45644);
nor UO_1727 (O_1727,N_47476,N_46333);
nand UO_1728 (O_1728,N_46561,N_47191);
nor UO_1729 (O_1729,N_49270,N_46691);
nand UO_1730 (O_1730,N_47469,N_46385);
and UO_1731 (O_1731,N_46384,N_47930);
or UO_1732 (O_1732,N_46326,N_49594);
nand UO_1733 (O_1733,N_46291,N_49009);
and UO_1734 (O_1734,N_49621,N_45098);
nor UO_1735 (O_1735,N_48885,N_45394);
nor UO_1736 (O_1736,N_47484,N_48773);
and UO_1737 (O_1737,N_48356,N_48371);
and UO_1738 (O_1738,N_49703,N_49523);
or UO_1739 (O_1739,N_48782,N_48938);
nand UO_1740 (O_1740,N_46010,N_48544);
nor UO_1741 (O_1741,N_45192,N_49562);
nand UO_1742 (O_1742,N_47088,N_45216);
or UO_1743 (O_1743,N_49728,N_47616);
nand UO_1744 (O_1744,N_46650,N_48714);
nand UO_1745 (O_1745,N_46229,N_45680);
and UO_1746 (O_1746,N_45328,N_49805);
xnor UO_1747 (O_1747,N_46884,N_49605);
nor UO_1748 (O_1748,N_48576,N_46225);
nand UO_1749 (O_1749,N_45598,N_47897);
nor UO_1750 (O_1750,N_45258,N_47192);
and UO_1751 (O_1751,N_47081,N_45608);
nand UO_1752 (O_1752,N_46308,N_46367);
and UO_1753 (O_1753,N_47663,N_48085);
xor UO_1754 (O_1754,N_45487,N_45956);
or UO_1755 (O_1755,N_45206,N_47091);
nand UO_1756 (O_1756,N_47233,N_49727);
xor UO_1757 (O_1757,N_45675,N_45178);
nor UO_1758 (O_1758,N_46028,N_49718);
nand UO_1759 (O_1759,N_46463,N_49167);
nand UO_1760 (O_1760,N_49698,N_45270);
xnor UO_1761 (O_1761,N_47999,N_48318);
and UO_1762 (O_1762,N_46409,N_47402);
nand UO_1763 (O_1763,N_48392,N_48820);
xnor UO_1764 (O_1764,N_47543,N_46823);
xnor UO_1765 (O_1765,N_46680,N_47181);
nand UO_1766 (O_1766,N_49451,N_49863);
nand UO_1767 (O_1767,N_45957,N_45840);
nor UO_1768 (O_1768,N_49707,N_48611);
or UO_1769 (O_1769,N_49339,N_45857);
nor UO_1770 (O_1770,N_47747,N_47817);
nand UO_1771 (O_1771,N_47831,N_48088);
or UO_1772 (O_1772,N_49160,N_46867);
nor UO_1773 (O_1773,N_45024,N_46030);
or UO_1774 (O_1774,N_47158,N_47279);
and UO_1775 (O_1775,N_49721,N_49773);
and UO_1776 (O_1776,N_45765,N_49255);
or UO_1777 (O_1777,N_46615,N_49052);
xnor UO_1778 (O_1778,N_47795,N_47446);
and UO_1779 (O_1779,N_45057,N_47605);
nand UO_1780 (O_1780,N_45954,N_45714);
nor UO_1781 (O_1781,N_48164,N_45531);
nor UO_1782 (O_1782,N_48823,N_48303);
and UO_1783 (O_1783,N_45875,N_47438);
nand UO_1784 (O_1784,N_49303,N_48181);
and UO_1785 (O_1785,N_49887,N_45151);
and UO_1786 (O_1786,N_46335,N_45917);
xnor UO_1787 (O_1787,N_45570,N_49564);
nand UO_1788 (O_1788,N_45111,N_46789);
nand UO_1789 (O_1789,N_45349,N_49150);
nor UO_1790 (O_1790,N_49333,N_46377);
nor UO_1791 (O_1791,N_46929,N_49710);
nand UO_1792 (O_1792,N_49251,N_47973);
or UO_1793 (O_1793,N_45828,N_45315);
nor UO_1794 (O_1794,N_46365,N_46054);
and UO_1795 (O_1795,N_49892,N_45684);
nor UO_1796 (O_1796,N_49450,N_47901);
nand UO_1797 (O_1797,N_45345,N_47184);
nand UO_1798 (O_1798,N_49608,N_49975);
or UO_1799 (O_1799,N_48805,N_46408);
nand UO_1800 (O_1800,N_48152,N_48971);
or UO_1801 (O_1801,N_49337,N_47065);
or UO_1802 (O_1802,N_45382,N_46178);
nand UO_1803 (O_1803,N_45944,N_46479);
nand UO_1804 (O_1804,N_46313,N_47873);
xor UO_1805 (O_1805,N_47998,N_48075);
nand UO_1806 (O_1806,N_48701,N_46382);
and UO_1807 (O_1807,N_46542,N_49625);
and UO_1808 (O_1808,N_47268,N_47523);
and UO_1809 (O_1809,N_47908,N_46622);
or UO_1810 (O_1810,N_47000,N_48615);
nor UO_1811 (O_1811,N_46378,N_49533);
xnor UO_1812 (O_1812,N_47774,N_48313);
and UO_1813 (O_1813,N_48268,N_49299);
nor UO_1814 (O_1814,N_49750,N_48074);
or UO_1815 (O_1815,N_47554,N_47954);
nor UO_1816 (O_1816,N_47503,N_49371);
nand UO_1817 (O_1817,N_45764,N_49820);
xor UO_1818 (O_1818,N_48430,N_46375);
nor UO_1819 (O_1819,N_47166,N_49392);
or UO_1820 (O_1820,N_45169,N_47704);
nand UO_1821 (O_1821,N_46725,N_47712);
or UO_1822 (O_1822,N_46391,N_46878);
nand UO_1823 (O_1823,N_45681,N_48135);
and UO_1824 (O_1824,N_49294,N_46960);
xnor UO_1825 (O_1825,N_48737,N_47855);
and UO_1826 (O_1826,N_47711,N_45927);
nor UO_1827 (O_1827,N_47719,N_47385);
nor UO_1828 (O_1828,N_45627,N_45848);
or UO_1829 (O_1829,N_46026,N_49068);
or UO_1830 (O_1830,N_47619,N_45010);
and UO_1831 (O_1831,N_48703,N_48184);
or UO_1832 (O_1832,N_48551,N_48445);
nand UO_1833 (O_1833,N_45301,N_47292);
and UO_1834 (O_1834,N_49457,N_49546);
or UO_1835 (O_1835,N_47896,N_45387);
or UO_1836 (O_1836,N_46452,N_49422);
nor UO_1837 (O_1837,N_45788,N_45682);
or UO_1838 (O_1838,N_48325,N_49646);
or UO_1839 (O_1839,N_46829,N_49045);
nand UO_1840 (O_1840,N_45021,N_48116);
or UO_1841 (O_1841,N_47525,N_46396);
or UO_1842 (O_1842,N_47550,N_46191);
xor UO_1843 (O_1843,N_46811,N_45407);
and UO_1844 (O_1844,N_49361,N_45250);
nand UO_1845 (O_1845,N_45906,N_45759);
nor UO_1846 (O_1846,N_45953,N_49939);
and UO_1847 (O_1847,N_47453,N_49199);
or UO_1848 (O_1848,N_49997,N_47502);
nand UO_1849 (O_1849,N_49561,N_46390);
nor UO_1850 (O_1850,N_45727,N_47260);
nor UO_1851 (O_1851,N_48007,N_48456);
nand UO_1852 (O_1852,N_47990,N_49991);
nor UO_1853 (O_1853,N_47339,N_46739);
nand UO_1854 (O_1854,N_45557,N_47411);
nor UO_1855 (O_1855,N_46402,N_46348);
nand UO_1856 (O_1856,N_47315,N_45415);
and UO_1857 (O_1857,N_49291,N_49896);
nand UO_1858 (O_1858,N_47082,N_48458);
nand UO_1859 (O_1859,N_47688,N_47624);
nand UO_1860 (O_1860,N_48958,N_46456);
nor UO_1861 (O_1861,N_45082,N_49406);
and UO_1862 (O_1862,N_45203,N_47777);
nor UO_1863 (O_1863,N_46016,N_45041);
or UO_1864 (O_1864,N_45825,N_47235);
xnor UO_1865 (O_1865,N_49310,N_45831);
nor UO_1866 (O_1866,N_48878,N_49297);
nand UO_1867 (O_1867,N_47674,N_46706);
nor UO_1868 (O_1868,N_48758,N_46640);
nand UO_1869 (O_1869,N_47353,N_46649);
or UO_1870 (O_1870,N_46870,N_46251);
xor UO_1871 (O_1871,N_46123,N_46177);
and UO_1872 (O_1872,N_45127,N_48936);
or UO_1873 (O_1873,N_48439,N_45123);
xnor UO_1874 (O_1874,N_45119,N_47317);
nor UO_1875 (O_1875,N_47785,N_45615);
and UO_1876 (O_1876,N_48887,N_46875);
nand UO_1877 (O_1877,N_45378,N_45979);
or UO_1878 (O_1878,N_49489,N_49679);
nand UO_1879 (O_1879,N_48554,N_48230);
nand UO_1880 (O_1880,N_49124,N_49668);
and UO_1881 (O_1881,N_46337,N_47080);
nand UO_1882 (O_1882,N_46963,N_47391);
or UO_1883 (O_1883,N_48808,N_46090);
xnor UO_1884 (O_1884,N_45635,N_45966);
or UO_1885 (O_1885,N_48335,N_46441);
and UO_1886 (O_1886,N_47336,N_49628);
or UO_1887 (O_1887,N_46756,N_45926);
nor UO_1888 (O_1888,N_46643,N_45887);
nor UO_1889 (O_1889,N_45190,N_47324);
nor UO_1890 (O_1890,N_45512,N_49030);
or UO_1891 (O_1891,N_45356,N_49641);
and UO_1892 (O_1892,N_48717,N_49223);
nor UO_1893 (O_1893,N_48987,N_49519);
nand UO_1894 (O_1894,N_48677,N_46449);
and UO_1895 (O_1895,N_46419,N_49704);
or UO_1896 (O_1896,N_45913,N_49335);
nor UO_1897 (O_1897,N_47028,N_45253);
xor UO_1898 (O_1898,N_49416,N_49850);
and UO_1899 (O_1899,N_45908,N_47111);
nor UO_1900 (O_1900,N_47947,N_47681);
or UO_1901 (O_1901,N_47175,N_48791);
nor UO_1902 (O_1902,N_46670,N_48709);
xor UO_1903 (O_1903,N_49362,N_48507);
nor UO_1904 (O_1904,N_47143,N_48624);
nand UO_1905 (O_1905,N_49089,N_49318);
xnor UO_1906 (O_1906,N_49243,N_47290);
or UO_1907 (O_1907,N_46392,N_46962);
and UO_1908 (O_1908,N_48962,N_49595);
and UO_1909 (O_1909,N_49568,N_45413);
nor UO_1910 (O_1910,N_45241,N_46285);
and UO_1911 (O_1911,N_47121,N_49996);
nand UO_1912 (O_1912,N_48560,N_45500);
nand UO_1913 (O_1913,N_45699,N_45458);
and UO_1914 (O_1914,N_47145,N_48693);
and UO_1915 (O_1915,N_47716,N_49824);
and UO_1916 (O_1916,N_47556,N_47744);
nor UO_1917 (O_1917,N_47966,N_47563);
nor UO_1918 (O_1918,N_46902,N_49328);
and UO_1919 (O_1919,N_48080,N_46269);
xor UO_1920 (O_1920,N_46105,N_45822);
nand UO_1921 (O_1921,N_49720,N_49031);
and UO_1922 (O_1922,N_45313,N_48065);
xor UO_1923 (O_1923,N_49948,N_49427);
nand UO_1924 (O_1924,N_47376,N_45625);
nand UO_1925 (O_1925,N_46571,N_46432);
nand UO_1926 (O_1926,N_48804,N_49029);
and UO_1927 (O_1927,N_45106,N_49035);
nor UO_1928 (O_1928,N_45393,N_47156);
nor UO_1929 (O_1929,N_46727,N_49764);
and UO_1930 (O_1930,N_46118,N_47019);
nand UO_1931 (O_1931,N_48542,N_46150);
or UO_1932 (O_1932,N_45775,N_45103);
nor UO_1933 (O_1933,N_45016,N_45280);
and UO_1934 (O_1934,N_48531,N_45886);
or UO_1935 (O_1935,N_47025,N_49286);
and UO_1936 (O_1936,N_49685,N_46460);
or UO_1937 (O_1937,N_45985,N_45934);
nand UO_1938 (O_1938,N_48113,N_48279);
nor UO_1939 (O_1939,N_49590,N_47367);
and UO_1940 (O_1940,N_48564,N_48929);
nor UO_1941 (O_1941,N_48029,N_49245);
xnor UO_1942 (O_1942,N_46128,N_45391);
and UO_1943 (O_1943,N_49020,N_47246);
or UO_1944 (O_1944,N_47309,N_45275);
nor UO_1945 (O_1945,N_49260,N_49148);
xor UO_1946 (O_1946,N_47107,N_46519);
nor UO_1947 (O_1947,N_48606,N_45536);
nor UO_1948 (O_1948,N_47806,N_49080);
or UO_1949 (O_1949,N_48783,N_46841);
and UO_1950 (O_1950,N_47985,N_45492);
and UO_1951 (O_1951,N_45397,N_46541);
or UO_1952 (O_1952,N_47656,N_48512);
nand UO_1953 (O_1953,N_45008,N_46533);
nand UO_1954 (O_1954,N_46992,N_45337);
and UO_1955 (O_1955,N_46209,N_47337);
xor UO_1956 (O_1956,N_49781,N_45838);
xor UO_1957 (O_1957,N_48294,N_45426);
nand UO_1958 (O_1958,N_48367,N_47969);
or UO_1959 (O_1959,N_47303,N_48794);
or UO_1960 (O_1960,N_45549,N_47426);
nor UO_1961 (O_1961,N_45972,N_48387);
nor UO_1962 (O_1962,N_48856,N_49806);
xor UO_1963 (O_1963,N_47221,N_49542);
nor UO_1964 (O_1964,N_47499,N_45361);
nor UO_1965 (O_1965,N_46861,N_47163);
nand UO_1966 (O_1966,N_48410,N_47904);
nor UO_1967 (O_1967,N_47551,N_48599);
nor UO_1968 (O_1968,N_49875,N_46197);
or UO_1969 (O_1969,N_48746,N_45364);
nor UO_1970 (O_1970,N_45968,N_45546);
or UO_1971 (O_1971,N_46152,N_46531);
and UO_1972 (O_1972,N_49285,N_48689);
xor UO_1973 (O_1973,N_49638,N_46592);
or UO_1974 (O_1974,N_47848,N_47539);
nor UO_1975 (O_1975,N_48195,N_48339);
and UO_1976 (O_1976,N_48666,N_49744);
xor UO_1977 (O_1977,N_49023,N_49300);
or UO_1978 (O_1978,N_49136,N_46433);
or UO_1979 (O_1979,N_48033,N_49209);
nand UO_1980 (O_1980,N_47043,N_46248);
nor UO_1981 (O_1981,N_49549,N_49420);
nor UO_1982 (O_1982,N_46164,N_45498);
xor UO_1983 (O_1983,N_45348,N_49421);
xnor UO_1984 (O_1984,N_45120,N_49649);
and UO_1985 (O_1985,N_49491,N_49653);
and UO_1986 (O_1986,N_48916,N_45329);
and UO_1987 (O_1987,N_45369,N_49179);
and UO_1988 (O_1988,N_47436,N_49752);
or UO_1989 (O_1989,N_49618,N_45205);
nand UO_1990 (O_1990,N_48124,N_45395);
nor UO_1991 (O_1991,N_47652,N_46144);
or UO_1992 (O_1992,N_46081,N_47629);
or UO_1993 (O_1993,N_45327,N_45237);
and UO_1994 (O_1994,N_47016,N_49428);
xor UO_1995 (O_1995,N_45343,N_47698);
and UO_1996 (O_1996,N_47837,N_46904);
or UO_1997 (O_1997,N_47200,N_49460);
nor UO_1998 (O_1998,N_47522,N_46654);
or UO_1999 (O_1999,N_47885,N_49814);
nand UO_2000 (O_2000,N_46954,N_49859);
xnor UO_2001 (O_2001,N_46761,N_46825);
nand UO_2002 (O_2002,N_46982,N_46736);
or UO_2003 (O_2003,N_45493,N_45342);
and UO_2004 (O_2004,N_48111,N_46236);
xnor UO_2005 (O_2005,N_49792,N_47792);
or UO_2006 (O_2006,N_45830,N_48724);
nor UO_2007 (O_2007,N_48875,N_45787);
or UO_2008 (O_2008,N_49527,N_47118);
or UO_2009 (O_2009,N_48067,N_46720);
xnor UO_2010 (O_2010,N_46961,N_47287);
and UO_2011 (O_2011,N_49749,N_48199);
and UO_2012 (O_2012,N_48097,N_47932);
nand UO_2013 (O_2013,N_49266,N_48571);
or UO_2014 (O_2014,N_48276,N_46129);
and UO_2015 (O_2015,N_46562,N_45808);
nor UO_2016 (O_2016,N_48694,N_45883);
or UO_2017 (O_2017,N_46953,N_46327);
nor UO_2018 (O_2018,N_49230,N_49109);
nor UO_2019 (O_2019,N_49591,N_46821);
nor UO_2020 (O_2020,N_46613,N_48886);
and UO_2021 (O_2021,N_47090,N_49659);
nand UO_2022 (O_2022,N_45193,N_47125);
or UO_2023 (O_2023,N_47517,N_49259);
nor UO_2024 (O_2024,N_48104,N_47335);
nor UO_2025 (O_2025,N_49236,N_49602);
nor UO_2026 (O_2026,N_49706,N_46798);
nor UO_2027 (O_2027,N_49856,N_46678);
or UO_2028 (O_2028,N_48869,N_45683);
and UO_2029 (O_2029,N_48484,N_49680);
nor UO_2030 (O_2030,N_48299,N_45437);
and UO_2031 (O_2031,N_45246,N_49612);
and UO_2032 (O_2032,N_49474,N_49214);
or UO_2033 (O_2033,N_49956,N_49190);
or UO_2034 (O_2034,N_47779,N_49772);
nand UO_2035 (O_2035,N_49193,N_46848);
xor UO_2036 (O_2036,N_45299,N_47886);
and UO_2037 (O_2037,N_45422,N_45180);
or UO_2038 (O_2038,N_48126,N_49487);
nor UO_2039 (O_2039,N_45457,N_47447);
and UO_2040 (O_2040,N_47506,N_48648);
nor UO_2041 (O_2041,N_46625,N_45641);
and UO_2042 (O_2042,N_47895,N_47599);
or UO_2043 (O_2043,N_46295,N_49987);
nand UO_2044 (O_2044,N_46096,N_46350);
nand UO_2045 (O_2045,N_45597,N_45463);
nand UO_2046 (O_2046,N_45058,N_45814);
nor UO_2047 (O_2047,N_48334,N_47898);
nor UO_2048 (O_2048,N_48233,N_45133);
and UO_2049 (O_2049,N_45918,N_48483);
nor UO_2050 (O_2050,N_46346,N_45796);
nand UO_2051 (O_2051,N_48188,N_48487);
or UO_2052 (O_2052,N_47709,N_48495);
or UO_2053 (O_2053,N_49326,N_48608);
or UO_2054 (O_2054,N_47079,N_45357);
and UO_2055 (O_2055,N_46989,N_47597);
and UO_2056 (O_2056,N_48057,N_48596);
nand UO_2057 (O_2057,N_47955,N_49121);
nand UO_2058 (O_2058,N_45620,N_45403);
nand UO_2059 (O_2059,N_47787,N_45080);
or UO_2060 (O_2060,N_49240,N_48610);
nor UO_2061 (O_2061,N_45143,N_45589);
nand UO_2062 (O_2062,N_46087,N_49895);
xnor UO_2063 (O_2063,N_48739,N_45842);
and UO_2064 (O_2064,N_45201,N_47172);
nor UO_2065 (O_2065,N_48591,N_46783);
nor UO_2066 (O_2066,N_46913,N_49355);
and UO_2067 (O_2067,N_47959,N_46709);
nor UO_2068 (O_2068,N_49993,N_46747);
nor UO_2069 (O_2069,N_49530,N_46159);
and UO_2070 (O_2070,N_45230,N_48601);
and UO_2071 (O_2071,N_48985,N_45820);
or UO_2072 (O_2072,N_49153,N_46120);
and UO_2073 (O_2073,N_45445,N_49084);
nand UO_2074 (O_2074,N_48613,N_45962);
and UO_2075 (O_2075,N_46809,N_48290);
nor UO_2076 (O_2076,N_47636,N_47768);
nand UO_2077 (O_2077,N_49701,N_46779);
nand UO_2078 (O_2078,N_46621,N_47800);
nand UO_2079 (O_2079,N_48370,N_46349);
nand UO_2080 (O_2080,N_45705,N_47224);
or UO_2081 (O_2081,N_45006,N_47607);
and UO_2082 (O_2082,N_48252,N_49585);
or UO_2083 (O_2083,N_47226,N_48742);
or UO_2084 (O_2084,N_46009,N_47006);
nand UO_2085 (O_2085,N_46689,N_47015);
nand UO_2086 (O_2086,N_49985,N_45656);
or UO_2087 (O_2087,N_45897,N_48752);
and UO_2088 (O_2088,N_49864,N_48779);
xnor UO_2089 (O_2089,N_45959,N_47086);
and UO_2090 (O_2090,N_45743,N_49128);
or UO_2091 (O_2091,N_49414,N_48767);
nor UO_2092 (O_2092,N_45870,N_47770);
nor UO_2093 (O_2093,N_45903,N_45379);
xor UO_2094 (O_2094,N_45623,N_47306);
nor UO_2095 (O_2095,N_45266,N_49182);
or UO_2096 (O_2096,N_46284,N_49932);
and UO_2097 (O_2097,N_49000,N_45318);
and UO_2098 (O_2098,N_49171,N_46180);
or UO_2099 (O_2099,N_45643,N_45844);
nand UO_2100 (O_2100,N_48117,N_45885);
and UO_2101 (O_2101,N_47710,N_46648);
and UO_2102 (O_2102,N_46876,N_49839);
and UO_2103 (O_2103,N_47900,N_48208);
nand UO_2104 (O_2104,N_49065,N_49980);
or UO_2105 (O_2105,N_46770,N_45708);
and UO_2106 (O_2106,N_46682,N_47689);
nand UO_2107 (O_2107,N_49583,N_49569);
nor UO_2108 (O_2108,N_48844,N_47811);
or UO_2109 (O_2109,N_46898,N_48158);
nor UO_2110 (O_2110,N_47444,N_47120);
xnor UO_2111 (O_2111,N_48407,N_49119);
and UO_2112 (O_2112,N_46300,N_49108);
nand UO_2113 (O_2113,N_46726,N_47643);
nand UO_2114 (O_2114,N_48421,N_46814);
or UO_2115 (O_2115,N_45654,N_49738);
nor UO_2116 (O_2116,N_46513,N_49700);
or UO_2117 (O_2117,N_47732,N_49571);
nand UO_2118 (O_2118,N_48423,N_48722);
and UO_2119 (O_2119,N_45790,N_48670);
nor UO_2120 (O_2120,N_47981,N_47001);
and UO_2121 (O_2121,N_49044,N_46093);
and UO_2122 (O_2122,N_46488,N_47461);
nand UO_2123 (O_2123,N_47977,N_46208);
and UO_2124 (O_2124,N_47611,N_45114);
xor UO_2125 (O_2125,N_46397,N_48780);
and UO_2126 (O_2126,N_49036,N_45398);
or UO_2127 (O_2127,N_48388,N_45789);
and UO_2128 (O_2128,N_45812,N_48357);
nand UO_2129 (O_2129,N_45056,N_45628);
nor UO_2130 (O_2130,N_47601,N_48136);
and UO_2131 (O_2131,N_49536,N_49917);
xor UO_2132 (O_2132,N_49088,N_45199);
nor UO_2133 (O_2133,N_49475,N_47211);
or UO_2134 (O_2134,N_49273,N_46246);
and UO_2135 (O_2135,N_47935,N_47325);
nand UO_2136 (O_2136,N_46828,N_45991);
nand UO_2137 (O_2137,N_48727,N_49078);
nor UO_2138 (O_2138,N_49233,N_49599);
or UO_2139 (O_2139,N_47618,N_46160);
or UO_2140 (O_2140,N_49534,N_47751);
xnor UO_2141 (O_2141,N_46237,N_47185);
xnor UO_2142 (O_2142,N_48172,N_49238);
nand UO_2143 (O_2143,N_46306,N_45679);
nand UO_2144 (O_2144,N_46858,N_46877);
nor UO_2145 (O_2145,N_47302,N_47534);
xor UO_2146 (O_2146,N_49482,N_45734);
and UO_2147 (O_2147,N_48450,N_45425);
nor UO_2148 (O_2148,N_47392,N_49937);
nand UO_2149 (O_2149,N_47139,N_48431);
nand UO_2150 (O_2150,N_46924,N_45449);
and UO_2151 (O_2151,N_46189,N_46056);
xor UO_2152 (O_2152,N_49872,N_45657);
and UO_2153 (O_2153,N_45858,N_49740);
xor UO_2154 (O_2154,N_47002,N_48516);
xnor UO_2155 (O_2155,N_46355,N_49083);
and UO_2156 (O_2156,N_47430,N_49579);
and UO_2157 (O_2157,N_46302,N_47229);
or UO_2158 (O_2158,N_48620,N_45179);
and UO_2159 (O_2159,N_49759,N_46558);
nor UO_2160 (O_2160,N_48159,N_48321);
nand UO_2161 (O_2161,N_48681,N_48659);
xor UO_2162 (O_2162,N_45561,N_47584);
or UO_2163 (O_2163,N_48915,N_46381);
and UO_2164 (O_2164,N_46891,N_45745);
nor UO_2165 (O_2165,N_45443,N_47136);
or UO_2166 (O_2166,N_45921,N_46866);
xnor UO_2167 (O_2167,N_49313,N_46359);
or UO_2168 (O_2168,N_48216,N_47384);
or UO_2169 (O_2169,N_47212,N_48981);
nand UO_2170 (O_2170,N_48850,N_45326);
or UO_2171 (O_2171,N_46794,N_45287);
or UO_2172 (O_2172,N_47938,N_46618);
nand UO_2173 (O_2173,N_49013,N_49213);
nand UO_2174 (O_2174,N_47741,N_47052);
and UO_2175 (O_2175,N_46830,N_49573);
or UO_2176 (O_2176,N_48692,N_47632);
and UO_2177 (O_2177,N_45878,N_47642);
or UO_2178 (O_2178,N_45490,N_48627);
xnor UO_2179 (O_2179,N_47717,N_49913);
or UO_2180 (O_2180,N_46318,N_49015);
and UO_2181 (O_2181,N_46751,N_47728);
and UO_2182 (O_2182,N_47805,N_46651);
and UO_2183 (O_2183,N_48798,N_46286);
or UO_2184 (O_2184,N_48210,N_47119);
nor UO_2185 (O_2185,N_46703,N_49943);
and UO_2186 (O_2186,N_45411,N_46115);
or UO_2187 (O_2187,N_48865,N_48069);
or UO_2188 (O_2188,N_49699,N_49965);
nand UO_2189 (O_2189,N_48801,N_49543);
nand UO_2190 (O_2190,N_45924,N_46366);
nand UO_2191 (O_2191,N_46612,N_45599);
or UO_2192 (O_2192,N_47833,N_49647);
xor UO_2193 (O_2193,N_49811,N_46403);
and UO_2194 (O_2194,N_46135,N_45741);
nand UO_2195 (O_2195,N_48634,N_48768);
nand UO_2196 (O_2196,N_45999,N_46551);
or UO_2197 (O_2197,N_49436,N_49974);
nand UO_2198 (O_2198,N_47928,N_48959);
nand UO_2199 (O_2199,N_46767,N_45096);
or UO_2200 (O_2200,N_49097,N_46762);
nand UO_2201 (O_2201,N_46064,N_49168);
or UO_2202 (O_2202,N_48876,N_48251);
nor UO_2203 (O_2203,N_46072,N_45161);
or UO_2204 (O_2204,N_49754,N_46277);
nand UO_2205 (O_2205,N_45851,N_46323);
and UO_2206 (O_2206,N_45186,N_45149);
xnor UO_2207 (O_2207,N_45780,N_48295);
nand UO_2208 (O_2208,N_48764,N_45686);
xor UO_2209 (O_2209,N_47213,N_48349);
nand UO_2210 (O_2210,N_46249,N_48710);
and UO_2211 (O_2211,N_49429,N_45419);
xor UO_2212 (O_2212,N_46532,N_47495);
or UO_2213 (O_2213,N_47271,N_46476);
nor UO_2214 (O_2214,N_47993,N_48604);
or UO_2215 (O_2215,N_45501,N_47035);
and UO_2216 (O_2216,N_49930,N_47053);
nand UO_2217 (O_2217,N_46094,N_46722);
nand UO_2218 (O_2218,N_46791,N_46617);
nand UO_2219 (O_2219,N_49175,N_49497);
nor UO_2220 (O_2220,N_47559,N_48082);
or UO_2221 (O_2221,N_49522,N_47307);
nand UO_2222 (O_2222,N_46820,N_48063);
nand UO_2223 (O_2223,N_46701,N_48066);
xor UO_2224 (O_2224,N_49057,N_45191);
nor UO_2225 (O_2225,N_49838,N_49118);
nor UO_2226 (O_2226,N_45933,N_49151);
nor UO_2227 (O_2227,N_46319,N_49778);
nor UO_2228 (O_2228,N_47578,N_47489);
and UO_2229 (O_2229,N_46203,N_47899);
nor UO_2230 (O_2230,N_49695,N_49317);
nor UO_2231 (O_2231,N_49405,N_46388);
and UO_2232 (O_2232,N_49909,N_48453);
and UO_2233 (O_2233,N_46467,N_48125);
nand UO_2234 (O_2234,N_47144,N_47931);
xor UO_2235 (O_2235,N_46429,N_48994);
xor UO_2236 (O_2236,N_49845,N_49552);
nand UO_2237 (O_2237,N_49090,N_47521);
and UO_2238 (O_2238,N_48864,N_49671);
nand UO_2239 (O_2239,N_47703,N_49876);
nor UO_2240 (O_2240,N_49836,N_49340);
nand UO_2241 (O_2241,N_48398,N_49998);
nor UO_2242 (O_2242,N_49769,N_47187);
nor UO_2243 (O_2243,N_45486,N_46714);
and UO_2244 (O_2244,N_45365,N_45718);
nand UO_2245 (O_2245,N_48037,N_45987);
nand UO_2246 (O_2246,N_46528,N_45937);
or UO_2247 (O_2247,N_46729,N_46872);
nand UO_2248 (O_2248,N_49911,N_49426);
nand UO_2249 (O_2249,N_49787,N_45377);
nor UO_2250 (O_2250,N_45588,N_49051);
and UO_2251 (O_2251,N_48023,N_45973);
and UO_2252 (O_2252,N_46944,N_46559);
nand UO_2253 (O_2253,N_48002,N_45670);
xnor UO_2254 (O_2254,N_47566,N_48131);
or UO_2255 (O_2255,N_49049,N_45606);
nor UO_2256 (O_2256,N_45303,N_47644);
nand UO_2257 (O_2257,N_48520,N_48792);
and UO_2258 (O_2258,N_46165,N_47468);
or UO_2259 (O_2259,N_47089,N_48513);
nor UO_2260 (O_2260,N_48454,N_45079);
nand UO_2261 (O_2261,N_48403,N_45900);
or UO_2262 (O_2262,N_46412,N_48983);
nor UO_2263 (O_2263,N_47012,N_48751);
nand UO_2264 (O_2264,N_45060,N_46594);
and UO_2265 (O_2265,N_48871,N_48738);
nand UO_2266 (O_2266,N_46438,N_45340);
xor UO_2267 (O_2267,N_45330,N_46742);
or UO_2268 (O_2268,N_47210,N_46322);
xnor UO_2269 (O_2269,N_49528,N_48822);
or UO_2270 (O_2270,N_46853,N_45837);
nand UO_2271 (O_2271,N_45171,N_46132);
nand UO_2272 (O_2272,N_47888,N_45554);
nor UO_2273 (O_2273,N_48532,N_49194);
and UO_2274 (O_2274,N_49785,N_47878);
nand UO_2275 (O_2275,N_45807,N_48147);
nor UO_2276 (O_2276,N_48405,N_45446);
or UO_2277 (O_2277,N_47842,N_46171);
nand UO_2278 (O_2278,N_46942,N_45712);
nor UO_2279 (O_2279,N_48744,N_46581);
or UO_2280 (O_2280,N_49982,N_45481);
and UO_2281 (O_2281,N_47413,N_48897);
or UO_2282 (O_2282,N_47057,N_48521);
and UO_2283 (O_2283,N_47911,N_47906);
nor UO_2284 (O_2284,N_47026,N_48004);
or UO_2285 (O_2285,N_49739,N_45661);
or UO_2286 (O_2286,N_49952,N_46484);
and UO_2287 (O_2287,N_45023,N_49898);
nor UO_2288 (O_2288,N_46524,N_49154);
nor UO_2289 (O_2289,N_47974,N_48219);
nand UO_2290 (O_2290,N_49192,N_46058);
nor UO_2291 (O_2291,N_48675,N_47513);
nor UO_2292 (O_2292,N_48863,N_46800);
nand UO_2293 (O_2293,N_46608,N_48190);
and UO_2294 (O_2294,N_46304,N_49741);
and UO_2295 (O_2295,N_47735,N_48397);
nand UO_2296 (O_2296,N_45638,N_49627);
and UO_2297 (O_2297,N_45824,N_46802);
nand UO_2298 (O_2298,N_49555,N_45958);
nand UO_2299 (O_2299,N_45465,N_49503);
nor UO_2300 (O_2300,N_48603,N_47008);
and UO_2301 (O_2301,N_45817,N_45863);
nand UO_2302 (O_2302,N_46634,N_46652);
or UO_2303 (O_2303,N_48406,N_46045);
nand UO_2304 (O_2304,N_48298,N_48616);
xnor UO_2305 (O_2305,N_46572,N_46750);
and UO_2306 (O_2306,N_49445,N_48167);
nand UO_2307 (O_2307,N_48493,N_47358);
xor UO_2308 (O_2308,N_46186,N_46149);
nand UO_2309 (O_2309,N_45066,N_46216);
xor UO_2310 (O_2310,N_47291,N_47603);
and UO_2311 (O_2311,N_45346,N_47509);
or UO_2312 (O_2312,N_45352,N_45579);
and UO_2313 (O_2313,N_46508,N_48362);
and UO_2314 (O_2314,N_47670,N_49377);
nand UO_2315 (O_2315,N_48118,N_49935);
nand UO_2316 (O_2316,N_45177,N_49283);
nand UO_2317 (O_2317,N_49058,N_49992);
and UO_2318 (O_2318,N_45688,N_47567);
and UO_2319 (O_2319,N_46997,N_46653);
nand UO_2320 (O_2320,N_47312,N_46737);
nor UO_2321 (O_2321,N_45517,N_45499);
nor UO_2322 (O_2322,N_47967,N_45819);
nand UO_2323 (O_2323,N_47803,N_48032);
and UO_2324 (O_2324,N_48042,N_49461);
and UO_2325 (O_2325,N_46224,N_45811);
nand UO_2326 (O_2326,N_49830,N_46748);
xor UO_2327 (O_2327,N_48436,N_49853);
nand UO_2328 (O_2328,N_45220,N_48635);
nor UO_2329 (O_2329,N_45374,N_49032);
xor UO_2330 (O_2330,N_49400,N_48843);
or UO_2331 (O_2331,N_46995,N_49812);
nand UO_2332 (O_2332,N_45404,N_45545);
nand UO_2333 (O_2333,N_49353,N_47135);
nand UO_2334 (O_2334,N_45800,N_46604);
and UO_2335 (O_2335,N_49402,N_46497);
or UO_2336 (O_2336,N_46312,N_46043);
nor UO_2337 (O_2337,N_47630,N_46266);
nand UO_2338 (O_2338,N_46760,N_49152);
xor UO_2339 (O_2339,N_47007,N_46228);
and UO_2340 (O_2340,N_45935,N_47961);
nand UO_2341 (O_2341,N_45285,N_49730);
or UO_2342 (O_2342,N_49995,N_45528);
or UO_2343 (O_2343,N_46451,N_48999);
and UO_2344 (O_2344,N_47234,N_48482);
nand UO_2345 (O_2345,N_45676,N_46671);
xor UO_2346 (O_2346,N_49765,N_48368);
nand UO_2347 (O_2347,N_46576,N_45665);
or UO_2348 (O_2348,N_46140,N_48175);
nor UO_2349 (O_2349,N_49620,N_49218);
nor UO_2350 (O_2350,N_47061,N_45054);
nand UO_2351 (O_2351,N_47537,N_48589);
nand UO_2352 (O_2352,N_46170,N_45740);
nand UO_2353 (O_2353,N_49081,N_48473);
nor UO_2354 (O_2354,N_49841,N_48952);
or UO_2355 (O_2355,N_45221,N_48672);
and UO_2356 (O_2356,N_47980,N_49395);
or UO_2357 (O_2357,N_47132,N_48731);
nand UO_2358 (O_2358,N_49717,N_49211);
or UO_2359 (O_2359,N_48455,N_46874);
nor UO_2360 (O_2360,N_46860,N_46444);
nor UO_2361 (O_2361,N_49354,N_45383);
xnor UO_2362 (O_2362,N_49606,N_47277);
or UO_2363 (O_2363,N_48386,N_45782);
nor UO_2364 (O_2364,N_49437,N_46288);
or UO_2365 (O_2365,N_45662,N_49978);
nand UO_2366 (O_2366,N_49560,N_48534);
nor UO_2367 (O_2367,N_48314,N_49095);
and UO_2368 (O_2368,N_45078,N_46505);
nor UO_2369 (O_2369,N_45593,N_47196);
or UO_2370 (O_2370,N_45219,N_45421);
or UO_2371 (O_2371,N_46765,N_47415);
and UO_2372 (O_2372,N_47270,N_49635);
nor UO_2373 (O_2373,N_49494,N_47418);
or UO_2374 (O_2374,N_45367,N_47791);
nor UO_2375 (O_2375,N_46628,N_45195);
nor UO_2376 (O_2376,N_49374,N_45470);
or UO_2377 (O_2377,N_49918,N_48209);
or UO_2378 (O_2378,N_48026,N_49115);
and UO_2379 (O_2379,N_49116,N_47929);
xor UO_2380 (O_2380,N_47769,N_45621);
or UO_2381 (O_2381,N_47369,N_46838);
or UO_2382 (O_2382,N_47372,N_46889);
nor UO_2383 (O_2383,N_45429,N_48921);
nand UO_2384 (O_2384,N_48194,N_46916);
nand UO_2385 (O_2385,N_46718,N_45767);
or UO_2386 (O_2386,N_45264,N_48480);
nand UO_2387 (O_2387,N_49141,N_47147);
nand UO_2388 (O_2388,N_49205,N_46936);
and UO_2389 (O_2389,N_49178,N_49358);
or UO_2390 (O_2390,N_46945,N_48997);
or UO_2391 (O_2391,N_49386,N_46011);
nor UO_2392 (O_2392,N_46719,N_45754);
or UO_2393 (O_2393,N_47678,N_45495);
nand UO_2394 (O_2394,N_47243,N_49736);
nand UO_2395 (O_2395,N_48047,N_49762);
nor UO_2396 (O_2396,N_48443,N_46398);
or UO_2397 (O_2397,N_49469,N_46758);
or UO_2398 (O_2398,N_49950,N_49472);
xnor UO_2399 (O_2399,N_48229,N_49761);
nand UO_2400 (O_2400,N_46527,N_47058);
or UO_2401 (O_2401,N_48382,N_47621);
and UO_2402 (O_2402,N_45135,N_47874);
nor UO_2403 (O_2403,N_49006,N_45004);
or UO_2404 (O_2404,N_49258,N_47600);
and UO_2405 (O_2405,N_47700,N_46759);
nand UO_2406 (O_2406,N_45992,N_46418);
or UO_2407 (O_2407,N_48287,N_47645);
nand UO_2408 (O_2408,N_45433,N_47810);
nand UO_2409 (O_2409,N_49208,N_48141);
and UO_2410 (O_2410,N_46461,N_45653);
or UO_2411 (O_2411,N_45769,N_47737);
and UO_2412 (O_2412,N_45074,N_46885);
nor UO_2413 (O_2413,N_48784,N_45904);
or UO_2414 (O_2414,N_47005,N_45227);
and UO_2415 (O_2415,N_46507,N_46262);
xor UO_2416 (O_2416,N_45538,N_49368);
and UO_2417 (O_2417,N_46597,N_45051);
or UO_2418 (O_2418,N_49586,N_45274);
nor UO_2419 (O_2419,N_49019,N_45967);
or UO_2420 (O_2420,N_45816,N_47836);
nor UO_2421 (O_2421,N_49456,N_46022);
nand UO_2422 (O_2422,N_49747,N_46919);
nor UO_2423 (O_2423,N_47982,N_45099);
or UO_2424 (O_2424,N_45132,N_48248);
and UO_2425 (O_2425,N_48927,N_49256);
nor UO_2426 (O_2426,N_47813,N_48428);
nor UO_2427 (O_2427,N_45234,N_45156);
and UO_2428 (O_2428,N_48091,N_47164);
or UO_2429 (O_2429,N_48933,N_45032);
xor UO_2430 (O_2430,N_49271,N_47481);
or UO_2431 (O_2431,N_46387,N_45511);
nand UO_2432 (O_2432,N_46529,N_48138);
and UO_2433 (O_2433,N_48932,N_49817);
nand UO_2434 (O_2434,N_49716,N_48134);
or UO_2435 (O_2435,N_46354,N_46371);
or UO_2436 (O_2436,N_45254,N_48166);
nand UO_2437 (O_2437,N_49770,N_49827);
or UO_2438 (O_2438,N_48288,N_45257);
nor UO_2439 (O_2439,N_49644,N_49164);
nand UO_2440 (O_2440,N_46588,N_49829);
and UO_2441 (O_2441,N_47818,N_49705);
nand UO_2442 (O_2442,N_46435,N_46520);
or UO_2443 (O_2443,N_45936,N_49064);
nand UO_2444 (O_2444,N_45872,N_46695);
and UO_2445 (O_2445,N_49893,N_48239);
and UO_2446 (O_2446,N_46025,N_49631);
and UO_2447 (O_2447,N_47382,N_46107);
xor UO_2448 (O_2448,N_45604,N_46584);
and UO_2449 (O_2449,N_45269,N_47216);
xor UO_2450 (O_2450,N_45785,N_47318);
nand UO_2451 (O_2451,N_47869,N_45965);
nand UO_2452 (O_2452,N_47696,N_46990);
or UO_2453 (O_2453,N_47480,N_47668);
nor UO_2454 (O_2454,N_48083,N_48449);
and UO_2455 (O_2455,N_47359,N_49369);
xor UO_2456 (O_2456,N_48993,N_46098);
xnor UO_2457 (O_2457,N_47910,N_45210);
nor UO_2458 (O_2458,N_48101,N_45198);
xnor UO_2459 (O_2459,N_45444,N_48377);
and UO_2460 (O_2460,N_45928,N_45779);
or UO_2461 (O_2461,N_49274,N_48924);
nand UO_2462 (O_2462,N_49480,N_46503);
xor UO_2463 (O_2463,N_46464,N_46445);
nor UO_2464 (O_2464,N_49485,N_46270);
xnor UO_2465 (O_2465,N_49623,N_46522);
or UO_2466 (O_2466,N_47462,N_45601);
and UO_2467 (O_2467,N_48338,N_46669);
nor UO_2468 (O_2468,N_47491,N_46930);
and UO_2469 (O_2469,N_49713,N_48732);
and UO_2470 (O_2470,N_45125,N_45482);
nand UO_2471 (O_2471,N_48676,N_46927);
or UO_2472 (O_2472,N_47096,N_49269);
nor UO_2473 (O_2473,N_49157,N_48812);
xor UO_2474 (O_2474,N_47108,N_48547);
nor UO_2475 (O_2475,N_45507,N_47868);
nor UO_2476 (O_2476,N_48957,N_45704);
and UO_2477 (O_2477,N_45440,N_46788);
or UO_2478 (O_2478,N_47056,N_49654);
and UO_2479 (O_2479,N_46166,N_48247);
and UO_2480 (O_2480,N_46184,N_47825);
or UO_2481 (O_2481,N_47573,N_48178);
or UO_2482 (O_2482,N_46846,N_48905);
nor UO_2483 (O_2483,N_45072,N_45583);
and UO_2484 (O_2484,N_45756,N_47634);
nor UO_2485 (O_2485,N_47265,N_46151);
and UO_2486 (O_2486,N_45696,N_48555);
xor UO_2487 (O_2487,N_48068,N_48759);
nor UO_2488 (O_2488,N_49722,N_48354);
or UO_2489 (O_2489,N_45503,N_45251);
nand UO_2490 (O_2490,N_47824,N_45895);
nand UO_2491 (O_2491,N_47783,N_46905);
or UO_2492 (O_2492,N_48360,N_46509);
and UO_2493 (O_2493,N_45930,N_45232);
or UO_2494 (O_2494,N_46975,N_45245);
nand UO_2495 (O_2495,N_49686,N_49860);
and UO_2496 (O_2496,N_47275,N_48100);
nand UO_2497 (O_2497,N_46038,N_48557);
nor UO_2498 (O_2498,N_48261,N_47639);
nand UO_2499 (O_2499,N_47604,N_48658);
nor UO_2500 (O_2500,N_49347,N_45310);
and UO_2501 (O_2501,N_47279,N_46580);
and UO_2502 (O_2502,N_48251,N_46416);
nor UO_2503 (O_2503,N_48621,N_45429);
nor UO_2504 (O_2504,N_49893,N_46028);
xnor UO_2505 (O_2505,N_45138,N_45022);
xor UO_2506 (O_2506,N_46758,N_48695);
or UO_2507 (O_2507,N_49729,N_45658);
or UO_2508 (O_2508,N_45964,N_45956);
xnor UO_2509 (O_2509,N_45875,N_46260);
nor UO_2510 (O_2510,N_45663,N_47324);
nand UO_2511 (O_2511,N_45144,N_46169);
nor UO_2512 (O_2512,N_48077,N_45078);
and UO_2513 (O_2513,N_47349,N_49538);
nand UO_2514 (O_2514,N_49381,N_49235);
and UO_2515 (O_2515,N_48623,N_49095);
xor UO_2516 (O_2516,N_45745,N_46511);
and UO_2517 (O_2517,N_49793,N_46403);
and UO_2518 (O_2518,N_48137,N_48407);
xor UO_2519 (O_2519,N_45672,N_49216);
nand UO_2520 (O_2520,N_46627,N_45228);
nand UO_2521 (O_2521,N_46958,N_49041);
nand UO_2522 (O_2522,N_49390,N_47887);
nand UO_2523 (O_2523,N_45741,N_48359);
or UO_2524 (O_2524,N_46490,N_45365);
and UO_2525 (O_2525,N_46898,N_47824);
nor UO_2526 (O_2526,N_45618,N_48217);
nor UO_2527 (O_2527,N_49333,N_48886);
or UO_2528 (O_2528,N_46677,N_49086);
nand UO_2529 (O_2529,N_48301,N_47181);
and UO_2530 (O_2530,N_47976,N_49448);
or UO_2531 (O_2531,N_45028,N_49809);
nor UO_2532 (O_2532,N_45282,N_48414);
or UO_2533 (O_2533,N_45397,N_47540);
or UO_2534 (O_2534,N_45080,N_46719);
or UO_2535 (O_2535,N_48336,N_48890);
or UO_2536 (O_2536,N_45079,N_49121);
or UO_2537 (O_2537,N_48991,N_49494);
nand UO_2538 (O_2538,N_46264,N_45083);
nand UO_2539 (O_2539,N_49736,N_48752);
nor UO_2540 (O_2540,N_49419,N_45087);
and UO_2541 (O_2541,N_46789,N_45797);
or UO_2542 (O_2542,N_45424,N_46975);
xnor UO_2543 (O_2543,N_45019,N_49841);
nand UO_2544 (O_2544,N_47206,N_47999);
or UO_2545 (O_2545,N_45665,N_45902);
nand UO_2546 (O_2546,N_48748,N_49959);
nand UO_2547 (O_2547,N_45674,N_46038);
xnor UO_2548 (O_2548,N_46214,N_47640);
and UO_2549 (O_2549,N_45140,N_47982);
xnor UO_2550 (O_2550,N_46320,N_48268);
nand UO_2551 (O_2551,N_48083,N_49478);
nor UO_2552 (O_2552,N_48498,N_49061);
nand UO_2553 (O_2553,N_47251,N_47777);
and UO_2554 (O_2554,N_49375,N_46997);
nand UO_2555 (O_2555,N_46396,N_49113);
nor UO_2556 (O_2556,N_49414,N_46512);
xnor UO_2557 (O_2557,N_45183,N_45059);
and UO_2558 (O_2558,N_49096,N_46742);
and UO_2559 (O_2559,N_46153,N_48246);
or UO_2560 (O_2560,N_47025,N_45137);
or UO_2561 (O_2561,N_49584,N_46399);
nor UO_2562 (O_2562,N_47189,N_49921);
nand UO_2563 (O_2563,N_48068,N_46904);
or UO_2564 (O_2564,N_49569,N_45584);
nor UO_2565 (O_2565,N_45228,N_49557);
nor UO_2566 (O_2566,N_45169,N_45671);
nor UO_2567 (O_2567,N_46109,N_45162);
nor UO_2568 (O_2568,N_46863,N_49959);
nor UO_2569 (O_2569,N_46224,N_48121);
xor UO_2570 (O_2570,N_47442,N_48791);
nand UO_2571 (O_2571,N_47550,N_46775);
and UO_2572 (O_2572,N_47806,N_46994);
nand UO_2573 (O_2573,N_47215,N_47673);
and UO_2574 (O_2574,N_47639,N_47742);
nor UO_2575 (O_2575,N_47165,N_46444);
xnor UO_2576 (O_2576,N_45807,N_45333);
nor UO_2577 (O_2577,N_47499,N_47867);
and UO_2578 (O_2578,N_45862,N_46872);
and UO_2579 (O_2579,N_49011,N_47720);
nor UO_2580 (O_2580,N_49832,N_49947);
and UO_2581 (O_2581,N_49430,N_46327);
nor UO_2582 (O_2582,N_46115,N_46534);
nor UO_2583 (O_2583,N_46929,N_48068);
nand UO_2584 (O_2584,N_49404,N_47850);
or UO_2585 (O_2585,N_45559,N_47438);
nand UO_2586 (O_2586,N_48253,N_45431);
or UO_2587 (O_2587,N_48310,N_49517);
and UO_2588 (O_2588,N_46654,N_45542);
or UO_2589 (O_2589,N_46755,N_46724);
and UO_2590 (O_2590,N_47513,N_45454);
nand UO_2591 (O_2591,N_47106,N_47041);
or UO_2592 (O_2592,N_49756,N_45664);
xnor UO_2593 (O_2593,N_49404,N_49626);
and UO_2594 (O_2594,N_49563,N_46951);
or UO_2595 (O_2595,N_47086,N_46511);
or UO_2596 (O_2596,N_46224,N_47659);
or UO_2597 (O_2597,N_48059,N_47767);
nor UO_2598 (O_2598,N_45222,N_45851);
nand UO_2599 (O_2599,N_47161,N_45138);
xnor UO_2600 (O_2600,N_45151,N_45353);
and UO_2601 (O_2601,N_49730,N_46623);
nor UO_2602 (O_2602,N_46102,N_48345);
nor UO_2603 (O_2603,N_45323,N_47746);
nand UO_2604 (O_2604,N_49761,N_46047);
nor UO_2605 (O_2605,N_46319,N_48459);
nor UO_2606 (O_2606,N_45053,N_45794);
or UO_2607 (O_2607,N_48012,N_45966);
or UO_2608 (O_2608,N_48521,N_49682);
nor UO_2609 (O_2609,N_49142,N_46827);
or UO_2610 (O_2610,N_47025,N_48711);
nand UO_2611 (O_2611,N_46705,N_47276);
nor UO_2612 (O_2612,N_47754,N_46726);
xor UO_2613 (O_2613,N_47745,N_45270);
nand UO_2614 (O_2614,N_46505,N_48488);
nor UO_2615 (O_2615,N_45114,N_49044);
and UO_2616 (O_2616,N_47040,N_46733);
nor UO_2617 (O_2617,N_48513,N_46942);
nor UO_2618 (O_2618,N_48475,N_47939);
xnor UO_2619 (O_2619,N_48997,N_47610);
xnor UO_2620 (O_2620,N_49270,N_48354);
nor UO_2621 (O_2621,N_47753,N_47678);
nand UO_2622 (O_2622,N_47571,N_49423);
and UO_2623 (O_2623,N_45960,N_45601);
or UO_2624 (O_2624,N_45586,N_47840);
nand UO_2625 (O_2625,N_46754,N_45742);
nand UO_2626 (O_2626,N_48802,N_48849);
or UO_2627 (O_2627,N_49394,N_45519);
nand UO_2628 (O_2628,N_46855,N_49613);
or UO_2629 (O_2629,N_45582,N_48535);
nand UO_2630 (O_2630,N_45518,N_49078);
xnor UO_2631 (O_2631,N_49974,N_45705);
or UO_2632 (O_2632,N_48078,N_48323);
and UO_2633 (O_2633,N_49351,N_45033);
nor UO_2634 (O_2634,N_48857,N_45262);
nor UO_2635 (O_2635,N_49083,N_47521);
nor UO_2636 (O_2636,N_48842,N_47740);
nand UO_2637 (O_2637,N_45356,N_45217);
or UO_2638 (O_2638,N_46469,N_49135);
and UO_2639 (O_2639,N_49540,N_45317);
or UO_2640 (O_2640,N_49976,N_46576);
nor UO_2641 (O_2641,N_49993,N_46913);
nand UO_2642 (O_2642,N_46088,N_46377);
nor UO_2643 (O_2643,N_45248,N_47270);
and UO_2644 (O_2644,N_47770,N_46430);
xor UO_2645 (O_2645,N_46046,N_47400);
nor UO_2646 (O_2646,N_49017,N_48450);
and UO_2647 (O_2647,N_45542,N_45119);
and UO_2648 (O_2648,N_45995,N_48853);
nor UO_2649 (O_2649,N_49199,N_45776);
nor UO_2650 (O_2650,N_49491,N_45002);
and UO_2651 (O_2651,N_48311,N_49567);
nand UO_2652 (O_2652,N_47518,N_49147);
or UO_2653 (O_2653,N_48254,N_45115);
xor UO_2654 (O_2654,N_47219,N_45292);
or UO_2655 (O_2655,N_45732,N_45127);
or UO_2656 (O_2656,N_47210,N_45038);
xnor UO_2657 (O_2657,N_48513,N_48391);
nor UO_2658 (O_2658,N_48561,N_45239);
nand UO_2659 (O_2659,N_45448,N_45711);
nand UO_2660 (O_2660,N_49081,N_46941);
or UO_2661 (O_2661,N_45376,N_45406);
nand UO_2662 (O_2662,N_48908,N_49071);
nor UO_2663 (O_2663,N_47085,N_48530);
nand UO_2664 (O_2664,N_48025,N_46228);
nand UO_2665 (O_2665,N_48971,N_46057);
nor UO_2666 (O_2666,N_48740,N_47961);
and UO_2667 (O_2667,N_47307,N_46782);
or UO_2668 (O_2668,N_48186,N_49239);
nand UO_2669 (O_2669,N_49058,N_48696);
and UO_2670 (O_2670,N_48953,N_47188);
or UO_2671 (O_2671,N_48925,N_47636);
nand UO_2672 (O_2672,N_49129,N_45954);
or UO_2673 (O_2673,N_47564,N_46517);
nand UO_2674 (O_2674,N_49936,N_49245);
or UO_2675 (O_2675,N_48647,N_48538);
or UO_2676 (O_2676,N_47100,N_48817);
and UO_2677 (O_2677,N_49780,N_48990);
xnor UO_2678 (O_2678,N_47330,N_45603);
nand UO_2679 (O_2679,N_45359,N_48223);
and UO_2680 (O_2680,N_49498,N_45541);
or UO_2681 (O_2681,N_47659,N_48626);
and UO_2682 (O_2682,N_47790,N_45426);
or UO_2683 (O_2683,N_46958,N_45532);
and UO_2684 (O_2684,N_49318,N_47681);
or UO_2685 (O_2685,N_47958,N_48126);
and UO_2686 (O_2686,N_49866,N_45277);
nand UO_2687 (O_2687,N_45887,N_47831);
and UO_2688 (O_2688,N_45490,N_47047);
and UO_2689 (O_2689,N_49607,N_48491);
nand UO_2690 (O_2690,N_47793,N_49877);
nor UO_2691 (O_2691,N_49331,N_48014);
xor UO_2692 (O_2692,N_49840,N_49186);
xor UO_2693 (O_2693,N_46957,N_46687);
nand UO_2694 (O_2694,N_48487,N_46853);
nand UO_2695 (O_2695,N_46765,N_46474);
and UO_2696 (O_2696,N_47357,N_46934);
and UO_2697 (O_2697,N_47139,N_48706);
nand UO_2698 (O_2698,N_49144,N_46463);
nor UO_2699 (O_2699,N_48746,N_46328);
or UO_2700 (O_2700,N_49020,N_47277);
xor UO_2701 (O_2701,N_48787,N_46872);
and UO_2702 (O_2702,N_48777,N_46300);
nor UO_2703 (O_2703,N_47864,N_45048);
xor UO_2704 (O_2704,N_48089,N_45016);
nor UO_2705 (O_2705,N_46852,N_46921);
nor UO_2706 (O_2706,N_46414,N_49444);
nor UO_2707 (O_2707,N_49691,N_47022);
xor UO_2708 (O_2708,N_47328,N_46149);
xnor UO_2709 (O_2709,N_47156,N_49036);
nor UO_2710 (O_2710,N_46282,N_49451);
nand UO_2711 (O_2711,N_48461,N_46448);
nand UO_2712 (O_2712,N_46908,N_48832);
and UO_2713 (O_2713,N_49714,N_45462);
nor UO_2714 (O_2714,N_45025,N_46596);
nor UO_2715 (O_2715,N_46093,N_47076);
and UO_2716 (O_2716,N_47792,N_47664);
nand UO_2717 (O_2717,N_49681,N_48864);
xor UO_2718 (O_2718,N_45878,N_47631);
nand UO_2719 (O_2719,N_46945,N_45481);
nor UO_2720 (O_2720,N_46944,N_47115);
nand UO_2721 (O_2721,N_48085,N_45040);
or UO_2722 (O_2722,N_47910,N_49245);
or UO_2723 (O_2723,N_45240,N_48517);
and UO_2724 (O_2724,N_48489,N_48027);
nor UO_2725 (O_2725,N_47015,N_49418);
nand UO_2726 (O_2726,N_45728,N_47997);
nor UO_2727 (O_2727,N_49887,N_45444);
xnor UO_2728 (O_2728,N_48910,N_48610);
nand UO_2729 (O_2729,N_48323,N_45945);
nor UO_2730 (O_2730,N_46986,N_47119);
nor UO_2731 (O_2731,N_46582,N_45857);
nand UO_2732 (O_2732,N_47147,N_46685);
and UO_2733 (O_2733,N_45355,N_49149);
or UO_2734 (O_2734,N_45146,N_45094);
nand UO_2735 (O_2735,N_47817,N_48450);
xor UO_2736 (O_2736,N_47479,N_48829);
nand UO_2737 (O_2737,N_49944,N_46928);
and UO_2738 (O_2738,N_45676,N_45980);
xor UO_2739 (O_2739,N_47935,N_47973);
or UO_2740 (O_2740,N_47570,N_48794);
or UO_2741 (O_2741,N_49693,N_45056);
nor UO_2742 (O_2742,N_48220,N_46023);
xnor UO_2743 (O_2743,N_46339,N_49052);
or UO_2744 (O_2744,N_46588,N_47614);
xnor UO_2745 (O_2745,N_49889,N_46991);
nor UO_2746 (O_2746,N_49345,N_45835);
nor UO_2747 (O_2747,N_49558,N_47230);
nand UO_2748 (O_2748,N_49782,N_49812);
nand UO_2749 (O_2749,N_49398,N_46915);
nor UO_2750 (O_2750,N_49772,N_48995);
or UO_2751 (O_2751,N_47537,N_49759);
or UO_2752 (O_2752,N_48723,N_48174);
and UO_2753 (O_2753,N_45782,N_47103);
nor UO_2754 (O_2754,N_49971,N_49615);
or UO_2755 (O_2755,N_47837,N_49304);
or UO_2756 (O_2756,N_45039,N_47619);
nor UO_2757 (O_2757,N_47112,N_45603);
nand UO_2758 (O_2758,N_45008,N_46248);
nand UO_2759 (O_2759,N_45746,N_48239);
nand UO_2760 (O_2760,N_47420,N_46457);
or UO_2761 (O_2761,N_45846,N_46954);
nand UO_2762 (O_2762,N_49857,N_45121);
and UO_2763 (O_2763,N_48467,N_48710);
nand UO_2764 (O_2764,N_47425,N_45358);
and UO_2765 (O_2765,N_49507,N_49731);
or UO_2766 (O_2766,N_47382,N_47507);
and UO_2767 (O_2767,N_48273,N_49888);
nand UO_2768 (O_2768,N_45829,N_46507);
and UO_2769 (O_2769,N_49357,N_49598);
nor UO_2770 (O_2770,N_47209,N_47139);
and UO_2771 (O_2771,N_47626,N_46603);
nand UO_2772 (O_2772,N_49202,N_46845);
and UO_2773 (O_2773,N_46043,N_47836);
nor UO_2774 (O_2774,N_47969,N_49321);
or UO_2775 (O_2775,N_46692,N_49952);
xor UO_2776 (O_2776,N_45601,N_46953);
or UO_2777 (O_2777,N_46099,N_49015);
nor UO_2778 (O_2778,N_46692,N_48727);
nand UO_2779 (O_2779,N_49209,N_49385);
nor UO_2780 (O_2780,N_46110,N_46052);
or UO_2781 (O_2781,N_49914,N_45896);
or UO_2782 (O_2782,N_49280,N_47785);
nor UO_2783 (O_2783,N_48846,N_47857);
and UO_2784 (O_2784,N_47037,N_47258);
and UO_2785 (O_2785,N_47201,N_49811);
nor UO_2786 (O_2786,N_47277,N_47920);
nor UO_2787 (O_2787,N_49068,N_47459);
or UO_2788 (O_2788,N_46096,N_48577);
and UO_2789 (O_2789,N_46310,N_49338);
xnor UO_2790 (O_2790,N_45686,N_45302);
and UO_2791 (O_2791,N_49506,N_48445);
and UO_2792 (O_2792,N_48149,N_48378);
nor UO_2793 (O_2793,N_47922,N_49933);
nor UO_2794 (O_2794,N_45146,N_46148);
nor UO_2795 (O_2795,N_45941,N_46459);
nor UO_2796 (O_2796,N_48814,N_46101);
nor UO_2797 (O_2797,N_46907,N_49330);
nand UO_2798 (O_2798,N_46399,N_48796);
xor UO_2799 (O_2799,N_46532,N_49144);
and UO_2800 (O_2800,N_48817,N_47155);
nor UO_2801 (O_2801,N_45083,N_49179);
xnor UO_2802 (O_2802,N_49232,N_49966);
xor UO_2803 (O_2803,N_47826,N_46732);
and UO_2804 (O_2804,N_46918,N_46204);
or UO_2805 (O_2805,N_46880,N_46645);
or UO_2806 (O_2806,N_49199,N_46915);
and UO_2807 (O_2807,N_47155,N_49684);
xor UO_2808 (O_2808,N_48186,N_47071);
nand UO_2809 (O_2809,N_47483,N_48273);
or UO_2810 (O_2810,N_46795,N_48128);
or UO_2811 (O_2811,N_49709,N_48223);
nand UO_2812 (O_2812,N_49818,N_45770);
xnor UO_2813 (O_2813,N_46023,N_46381);
nand UO_2814 (O_2814,N_45869,N_48037);
xor UO_2815 (O_2815,N_45761,N_45158);
nand UO_2816 (O_2816,N_48427,N_45459);
nand UO_2817 (O_2817,N_46149,N_46875);
nor UO_2818 (O_2818,N_47153,N_46017);
and UO_2819 (O_2819,N_46985,N_49953);
nand UO_2820 (O_2820,N_46426,N_48477);
and UO_2821 (O_2821,N_46882,N_49000);
or UO_2822 (O_2822,N_45588,N_48372);
xnor UO_2823 (O_2823,N_45377,N_46566);
nand UO_2824 (O_2824,N_48633,N_45938);
nand UO_2825 (O_2825,N_45598,N_48119);
and UO_2826 (O_2826,N_47170,N_48866);
or UO_2827 (O_2827,N_46447,N_49396);
nor UO_2828 (O_2828,N_48926,N_49688);
xnor UO_2829 (O_2829,N_45139,N_46792);
or UO_2830 (O_2830,N_46655,N_48121);
nor UO_2831 (O_2831,N_47906,N_48270);
or UO_2832 (O_2832,N_48278,N_48440);
or UO_2833 (O_2833,N_49563,N_49092);
and UO_2834 (O_2834,N_47759,N_48438);
and UO_2835 (O_2835,N_49217,N_45975);
nor UO_2836 (O_2836,N_46191,N_47304);
nor UO_2837 (O_2837,N_46663,N_47613);
nor UO_2838 (O_2838,N_47105,N_49528);
or UO_2839 (O_2839,N_46881,N_49805);
or UO_2840 (O_2840,N_46581,N_48728);
nor UO_2841 (O_2841,N_45359,N_46857);
nor UO_2842 (O_2842,N_47936,N_47323);
or UO_2843 (O_2843,N_48761,N_46776);
xnor UO_2844 (O_2844,N_46790,N_49412);
or UO_2845 (O_2845,N_49024,N_49521);
or UO_2846 (O_2846,N_46537,N_46163);
or UO_2847 (O_2847,N_47768,N_48279);
and UO_2848 (O_2848,N_49574,N_49638);
and UO_2849 (O_2849,N_46201,N_47340);
and UO_2850 (O_2850,N_49743,N_48870);
nor UO_2851 (O_2851,N_47620,N_46306);
xor UO_2852 (O_2852,N_45369,N_45713);
nand UO_2853 (O_2853,N_47861,N_47476);
xnor UO_2854 (O_2854,N_45992,N_46050);
nand UO_2855 (O_2855,N_47844,N_45560);
or UO_2856 (O_2856,N_48717,N_46734);
and UO_2857 (O_2857,N_46906,N_48883);
or UO_2858 (O_2858,N_48939,N_48696);
nand UO_2859 (O_2859,N_46979,N_45847);
nand UO_2860 (O_2860,N_47126,N_47790);
nor UO_2861 (O_2861,N_49117,N_45100);
or UO_2862 (O_2862,N_46300,N_46405);
nor UO_2863 (O_2863,N_46533,N_47947);
and UO_2864 (O_2864,N_47846,N_46794);
and UO_2865 (O_2865,N_48315,N_48978);
nor UO_2866 (O_2866,N_47906,N_47328);
or UO_2867 (O_2867,N_49493,N_49473);
nor UO_2868 (O_2868,N_46137,N_49194);
nor UO_2869 (O_2869,N_48514,N_45512);
or UO_2870 (O_2870,N_47143,N_49604);
nor UO_2871 (O_2871,N_47350,N_46081);
or UO_2872 (O_2872,N_49771,N_46451);
xor UO_2873 (O_2873,N_46710,N_49367);
and UO_2874 (O_2874,N_47499,N_47035);
and UO_2875 (O_2875,N_48518,N_49304);
nand UO_2876 (O_2876,N_47366,N_46255);
nand UO_2877 (O_2877,N_46876,N_49005);
xor UO_2878 (O_2878,N_47704,N_45336);
nand UO_2879 (O_2879,N_47874,N_47174);
and UO_2880 (O_2880,N_47040,N_46636);
nor UO_2881 (O_2881,N_45498,N_48692);
or UO_2882 (O_2882,N_46736,N_49037);
or UO_2883 (O_2883,N_49885,N_49221);
or UO_2884 (O_2884,N_45477,N_49335);
xor UO_2885 (O_2885,N_49678,N_48521);
or UO_2886 (O_2886,N_49074,N_45104);
or UO_2887 (O_2887,N_49910,N_45994);
nor UO_2888 (O_2888,N_45007,N_49031);
nand UO_2889 (O_2889,N_47680,N_46206);
and UO_2890 (O_2890,N_47598,N_45166);
and UO_2891 (O_2891,N_45764,N_49622);
nand UO_2892 (O_2892,N_46192,N_49353);
nor UO_2893 (O_2893,N_45062,N_49965);
and UO_2894 (O_2894,N_49857,N_47507);
xor UO_2895 (O_2895,N_45930,N_49783);
and UO_2896 (O_2896,N_48402,N_47652);
and UO_2897 (O_2897,N_49533,N_49634);
and UO_2898 (O_2898,N_47387,N_46178);
xnor UO_2899 (O_2899,N_45390,N_49558);
and UO_2900 (O_2900,N_49804,N_49836);
nor UO_2901 (O_2901,N_45651,N_48963);
nor UO_2902 (O_2902,N_47027,N_47179);
nand UO_2903 (O_2903,N_47578,N_46141);
nor UO_2904 (O_2904,N_49535,N_45675);
nand UO_2905 (O_2905,N_45598,N_47766);
nor UO_2906 (O_2906,N_46419,N_49311);
nand UO_2907 (O_2907,N_45294,N_45120);
nor UO_2908 (O_2908,N_48048,N_46442);
nor UO_2909 (O_2909,N_45635,N_47632);
or UO_2910 (O_2910,N_46626,N_45963);
and UO_2911 (O_2911,N_45509,N_48885);
nand UO_2912 (O_2912,N_46929,N_48747);
nor UO_2913 (O_2913,N_46888,N_46977);
and UO_2914 (O_2914,N_46769,N_45427);
nand UO_2915 (O_2915,N_46591,N_47076);
and UO_2916 (O_2916,N_47398,N_48081);
nand UO_2917 (O_2917,N_47803,N_47036);
xnor UO_2918 (O_2918,N_48732,N_48329);
nor UO_2919 (O_2919,N_46106,N_47729);
or UO_2920 (O_2920,N_45211,N_49732);
xnor UO_2921 (O_2921,N_49455,N_47656);
nor UO_2922 (O_2922,N_47657,N_45138);
and UO_2923 (O_2923,N_49576,N_47142);
xor UO_2924 (O_2924,N_48375,N_45858);
nand UO_2925 (O_2925,N_49855,N_47674);
and UO_2926 (O_2926,N_45742,N_45224);
and UO_2927 (O_2927,N_45242,N_45482);
and UO_2928 (O_2928,N_46873,N_46864);
nor UO_2929 (O_2929,N_48042,N_47131);
nand UO_2930 (O_2930,N_47369,N_49599);
nand UO_2931 (O_2931,N_45139,N_46633);
nor UO_2932 (O_2932,N_45102,N_45982);
nand UO_2933 (O_2933,N_48802,N_49895);
nor UO_2934 (O_2934,N_46971,N_46706);
or UO_2935 (O_2935,N_46654,N_47744);
nand UO_2936 (O_2936,N_45208,N_47231);
nand UO_2937 (O_2937,N_49975,N_49239);
nor UO_2938 (O_2938,N_49839,N_47479);
nand UO_2939 (O_2939,N_46542,N_48471);
nand UO_2940 (O_2940,N_49727,N_45954);
nor UO_2941 (O_2941,N_47150,N_47077);
nor UO_2942 (O_2942,N_48865,N_46731);
nand UO_2943 (O_2943,N_48001,N_46822);
nand UO_2944 (O_2944,N_49840,N_46949);
and UO_2945 (O_2945,N_49993,N_48969);
nor UO_2946 (O_2946,N_48789,N_48909);
or UO_2947 (O_2947,N_49295,N_46827);
or UO_2948 (O_2948,N_47801,N_49562);
or UO_2949 (O_2949,N_48093,N_46859);
nand UO_2950 (O_2950,N_49485,N_48525);
nand UO_2951 (O_2951,N_48904,N_49565);
nand UO_2952 (O_2952,N_47936,N_48816);
and UO_2953 (O_2953,N_49252,N_46427);
nand UO_2954 (O_2954,N_46819,N_45783);
nor UO_2955 (O_2955,N_47589,N_46750);
nand UO_2956 (O_2956,N_45378,N_46539);
nor UO_2957 (O_2957,N_49138,N_48866);
and UO_2958 (O_2958,N_48224,N_46601);
or UO_2959 (O_2959,N_48746,N_47390);
nor UO_2960 (O_2960,N_48931,N_49360);
or UO_2961 (O_2961,N_47800,N_49571);
xor UO_2962 (O_2962,N_48126,N_48335);
or UO_2963 (O_2963,N_48262,N_48674);
nor UO_2964 (O_2964,N_47305,N_47183);
and UO_2965 (O_2965,N_47118,N_47208);
xnor UO_2966 (O_2966,N_48671,N_45148);
or UO_2967 (O_2967,N_47771,N_46089);
and UO_2968 (O_2968,N_46827,N_48871);
xnor UO_2969 (O_2969,N_46986,N_48215);
and UO_2970 (O_2970,N_47961,N_49288);
and UO_2971 (O_2971,N_47438,N_45927);
xnor UO_2972 (O_2972,N_47309,N_47076);
nand UO_2973 (O_2973,N_48038,N_49678);
nor UO_2974 (O_2974,N_46273,N_45560);
nand UO_2975 (O_2975,N_45077,N_47043);
xor UO_2976 (O_2976,N_46418,N_49664);
nor UO_2977 (O_2977,N_46495,N_45064);
nand UO_2978 (O_2978,N_46412,N_46520);
nand UO_2979 (O_2979,N_46791,N_47364);
or UO_2980 (O_2980,N_45457,N_45546);
or UO_2981 (O_2981,N_49900,N_47261);
xnor UO_2982 (O_2982,N_49370,N_48674);
nor UO_2983 (O_2983,N_49972,N_48054);
or UO_2984 (O_2984,N_49105,N_49222);
or UO_2985 (O_2985,N_45951,N_49866);
or UO_2986 (O_2986,N_48169,N_47195);
nor UO_2987 (O_2987,N_49726,N_48226);
nor UO_2988 (O_2988,N_47624,N_49004);
or UO_2989 (O_2989,N_48062,N_47140);
nor UO_2990 (O_2990,N_48592,N_47700);
nor UO_2991 (O_2991,N_48142,N_46916);
or UO_2992 (O_2992,N_47845,N_46673);
and UO_2993 (O_2993,N_49491,N_45679);
or UO_2994 (O_2994,N_47242,N_48902);
or UO_2995 (O_2995,N_45441,N_48840);
and UO_2996 (O_2996,N_48220,N_46723);
or UO_2997 (O_2997,N_45655,N_47418);
nand UO_2998 (O_2998,N_49057,N_48729);
xor UO_2999 (O_2999,N_47277,N_46213);
and UO_3000 (O_3000,N_47121,N_49126);
nor UO_3001 (O_3001,N_49100,N_49348);
and UO_3002 (O_3002,N_47832,N_45264);
and UO_3003 (O_3003,N_46569,N_46819);
nor UO_3004 (O_3004,N_49838,N_49880);
or UO_3005 (O_3005,N_48349,N_48748);
and UO_3006 (O_3006,N_48829,N_49039);
nand UO_3007 (O_3007,N_46579,N_47168);
nor UO_3008 (O_3008,N_48248,N_48186);
nor UO_3009 (O_3009,N_46017,N_46919);
nand UO_3010 (O_3010,N_49785,N_49117);
or UO_3011 (O_3011,N_49188,N_49214);
and UO_3012 (O_3012,N_49415,N_45902);
and UO_3013 (O_3013,N_45869,N_45573);
nand UO_3014 (O_3014,N_45408,N_45961);
or UO_3015 (O_3015,N_46103,N_45937);
and UO_3016 (O_3016,N_45635,N_49035);
or UO_3017 (O_3017,N_49211,N_49112);
and UO_3018 (O_3018,N_45925,N_48445);
or UO_3019 (O_3019,N_47237,N_47389);
or UO_3020 (O_3020,N_49609,N_49762);
and UO_3021 (O_3021,N_48041,N_49005);
and UO_3022 (O_3022,N_45176,N_45267);
or UO_3023 (O_3023,N_48170,N_49050);
nand UO_3024 (O_3024,N_45244,N_49317);
or UO_3025 (O_3025,N_48366,N_47520);
nand UO_3026 (O_3026,N_47899,N_48932);
xnor UO_3027 (O_3027,N_47071,N_46033);
or UO_3028 (O_3028,N_46316,N_47839);
xnor UO_3029 (O_3029,N_47265,N_49838);
nor UO_3030 (O_3030,N_47623,N_47163);
nand UO_3031 (O_3031,N_49659,N_47476);
or UO_3032 (O_3032,N_45387,N_49593);
nor UO_3033 (O_3033,N_48062,N_46328);
and UO_3034 (O_3034,N_47977,N_48201);
nor UO_3035 (O_3035,N_48937,N_48821);
or UO_3036 (O_3036,N_45491,N_48266);
or UO_3037 (O_3037,N_49456,N_45484);
and UO_3038 (O_3038,N_47958,N_45316);
and UO_3039 (O_3039,N_47088,N_45519);
or UO_3040 (O_3040,N_46884,N_45819);
or UO_3041 (O_3041,N_48355,N_49676);
or UO_3042 (O_3042,N_48374,N_48190);
nand UO_3043 (O_3043,N_46585,N_45266);
or UO_3044 (O_3044,N_45614,N_49942);
nand UO_3045 (O_3045,N_45742,N_45585);
nor UO_3046 (O_3046,N_49557,N_47074);
nand UO_3047 (O_3047,N_47561,N_46078);
nand UO_3048 (O_3048,N_48958,N_49095);
and UO_3049 (O_3049,N_45882,N_47482);
nand UO_3050 (O_3050,N_47387,N_48538);
nor UO_3051 (O_3051,N_48330,N_46616);
xor UO_3052 (O_3052,N_46159,N_48199);
and UO_3053 (O_3053,N_48965,N_47407);
xnor UO_3054 (O_3054,N_46319,N_46444);
or UO_3055 (O_3055,N_46572,N_49161);
and UO_3056 (O_3056,N_47589,N_46026);
and UO_3057 (O_3057,N_49470,N_45305);
nor UO_3058 (O_3058,N_47713,N_49267);
nand UO_3059 (O_3059,N_45701,N_45428);
nor UO_3060 (O_3060,N_49810,N_49421);
or UO_3061 (O_3061,N_48208,N_49716);
nand UO_3062 (O_3062,N_47475,N_48936);
xor UO_3063 (O_3063,N_47939,N_48305);
or UO_3064 (O_3064,N_47556,N_49066);
nand UO_3065 (O_3065,N_49421,N_46683);
and UO_3066 (O_3066,N_47457,N_49399);
and UO_3067 (O_3067,N_47409,N_46098);
and UO_3068 (O_3068,N_49200,N_45560);
nand UO_3069 (O_3069,N_45605,N_49176);
nor UO_3070 (O_3070,N_47853,N_47444);
and UO_3071 (O_3071,N_47637,N_45346);
or UO_3072 (O_3072,N_49748,N_48708);
nor UO_3073 (O_3073,N_46193,N_45931);
nor UO_3074 (O_3074,N_49537,N_45911);
or UO_3075 (O_3075,N_48662,N_48043);
or UO_3076 (O_3076,N_49098,N_47501);
xor UO_3077 (O_3077,N_48234,N_46458);
and UO_3078 (O_3078,N_49373,N_45290);
and UO_3079 (O_3079,N_45898,N_46706);
nor UO_3080 (O_3080,N_49531,N_49355);
and UO_3081 (O_3081,N_45528,N_45220);
and UO_3082 (O_3082,N_45502,N_49464);
or UO_3083 (O_3083,N_48508,N_47116);
nor UO_3084 (O_3084,N_49009,N_47326);
or UO_3085 (O_3085,N_48550,N_46653);
nor UO_3086 (O_3086,N_49190,N_49016);
nor UO_3087 (O_3087,N_49877,N_49396);
and UO_3088 (O_3088,N_47829,N_48491);
and UO_3089 (O_3089,N_45854,N_45231);
nand UO_3090 (O_3090,N_47821,N_48372);
xnor UO_3091 (O_3091,N_47979,N_48341);
and UO_3092 (O_3092,N_45589,N_48180);
and UO_3093 (O_3093,N_46642,N_48106);
nand UO_3094 (O_3094,N_45776,N_45111);
and UO_3095 (O_3095,N_46158,N_45993);
or UO_3096 (O_3096,N_46629,N_49384);
and UO_3097 (O_3097,N_46675,N_47806);
nor UO_3098 (O_3098,N_46852,N_46492);
and UO_3099 (O_3099,N_45214,N_47126);
nor UO_3100 (O_3100,N_49539,N_49356);
nand UO_3101 (O_3101,N_45073,N_49918);
and UO_3102 (O_3102,N_48510,N_48569);
nand UO_3103 (O_3103,N_47689,N_48930);
and UO_3104 (O_3104,N_49466,N_49458);
and UO_3105 (O_3105,N_49829,N_49107);
nor UO_3106 (O_3106,N_49110,N_49027);
or UO_3107 (O_3107,N_45391,N_46739);
or UO_3108 (O_3108,N_47294,N_45361);
xnor UO_3109 (O_3109,N_45094,N_49087);
xnor UO_3110 (O_3110,N_47166,N_47416);
nand UO_3111 (O_3111,N_47186,N_48287);
and UO_3112 (O_3112,N_45404,N_49613);
nor UO_3113 (O_3113,N_46453,N_47832);
nand UO_3114 (O_3114,N_47270,N_49762);
nand UO_3115 (O_3115,N_47024,N_45074);
or UO_3116 (O_3116,N_49456,N_48797);
and UO_3117 (O_3117,N_45697,N_46078);
and UO_3118 (O_3118,N_46042,N_49410);
or UO_3119 (O_3119,N_47400,N_47929);
nand UO_3120 (O_3120,N_47366,N_46709);
and UO_3121 (O_3121,N_49623,N_49650);
and UO_3122 (O_3122,N_46637,N_47841);
nor UO_3123 (O_3123,N_45976,N_45709);
or UO_3124 (O_3124,N_45526,N_46721);
and UO_3125 (O_3125,N_45015,N_46883);
and UO_3126 (O_3126,N_46466,N_49804);
nand UO_3127 (O_3127,N_46629,N_49120);
nor UO_3128 (O_3128,N_45234,N_48998);
and UO_3129 (O_3129,N_45799,N_48483);
nor UO_3130 (O_3130,N_48248,N_46489);
and UO_3131 (O_3131,N_45751,N_49733);
and UO_3132 (O_3132,N_47926,N_45766);
nor UO_3133 (O_3133,N_45743,N_45627);
nand UO_3134 (O_3134,N_48907,N_46967);
xor UO_3135 (O_3135,N_48700,N_45005);
or UO_3136 (O_3136,N_48821,N_46092);
nor UO_3137 (O_3137,N_45060,N_46830);
or UO_3138 (O_3138,N_48632,N_45805);
nor UO_3139 (O_3139,N_47648,N_49211);
and UO_3140 (O_3140,N_48480,N_48574);
or UO_3141 (O_3141,N_46730,N_45270);
and UO_3142 (O_3142,N_46759,N_45249);
and UO_3143 (O_3143,N_46871,N_49112);
nor UO_3144 (O_3144,N_46870,N_46185);
nand UO_3145 (O_3145,N_48388,N_47834);
or UO_3146 (O_3146,N_45837,N_48650);
nor UO_3147 (O_3147,N_46551,N_47272);
and UO_3148 (O_3148,N_49305,N_45666);
xnor UO_3149 (O_3149,N_46277,N_46137);
nor UO_3150 (O_3150,N_45154,N_49374);
nand UO_3151 (O_3151,N_48816,N_48389);
xnor UO_3152 (O_3152,N_48530,N_45815);
nor UO_3153 (O_3153,N_46917,N_46409);
nand UO_3154 (O_3154,N_49642,N_47065);
or UO_3155 (O_3155,N_46549,N_47001);
nand UO_3156 (O_3156,N_47816,N_46613);
nand UO_3157 (O_3157,N_45105,N_49526);
and UO_3158 (O_3158,N_48723,N_47315);
and UO_3159 (O_3159,N_45331,N_49241);
nand UO_3160 (O_3160,N_47129,N_45703);
nor UO_3161 (O_3161,N_48930,N_46414);
nor UO_3162 (O_3162,N_46874,N_46990);
and UO_3163 (O_3163,N_49857,N_47403);
xor UO_3164 (O_3164,N_48658,N_48315);
nand UO_3165 (O_3165,N_46955,N_48606);
nor UO_3166 (O_3166,N_46774,N_45732);
xor UO_3167 (O_3167,N_49460,N_46685);
nor UO_3168 (O_3168,N_46909,N_45312);
nor UO_3169 (O_3169,N_48560,N_49373);
or UO_3170 (O_3170,N_46087,N_47706);
nor UO_3171 (O_3171,N_45566,N_49051);
nand UO_3172 (O_3172,N_49097,N_46967);
nor UO_3173 (O_3173,N_45930,N_45972);
nor UO_3174 (O_3174,N_47890,N_49657);
or UO_3175 (O_3175,N_45030,N_49792);
and UO_3176 (O_3176,N_45825,N_45129);
or UO_3177 (O_3177,N_47228,N_46082);
nand UO_3178 (O_3178,N_48169,N_47694);
or UO_3179 (O_3179,N_45513,N_49627);
nor UO_3180 (O_3180,N_49949,N_46136);
nor UO_3181 (O_3181,N_45286,N_48158);
nor UO_3182 (O_3182,N_48876,N_47682);
or UO_3183 (O_3183,N_45740,N_45585);
nor UO_3184 (O_3184,N_47867,N_47290);
and UO_3185 (O_3185,N_45829,N_46900);
or UO_3186 (O_3186,N_46785,N_49229);
or UO_3187 (O_3187,N_46313,N_49281);
nor UO_3188 (O_3188,N_46800,N_48281);
or UO_3189 (O_3189,N_45100,N_48554);
and UO_3190 (O_3190,N_48231,N_48474);
xnor UO_3191 (O_3191,N_49564,N_45560);
and UO_3192 (O_3192,N_46371,N_46653);
nand UO_3193 (O_3193,N_47258,N_45460);
nand UO_3194 (O_3194,N_46731,N_46103);
nor UO_3195 (O_3195,N_46376,N_46023);
or UO_3196 (O_3196,N_49885,N_47077);
or UO_3197 (O_3197,N_45690,N_46335);
or UO_3198 (O_3198,N_47678,N_48861);
nor UO_3199 (O_3199,N_47028,N_46207);
or UO_3200 (O_3200,N_49556,N_45320);
xnor UO_3201 (O_3201,N_48622,N_46909);
nor UO_3202 (O_3202,N_49990,N_48481);
and UO_3203 (O_3203,N_47594,N_46417);
and UO_3204 (O_3204,N_45591,N_45525);
or UO_3205 (O_3205,N_49961,N_49136);
and UO_3206 (O_3206,N_48754,N_46871);
and UO_3207 (O_3207,N_47081,N_45346);
nor UO_3208 (O_3208,N_49966,N_48109);
nor UO_3209 (O_3209,N_48793,N_48934);
nand UO_3210 (O_3210,N_49428,N_47060);
and UO_3211 (O_3211,N_48909,N_49048);
nor UO_3212 (O_3212,N_47813,N_46303);
or UO_3213 (O_3213,N_46855,N_49460);
or UO_3214 (O_3214,N_47235,N_45964);
nor UO_3215 (O_3215,N_46670,N_46303);
nor UO_3216 (O_3216,N_45019,N_47342);
or UO_3217 (O_3217,N_45428,N_49339);
or UO_3218 (O_3218,N_49424,N_46811);
or UO_3219 (O_3219,N_46831,N_46886);
nand UO_3220 (O_3220,N_45480,N_47734);
xor UO_3221 (O_3221,N_46953,N_45784);
or UO_3222 (O_3222,N_48025,N_49319);
xnor UO_3223 (O_3223,N_49633,N_48139);
nor UO_3224 (O_3224,N_48291,N_46192);
and UO_3225 (O_3225,N_48732,N_46091);
nor UO_3226 (O_3226,N_48269,N_45222);
xor UO_3227 (O_3227,N_45259,N_46784);
and UO_3228 (O_3228,N_48609,N_46342);
xor UO_3229 (O_3229,N_46554,N_49401);
or UO_3230 (O_3230,N_49053,N_46611);
xnor UO_3231 (O_3231,N_48411,N_48935);
nand UO_3232 (O_3232,N_46421,N_46496);
or UO_3233 (O_3233,N_47755,N_45953);
nor UO_3234 (O_3234,N_46164,N_49532);
nand UO_3235 (O_3235,N_45140,N_46914);
and UO_3236 (O_3236,N_48386,N_46508);
nor UO_3237 (O_3237,N_45303,N_49350);
or UO_3238 (O_3238,N_48789,N_47791);
nor UO_3239 (O_3239,N_48029,N_47614);
and UO_3240 (O_3240,N_49943,N_48587);
nand UO_3241 (O_3241,N_49305,N_47541);
nand UO_3242 (O_3242,N_49381,N_45249);
or UO_3243 (O_3243,N_49338,N_45639);
or UO_3244 (O_3244,N_47159,N_45537);
nand UO_3245 (O_3245,N_48150,N_47229);
and UO_3246 (O_3246,N_45995,N_45718);
or UO_3247 (O_3247,N_46480,N_46582);
nand UO_3248 (O_3248,N_45261,N_46945);
nor UO_3249 (O_3249,N_49644,N_48309);
nor UO_3250 (O_3250,N_46271,N_49796);
xnor UO_3251 (O_3251,N_47005,N_47792);
or UO_3252 (O_3252,N_47422,N_47438);
or UO_3253 (O_3253,N_49194,N_49415);
or UO_3254 (O_3254,N_47972,N_45745);
or UO_3255 (O_3255,N_48506,N_49990);
or UO_3256 (O_3256,N_49682,N_46465);
xor UO_3257 (O_3257,N_48562,N_48781);
nor UO_3258 (O_3258,N_49930,N_48940);
and UO_3259 (O_3259,N_45673,N_45630);
nor UO_3260 (O_3260,N_48400,N_47070);
nor UO_3261 (O_3261,N_47314,N_46789);
nor UO_3262 (O_3262,N_45643,N_46892);
nor UO_3263 (O_3263,N_48601,N_47728);
nand UO_3264 (O_3264,N_45667,N_45517);
and UO_3265 (O_3265,N_47235,N_46857);
nor UO_3266 (O_3266,N_45777,N_46629);
nor UO_3267 (O_3267,N_49617,N_47363);
nor UO_3268 (O_3268,N_49009,N_48044);
nor UO_3269 (O_3269,N_48626,N_46913);
nand UO_3270 (O_3270,N_46428,N_46496);
and UO_3271 (O_3271,N_47417,N_46744);
nand UO_3272 (O_3272,N_45027,N_45729);
nand UO_3273 (O_3273,N_48215,N_49325);
xnor UO_3274 (O_3274,N_47394,N_48355);
nand UO_3275 (O_3275,N_45177,N_46615);
nor UO_3276 (O_3276,N_49394,N_46865);
nor UO_3277 (O_3277,N_47608,N_45127);
nand UO_3278 (O_3278,N_45918,N_47525);
and UO_3279 (O_3279,N_48823,N_47007);
and UO_3280 (O_3280,N_45339,N_48683);
nor UO_3281 (O_3281,N_47102,N_49377);
or UO_3282 (O_3282,N_48264,N_47870);
nor UO_3283 (O_3283,N_49121,N_46596);
and UO_3284 (O_3284,N_48972,N_47763);
and UO_3285 (O_3285,N_47533,N_45137);
nor UO_3286 (O_3286,N_45563,N_45469);
or UO_3287 (O_3287,N_48220,N_47592);
nand UO_3288 (O_3288,N_46093,N_47340);
nand UO_3289 (O_3289,N_48945,N_47003);
or UO_3290 (O_3290,N_47886,N_47751);
and UO_3291 (O_3291,N_47498,N_48579);
nand UO_3292 (O_3292,N_47576,N_45640);
or UO_3293 (O_3293,N_47245,N_47881);
and UO_3294 (O_3294,N_48007,N_49451);
xor UO_3295 (O_3295,N_48200,N_47293);
nand UO_3296 (O_3296,N_48146,N_47507);
nor UO_3297 (O_3297,N_47645,N_45088);
nor UO_3298 (O_3298,N_45310,N_45379);
xnor UO_3299 (O_3299,N_45685,N_48473);
and UO_3300 (O_3300,N_45141,N_48744);
and UO_3301 (O_3301,N_49073,N_46664);
and UO_3302 (O_3302,N_47701,N_48573);
or UO_3303 (O_3303,N_47380,N_48812);
or UO_3304 (O_3304,N_49566,N_45973);
nor UO_3305 (O_3305,N_49142,N_45102);
and UO_3306 (O_3306,N_45158,N_46262);
nor UO_3307 (O_3307,N_49806,N_49067);
or UO_3308 (O_3308,N_48563,N_49402);
and UO_3309 (O_3309,N_48406,N_46047);
and UO_3310 (O_3310,N_48769,N_46530);
nor UO_3311 (O_3311,N_45938,N_49625);
and UO_3312 (O_3312,N_47259,N_45845);
or UO_3313 (O_3313,N_48540,N_48220);
nor UO_3314 (O_3314,N_47220,N_47462);
nand UO_3315 (O_3315,N_49682,N_46824);
or UO_3316 (O_3316,N_45896,N_46859);
xnor UO_3317 (O_3317,N_47228,N_49528);
nor UO_3318 (O_3318,N_47640,N_45995);
nor UO_3319 (O_3319,N_48692,N_47047);
nor UO_3320 (O_3320,N_46009,N_46331);
nor UO_3321 (O_3321,N_48765,N_46892);
or UO_3322 (O_3322,N_45518,N_48241);
nor UO_3323 (O_3323,N_47737,N_48672);
or UO_3324 (O_3324,N_47865,N_45747);
and UO_3325 (O_3325,N_48839,N_49679);
nand UO_3326 (O_3326,N_45115,N_45679);
or UO_3327 (O_3327,N_49683,N_47925);
nand UO_3328 (O_3328,N_49495,N_47822);
or UO_3329 (O_3329,N_46267,N_47574);
or UO_3330 (O_3330,N_46874,N_46096);
or UO_3331 (O_3331,N_47668,N_47368);
or UO_3332 (O_3332,N_45175,N_47656);
and UO_3333 (O_3333,N_48822,N_48907);
and UO_3334 (O_3334,N_49423,N_48487);
or UO_3335 (O_3335,N_49892,N_45522);
nand UO_3336 (O_3336,N_46564,N_45578);
nor UO_3337 (O_3337,N_45884,N_45084);
and UO_3338 (O_3338,N_46057,N_49466);
and UO_3339 (O_3339,N_45378,N_46112);
nand UO_3340 (O_3340,N_45658,N_46597);
or UO_3341 (O_3341,N_46015,N_46746);
nand UO_3342 (O_3342,N_46481,N_49183);
and UO_3343 (O_3343,N_48574,N_45247);
or UO_3344 (O_3344,N_48203,N_47727);
nand UO_3345 (O_3345,N_47113,N_48413);
or UO_3346 (O_3346,N_46538,N_48750);
or UO_3347 (O_3347,N_45908,N_47835);
nand UO_3348 (O_3348,N_46757,N_47103);
nor UO_3349 (O_3349,N_49036,N_45448);
nor UO_3350 (O_3350,N_45580,N_46067);
or UO_3351 (O_3351,N_48752,N_47853);
or UO_3352 (O_3352,N_47986,N_47715);
or UO_3353 (O_3353,N_46962,N_47235);
nand UO_3354 (O_3354,N_47988,N_46082);
and UO_3355 (O_3355,N_47692,N_45294);
or UO_3356 (O_3356,N_49829,N_45873);
or UO_3357 (O_3357,N_46610,N_48554);
and UO_3358 (O_3358,N_47161,N_48939);
nor UO_3359 (O_3359,N_45879,N_45350);
nand UO_3360 (O_3360,N_47096,N_48382);
or UO_3361 (O_3361,N_47070,N_45948);
nor UO_3362 (O_3362,N_48750,N_49179);
and UO_3363 (O_3363,N_47144,N_45931);
nand UO_3364 (O_3364,N_49027,N_46203);
nand UO_3365 (O_3365,N_49939,N_49278);
and UO_3366 (O_3366,N_48421,N_46578);
nand UO_3367 (O_3367,N_49631,N_47393);
or UO_3368 (O_3368,N_45069,N_46999);
and UO_3369 (O_3369,N_46898,N_46968);
nor UO_3370 (O_3370,N_45759,N_48251);
or UO_3371 (O_3371,N_47397,N_45404);
or UO_3372 (O_3372,N_49693,N_45349);
or UO_3373 (O_3373,N_45549,N_49219);
and UO_3374 (O_3374,N_48880,N_46155);
and UO_3375 (O_3375,N_45328,N_48878);
and UO_3376 (O_3376,N_49705,N_46260);
or UO_3377 (O_3377,N_45071,N_45641);
or UO_3378 (O_3378,N_49895,N_49719);
and UO_3379 (O_3379,N_46238,N_46842);
and UO_3380 (O_3380,N_45181,N_49157);
nor UO_3381 (O_3381,N_47236,N_48509);
nand UO_3382 (O_3382,N_46337,N_47827);
nand UO_3383 (O_3383,N_46019,N_48518);
and UO_3384 (O_3384,N_49892,N_49042);
nand UO_3385 (O_3385,N_45394,N_49198);
xor UO_3386 (O_3386,N_46939,N_46574);
and UO_3387 (O_3387,N_45272,N_47222);
or UO_3388 (O_3388,N_47945,N_45042);
nor UO_3389 (O_3389,N_48696,N_46436);
xnor UO_3390 (O_3390,N_45277,N_48080);
and UO_3391 (O_3391,N_49760,N_45892);
nand UO_3392 (O_3392,N_47008,N_49914);
nand UO_3393 (O_3393,N_45223,N_49926);
nand UO_3394 (O_3394,N_45241,N_46255);
nand UO_3395 (O_3395,N_46667,N_45964);
nor UO_3396 (O_3396,N_47731,N_46979);
nor UO_3397 (O_3397,N_45498,N_48803);
xor UO_3398 (O_3398,N_46450,N_45415);
xnor UO_3399 (O_3399,N_45986,N_49795);
nand UO_3400 (O_3400,N_49855,N_48262);
and UO_3401 (O_3401,N_46518,N_45300);
nor UO_3402 (O_3402,N_49084,N_47254);
and UO_3403 (O_3403,N_45007,N_47372);
or UO_3404 (O_3404,N_48009,N_47663);
nor UO_3405 (O_3405,N_46014,N_48813);
nand UO_3406 (O_3406,N_48550,N_47509);
nand UO_3407 (O_3407,N_49792,N_47359);
xor UO_3408 (O_3408,N_46281,N_45921);
or UO_3409 (O_3409,N_47233,N_46382);
or UO_3410 (O_3410,N_46741,N_45574);
or UO_3411 (O_3411,N_47036,N_46019);
xor UO_3412 (O_3412,N_45188,N_47483);
nor UO_3413 (O_3413,N_45163,N_49192);
and UO_3414 (O_3414,N_49634,N_46933);
or UO_3415 (O_3415,N_47508,N_47600);
nor UO_3416 (O_3416,N_48897,N_48210);
nand UO_3417 (O_3417,N_48258,N_49277);
nor UO_3418 (O_3418,N_49743,N_49396);
or UO_3419 (O_3419,N_48673,N_48653);
nand UO_3420 (O_3420,N_45630,N_46972);
and UO_3421 (O_3421,N_47308,N_45555);
xor UO_3422 (O_3422,N_48568,N_48848);
and UO_3423 (O_3423,N_45750,N_45338);
and UO_3424 (O_3424,N_47461,N_47867);
nand UO_3425 (O_3425,N_47636,N_45728);
nor UO_3426 (O_3426,N_48787,N_48992);
and UO_3427 (O_3427,N_45465,N_46431);
or UO_3428 (O_3428,N_49703,N_49300);
xnor UO_3429 (O_3429,N_48912,N_46823);
and UO_3430 (O_3430,N_48032,N_45609);
nand UO_3431 (O_3431,N_47641,N_45667);
nor UO_3432 (O_3432,N_47628,N_47024);
or UO_3433 (O_3433,N_49895,N_45281);
nor UO_3434 (O_3434,N_47393,N_48761);
and UO_3435 (O_3435,N_45479,N_46162);
nand UO_3436 (O_3436,N_46472,N_45013);
nand UO_3437 (O_3437,N_46827,N_48165);
and UO_3438 (O_3438,N_46506,N_45629);
xnor UO_3439 (O_3439,N_47637,N_49202);
or UO_3440 (O_3440,N_46103,N_45095);
nand UO_3441 (O_3441,N_49677,N_48046);
nor UO_3442 (O_3442,N_48397,N_49913);
nand UO_3443 (O_3443,N_49203,N_49514);
nor UO_3444 (O_3444,N_47555,N_49979);
and UO_3445 (O_3445,N_45986,N_47923);
and UO_3446 (O_3446,N_48757,N_48321);
or UO_3447 (O_3447,N_46895,N_46544);
or UO_3448 (O_3448,N_48464,N_49413);
and UO_3449 (O_3449,N_45164,N_46890);
or UO_3450 (O_3450,N_48555,N_45089);
nor UO_3451 (O_3451,N_49241,N_47131);
or UO_3452 (O_3452,N_48474,N_48664);
nand UO_3453 (O_3453,N_45550,N_48864);
nor UO_3454 (O_3454,N_49059,N_48991);
nor UO_3455 (O_3455,N_45089,N_49496);
or UO_3456 (O_3456,N_47462,N_48896);
nor UO_3457 (O_3457,N_47916,N_47184);
xor UO_3458 (O_3458,N_47716,N_48267);
nor UO_3459 (O_3459,N_47319,N_47616);
nor UO_3460 (O_3460,N_47158,N_47528);
nor UO_3461 (O_3461,N_47769,N_48496);
nand UO_3462 (O_3462,N_48540,N_49589);
nand UO_3463 (O_3463,N_45945,N_46889);
nand UO_3464 (O_3464,N_49388,N_48142);
and UO_3465 (O_3465,N_47146,N_48237);
nor UO_3466 (O_3466,N_45213,N_46505);
nand UO_3467 (O_3467,N_47463,N_47286);
and UO_3468 (O_3468,N_49957,N_47295);
nor UO_3469 (O_3469,N_48957,N_48503);
nand UO_3470 (O_3470,N_46332,N_47081);
and UO_3471 (O_3471,N_48808,N_48805);
or UO_3472 (O_3472,N_47153,N_47757);
nor UO_3473 (O_3473,N_48740,N_49354);
and UO_3474 (O_3474,N_45635,N_49082);
or UO_3475 (O_3475,N_49998,N_49482);
or UO_3476 (O_3476,N_48006,N_45265);
nand UO_3477 (O_3477,N_46560,N_47159);
nor UO_3478 (O_3478,N_45666,N_48927);
or UO_3479 (O_3479,N_46932,N_45323);
and UO_3480 (O_3480,N_45051,N_45030);
and UO_3481 (O_3481,N_45577,N_48872);
nand UO_3482 (O_3482,N_47718,N_47116);
xor UO_3483 (O_3483,N_48319,N_46287);
nand UO_3484 (O_3484,N_45421,N_46175);
nor UO_3485 (O_3485,N_47423,N_49824);
or UO_3486 (O_3486,N_48219,N_48738);
and UO_3487 (O_3487,N_49328,N_46057);
nor UO_3488 (O_3488,N_47397,N_47525);
or UO_3489 (O_3489,N_45989,N_48251);
nand UO_3490 (O_3490,N_49618,N_49960);
xnor UO_3491 (O_3491,N_48758,N_45514);
nor UO_3492 (O_3492,N_47626,N_49366);
xnor UO_3493 (O_3493,N_46639,N_46783);
nand UO_3494 (O_3494,N_45114,N_47145);
xnor UO_3495 (O_3495,N_47495,N_49647);
nor UO_3496 (O_3496,N_49675,N_49793);
nor UO_3497 (O_3497,N_48284,N_48034);
nor UO_3498 (O_3498,N_45459,N_48918);
nor UO_3499 (O_3499,N_45742,N_45432);
nand UO_3500 (O_3500,N_46762,N_47217);
or UO_3501 (O_3501,N_45751,N_45108);
nand UO_3502 (O_3502,N_47775,N_49354);
or UO_3503 (O_3503,N_45687,N_46464);
nand UO_3504 (O_3504,N_48840,N_47836);
and UO_3505 (O_3505,N_49015,N_48495);
or UO_3506 (O_3506,N_46411,N_47809);
nand UO_3507 (O_3507,N_45110,N_47138);
and UO_3508 (O_3508,N_48933,N_47060);
nand UO_3509 (O_3509,N_45936,N_47552);
nor UO_3510 (O_3510,N_45791,N_46457);
nor UO_3511 (O_3511,N_45858,N_49210);
or UO_3512 (O_3512,N_47100,N_48492);
nor UO_3513 (O_3513,N_46487,N_46770);
and UO_3514 (O_3514,N_47936,N_46964);
nand UO_3515 (O_3515,N_49614,N_46047);
nor UO_3516 (O_3516,N_47047,N_48876);
xor UO_3517 (O_3517,N_46840,N_47571);
nor UO_3518 (O_3518,N_47953,N_47031);
nand UO_3519 (O_3519,N_46293,N_46893);
or UO_3520 (O_3520,N_47309,N_46583);
and UO_3521 (O_3521,N_46747,N_47850);
and UO_3522 (O_3522,N_46024,N_48876);
and UO_3523 (O_3523,N_46575,N_48308);
nand UO_3524 (O_3524,N_45328,N_49280);
nor UO_3525 (O_3525,N_46935,N_49676);
nor UO_3526 (O_3526,N_47554,N_47445);
nand UO_3527 (O_3527,N_49787,N_46622);
and UO_3528 (O_3528,N_46062,N_46618);
nor UO_3529 (O_3529,N_48189,N_47676);
xor UO_3530 (O_3530,N_47757,N_47633);
xnor UO_3531 (O_3531,N_45626,N_47306);
nor UO_3532 (O_3532,N_49631,N_46340);
or UO_3533 (O_3533,N_47062,N_47794);
or UO_3534 (O_3534,N_49311,N_45949);
nor UO_3535 (O_3535,N_48845,N_48586);
or UO_3536 (O_3536,N_46017,N_45572);
nor UO_3537 (O_3537,N_46934,N_49229);
and UO_3538 (O_3538,N_46291,N_46951);
nor UO_3539 (O_3539,N_45037,N_45832);
nand UO_3540 (O_3540,N_46044,N_45483);
and UO_3541 (O_3541,N_46052,N_46323);
and UO_3542 (O_3542,N_49752,N_45164);
and UO_3543 (O_3543,N_45088,N_48905);
or UO_3544 (O_3544,N_48598,N_49568);
nor UO_3545 (O_3545,N_48955,N_45380);
or UO_3546 (O_3546,N_46809,N_48236);
or UO_3547 (O_3547,N_46218,N_47174);
or UO_3548 (O_3548,N_45321,N_45641);
nor UO_3549 (O_3549,N_47296,N_48514);
nand UO_3550 (O_3550,N_46411,N_49967);
nand UO_3551 (O_3551,N_46550,N_49322);
nor UO_3552 (O_3552,N_48836,N_46294);
and UO_3553 (O_3553,N_47298,N_47727);
nand UO_3554 (O_3554,N_46478,N_46332);
and UO_3555 (O_3555,N_45305,N_49349);
nor UO_3556 (O_3556,N_45113,N_47802);
nor UO_3557 (O_3557,N_48611,N_47830);
nand UO_3558 (O_3558,N_48964,N_49385);
and UO_3559 (O_3559,N_46708,N_49165);
xnor UO_3560 (O_3560,N_48527,N_47763);
nor UO_3561 (O_3561,N_46120,N_48646);
or UO_3562 (O_3562,N_45081,N_47263);
and UO_3563 (O_3563,N_45340,N_45727);
xnor UO_3564 (O_3564,N_49727,N_49411);
nor UO_3565 (O_3565,N_47348,N_45426);
nand UO_3566 (O_3566,N_48729,N_46017);
or UO_3567 (O_3567,N_46365,N_45161);
and UO_3568 (O_3568,N_48138,N_45280);
nand UO_3569 (O_3569,N_49735,N_46991);
and UO_3570 (O_3570,N_49055,N_49891);
and UO_3571 (O_3571,N_46015,N_46020);
and UO_3572 (O_3572,N_45594,N_49696);
or UO_3573 (O_3573,N_45983,N_48984);
and UO_3574 (O_3574,N_49938,N_45233);
nand UO_3575 (O_3575,N_49992,N_47963);
xnor UO_3576 (O_3576,N_47612,N_47347);
and UO_3577 (O_3577,N_49784,N_49018);
nand UO_3578 (O_3578,N_46578,N_45630);
and UO_3579 (O_3579,N_46130,N_49233);
or UO_3580 (O_3580,N_47356,N_45966);
or UO_3581 (O_3581,N_46709,N_48317);
and UO_3582 (O_3582,N_45507,N_46711);
xnor UO_3583 (O_3583,N_49253,N_48148);
nand UO_3584 (O_3584,N_49357,N_46854);
nor UO_3585 (O_3585,N_49735,N_47690);
or UO_3586 (O_3586,N_48724,N_45835);
and UO_3587 (O_3587,N_48308,N_45738);
nand UO_3588 (O_3588,N_47558,N_49558);
xor UO_3589 (O_3589,N_46805,N_49859);
or UO_3590 (O_3590,N_45142,N_48955);
and UO_3591 (O_3591,N_47243,N_47277);
and UO_3592 (O_3592,N_47228,N_47172);
nor UO_3593 (O_3593,N_46050,N_48318);
nor UO_3594 (O_3594,N_49695,N_48672);
xnor UO_3595 (O_3595,N_46960,N_46816);
xnor UO_3596 (O_3596,N_49365,N_45991);
nand UO_3597 (O_3597,N_47805,N_47709);
nand UO_3598 (O_3598,N_47247,N_45038);
nand UO_3599 (O_3599,N_46235,N_47993);
nor UO_3600 (O_3600,N_48824,N_48134);
and UO_3601 (O_3601,N_47574,N_47883);
nor UO_3602 (O_3602,N_48440,N_47333);
or UO_3603 (O_3603,N_49485,N_49714);
or UO_3604 (O_3604,N_48067,N_48696);
or UO_3605 (O_3605,N_46436,N_49634);
xnor UO_3606 (O_3606,N_47355,N_49591);
or UO_3607 (O_3607,N_45746,N_47586);
or UO_3608 (O_3608,N_46904,N_47909);
or UO_3609 (O_3609,N_48824,N_48828);
nand UO_3610 (O_3610,N_49480,N_49893);
or UO_3611 (O_3611,N_47783,N_46677);
xnor UO_3612 (O_3612,N_48023,N_49103);
or UO_3613 (O_3613,N_48252,N_49810);
nor UO_3614 (O_3614,N_46448,N_48591);
or UO_3615 (O_3615,N_47751,N_48464);
or UO_3616 (O_3616,N_47569,N_46034);
or UO_3617 (O_3617,N_48308,N_49241);
or UO_3618 (O_3618,N_47358,N_45333);
or UO_3619 (O_3619,N_49224,N_47019);
nand UO_3620 (O_3620,N_45107,N_49483);
or UO_3621 (O_3621,N_45736,N_47921);
nand UO_3622 (O_3622,N_49557,N_46398);
nor UO_3623 (O_3623,N_48289,N_46857);
and UO_3624 (O_3624,N_46898,N_47577);
nor UO_3625 (O_3625,N_47497,N_47422);
or UO_3626 (O_3626,N_46888,N_46544);
nand UO_3627 (O_3627,N_45567,N_49522);
or UO_3628 (O_3628,N_49423,N_46471);
or UO_3629 (O_3629,N_46659,N_48859);
or UO_3630 (O_3630,N_45352,N_45161);
xor UO_3631 (O_3631,N_46700,N_45699);
and UO_3632 (O_3632,N_47818,N_45970);
nor UO_3633 (O_3633,N_47428,N_48262);
xor UO_3634 (O_3634,N_47065,N_46333);
or UO_3635 (O_3635,N_46734,N_48968);
nor UO_3636 (O_3636,N_49220,N_49620);
nand UO_3637 (O_3637,N_45890,N_49672);
nor UO_3638 (O_3638,N_45413,N_48838);
xor UO_3639 (O_3639,N_46236,N_47952);
and UO_3640 (O_3640,N_45306,N_46103);
nor UO_3641 (O_3641,N_48687,N_47423);
or UO_3642 (O_3642,N_49710,N_46019);
nand UO_3643 (O_3643,N_47197,N_47226);
nand UO_3644 (O_3644,N_46312,N_46887);
nor UO_3645 (O_3645,N_48485,N_45010);
nor UO_3646 (O_3646,N_45649,N_47771);
or UO_3647 (O_3647,N_48946,N_47795);
nand UO_3648 (O_3648,N_49307,N_45266);
nor UO_3649 (O_3649,N_49345,N_47779);
and UO_3650 (O_3650,N_45887,N_48046);
or UO_3651 (O_3651,N_49910,N_49413);
xnor UO_3652 (O_3652,N_45008,N_48018);
nor UO_3653 (O_3653,N_49277,N_48013);
nand UO_3654 (O_3654,N_47727,N_48478);
nor UO_3655 (O_3655,N_45595,N_49633);
nor UO_3656 (O_3656,N_47068,N_47073);
and UO_3657 (O_3657,N_49519,N_46677);
and UO_3658 (O_3658,N_48698,N_47685);
nand UO_3659 (O_3659,N_45439,N_47751);
xnor UO_3660 (O_3660,N_46416,N_48178);
or UO_3661 (O_3661,N_48777,N_49344);
nor UO_3662 (O_3662,N_49170,N_49702);
nand UO_3663 (O_3663,N_48081,N_48576);
or UO_3664 (O_3664,N_46149,N_46072);
or UO_3665 (O_3665,N_47848,N_48796);
xor UO_3666 (O_3666,N_47749,N_47229);
and UO_3667 (O_3667,N_47621,N_45208);
or UO_3668 (O_3668,N_45684,N_46229);
nand UO_3669 (O_3669,N_45782,N_47314);
and UO_3670 (O_3670,N_48567,N_49657);
nor UO_3671 (O_3671,N_48714,N_48264);
and UO_3672 (O_3672,N_46424,N_47606);
nor UO_3673 (O_3673,N_45130,N_49132);
nand UO_3674 (O_3674,N_49647,N_49998);
and UO_3675 (O_3675,N_45396,N_46255);
nand UO_3676 (O_3676,N_48117,N_48619);
or UO_3677 (O_3677,N_46093,N_47366);
nor UO_3678 (O_3678,N_49506,N_48898);
nor UO_3679 (O_3679,N_47249,N_46254);
and UO_3680 (O_3680,N_49077,N_49334);
nor UO_3681 (O_3681,N_48547,N_48947);
nor UO_3682 (O_3682,N_47541,N_48853);
and UO_3683 (O_3683,N_48287,N_47462);
nor UO_3684 (O_3684,N_46914,N_49284);
or UO_3685 (O_3685,N_47439,N_47909);
nor UO_3686 (O_3686,N_46225,N_48808);
nor UO_3687 (O_3687,N_45757,N_45214);
nor UO_3688 (O_3688,N_48382,N_49200);
nand UO_3689 (O_3689,N_49582,N_47352);
or UO_3690 (O_3690,N_49643,N_46253);
or UO_3691 (O_3691,N_46801,N_48994);
and UO_3692 (O_3692,N_47869,N_46559);
or UO_3693 (O_3693,N_46455,N_47875);
and UO_3694 (O_3694,N_46145,N_45158);
xnor UO_3695 (O_3695,N_48347,N_45842);
or UO_3696 (O_3696,N_45518,N_48028);
and UO_3697 (O_3697,N_49530,N_47054);
nand UO_3698 (O_3698,N_49611,N_46448);
nand UO_3699 (O_3699,N_46283,N_45179);
nor UO_3700 (O_3700,N_47185,N_49534);
or UO_3701 (O_3701,N_49430,N_45085);
nor UO_3702 (O_3702,N_48066,N_46343);
nand UO_3703 (O_3703,N_46723,N_47641);
and UO_3704 (O_3704,N_48460,N_48798);
and UO_3705 (O_3705,N_48525,N_49578);
or UO_3706 (O_3706,N_46951,N_49967);
nor UO_3707 (O_3707,N_47145,N_45774);
nor UO_3708 (O_3708,N_46058,N_47869);
and UO_3709 (O_3709,N_45983,N_47679);
nand UO_3710 (O_3710,N_48316,N_47123);
or UO_3711 (O_3711,N_46931,N_47508);
nor UO_3712 (O_3712,N_48954,N_46144);
nand UO_3713 (O_3713,N_45393,N_47329);
nand UO_3714 (O_3714,N_46696,N_47514);
xnor UO_3715 (O_3715,N_45347,N_46338);
nor UO_3716 (O_3716,N_49634,N_47879);
nand UO_3717 (O_3717,N_49441,N_49259);
nor UO_3718 (O_3718,N_49064,N_45433);
nand UO_3719 (O_3719,N_48600,N_46491);
or UO_3720 (O_3720,N_46088,N_49025);
xnor UO_3721 (O_3721,N_45762,N_49606);
or UO_3722 (O_3722,N_45431,N_48920);
nor UO_3723 (O_3723,N_48287,N_49933);
or UO_3724 (O_3724,N_46908,N_47795);
and UO_3725 (O_3725,N_47938,N_46103);
nand UO_3726 (O_3726,N_49522,N_45800);
and UO_3727 (O_3727,N_45933,N_47230);
or UO_3728 (O_3728,N_49685,N_45876);
nor UO_3729 (O_3729,N_46015,N_48503);
nand UO_3730 (O_3730,N_49157,N_45514);
nor UO_3731 (O_3731,N_49691,N_49362);
or UO_3732 (O_3732,N_46067,N_47723);
nor UO_3733 (O_3733,N_47463,N_48152);
xnor UO_3734 (O_3734,N_46632,N_49040);
and UO_3735 (O_3735,N_48497,N_45411);
nor UO_3736 (O_3736,N_49708,N_47016);
and UO_3737 (O_3737,N_49970,N_46711);
nand UO_3738 (O_3738,N_48379,N_46053);
xnor UO_3739 (O_3739,N_45983,N_46861);
and UO_3740 (O_3740,N_48465,N_48323);
and UO_3741 (O_3741,N_45107,N_47030);
or UO_3742 (O_3742,N_47048,N_46049);
nor UO_3743 (O_3743,N_49759,N_47496);
nor UO_3744 (O_3744,N_45044,N_48272);
and UO_3745 (O_3745,N_46415,N_45418);
and UO_3746 (O_3746,N_46411,N_45819);
nand UO_3747 (O_3747,N_48323,N_47967);
nor UO_3748 (O_3748,N_49768,N_47608);
nand UO_3749 (O_3749,N_45908,N_48349);
nand UO_3750 (O_3750,N_45813,N_46983);
nor UO_3751 (O_3751,N_49927,N_46679);
nor UO_3752 (O_3752,N_49222,N_49435);
xor UO_3753 (O_3753,N_49294,N_46829);
xor UO_3754 (O_3754,N_49461,N_45198);
nand UO_3755 (O_3755,N_46630,N_49783);
nor UO_3756 (O_3756,N_45954,N_49125);
nor UO_3757 (O_3757,N_49418,N_49846);
and UO_3758 (O_3758,N_49250,N_47581);
and UO_3759 (O_3759,N_49384,N_45273);
nand UO_3760 (O_3760,N_48056,N_49754);
nor UO_3761 (O_3761,N_47205,N_49059);
or UO_3762 (O_3762,N_45899,N_47064);
nor UO_3763 (O_3763,N_47454,N_47550);
nor UO_3764 (O_3764,N_45467,N_49496);
nor UO_3765 (O_3765,N_47405,N_49387);
or UO_3766 (O_3766,N_48028,N_49388);
nand UO_3767 (O_3767,N_49887,N_49945);
or UO_3768 (O_3768,N_48517,N_45430);
nand UO_3769 (O_3769,N_47776,N_49610);
nand UO_3770 (O_3770,N_49335,N_49713);
nand UO_3771 (O_3771,N_49301,N_45180);
or UO_3772 (O_3772,N_48309,N_48690);
nor UO_3773 (O_3773,N_49446,N_48413);
or UO_3774 (O_3774,N_45148,N_48504);
xor UO_3775 (O_3775,N_46338,N_47427);
nor UO_3776 (O_3776,N_49072,N_49399);
or UO_3777 (O_3777,N_45779,N_48589);
or UO_3778 (O_3778,N_46984,N_46847);
and UO_3779 (O_3779,N_47481,N_48989);
nor UO_3780 (O_3780,N_47543,N_45136);
nand UO_3781 (O_3781,N_48127,N_47524);
or UO_3782 (O_3782,N_47339,N_45150);
nand UO_3783 (O_3783,N_45170,N_48653);
nand UO_3784 (O_3784,N_48503,N_45707);
xor UO_3785 (O_3785,N_46461,N_48290);
or UO_3786 (O_3786,N_47498,N_48412);
and UO_3787 (O_3787,N_47288,N_47453);
nor UO_3788 (O_3788,N_49418,N_48662);
and UO_3789 (O_3789,N_48914,N_47332);
nor UO_3790 (O_3790,N_49053,N_49383);
nor UO_3791 (O_3791,N_49840,N_49311);
and UO_3792 (O_3792,N_45744,N_48434);
and UO_3793 (O_3793,N_48972,N_48942);
nor UO_3794 (O_3794,N_49405,N_46400);
nand UO_3795 (O_3795,N_47954,N_47427);
nand UO_3796 (O_3796,N_45801,N_48941);
and UO_3797 (O_3797,N_48541,N_46598);
and UO_3798 (O_3798,N_47270,N_49081);
and UO_3799 (O_3799,N_46874,N_49076);
nand UO_3800 (O_3800,N_45476,N_49253);
nor UO_3801 (O_3801,N_49933,N_48531);
or UO_3802 (O_3802,N_49362,N_45914);
nand UO_3803 (O_3803,N_45658,N_49466);
nand UO_3804 (O_3804,N_45946,N_46309);
xor UO_3805 (O_3805,N_46901,N_46618);
nor UO_3806 (O_3806,N_47114,N_45260);
and UO_3807 (O_3807,N_45914,N_47398);
nor UO_3808 (O_3808,N_48807,N_49223);
or UO_3809 (O_3809,N_49777,N_49603);
nand UO_3810 (O_3810,N_49386,N_45632);
or UO_3811 (O_3811,N_47848,N_49032);
nor UO_3812 (O_3812,N_49793,N_48632);
and UO_3813 (O_3813,N_49759,N_49309);
or UO_3814 (O_3814,N_46150,N_47292);
nor UO_3815 (O_3815,N_47253,N_47727);
and UO_3816 (O_3816,N_45938,N_48914);
or UO_3817 (O_3817,N_49748,N_47900);
nand UO_3818 (O_3818,N_48238,N_48756);
or UO_3819 (O_3819,N_45740,N_47891);
or UO_3820 (O_3820,N_49002,N_49903);
and UO_3821 (O_3821,N_46269,N_48708);
nor UO_3822 (O_3822,N_47785,N_45369);
or UO_3823 (O_3823,N_49993,N_46807);
or UO_3824 (O_3824,N_45925,N_47281);
and UO_3825 (O_3825,N_47725,N_49657);
nand UO_3826 (O_3826,N_49708,N_49912);
and UO_3827 (O_3827,N_46893,N_47345);
or UO_3828 (O_3828,N_45453,N_47820);
or UO_3829 (O_3829,N_45175,N_47909);
xor UO_3830 (O_3830,N_49773,N_47967);
and UO_3831 (O_3831,N_46206,N_47806);
xnor UO_3832 (O_3832,N_49274,N_47331);
nand UO_3833 (O_3833,N_48980,N_49153);
or UO_3834 (O_3834,N_49503,N_49342);
xnor UO_3835 (O_3835,N_45826,N_47374);
nand UO_3836 (O_3836,N_46622,N_49790);
and UO_3837 (O_3837,N_49966,N_48730);
nor UO_3838 (O_3838,N_46690,N_48291);
nor UO_3839 (O_3839,N_45437,N_48451);
xor UO_3840 (O_3840,N_46063,N_46824);
xnor UO_3841 (O_3841,N_45803,N_46531);
nand UO_3842 (O_3842,N_47599,N_45022);
or UO_3843 (O_3843,N_47730,N_45321);
and UO_3844 (O_3844,N_47232,N_48057);
nor UO_3845 (O_3845,N_45369,N_46246);
nand UO_3846 (O_3846,N_49541,N_48247);
xnor UO_3847 (O_3847,N_45944,N_45938);
nor UO_3848 (O_3848,N_47352,N_49392);
and UO_3849 (O_3849,N_49222,N_45382);
or UO_3850 (O_3850,N_45737,N_48874);
or UO_3851 (O_3851,N_48227,N_49062);
and UO_3852 (O_3852,N_48397,N_45002);
nor UO_3853 (O_3853,N_45253,N_47986);
and UO_3854 (O_3854,N_47424,N_49776);
or UO_3855 (O_3855,N_46080,N_49841);
or UO_3856 (O_3856,N_48453,N_49798);
or UO_3857 (O_3857,N_46213,N_45723);
nand UO_3858 (O_3858,N_45220,N_45675);
or UO_3859 (O_3859,N_49539,N_47986);
nand UO_3860 (O_3860,N_45908,N_45914);
or UO_3861 (O_3861,N_49721,N_45919);
nand UO_3862 (O_3862,N_45289,N_46483);
nor UO_3863 (O_3863,N_49616,N_45748);
and UO_3864 (O_3864,N_48014,N_47241);
or UO_3865 (O_3865,N_48697,N_45369);
or UO_3866 (O_3866,N_49735,N_47013);
nand UO_3867 (O_3867,N_45567,N_49128);
or UO_3868 (O_3868,N_48224,N_49114);
nor UO_3869 (O_3869,N_46954,N_46634);
nand UO_3870 (O_3870,N_49131,N_46837);
or UO_3871 (O_3871,N_46264,N_47865);
nand UO_3872 (O_3872,N_47682,N_48898);
nor UO_3873 (O_3873,N_45747,N_45942);
nor UO_3874 (O_3874,N_47845,N_45158);
nor UO_3875 (O_3875,N_49098,N_47544);
nor UO_3876 (O_3876,N_45520,N_47716);
or UO_3877 (O_3877,N_49058,N_48100);
nand UO_3878 (O_3878,N_49237,N_47039);
or UO_3879 (O_3879,N_48213,N_46663);
nor UO_3880 (O_3880,N_49571,N_49016);
or UO_3881 (O_3881,N_47577,N_45813);
and UO_3882 (O_3882,N_47969,N_47362);
or UO_3883 (O_3883,N_46065,N_47132);
or UO_3884 (O_3884,N_48225,N_45075);
or UO_3885 (O_3885,N_46735,N_46313);
or UO_3886 (O_3886,N_45182,N_49050);
or UO_3887 (O_3887,N_48563,N_45685);
nor UO_3888 (O_3888,N_47765,N_45328);
nor UO_3889 (O_3889,N_47114,N_48100);
nand UO_3890 (O_3890,N_49257,N_48969);
or UO_3891 (O_3891,N_45947,N_49248);
or UO_3892 (O_3892,N_47115,N_49868);
nand UO_3893 (O_3893,N_46286,N_46886);
nand UO_3894 (O_3894,N_48721,N_47952);
nor UO_3895 (O_3895,N_46256,N_47694);
or UO_3896 (O_3896,N_49417,N_46843);
and UO_3897 (O_3897,N_46586,N_48219);
xor UO_3898 (O_3898,N_45304,N_46528);
nor UO_3899 (O_3899,N_47899,N_46386);
and UO_3900 (O_3900,N_46942,N_45056);
xor UO_3901 (O_3901,N_48725,N_48416);
or UO_3902 (O_3902,N_45867,N_46815);
nor UO_3903 (O_3903,N_49941,N_46761);
and UO_3904 (O_3904,N_45021,N_48559);
nand UO_3905 (O_3905,N_48983,N_45622);
nor UO_3906 (O_3906,N_49995,N_47804);
or UO_3907 (O_3907,N_45970,N_48477);
or UO_3908 (O_3908,N_48445,N_49524);
and UO_3909 (O_3909,N_49309,N_48641);
and UO_3910 (O_3910,N_49471,N_47581);
nand UO_3911 (O_3911,N_47848,N_46272);
xnor UO_3912 (O_3912,N_46165,N_45792);
or UO_3913 (O_3913,N_45537,N_47074);
or UO_3914 (O_3914,N_45744,N_45559);
and UO_3915 (O_3915,N_46413,N_48633);
nor UO_3916 (O_3916,N_45610,N_45636);
nor UO_3917 (O_3917,N_47156,N_47731);
or UO_3918 (O_3918,N_46041,N_48215);
nor UO_3919 (O_3919,N_49163,N_48850);
nand UO_3920 (O_3920,N_46818,N_48436);
nand UO_3921 (O_3921,N_45952,N_48367);
nor UO_3922 (O_3922,N_48874,N_49408);
xor UO_3923 (O_3923,N_48001,N_49462);
nand UO_3924 (O_3924,N_45575,N_49160);
nor UO_3925 (O_3925,N_49624,N_47460);
or UO_3926 (O_3926,N_45806,N_48957);
or UO_3927 (O_3927,N_49727,N_47821);
xor UO_3928 (O_3928,N_48494,N_47495);
nand UO_3929 (O_3929,N_48384,N_47545);
nor UO_3930 (O_3930,N_47682,N_46800);
nand UO_3931 (O_3931,N_47058,N_45208);
and UO_3932 (O_3932,N_46781,N_47862);
or UO_3933 (O_3933,N_49200,N_45543);
or UO_3934 (O_3934,N_46949,N_46470);
or UO_3935 (O_3935,N_45414,N_46324);
nand UO_3936 (O_3936,N_46559,N_49059);
nor UO_3937 (O_3937,N_48552,N_45526);
and UO_3938 (O_3938,N_47424,N_46041);
nor UO_3939 (O_3939,N_47248,N_45108);
and UO_3940 (O_3940,N_47358,N_49061);
and UO_3941 (O_3941,N_48617,N_47838);
or UO_3942 (O_3942,N_47099,N_45932);
and UO_3943 (O_3943,N_45475,N_49690);
or UO_3944 (O_3944,N_46618,N_48725);
nor UO_3945 (O_3945,N_45161,N_45206);
nor UO_3946 (O_3946,N_47915,N_48097);
and UO_3947 (O_3947,N_49106,N_45915);
nand UO_3948 (O_3948,N_49341,N_47159);
nor UO_3949 (O_3949,N_47525,N_49465);
nand UO_3950 (O_3950,N_46481,N_48228);
nor UO_3951 (O_3951,N_46448,N_48592);
nor UO_3952 (O_3952,N_47242,N_45283);
or UO_3953 (O_3953,N_49994,N_48079);
nand UO_3954 (O_3954,N_46677,N_46832);
nor UO_3955 (O_3955,N_46555,N_46569);
and UO_3956 (O_3956,N_49520,N_47012);
nand UO_3957 (O_3957,N_48694,N_47518);
nand UO_3958 (O_3958,N_49020,N_46319);
and UO_3959 (O_3959,N_49307,N_45087);
nor UO_3960 (O_3960,N_48853,N_45301);
xor UO_3961 (O_3961,N_48889,N_48929);
nor UO_3962 (O_3962,N_48363,N_45258);
and UO_3963 (O_3963,N_47651,N_48850);
or UO_3964 (O_3964,N_46778,N_48356);
xnor UO_3965 (O_3965,N_47886,N_48264);
xor UO_3966 (O_3966,N_48738,N_49427);
or UO_3967 (O_3967,N_46047,N_47649);
nor UO_3968 (O_3968,N_49088,N_45543);
or UO_3969 (O_3969,N_47718,N_46989);
or UO_3970 (O_3970,N_47115,N_49547);
nand UO_3971 (O_3971,N_47428,N_46482);
nor UO_3972 (O_3972,N_45979,N_45375);
or UO_3973 (O_3973,N_49833,N_49499);
nand UO_3974 (O_3974,N_49561,N_45126);
nor UO_3975 (O_3975,N_46681,N_46923);
xnor UO_3976 (O_3976,N_45750,N_45765);
xnor UO_3977 (O_3977,N_48710,N_48277);
nor UO_3978 (O_3978,N_47951,N_45023);
nor UO_3979 (O_3979,N_48542,N_48945);
or UO_3980 (O_3980,N_45991,N_45168);
nor UO_3981 (O_3981,N_46730,N_49160);
or UO_3982 (O_3982,N_49498,N_48439);
nor UO_3983 (O_3983,N_49252,N_46999);
or UO_3984 (O_3984,N_48197,N_49223);
or UO_3985 (O_3985,N_46942,N_49992);
and UO_3986 (O_3986,N_46757,N_45014);
xor UO_3987 (O_3987,N_49654,N_47596);
nor UO_3988 (O_3988,N_46114,N_49220);
and UO_3989 (O_3989,N_46010,N_47750);
nor UO_3990 (O_3990,N_49550,N_49887);
nand UO_3991 (O_3991,N_47292,N_46644);
nand UO_3992 (O_3992,N_49747,N_47574);
or UO_3993 (O_3993,N_48203,N_47668);
or UO_3994 (O_3994,N_45254,N_48686);
nand UO_3995 (O_3995,N_48354,N_48996);
and UO_3996 (O_3996,N_48491,N_46460);
nor UO_3997 (O_3997,N_47762,N_47788);
xnor UO_3998 (O_3998,N_48411,N_49450);
nor UO_3999 (O_3999,N_49282,N_45784);
and UO_4000 (O_4000,N_45629,N_49128);
or UO_4001 (O_4001,N_45005,N_45542);
xor UO_4002 (O_4002,N_46857,N_47356);
nand UO_4003 (O_4003,N_45881,N_47990);
xor UO_4004 (O_4004,N_49311,N_48390);
nand UO_4005 (O_4005,N_45948,N_47167);
and UO_4006 (O_4006,N_45655,N_47617);
or UO_4007 (O_4007,N_47236,N_45170);
nor UO_4008 (O_4008,N_46726,N_48905);
or UO_4009 (O_4009,N_47758,N_47673);
nand UO_4010 (O_4010,N_46676,N_47909);
and UO_4011 (O_4011,N_47602,N_46462);
nand UO_4012 (O_4012,N_49054,N_49093);
or UO_4013 (O_4013,N_47760,N_45034);
and UO_4014 (O_4014,N_48539,N_45435);
and UO_4015 (O_4015,N_45688,N_47411);
nor UO_4016 (O_4016,N_47028,N_47135);
and UO_4017 (O_4017,N_49425,N_45731);
and UO_4018 (O_4018,N_49362,N_45582);
or UO_4019 (O_4019,N_49342,N_45131);
and UO_4020 (O_4020,N_45304,N_48778);
or UO_4021 (O_4021,N_45995,N_47111);
or UO_4022 (O_4022,N_46512,N_45809);
or UO_4023 (O_4023,N_46859,N_47329);
and UO_4024 (O_4024,N_48299,N_49328);
nor UO_4025 (O_4025,N_45892,N_45789);
nor UO_4026 (O_4026,N_47482,N_47526);
nor UO_4027 (O_4027,N_46254,N_46116);
xor UO_4028 (O_4028,N_46339,N_49370);
and UO_4029 (O_4029,N_47718,N_49978);
or UO_4030 (O_4030,N_46597,N_45909);
nand UO_4031 (O_4031,N_47450,N_47710);
nor UO_4032 (O_4032,N_48239,N_47590);
and UO_4033 (O_4033,N_46102,N_49478);
nand UO_4034 (O_4034,N_47232,N_49763);
nand UO_4035 (O_4035,N_49137,N_46440);
nand UO_4036 (O_4036,N_48484,N_48304);
nor UO_4037 (O_4037,N_47473,N_46154);
or UO_4038 (O_4038,N_45267,N_46459);
nand UO_4039 (O_4039,N_46213,N_45456);
nand UO_4040 (O_4040,N_49470,N_48543);
or UO_4041 (O_4041,N_49472,N_48140);
nand UO_4042 (O_4042,N_48601,N_45653);
and UO_4043 (O_4043,N_49667,N_47157);
nor UO_4044 (O_4044,N_46321,N_46284);
nand UO_4045 (O_4045,N_45550,N_47060);
nor UO_4046 (O_4046,N_48429,N_48944);
nand UO_4047 (O_4047,N_45795,N_45333);
and UO_4048 (O_4048,N_48263,N_46411);
and UO_4049 (O_4049,N_49297,N_49851);
or UO_4050 (O_4050,N_45822,N_45292);
nand UO_4051 (O_4051,N_47699,N_46059);
xor UO_4052 (O_4052,N_45424,N_47922);
or UO_4053 (O_4053,N_45117,N_47307);
nor UO_4054 (O_4054,N_46617,N_47304);
and UO_4055 (O_4055,N_47242,N_47975);
nand UO_4056 (O_4056,N_45984,N_47041);
nor UO_4057 (O_4057,N_48337,N_48702);
nor UO_4058 (O_4058,N_49880,N_45421);
nor UO_4059 (O_4059,N_48902,N_49966);
nand UO_4060 (O_4060,N_49987,N_45989);
nand UO_4061 (O_4061,N_46913,N_48581);
and UO_4062 (O_4062,N_45526,N_47861);
nor UO_4063 (O_4063,N_45758,N_46876);
or UO_4064 (O_4064,N_47226,N_45234);
nor UO_4065 (O_4065,N_48278,N_45887);
nand UO_4066 (O_4066,N_47982,N_49991);
nor UO_4067 (O_4067,N_46205,N_46435);
nand UO_4068 (O_4068,N_46572,N_45174);
nor UO_4069 (O_4069,N_46466,N_48598);
or UO_4070 (O_4070,N_49643,N_47820);
nor UO_4071 (O_4071,N_45804,N_45618);
and UO_4072 (O_4072,N_48861,N_48645);
or UO_4073 (O_4073,N_45398,N_46746);
and UO_4074 (O_4074,N_45685,N_49249);
and UO_4075 (O_4075,N_47371,N_48322);
nand UO_4076 (O_4076,N_47282,N_48793);
nand UO_4077 (O_4077,N_48509,N_48042);
nand UO_4078 (O_4078,N_49457,N_48770);
and UO_4079 (O_4079,N_46429,N_48213);
nor UO_4080 (O_4080,N_46724,N_48684);
nand UO_4081 (O_4081,N_49233,N_48255);
and UO_4082 (O_4082,N_49358,N_48935);
nand UO_4083 (O_4083,N_46236,N_49356);
and UO_4084 (O_4084,N_45085,N_49172);
nor UO_4085 (O_4085,N_47109,N_49447);
or UO_4086 (O_4086,N_45912,N_48819);
or UO_4087 (O_4087,N_49074,N_47970);
nand UO_4088 (O_4088,N_46887,N_45901);
nand UO_4089 (O_4089,N_45229,N_45088);
nand UO_4090 (O_4090,N_48833,N_45218);
or UO_4091 (O_4091,N_45461,N_47177);
nand UO_4092 (O_4092,N_48932,N_49420);
xnor UO_4093 (O_4093,N_45364,N_49209);
nand UO_4094 (O_4094,N_46286,N_45418);
xor UO_4095 (O_4095,N_49374,N_46456);
nand UO_4096 (O_4096,N_45185,N_45354);
nor UO_4097 (O_4097,N_46877,N_47167);
or UO_4098 (O_4098,N_48361,N_48473);
nand UO_4099 (O_4099,N_46850,N_48838);
or UO_4100 (O_4100,N_46842,N_46650);
nor UO_4101 (O_4101,N_47434,N_45046);
or UO_4102 (O_4102,N_46496,N_45683);
nor UO_4103 (O_4103,N_45326,N_46360);
or UO_4104 (O_4104,N_48600,N_48809);
and UO_4105 (O_4105,N_49179,N_46067);
or UO_4106 (O_4106,N_45504,N_48757);
or UO_4107 (O_4107,N_45548,N_49496);
and UO_4108 (O_4108,N_49824,N_46467);
nand UO_4109 (O_4109,N_48662,N_48392);
nand UO_4110 (O_4110,N_46208,N_48712);
xor UO_4111 (O_4111,N_46526,N_47646);
nor UO_4112 (O_4112,N_45137,N_48288);
nand UO_4113 (O_4113,N_46093,N_47707);
xor UO_4114 (O_4114,N_47579,N_47320);
nor UO_4115 (O_4115,N_48677,N_47655);
nor UO_4116 (O_4116,N_48551,N_46321);
or UO_4117 (O_4117,N_45022,N_45029);
xor UO_4118 (O_4118,N_45352,N_45328);
nand UO_4119 (O_4119,N_45602,N_48699);
nand UO_4120 (O_4120,N_47399,N_48296);
nor UO_4121 (O_4121,N_46568,N_45799);
nand UO_4122 (O_4122,N_48406,N_46869);
nand UO_4123 (O_4123,N_45122,N_48364);
or UO_4124 (O_4124,N_49546,N_49666);
nand UO_4125 (O_4125,N_47664,N_49280);
nand UO_4126 (O_4126,N_46933,N_45060);
and UO_4127 (O_4127,N_49414,N_48934);
nor UO_4128 (O_4128,N_45699,N_48025);
nand UO_4129 (O_4129,N_48555,N_46120);
nand UO_4130 (O_4130,N_45411,N_49285);
and UO_4131 (O_4131,N_48466,N_48659);
xor UO_4132 (O_4132,N_49112,N_48812);
xor UO_4133 (O_4133,N_45629,N_48943);
or UO_4134 (O_4134,N_46770,N_45262);
nor UO_4135 (O_4135,N_47889,N_46065);
and UO_4136 (O_4136,N_45508,N_48762);
nor UO_4137 (O_4137,N_48324,N_48978);
xnor UO_4138 (O_4138,N_45254,N_48235);
or UO_4139 (O_4139,N_46388,N_47445);
nand UO_4140 (O_4140,N_46051,N_49918);
nor UO_4141 (O_4141,N_46104,N_47500);
nor UO_4142 (O_4142,N_48304,N_45998);
nor UO_4143 (O_4143,N_47664,N_49370);
and UO_4144 (O_4144,N_46122,N_49508);
nand UO_4145 (O_4145,N_46400,N_49488);
xnor UO_4146 (O_4146,N_47412,N_47852);
or UO_4147 (O_4147,N_45081,N_48286);
nand UO_4148 (O_4148,N_49962,N_45070);
nand UO_4149 (O_4149,N_47234,N_46798);
nor UO_4150 (O_4150,N_45723,N_48189);
nand UO_4151 (O_4151,N_49156,N_46168);
nor UO_4152 (O_4152,N_48697,N_49706);
nor UO_4153 (O_4153,N_49903,N_48186);
and UO_4154 (O_4154,N_49360,N_46276);
nor UO_4155 (O_4155,N_49143,N_46801);
nand UO_4156 (O_4156,N_45160,N_48703);
and UO_4157 (O_4157,N_49506,N_48924);
or UO_4158 (O_4158,N_47717,N_48829);
nor UO_4159 (O_4159,N_45532,N_49388);
nor UO_4160 (O_4160,N_49619,N_49959);
and UO_4161 (O_4161,N_46062,N_49378);
nor UO_4162 (O_4162,N_48852,N_46126);
or UO_4163 (O_4163,N_45717,N_45405);
and UO_4164 (O_4164,N_48289,N_45916);
and UO_4165 (O_4165,N_49049,N_45151);
and UO_4166 (O_4166,N_48532,N_45743);
xnor UO_4167 (O_4167,N_48503,N_47395);
nor UO_4168 (O_4168,N_48123,N_48972);
and UO_4169 (O_4169,N_45222,N_48391);
and UO_4170 (O_4170,N_46504,N_46910);
nand UO_4171 (O_4171,N_46777,N_47984);
xnor UO_4172 (O_4172,N_48250,N_49202);
or UO_4173 (O_4173,N_49066,N_48625);
nand UO_4174 (O_4174,N_46856,N_47129);
nor UO_4175 (O_4175,N_48494,N_49895);
nand UO_4176 (O_4176,N_48808,N_47719);
nand UO_4177 (O_4177,N_45154,N_46052);
nand UO_4178 (O_4178,N_45791,N_49812);
nand UO_4179 (O_4179,N_49339,N_45544);
or UO_4180 (O_4180,N_47023,N_45358);
or UO_4181 (O_4181,N_48878,N_47694);
nand UO_4182 (O_4182,N_47824,N_47617);
nor UO_4183 (O_4183,N_45619,N_46769);
or UO_4184 (O_4184,N_47148,N_46674);
and UO_4185 (O_4185,N_49878,N_49726);
and UO_4186 (O_4186,N_45569,N_49320);
nand UO_4187 (O_4187,N_46639,N_45784);
nor UO_4188 (O_4188,N_45556,N_48018);
nand UO_4189 (O_4189,N_49184,N_48051);
or UO_4190 (O_4190,N_49334,N_46832);
or UO_4191 (O_4191,N_47739,N_46758);
and UO_4192 (O_4192,N_47781,N_45312);
nand UO_4193 (O_4193,N_46566,N_46641);
xor UO_4194 (O_4194,N_48872,N_48873);
nor UO_4195 (O_4195,N_46111,N_48335);
and UO_4196 (O_4196,N_47019,N_46770);
xnor UO_4197 (O_4197,N_46052,N_47981);
nand UO_4198 (O_4198,N_49934,N_45361);
nand UO_4199 (O_4199,N_46251,N_47988);
and UO_4200 (O_4200,N_49627,N_46483);
nand UO_4201 (O_4201,N_45512,N_46969);
or UO_4202 (O_4202,N_49518,N_46846);
nand UO_4203 (O_4203,N_46012,N_49867);
or UO_4204 (O_4204,N_46745,N_47907);
nand UO_4205 (O_4205,N_49263,N_49109);
and UO_4206 (O_4206,N_48723,N_46538);
and UO_4207 (O_4207,N_47615,N_45780);
or UO_4208 (O_4208,N_49718,N_47208);
or UO_4209 (O_4209,N_45841,N_48569);
or UO_4210 (O_4210,N_46343,N_46225);
nand UO_4211 (O_4211,N_47537,N_49769);
nor UO_4212 (O_4212,N_47786,N_47627);
and UO_4213 (O_4213,N_48029,N_46494);
nand UO_4214 (O_4214,N_46550,N_45847);
or UO_4215 (O_4215,N_45719,N_46837);
xnor UO_4216 (O_4216,N_47853,N_47518);
xnor UO_4217 (O_4217,N_49237,N_45213);
nand UO_4218 (O_4218,N_46986,N_47197);
or UO_4219 (O_4219,N_46892,N_46338);
and UO_4220 (O_4220,N_46182,N_47373);
nand UO_4221 (O_4221,N_49716,N_49441);
nor UO_4222 (O_4222,N_46319,N_48968);
xnor UO_4223 (O_4223,N_48093,N_49595);
or UO_4224 (O_4224,N_48329,N_48513);
xnor UO_4225 (O_4225,N_47476,N_48749);
nor UO_4226 (O_4226,N_46837,N_49448);
nand UO_4227 (O_4227,N_48723,N_49130);
xor UO_4228 (O_4228,N_46501,N_47375);
nor UO_4229 (O_4229,N_45151,N_47853);
or UO_4230 (O_4230,N_49911,N_49604);
and UO_4231 (O_4231,N_46736,N_48230);
nand UO_4232 (O_4232,N_47774,N_48855);
nor UO_4233 (O_4233,N_45095,N_48019);
or UO_4234 (O_4234,N_49923,N_48756);
nor UO_4235 (O_4235,N_45533,N_47005);
and UO_4236 (O_4236,N_47060,N_45075);
xor UO_4237 (O_4237,N_48765,N_46783);
nor UO_4238 (O_4238,N_46266,N_47544);
nand UO_4239 (O_4239,N_48618,N_46725);
xnor UO_4240 (O_4240,N_47178,N_49138);
or UO_4241 (O_4241,N_49943,N_49699);
nand UO_4242 (O_4242,N_45544,N_48329);
and UO_4243 (O_4243,N_49584,N_49517);
nand UO_4244 (O_4244,N_48709,N_48466);
and UO_4245 (O_4245,N_45385,N_47979);
and UO_4246 (O_4246,N_48828,N_45188);
and UO_4247 (O_4247,N_48190,N_48966);
and UO_4248 (O_4248,N_49712,N_49318);
and UO_4249 (O_4249,N_45760,N_49039);
and UO_4250 (O_4250,N_45753,N_47354);
and UO_4251 (O_4251,N_46151,N_49240);
and UO_4252 (O_4252,N_46517,N_49381);
nand UO_4253 (O_4253,N_46903,N_49665);
or UO_4254 (O_4254,N_48389,N_46181);
nand UO_4255 (O_4255,N_45958,N_45678);
nand UO_4256 (O_4256,N_45274,N_45618);
nor UO_4257 (O_4257,N_46177,N_47455);
and UO_4258 (O_4258,N_49214,N_45409);
or UO_4259 (O_4259,N_45561,N_46516);
and UO_4260 (O_4260,N_45667,N_45459);
nor UO_4261 (O_4261,N_46692,N_45249);
nand UO_4262 (O_4262,N_46345,N_49968);
xor UO_4263 (O_4263,N_47522,N_48682);
or UO_4264 (O_4264,N_48904,N_45927);
xor UO_4265 (O_4265,N_47398,N_46630);
nor UO_4266 (O_4266,N_47201,N_48472);
nand UO_4267 (O_4267,N_46090,N_46626);
nand UO_4268 (O_4268,N_47978,N_46500);
nand UO_4269 (O_4269,N_45707,N_48412);
or UO_4270 (O_4270,N_49371,N_48051);
nand UO_4271 (O_4271,N_46477,N_49452);
or UO_4272 (O_4272,N_48727,N_49083);
and UO_4273 (O_4273,N_45677,N_47491);
or UO_4274 (O_4274,N_48057,N_48816);
nor UO_4275 (O_4275,N_45643,N_46182);
xnor UO_4276 (O_4276,N_46947,N_49352);
nor UO_4277 (O_4277,N_47929,N_47175);
and UO_4278 (O_4278,N_46320,N_48445);
and UO_4279 (O_4279,N_45395,N_47969);
and UO_4280 (O_4280,N_45447,N_47119);
nor UO_4281 (O_4281,N_49875,N_47062);
nor UO_4282 (O_4282,N_49885,N_49926);
or UO_4283 (O_4283,N_47188,N_49121);
or UO_4284 (O_4284,N_49595,N_49955);
nand UO_4285 (O_4285,N_45091,N_49015);
xor UO_4286 (O_4286,N_47116,N_48818);
and UO_4287 (O_4287,N_49316,N_49456);
and UO_4288 (O_4288,N_46744,N_47636);
or UO_4289 (O_4289,N_47650,N_49676);
and UO_4290 (O_4290,N_45054,N_45596);
and UO_4291 (O_4291,N_48184,N_49639);
and UO_4292 (O_4292,N_49153,N_45140);
or UO_4293 (O_4293,N_45831,N_46927);
and UO_4294 (O_4294,N_46526,N_47687);
xnor UO_4295 (O_4295,N_47679,N_47263);
or UO_4296 (O_4296,N_48967,N_48528);
nor UO_4297 (O_4297,N_45510,N_48806);
nor UO_4298 (O_4298,N_49100,N_47043);
nand UO_4299 (O_4299,N_46684,N_46712);
and UO_4300 (O_4300,N_45639,N_49726);
nand UO_4301 (O_4301,N_47460,N_45271);
or UO_4302 (O_4302,N_45685,N_45295);
and UO_4303 (O_4303,N_49567,N_48089);
nor UO_4304 (O_4304,N_46699,N_46782);
or UO_4305 (O_4305,N_47760,N_49847);
nor UO_4306 (O_4306,N_48908,N_46457);
and UO_4307 (O_4307,N_46402,N_49698);
or UO_4308 (O_4308,N_46527,N_49650);
and UO_4309 (O_4309,N_49757,N_47878);
or UO_4310 (O_4310,N_45315,N_49968);
and UO_4311 (O_4311,N_45068,N_47422);
xor UO_4312 (O_4312,N_46622,N_49139);
nor UO_4313 (O_4313,N_46364,N_48544);
xnor UO_4314 (O_4314,N_49811,N_47991);
xor UO_4315 (O_4315,N_47395,N_46957);
or UO_4316 (O_4316,N_47896,N_46995);
or UO_4317 (O_4317,N_45557,N_48120);
nand UO_4318 (O_4318,N_47059,N_45194);
or UO_4319 (O_4319,N_47411,N_48224);
or UO_4320 (O_4320,N_49762,N_49295);
xor UO_4321 (O_4321,N_45019,N_46186);
nand UO_4322 (O_4322,N_49732,N_48112);
nand UO_4323 (O_4323,N_47301,N_49746);
and UO_4324 (O_4324,N_45608,N_49569);
or UO_4325 (O_4325,N_45769,N_49588);
nor UO_4326 (O_4326,N_45894,N_47323);
nand UO_4327 (O_4327,N_48191,N_48657);
nor UO_4328 (O_4328,N_46326,N_46941);
nor UO_4329 (O_4329,N_46593,N_49924);
nand UO_4330 (O_4330,N_46766,N_47954);
xnor UO_4331 (O_4331,N_46986,N_46002);
nand UO_4332 (O_4332,N_45401,N_46833);
nor UO_4333 (O_4333,N_48436,N_45103);
nor UO_4334 (O_4334,N_46353,N_48888);
and UO_4335 (O_4335,N_48393,N_49233);
xor UO_4336 (O_4336,N_46290,N_45676);
nand UO_4337 (O_4337,N_48985,N_47769);
and UO_4338 (O_4338,N_47426,N_45686);
xor UO_4339 (O_4339,N_48483,N_46016);
nand UO_4340 (O_4340,N_49117,N_49397);
or UO_4341 (O_4341,N_45735,N_47924);
nand UO_4342 (O_4342,N_45409,N_48438);
nor UO_4343 (O_4343,N_48323,N_45319);
and UO_4344 (O_4344,N_49337,N_46971);
or UO_4345 (O_4345,N_45298,N_47276);
or UO_4346 (O_4346,N_49982,N_45790);
nand UO_4347 (O_4347,N_49591,N_49907);
and UO_4348 (O_4348,N_46672,N_47215);
nand UO_4349 (O_4349,N_46923,N_47392);
nand UO_4350 (O_4350,N_47271,N_45021);
nor UO_4351 (O_4351,N_47809,N_46912);
nor UO_4352 (O_4352,N_49594,N_46460);
nand UO_4353 (O_4353,N_49942,N_48770);
or UO_4354 (O_4354,N_46068,N_46826);
nand UO_4355 (O_4355,N_49657,N_46235);
and UO_4356 (O_4356,N_45274,N_46917);
and UO_4357 (O_4357,N_46628,N_45554);
nor UO_4358 (O_4358,N_46214,N_47520);
and UO_4359 (O_4359,N_48175,N_49939);
or UO_4360 (O_4360,N_49699,N_46795);
nand UO_4361 (O_4361,N_45500,N_46763);
xor UO_4362 (O_4362,N_47910,N_48728);
nand UO_4363 (O_4363,N_48928,N_47726);
or UO_4364 (O_4364,N_45723,N_46146);
and UO_4365 (O_4365,N_45891,N_47794);
nand UO_4366 (O_4366,N_45523,N_47202);
nor UO_4367 (O_4367,N_46339,N_48058);
nand UO_4368 (O_4368,N_47886,N_48348);
and UO_4369 (O_4369,N_47947,N_47687);
and UO_4370 (O_4370,N_45340,N_47734);
nand UO_4371 (O_4371,N_45210,N_48529);
and UO_4372 (O_4372,N_47790,N_48392);
and UO_4373 (O_4373,N_49669,N_46353);
nor UO_4374 (O_4374,N_46764,N_49438);
nand UO_4375 (O_4375,N_45177,N_46428);
nor UO_4376 (O_4376,N_45766,N_48234);
xor UO_4377 (O_4377,N_48464,N_47825);
xnor UO_4378 (O_4378,N_46627,N_46331);
and UO_4379 (O_4379,N_48252,N_47333);
nand UO_4380 (O_4380,N_45285,N_48396);
xor UO_4381 (O_4381,N_49386,N_47323);
or UO_4382 (O_4382,N_49715,N_46025);
nand UO_4383 (O_4383,N_46798,N_47707);
nand UO_4384 (O_4384,N_46247,N_49173);
nand UO_4385 (O_4385,N_45233,N_49590);
and UO_4386 (O_4386,N_48466,N_45874);
or UO_4387 (O_4387,N_45064,N_47569);
or UO_4388 (O_4388,N_46968,N_45456);
xnor UO_4389 (O_4389,N_47659,N_45570);
or UO_4390 (O_4390,N_47411,N_48849);
and UO_4391 (O_4391,N_45661,N_49186);
nand UO_4392 (O_4392,N_48636,N_46742);
or UO_4393 (O_4393,N_46267,N_48875);
nand UO_4394 (O_4394,N_48594,N_49654);
nand UO_4395 (O_4395,N_46665,N_48507);
nand UO_4396 (O_4396,N_49858,N_49635);
and UO_4397 (O_4397,N_46593,N_47035);
xnor UO_4398 (O_4398,N_46050,N_48335);
and UO_4399 (O_4399,N_48527,N_46040);
nor UO_4400 (O_4400,N_45748,N_46642);
nand UO_4401 (O_4401,N_47701,N_48033);
or UO_4402 (O_4402,N_46759,N_47481);
or UO_4403 (O_4403,N_45630,N_45666);
nand UO_4404 (O_4404,N_46882,N_45622);
nor UO_4405 (O_4405,N_45476,N_46638);
nor UO_4406 (O_4406,N_46942,N_48995);
or UO_4407 (O_4407,N_47560,N_49682);
and UO_4408 (O_4408,N_48670,N_49523);
nor UO_4409 (O_4409,N_47976,N_48595);
and UO_4410 (O_4410,N_49896,N_46174);
or UO_4411 (O_4411,N_46295,N_47675);
nand UO_4412 (O_4412,N_47059,N_49051);
or UO_4413 (O_4413,N_48824,N_47680);
and UO_4414 (O_4414,N_46079,N_45989);
nor UO_4415 (O_4415,N_49666,N_47113);
nor UO_4416 (O_4416,N_45222,N_48285);
or UO_4417 (O_4417,N_48621,N_47212);
nor UO_4418 (O_4418,N_47469,N_45194);
nor UO_4419 (O_4419,N_45096,N_49619);
nand UO_4420 (O_4420,N_46680,N_45128);
nor UO_4421 (O_4421,N_49548,N_46810);
xor UO_4422 (O_4422,N_46674,N_46042);
nand UO_4423 (O_4423,N_45937,N_45625);
and UO_4424 (O_4424,N_46187,N_47745);
and UO_4425 (O_4425,N_47594,N_47639);
nor UO_4426 (O_4426,N_49029,N_47539);
nor UO_4427 (O_4427,N_46331,N_47029);
or UO_4428 (O_4428,N_45207,N_46099);
nand UO_4429 (O_4429,N_49201,N_45991);
nor UO_4430 (O_4430,N_47088,N_49391);
xnor UO_4431 (O_4431,N_46258,N_46640);
nor UO_4432 (O_4432,N_49236,N_46902);
nand UO_4433 (O_4433,N_49286,N_45819);
nor UO_4434 (O_4434,N_46070,N_47414);
nand UO_4435 (O_4435,N_46016,N_48003);
or UO_4436 (O_4436,N_49821,N_45345);
or UO_4437 (O_4437,N_49936,N_48647);
nor UO_4438 (O_4438,N_49035,N_45473);
nand UO_4439 (O_4439,N_45185,N_45205);
xnor UO_4440 (O_4440,N_45058,N_47361);
nor UO_4441 (O_4441,N_48803,N_45977);
nor UO_4442 (O_4442,N_49209,N_45660);
nor UO_4443 (O_4443,N_48941,N_46025);
and UO_4444 (O_4444,N_49509,N_46658);
or UO_4445 (O_4445,N_46814,N_48853);
nand UO_4446 (O_4446,N_45647,N_46724);
and UO_4447 (O_4447,N_45269,N_47292);
nor UO_4448 (O_4448,N_49464,N_49465);
and UO_4449 (O_4449,N_48262,N_46014);
and UO_4450 (O_4450,N_48643,N_46530);
nand UO_4451 (O_4451,N_46154,N_48105);
and UO_4452 (O_4452,N_49509,N_47234);
and UO_4453 (O_4453,N_48377,N_45800);
or UO_4454 (O_4454,N_47093,N_46683);
nor UO_4455 (O_4455,N_45701,N_47212);
or UO_4456 (O_4456,N_46404,N_49440);
xor UO_4457 (O_4457,N_48092,N_47114);
xor UO_4458 (O_4458,N_47492,N_48761);
nor UO_4459 (O_4459,N_49407,N_46262);
nor UO_4460 (O_4460,N_49153,N_45953);
xnor UO_4461 (O_4461,N_49074,N_47194);
and UO_4462 (O_4462,N_46519,N_46969);
and UO_4463 (O_4463,N_47256,N_46895);
and UO_4464 (O_4464,N_45814,N_49004);
or UO_4465 (O_4465,N_47361,N_49215);
or UO_4466 (O_4466,N_46647,N_49527);
nand UO_4467 (O_4467,N_49032,N_47333);
or UO_4468 (O_4468,N_45134,N_46492);
nor UO_4469 (O_4469,N_47156,N_46097);
xor UO_4470 (O_4470,N_46279,N_45632);
nor UO_4471 (O_4471,N_48480,N_48709);
or UO_4472 (O_4472,N_47664,N_48922);
nand UO_4473 (O_4473,N_46134,N_48076);
xnor UO_4474 (O_4474,N_49230,N_47355);
or UO_4475 (O_4475,N_46553,N_46181);
nand UO_4476 (O_4476,N_47469,N_47902);
or UO_4477 (O_4477,N_49614,N_48226);
and UO_4478 (O_4478,N_45166,N_48669);
nor UO_4479 (O_4479,N_47558,N_47061);
nor UO_4480 (O_4480,N_46978,N_47611);
xnor UO_4481 (O_4481,N_46879,N_45057);
nand UO_4482 (O_4482,N_45620,N_49845);
xnor UO_4483 (O_4483,N_49209,N_45994);
nor UO_4484 (O_4484,N_47720,N_46705);
or UO_4485 (O_4485,N_46624,N_47246);
nor UO_4486 (O_4486,N_46017,N_49491);
and UO_4487 (O_4487,N_48954,N_46884);
nor UO_4488 (O_4488,N_49263,N_49296);
and UO_4489 (O_4489,N_49756,N_45167);
or UO_4490 (O_4490,N_49778,N_47251);
nand UO_4491 (O_4491,N_45858,N_49350);
nor UO_4492 (O_4492,N_46362,N_48264);
nor UO_4493 (O_4493,N_49939,N_46511);
xnor UO_4494 (O_4494,N_47036,N_48842);
xnor UO_4495 (O_4495,N_46423,N_47749);
nand UO_4496 (O_4496,N_49904,N_46691);
nand UO_4497 (O_4497,N_46926,N_48848);
or UO_4498 (O_4498,N_47363,N_48519);
xor UO_4499 (O_4499,N_45524,N_45424);
and UO_4500 (O_4500,N_46400,N_46729);
and UO_4501 (O_4501,N_48359,N_47901);
or UO_4502 (O_4502,N_45572,N_46622);
nand UO_4503 (O_4503,N_48828,N_47883);
nor UO_4504 (O_4504,N_47151,N_46422);
and UO_4505 (O_4505,N_48508,N_46753);
or UO_4506 (O_4506,N_46611,N_48883);
and UO_4507 (O_4507,N_45993,N_45927);
nor UO_4508 (O_4508,N_45844,N_46972);
or UO_4509 (O_4509,N_46916,N_45293);
or UO_4510 (O_4510,N_47639,N_45020);
nor UO_4511 (O_4511,N_47549,N_47715);
nor UO_4512 (O_4512,N_46553,N_46572);
nand UO_4513 (O_4513,N_49481,N_46777);
nand UO_4514 (O_4514,N_46765,N_48106);
xor UO_4515 (O_4515,N_45106,N_49313);
and UO_4516 (O_4516,N_47914,N_48392);
and UO_4517 (O_4517,N_47885,N_48006);
nor UO_4518 (O_4518,N_49764,N_45258);
or UO_4519 (O_4519,N_48738,N_49805);
and UO_4520 (O_4520,N_45117,N_46634);
nor UO_4521 (O_4521,N_47052,N_46434);
nor UO_4522 (O_4522,N_45103,N_49548);
or UO_4523 (O_4523,N_49654,N_48631);
or UO_4524 (O_4524,N_47746,N_47578);
or UO_4525 (O_4525,N_49733,N_45515);
nand UO_4526 (O_4526,N_48504,N_45396);
and UO_4527 (O_4527,N_49636,N_48197);
or UO_4528 (O_4528,N_49478,N_48326);
xnor UO_4529 (O_4529,N_46902,N_45423);
nand UO_4530 (O_4530,N_48389,N_45152);
nand UO_4531 (O_4531,N_45010,N_46277);
nor UO_4532 (O_4532,N_46046,N_45342);
nor UO_4533 (O_4533,N_46684,N_47109);
and UO_4534 (O_4534,N_47526,N_46044);
nand UO_4535 (O_4535,N_49477,N_45317);
nor UO_4536 (O_4536,N_48502,N_46486);
and UO_4537 (O_4537,N_48716,N_46085);
or UO_4538 (O_4538,N_49701,N_47202);
nand UO_4539 (O_4539,N_48774,N_49067);
nor UO_4540 (O_4540,N_49384,N_47151);
xor UO_4541 (O_4541,N_47689,N_46823);
nor UO_4542 (O_4542,N_47641,N_48558);
or UO_4543 (O_4543,N_46957,N_45582);
nand UO_4544 (O_4544,N_48115,N_45253);
and UO_4545 (O_4545,N_49162,N_47274);
nand UO_4546 (O_4546,N_46875,N_49045);
nor UO_4547 (O_4547,N_45894,N_47747);
nand UO_4548 (O_4548,N_45259,N_48218);
or UO_4549 (O_4549,N_49200,N_45746);
nor UO_4550 (O_4550,N_45218,N_49280);
or UO_4551 (O_4551,N_48133,N_49079);
nand UO_4552 (O_4552,N_46494,N_49645);
nor UO_4553 (O_4553,N_48309,N_46615);
xor UO_4554 (O_4554,N_48494,N_49133);
or UO_4555 (O_4555,N_47570,N_45382);
or UO_4556 (O_4556,N_48769,N_47745);
nand UO_4557 (O_4557,N_46602,N_45368);
nand UO_4558 (O_4558,N_47091,N_49598);
and UO_4559 (O_4559,N_48842,N_49958);
and UO_4560 (O_4560,N_45842,N_49607);
or UO_4561 (O_4561,N_49761,N_49507);
or UO_4562 (O_4562,N_45481,N_46637);
nand UO_4563 (O_4563,N_49919,N_47991);
nand UO_4564 (O_4564,N_45796,N_48469);
or UO_4565 (O_4565,N_48794,N_48904);
xnor UO_4566 (O_4566,N_49678,N_47838);
and UO_4567 (O_4567,N_48276,N_47531);
and UO_4568 (O_4568,N_46512,N_45402);
nor UO_4569 (O_4569,N_47058,N_47324);
xnor UO_4570 (O_4570,N_49969,N_49526);
xnor UO_4571 (O_4571,N_48323,N_49117);
and UO_4572 (O_4572,N_48975,N_47954);
nand UO_4573 (O_4573,N_49139,N_47837);
nand UO_4574 (O_4574,N_46643,N_47857);
nand UO_4575 (O_4575,N_49517,N_48743);
or UO_4576 (O_4576,N_47453,N_48824);
nand UO_4577 (O_4577,N_47654,N_47173);
nand UO_4578 (O_4578,N_48120,N_45251);
nand UO_4579 (O_4579,N_45432,N_47749);
nand UO_4580 (O_4580,N_47361,N_45363);
nor UO_4581 (O_4581,N_49155,N_45604);
nor UO_4582 (O_4582,N_45776,N_48308);
and UO_4583 (O_4583,N_49985,N_45245);
nor UO_4584 (O_4584,N_49969,N_48100);
and UO_4585 (O_4585,N_47897,N_46005);
and UO_4586 (O_4586,N_45211,N_45618);
or UO_4587 (O_4587,N_45812,N_49072);
and UO_4588 (O_4588,N_49145,N_45594);
nor UO_4589 (O_4589,N_49999,N_48179);
and UO_4590 (O_4590,N_49187,N_45393);
xnor UO_4591 (O_4591,N_49579,N_45208);
nor UO_4592 (O_4592,N_45613,N_47505);
nand UO_4593 (O_4593,N_47967,N_49012);
and UO_4594 (O_4594,N_48460,N_46200);
nand UO_4595 (O_4595,N_49647,N_46975);
nand UO_4596 (O_4596,N_49869,N_46011);
nor UO_4597 (O_4597,N_45135,N_47573);
and UO_4598 (O_4598,N_48808,N_45798);
nand UO_4599 (O_4599,N_49699,N_47865);
or UO_4600 (O_4600,N_48999,N_48939);
or UO_4601 (O_4601,N_48878,N_49009);
nor UO_4602 (O_4602,N_48712,N_48443);
nor UO_4603 (O_4603,N_48628,N_49510);
or UO_4604 (O_4604,N_45649,N_45871);
nand UO_4605 (O_4605,N_49411,N_45325);
or UO_4606 (O_4606,N_48727,N_46419);
nand UO_4607 (O_4607,N_48962,N_45853);
nor UO_4608 (O_4608,N_48412,N_47810);
and UO_4609 (O_4609,N_45414,N_46914);
nor UO_4610 (O_4610,N_47901,N_48475);
nor UO_4611 (O_4611,N_48085,N_46962);
and UO_4612 (O_4612,N_46503,N_48035);
nand UO_4613 (O_4613,N_45431,N_45851);
nand UO_4614 (O_4614,N_47526,N_49528);
and UO_4615 (O_4615,N_49977,N_47949);
xor UO_4616 (O_4616,N_45857,N_46236);
and UO_4617 (O_4617,N_45323,N_47621);
nand UO_4618 (O_4618,N_48760,N_46588);
nor UO_4619 (O_4619,N_49042,N_48750);
or UO_4620 (O_4620,N_49158,N_47081);
nand UO_4621 (O_4621,N_47823,N_48251);
or UO_4622 (O_4622,N_46584,N_49135);
nand UO_4623 (O_4623,N_45270,N_48651);
nand UO_4624 (O_4624,N_47132,N_46900);
or UO_4625 (O_4625,N_47750,N_49627);
nor UO_4626 (O_4626,N_45344,N_47222);
nor UO_4627 (O_4627,N_45242,N_49162);
nand UO_4628 (O_4628,N_48011,N_47198);
nor UO_4629 (O_4629,N_49722,N_45792);
nor UO_4630 (O_4630,N_45246,N_45166);
xnor UO_4631 (O_4631,N_45723,N_48353);
xor UO_4632 (O_4632,N_46509,N_49467);
and UO_4633 (O_4633,N_47340,N_46740);
or UO_4634 (O_4634,N_45677,N_47878);
xor UO_4635 (O_4635,N_48842,N_49340);
nor UO_4636 (O_4636,N_45449,N_47394);
nor UO_4637 (O_4637,N_46253,N_49164);
nand UO_4638 (O_4638,N_49523,N_49648);
nor UO_4639 (O_4639,N_48315,N_48481);
nand UO_4640 (O_4640,N_49722,N_45888);
nand UO_4641 (O_4641,N_47871,N_48927);
and UO_4642 (O_4642,N_45668,N_48563);
nand UO_4643 (O_4643,N_45687,N_49905);
and UO_4644 (O_4644,N_46286,N_45041);
or UO_4645 (O_4645,N_46798,N_45217);
xor UO_4646 (O_4646,N_48722,N_45918);
xor UO_4647 (O_4647,N_46904,N_48556);
and UO_4648 (O_4648,N_49279,N_48816);
and UO_4649 (O_4649,N_46936,N_47903);
nand UO_4650 (O_4650,N_47837,N_47944);
or UO_4651 (O_4651,N_45059,N_48733);
and UO_4652 (O_4652,N_47974,N_45702);
and UO_4653 (O_4653,N_48719,N_47805);
nand UO_4654 (O_4654,N_45952,N_47478);
or UO_4655 (O_4655,N_47940,N_47666);
or UO_4656 (O_4656,N_46301,N_46177);
and UO_4657 (O_4657,N_47333,N_45368);
and UO_4658 (O_4658,N_48278,N_48993);
or UO_4659 (O_4659,N_47630,N_47040);
xnor UO_4660 (O_4660,N_48881,N_48719);
nor UO_4661 (O_4661,N_46777,N_46035);
nand UO_4662 (O_4662,N_49148,N_46202);
xnor UO_4663 (O_4663,N_46060,N_45577);
or UO_4664 (O_4664,N_49086,N_48856);
or UO_4665 (O_4665,N_46342,N_49164);
or UO_4666 (O_4666,N_49864,N_46474);
nor UO_4667 (O_4667,N_45402,N_45846);
or UO_4668 (O_4668,N_46223,N_46241);
xor UO_4669 (O_4669,N_49762,N_47350);
or UO_4670 (O_4670,N_47066,N_45446);
xnor UO_4671 (O_4671,N_46356,N_45951);
or UO_4672 (O_4672,N_45197,N_46171);
or UO_4673 (O_4673,N_49944,N_48492);
and UO_4674 (O_4674,N_46176,N_47537);
nor UO_4675 (O_4675,N_46255,N_45645);
and UO_4676 (O_4676,N_45858,N_45150);
nor UO_4677 (O_4677,N_46060,N_49885);
and UO_4678 (O_4678,N_47869,N_45213);
and UO_4679 (O_4679,N_47906,N_45444);
nor UO_4680 (O_4680,N_49377,N_45291);
or UO_4681 (O_4681,N_49779,N_49352);
nor UO_4682 (O_4682,N_48045,N_46906);
and UO_4683 (O_4683,N_49039,N_48637);
and UO_4684 (O_4684,N_49312,N_45556);
and UO_4685 (O_4685,N_48420,N_48426);
nand UO_4686 (O_4686,N_49895,N_48267);
nor UO_4687 (O_4687,N_45054,N_48638);
nor UO_4688 (O_4688,N_46144,N_48027);
or UO_4689 (O_4689,N_47245,N_46375);
and UO_4690 (O_4690,N_48153,N_47233);
and UO_4691 (O_4691,N_47966,N_47207);
nand UO_4692 (O_4692,N_47003,N_46287);
and UO_4693 (O_4693,N_49804,N_47802);
or UO_4694 (O_4694,N_48022,N_45858);
nand UO_4695 (O_4695,N_49962,N_49982);
or UO_4696 (O_4696,N_46838,N_49423);
nand UO_4697 (O_4697,N_45834,N_45737);
or UO_4698 (O_4698,N_48682,N_46281);
and UO_4699 (O_4699,N_46187,N_46494);
nand UO_4700 (O_4700,N_48441,N_46532);
or UO_4701 (O_4701,N_45203,N_47671);
nand UO_4702 (O_4702,N_48170,N_47764);
or UO_4703 (O_4703,N_48729,N_47850);
nor UO_4704 (O_4704,N_48660,N_48548);
nor UO_4705 (O_4705,N_45286,N_48775);
nand UO_4706 (O_4706,N_48015,N_47177);
or UO_4707 (O_4707,N_49216,N_49036);
or UO_4708 (O_4708,N_49408,N_46362);
or UO_4709 (O_4709,N_49525,N_48144);
or UO_4710 (O_4710,N_49398,N_46221);
and UO_4711 (O_4711,N_49604,N_49950);
nor UO_4712 (O_4712,N_45728,N_47260);
and UO_4713 (O_4713,N_49300,N_45293);
nand UO_4714 (O_4714,N_46603,N_49419);
xor UO_4715 (O_4715,N_48553,N_49998);
nor UO_4716 (O_4716,N_45854,N_45623);
nor UO_4717 (O_4717,N_47726,N_45932);
nor UO_4718 (O_4718,N_49590,N_49541);
nand UO_4719 (O_4719,N_46124,N_46079);
or UO_4720 (O_4720,N_48125,N_48013);
or UO_4721 (O_4721,N_46062,N_47614);
nor UO_4722 (O_4722,N_45822,N_46329);
nand UO_4723 (O_4723,N_47140,N_47385);
or UO_4724 (O_4724,N_49022,N_47678);
and UO_4725 (O_4725,N_47924,N_47375);
nor UO_4726 (O_4726,N_47561,N_45265);
or UO_4727 (O_4727,N_47890,N_48103);
and UO_4728 (O_4728,N_45206,N_48515);
and UO_4729 (O_4729,N_48379,N_45241);
nor UO_4730 (O_4730,N_46053,N_46763);
and UO_4731 (O_4731,N_48750,N_46624);
or UO_4732 (O_4732,N_49515,N_49926);
nor UO_4733 (O_4733,N_49502,N_48073);
or UO_4734 (O_4734,N_46881,N_45303);
nor UO_4735 (O_4735,N_47341,N_46322);
or UO_4736 (O_4736,N_48287,N_46065);
and UO_4737 (O_4737,N_48288,N_47220);
nand UO_4738 (O_4738,N_48717,N_45346);
or UO_4739 (O_4739,N_48337,N_45376);
or UO_4740 (O_4740,N_48549,N_48985);
and UO_4741 (O_4741,N_47217,N_47476);
and UO_4742 (O_4742,N_49247,N_45621);
nor UO_4743 (O_4743,N_47052,N_46178);
xnor UO_4744 (O_4744,N_48656,N_49977);
nand UO_4745 (O_4745,N_45388,N_47827);
and UO_4746 (O_4746,N_48007,N_46837);
nor UO_4747 (O_4747,N_48449,N_47343);
nor UO_4748 (O_4748,N_49295,N_48895);
nand UO_4749 (O_4749,N_48798,N_46778);
nand UO_4750 (O_4750,N_45398,N_47510);
xnor UO_4751 (O_4751,N_46940,N_49700);
xor UO_4752 (O_4752,N_45751,N_49903);
nand UO_4753 (O_4753,N_47985,N_45999);
xnor UO_4754 (O_4754,N_49275,N_49256);
nor UO_4755 (O_4755,N_46138,N_45243);
or UO_4756 (O_4756,N_48442,N_48839);
or UO_4757 (O_4757,N_49853,N_47366);
and UO_4758 (O_4758,N_49828,N_45318);
nand UO_4759 (O_4759,N_45938,N_49723);
and UO_4760 (O_4760,N_47072,N_49391);
nand UO_4761 (O_4761,N_49569,N_46969);
and UO_4762 (O_4762,N_46117,N_48657);
nand UO_4763 (O_4763,N_49688,N_48985);
nand UO_4764 (O_4764,N_47122,N_45251);
and UO_4765 (O_4765,N_49497,N_45822);
nor UO_4766 (O_4766,N_45737,N_48462);
and UO_4767 (O_4767,N_48190,N_46962);
nor UO_4768 (O_4768,N_48518,N_49079);
nor UO_4769 (O_4769,N_48522,N_47381);
nor UO_4770 (O_4770,N_46733,N_49267);
nand UO_4771 (O_4771,N_48237,N_47046);
or UO_4772 (O_4772,N_45370,N_45314);
nand UO_4773 (O_4773,N_48837,N_46304);
nor UO_4774 (O_4774,N_47313,N_48979);
or UO_4775 (O_4775,N_49528,N_46491);
nor UO_4776 (O_4776,N_46458,N_47114);
or UO_4777 (O_4777,N_46185,N_48526);
or UO_4778 (O_4778,N_48725,N_48227);
nand UO_4779 (O_4779,N_49217,N_45943);
nor UO_4780 (O_4780,N_49273,N_46106);
and UO_4781 (O_4781,N_48079,N_49827);
and UO_4782 (O_4782,N_48891,N_47148);
and UO_4783 (O_4783,N_47905,N_48317);
and UO_4784 (O_4784,N_49036,N_45250);
nand UO_4785 (O_4785,N_49012,N_46508);
nor UO_4786 (O_4786,N_47936,N_47946);
nand UO_4787 (O_4787,N_47660,N_48375);
or UO_4788 (O_4788,N_46117,N_47061);
and UO_4789 (O_4789,N_48549,N_46875);
nor UO_4790 (O_4790,N_49207,N_49410);
nor UO_4791 (O_4791,N_45428,N_47250);
nor UO_4792 (O_4792,N_45475,N_45471);
or UO_4793 (O_4793,N_46337,N_47970);
or UO_4794 (O_4794,N_49028,N_46252);
nand UO_4795 (O_4795,N_48500,N_45346);
nor UO_4796 (O_4796,N_46020,N_47978);
xnor UO_4797 (O_4797,N_46137,N_46466);
and UO_4798 (O_4798,N_46138,N_49556);
or UO_4799 (O_4799,N_47570,N_48726);
xnor UO_4800 (O_4800,N_49020,N_48210);
xor UO_4801 (O_4801,N_48485,N_49523);
nand UO_4802 (O_4802,N_47037,N_46461);
xor UO_4803 (O_4803,N_48973,N_46567);
nor UO_4804 (O_4804,N_46377,N_49876);
and UO_4805 (O_4805,N_46501,N_48060);
nor UO_4806 (O_4806,N_47996,N_45042);
nand UO_4807 (O_4807,N_49533,N_47663);
nand UO_4808 (O_4808,N_46399,N_46046);
nand UO_4809 (O_4809,N_47985,N_49792);
or UO_4810 (O_4810,N_45175,N_48609);
xor UO_4811 (O_4811,N_46500,N_46708);
or UO_4812 (O_4812,N_49442,N_48235);
nand UO_4813 (O_4813,N_46266,N_47464);
xnor UO_4814 (O_4814,N_48570,N_45751);
and UO_4815 (O_4815,N_45498,N_45673);
nor UO_4816 (O_4816,N_46627,N_46258);
or UO_4817 (O_4817,N_46804,N_45718);
xor UO_4818 (O_4818,N_49746,N_46709);
nand UO_4819 (O_4819,N_46635,N_45177);
nor UO_4820 (O_4820,N_46184,N_46555);
nor UO_4821 (O_4821,N_49159,N_49467);
and UO_4822 (O_4822,N_47379,N_48399);
and UO_4823 (O_4823,N_45844,N_48574);
or UO_4824 (O_4824,N_48800,N_48627);
nand UO_4825 (O_4825,N_47029,N_46217);
nor UO_4826 (O_4826,N_45181,N_49009);
xor UO_4827 (O_4827,N_48832,N_47203);
nor UO_4828 (O_4828,N_47794,N_48546);
xor UO_4829 (O_4829,N_48421,N_49145);
xnor UO_4830 (O_4830,N_48010,N_46633);
nand UO_4831 (O_4831,N_49062,N_46075);
nand UO_4832 (O_4832,N_45251,N_49076);
and UO_4833 (O_4833,N_46300,N_48625);
and UO_4834 (O_4834,N_47674,N_45560);
nand UO_4835 (O_4835,N_46449,N_49637);
and UO_4836 (O_4836,N_46891,N_45605);
and UO_4837 (O_4837,N_49299,N_49297);
nor UO_4838 (O_4838,N_46651,N_46662);
and UO_4839 (O_4839,N_45705,N_45987);
or UO_4840 (O_4840,N_47169,N_45649);
or UO_4841 (O_4841,N_45906,N_49804);
xor UO_4842 (O_4842,N_47262,N_46246);
nand UO_4843 (O_4843,N_46735,N_45202);
and UO_4844 (O_4844,N_49718,N_48540);
or UO_4845 (O_4845,N_49723,N_47648);
nor UO_4846 (O_4846,N_47755,N_47243);
and UO_4847 (O_4847,N_48479,N_49395);
and UO_4848 (O_4848,N_45161,N_46290);
or UO_4849 (O_4849,N_47893,N_45141);
nand UO_4850 (O_4850,N_46777,N_49628);
and UO_4851 (O_4851,N_49720,N_49851);
or UO_4852 (O_4852,N_47459,N_48977);
nor UO_4853 (O_4853,N_45112,N_45271);
or UO_4854 (O_4854,N_49003,N_46371);
nor UO_4855 (O_4855,N_48771,N_48562);
and UO_4856 (O_4856,N_46722,N_49357);
nand UO_4857 (O_4857,N_46411,N_48655);
nand UO_4858 (O_4858,N_46011,N_49243);
nand UO_4859 (O_4859,N_46190,N_48276);
nor UO_4860 (O_4860,N_48057,N_46456);
or UO_4861 (O_4861,N_48755,N_48575);
nand UO_4862 (O_4862,N_48440,N_48393);
nand UO_4863 (O_4863,N_47827,N_47145);
nor UO_4864 (O_4864,N_46572,N_48307);
nand UO_4865 (O_4865,N_49627,N_45497);
xor UO_4866 (O_4866,N_45416,N_46272);
nand UO_4867 (O_4867,N_46440,N_46766);
xor UO_4868 (O_4868,N_47012,N_48110);
nor UO_4869 (O_4869,N_49030,N_45338);
nand UO_4870 (O_4870,N_49370,N_49437);
or UO_4871 (O_4871,N_45182,N_45185);
and UO_4872 (O_4872,N_47616,N_48189);
and UO_4873 (O_4873,N_45948,N_45366);
nor UO_4874 (O_4874,N_48947,N_45190);
nand UO_4875 (O_4875,N_49806,N_47194);
nand UO_4876 (O_4876,N_47812,N_45580);
nand UO_4877 (O_4877,N_48936,N_45873);
and UO_4878 (O_4878,N_45153,N_45871);
nor UO_4879 (O_4879,N_46977,N_49644);
nand UO_4880 (O_4880,N_46808,N_47033);
or UO_4881 (O_4881,N_49367,N_46930);
or UO_4882 (O_4882,N_48858,N_46480);
xnor UO_4883 (O_4883,N_46489,N_45288);
or UO_4884 (O_4884,N_45771,N_49220);
nor UO_4885 (O_4885,N_48585,N_48139);
or UO_4886 (O_4886,N_45406,N_49153);
and UO_4887 (O_4887,N_47542,N_48016);
and UO_4888 (O_4888,N_47359,N_46915);
or UO_4889 (O_4889,N_47121,N_49472);
nor UO_4890 (O_4890,N_49959,N_47753);
xnor UO_4891 (O_4891,N_46460,N_45123);
nand UO_4892 (O_4892,N_49011,N_46449);
and UO_4893 (O_4893,N_46749,N_45850);
nor UO_4894 (O_4894,N_46584,N_45234);
nand UO_4895 (O_4895,N_49117,N_47524);
and UO_4896 (O_4896,N_45839,N_46332);
nand UO_4897 (O_4897,N_48446,N_45387);
nor UO_4898 (O_4898,N_48976,N_46552);
nand UO_4899 (O_4899,N_48855,N_46860);
or UO_4900 (O_4900,N_49915,N_48427);
nor UO_4901 (O_4901,N_45730,N_47327);
and UO_4902 (O_4902,N_49190,N_45545);
nand UO_4903 (O_4903,N_48293,N_46893);
and UO_4904 (O_4904,N_49555,N_45278);
xor UO_4905 (O_4905,N_48318,N_46694);
xor UO_4906 (O_4906,N_47529,N_46892);
and UO_4907 (O_4907,N_48851,N_47090);
xor UO_4908 (O_4908,N_49015,N_49048);
or UO_4909 (O_4909,N_46143,N_49106);
or UO_4910 (O_4910,N_46320,N_48190);
xnor UO_4911 (O_4911,N_48191,N_45702);
xor UO_4912 (O_4912,N_46261,N_46072);
nor UO_4913 (O_4913,N_48847,N_45346);
nor UO_4914 (O_4914,N_46488,N_49627);
xnor UO_4915 (O_4915,N_48288,N_46780);
or UO_4916 (O_4916,N_47523,N_45350);
nor UO_4917 (O_4917,N_45781,N_48415);
and UO_4918 (O_4918,N_49423,N_46491);
nand UO_4919 (O_4919,N_49965,N_48020);
or UO_4920 (O_4920,N_46735,N_48331);
nor UO_4921 (O_4921,N_45364,N_47507);
nor UO_4922 (O_4922,N_48811,N_49591);
nand UO_4923 (O_4923,N_48628,N_48794);
nand UO_4924 (O_4924,N_49411,N_45757);
nand UO_4925 (O_4925,N_48625,N_47381);
and UO_4926 (O_4926,N_45973,N_47990);
nor UO_4927 (O_4927,N_49799,N_48526);
nor UO_4928 (O_4928,N_46077,N_45310);
and UO_4929 (O_4929,N_47539,N_45326);
nand UO_4930 (O_4930,N_46594,N_48502);
nor UO_4931 (O_4931,N_49151,N_45405);
and UO_4932 (O_4932,N_46199,N_49794);
and UO_4933 (O_4933,N_46884,N_47368);
nand UO_4934 (O_4934,N_49287,N_47340);
nor UO_4935 (O_4935,N_46997,N_48338);
or UO_4936 (O_4936,N_48998,N_49858);
or UO_4937 (O_4937,N_48205,N_46350);
and UO_4938 (O_4938,N_49697,N_45194);
nor UO_4939 (O_4939,N_45127,N_47958);
and UO_4940 (O_4940,N_47622,N_45982);
nor UO_4941 (O_4941,N_47519,N_45823);
or UO_4942 (O_4942,N_47779,N_48579);
nand UO_4943 (O_4943,N_48924,N_47810);
or UO_4944 (O_4944,N_47222,N_46545);
or UO_4945 (O_4945,N_46712,N_45624);
nand UO_4946 (O_4946,N_46424,N_49988);
or UO_4947 (O_4947,N_48746,N_45416);
or UO_4948 (O_4948,N_46338,N_48664);
and UO_4949 (O_4949,N_49891,N_45657);
and UO_4950 (O_4950,N_46067,N_45961);
and UO_4951 (O_4951,N_49839,N_47783);
and UO_4952 (O_4952,N_48629,N_49548);
or UO_4953 (O_4953,N_46036,N_47199);
nand UO_4954 (O_4954,N_49993,N_46881);
or UO_4955 (O_4955,N_49754,N_49888);
or UO_4956 (O_4956,N_47203,N_48927);
nor UO_4957 (O_4957,N_46731,N_47762);
or UO_4958 (O_4958,N_49254,N_49116);
xor UO_4959 (O_4959,N_49756,N_47765);
nand UO_4960 (O_4960,N_47666,N_47836);
nor UO_4961 (O_4961,N_46479,N_49936);
nor UO_4962 (O_4962,N_47921,N_45359);
nor UO_4963 (O_4963,N_48207,N_45904);
or UO_4964 (O_4964,N_46751,N_48959);
nand UO_4965 (O_4965,N_47287,N_49237);
nor UO_4966 (O_4966,N_49899,N_47044);
nor UO_4967 (O_4967,N_49246,N_46530);
nor UO_4968 (O_4968,N_47898,N_48481);
xnor UO_4969 (O_4969,N_46551,N_46009);
nand UO_4970 (O_4970,N_45632,N_46901);
and UO_4971 (O_4971,N_49672,N_47806);
nand UO_4972 (O_4972,N_48464,N_49710);
or UO_4973 (O_4973,N_47264,N_47949);
or UO_4974 (O_4974,N_45001,N_47819);
or UO_4975 (O_4975,N_47105,N_49675);
or UO_4976 (O_4976,N_45352,N_46823);
and UO_4977 (O_4977,N_45309,N_46043);
nand UO_4978 (O_4978,N_47967,N_46054);
nand UO_4979 (O_4979,N_45259,N_47635);
nor UO_4980 (O_4980,N_48192,N_47652);
and UO_4981 (O_4981,N_48978,N_48430);
nand UO_4982 (O_4982,N_49337,N_46675);
xor UO_4983 (O_4983,N_45481,N_46052);
nor UO_4984 (O_4984,N_45313,N_45968);
nor UO_4985 (O_4985,N_46748,N_47630);
and UO_4986 (O_4986,N_46531,N_49781);
nand UO_4987 (O_4987,N_46741,N_49999);
or UO_4988 (O_4988,N_47501,N_45513);
or UO_4989 (O_4989,N_49942,N_48237);
and UO_4990 (O_4990,N_46532,N_48731);
nor UO_4991 (O_4991,N_47760,N_49445);
and UO_4992 (O_4992,N_48299,N_49825);
nor UO_4993 (O_4993,N_46613,N_49017);
or UO_4994 (O_4994,N_48162,N_47016);
nand UO_4995 (O_4995,N_49684,N_45850);
and UO_4996 (O_4996,N_45430,N_45485);
and UO_4997 (O_4997,N_47362,N_47373);
and UO_4998 (O_4998,N_46464,N_46138);
and UO_4999 (O_4999,N_49274,N_48474);
endmodule