module basic_1000_10000_1500_20_levels_5xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
and U0 (N_0,In_501,In_111);
nand U1 (N_1,In_188,In_230);
and U2 (N_2,In_876,In_517);
and U3 (N_3,In_438,In_778);
or U4 (N_4,In_931,In_995);
and U5 (N_5,In_108,In_201);
nor U6 (N_6,In_270,In_71);
nand U7 (N_7,In_489,In_790);
or U8 (N_8,In_616,In_533);
xor U9 (N_9,In_179,In_804);
nand U10 (N_10,In_635,In_37);
xor U11 (N_11,In_6,In_186);
nor U12 (N_12,In_828,In_996);
and U13 (N_13,In_519,In_877);
nand U14 (N_14,In_624,In_194);
or U15 (N_15,In_477,In_861);
or U16 (N_16,In_484,In_520);
nand U17 (N_17,In_391,In_286);
and U18 (N_18,In_18,In_570);
and U19 (N_19,In_394,In_76);
nand U20 (N_20,In_573,In_531);
and U21 (N_21,In_219,In_26);
and U22 (N_22,In_283,In_120);
or U23 (N_23,In_740,In_96);
or U24 (N_24,In_481,In_572);
nor U25 (N_25,In_408,In_374);
nand U26 (N_26,In_504,In_248);
nand U27 (N_27,In_850,In_918);
xnor U28 (N_28,In_537,In_817);
and U29 (N_29,In_310,In_753);
nor U30 (N_30,In_147,In_524);
and U31 (N_31,In_898,In_433);
nand U32 (N_32,In_767,In_422);
nor U33 (N_33,In_508,In_991);
nor U34 (N_34,In_428,In_264);
or U35 (N_35,In_739,In_676);
nor U36 (N_36,In_540,In_378);
nor U37 (N_37,In_290,In_172);
xor U38 (N_38,In_759,In_278);
and U39 (N_39,In_687,In_254);
nand U40 (N_40,In_69,In_605);
nand U41 (N_41,In_403,In_232);
nand U42 (N_42,In_471,In_858);
or U43 (N_43,In_122,In_192);
nor U44 (N_44,In_937,In_947);
or U45 (N_45,In_217,In_810);
nor U46 (N_46,In_466,In_974);
or U47 (N_47,In_480,In_284);
and U48 (N_48,In_765,In_72);
or U49 (N_49,In_240,In_648);
nor U50 (N_50,In_855,In_314);
nand U51 (N_51,In_27,In_756);
xor U52 (N_52,In_620,In_157);
and U53 (N_53,In_338,In_706);
or U54 (N_54,In_46,In_460);
nand U55 (N_55,In_574,In_784);
and U56 (N_56,In_358,In_972);
and U57 (N_57,In_981,In_672);
and U58 (N_58,In_594,In_214);
xor U59 (N_59,In_900,In_293);
xor U60 (N_60,In_993,In_780);
or U61 (N_61,In_805,In_811);
xor U62 (N_62,In_277,In_450);
nor U63 (N_63,In_306,In_137);
and U64 (N_64,In_545,In_838);
or U65 (N_65,In_532,In_603);
and U66 (N_66,In_614,In_48);
nor U67 (N_67,In_109,In_643);
nand U68 (N_68,In_239,In_81);
nand U69 (N_69,In_263,In_772);
or U70 (N_70,In_39,In_365);
nor U71 (N_71,In_255,In_454);
xnor U72 (N_72,In_329,In_198);
or U73 (N_73,In_802,In_853);
nor U74 (N_74,In_300,In_766);
nor U75 (N_75,In_395,In_190);
and U76 (N_76,In_500,In_177);
nand U77 (N_77,In_813,In_667);
or U78 (N_78,In_102,In_820);
and U79 (N_79,In_328,In_985);
and U80 (N_80,In_384,In_11);
and U81 (N_81,In_116,In_758);
nand U82 (N_82,In_912,In_410);
and U83 (N_83,In_13,In_237);
and U84 (N_84,In_875,In_640);
and U85 (N_85,In_107,In_146);
nor U86 (N_86,In_138,In_722);
nand U87 (N_87,In_982,In_854);
nand U88 (N_88,In_266,In_337);
and U89 (N_89,In_692,In_274);
or U90 (N_90,In_970,In_564);
and U91 (N_91,In_407,In_65);
or U92 (N_92,In_521,In_807);
nor U93 (N_93,In_835,In_461);
and U94 (N_94,In_24,In_720);
or U95 (N_95,In_741,In_78);
xor U96 (N_96,In_404,In_843);
or U97 (N_97,In_690,In_942);
or U98 (N_98,In_886,In_117);
and U99 (N_99,In_431,In_891);
and U100 (N_100,In_356,In_375);
nand U101 (N_101,In_303,In_389);
or U102 (N_102,In_934,In_355);
or U103 (N_103,In_381,In_79);
and U104 (N_104,In_650,In_400);
or U105 (N_105,In_150,In_644);
and U106 (N_106,In_344,In_7);
xnor U107 (N_107,In_983,In_830);
nor U108 (N_108,In_556,In_724);
nor U109 (N_109,In_241,In_615);
or U110 (N_110,In_144,In_599);
nor U111 (N_111,In_353,In_253);
and U112 (N_112,In_244,In_304);
nand U113 (N_113,In_448,In_215);
nor U114 (N_114,In_485,In_60);
and U115 (N_115,In_459,In_536);
or U116 (N_116,In_955,In_131);
nor U117 (N_117,In_326,In_617);
nand U118 (N_118,In_658,In_630);
and U119 (N_119,In_362,In_806);
nand U120 (N_120,In_246,In_622);
nand U121 (N_121,In_213,In_771);
and U122 (N_122,In_625,In_307);
or U123 (N_123,In_135,In_915);
xor U124 (N_124,In_357,In_867);
or U125 (N_125,In_323,In_827);
nand U126 (N_126,In_354,In_693);
xor U127 (N_127,In_231,In_161);
and U128 (N_128,In_997,In_350);
and U129 (N_129,In_604,In_833);
nand U130 (N_130,In_197,In_289);
xor U131 (N_131,In_52,In_718);
nor U132 (N_132,In_542,In_467);
xnor U133 (N_133,In_799,In_364);
and U134 (N_134,In_969,In_429);
or U135 (N_135,In_779,In_265);
and U136 (N_136,In_941,In_469);
xnor U137 (N_137,In_530,In_988);
nor U138 (N_138,In_68,In_414);
xor U139 (N_139,In_619,In_539);
nand U140 (N_140,In_607,In_697);
and U141 (N_141,In_41,In_881);
nand U142 (N_142,In_57,In_346);
and U143 (N_143,In_954,In_800);
nand U144 (N_144,In_583,In_923);
or U145 (N_145,In_200,In_966);
and U146 (N_146,In_924,In_751);
nand U147 (N_147,In_432,In_888);
nand U148 (N_148,In_38,In_309);
nor U149 (N_149,In_476,In_869);
nand U150 (N_150,In_348,In_401);
and U151 (N_151,In_787,In_294);
or U152 (N_152,In_322,In_960);
or U153 (N_153,In_773,In_872);
nand U154 (N_154,In_535,In_297);
xnor U155 (N_155,In_575,In_761);
nand U156 (N_156,In_848,In_268);
and U157 (N_157,In_950,In_93);
nand U158 (N_158,In_863,In_791);
xor U159 (N_159,In_725,In_12);
nor U160 (N_160,In_19,In_158);
and U161 (N_161,In_977,In_45);
or U162 (N_162,In_698,In_238);
or U163 (N_163,In_713,In_503);
and U164 (N_164,In_701,In_785);
nand U165 (N_165,In_124,In_170);
nor U166 (N_166,In_451,In_409);
nor U167 (N_167,In_475,In_700);
nand U168 (N_168,In_973,In_957);
nor U169 (N_169,In_153,In_180);
and U170 (N_170,In_525,In_97);
xnor U171 (N_171,In_171,In_491);
and U172 (N_172,In_351,In_9);
nor U173 (N_173,In_16,In_708);
nor U174 (N_174,In_203,In_516);
nor U175 (N_175,In_175,In_112);
and U176 (N_176,In_435,In_205);
and U177 (N_177,In_465,In_664);
or U178 (N_178,In_449,In_398);
or U179 (N_179,In_482,In_638);
xor U180 (N_180,In_225,In_506);
xnor U181 (N_181,In_49,In_84);
nor U182 (N_182,In_557,In_296);
nor U183 (N_183,In_383,In_627);
and U184 (N_184,In_814,In_749);
and U185 (N_185,In_932,In_94);
and U186 (N_186,In_308,In_544);
nor U187 (N_187,In_498,In_14);
nor U188 (N_188,In_686,In_757);
xnor U189 (N_189,In_665,In_699);
nand U190 (N_190,In_486,In_818);
xor U191 (N_191,In_4,In_669);
and U192 (N_192,In_56,In_427);
nor U193 (N_193,In_752,In_986);
nor U194 (N_194,In_34,In_457);
nor U195 (N_195,In_373,In_889);
nor U196 (N_196,In_430,In_420);
nand U197 (N_197,In_559,In_515);
or U198 (N_198,In_563,In_971);
nor U199 (N_199,In_98,In_512);
and U200 (N_200,In_642,In_55);
nand U201 (N_201,In_865,In_839);
or U202 (N_202,In_141,In_943);
or U203 (N_203,In_837,In_893);
or U204 (N_204,In_242,In_866);
nand U205 (N_205,In_319,In_793);
and U206 (N_206,In_914,In_589);
and U207 (N_207,In_396,In_577);
or U208 (N_208,In_815,In_887);
nand U209 (N_209,In_376,In_377);
and U210 (N_210,In_682,In_361);
and U211 (N_211,In_788,In_714);
and U212 (N_212,In_149,In_458);
or U213 (N_213,In_646,In_490);
nor U214 (N_214,In_317,In_281);
or U215 (N_215,In_597,In_250);
or U216 (N_216,In_5,In_495);
nand U217 (N_217,In_769,In_656);
xnor U218 (N_218,In_321,In_100);
nand U219 (N_219,In_1,In_655);
and U220 (N_220,In_110,In_909);
and U221 (N_221,In_940,In_154);
or U222 (N_222,In_152,In_908);
or U223 (N_223,In_743,In_202);
and U224 (N_224,In_593,In_226);
nor U225 (N_225,In_132,In_77);
nand U226 (N_226,In_185,In_663);
or U227 (N_227,In_582,In_155);
nor U228 (N_228,In_312,In_590);
nand U229 (N_229,In_511,In_978);
xnor U230 (N_230,In_808,In_823);
nor U231 (N_231,In_261,In_21);
or U232 (N_232,In_862,In_474);
nor U233 (N_233,In_975,In_212);
or U234 (N_234,In_683,In_812);
and U235 (N_235,In_412,In_731);
nor U236 (N_236,In_846,In_101);
and U237 (N_237,In_387,In_426);
nand U238 (N_238,In_632,In_796);
or U239 (N_239,In_847,In_236);
nand U240 (N_240,In_935,In_229);
nand U241 (N_241,In_874,In_316);
nand U242 (N_242,In_927,In_273);
nor U243 (N_243,In_845,In_330);
and U244 (N_244,In_195,In_445);
nor U245 (N_245,In_390,In_671);
nor U246 (N_246,In_775,In_159);
and U247 (N_247,In_528,In_762);
or U248 (N_248,In_715,In_189);
nand U249 (N_249,In_911,In_167);
or U250 (N_250,In_860,In_726);
nor U251 (N_251,In_613,In_952);
nand U252 (N_252,In_781,In_89);
nand U253 (N_253,In_191,In_82);
and U254 (N_254,In_32,In_803);
or U255 (N_255,In_998,In_629);
and U256 (N_256,In_43,In_372);
or U257 (N_257,In_456,In_140);
nor U258 (N_258,In_473,In_178);
and U259 (N_259,In_505,In_600);
nand U260 (N_260,In_88,In_251);
and U261 (N_261,In_29,In_857);
and U262 (N_262,In_782,In_989);
nor U263 (N_263,In_35,In_134);
nand U264 (N_264,In_976,In_568);
nor U265 (N_265,In_962,In_606);
or U266 (N_266,In_113,In_645);
nand U267 (N_267,In_369,In_580);
or U268 (N_268,In_335,In_86);
or U269 (N_269,In_841,In_340);
nor U270 (N_270,In_562,In_143);
or U271 (N_271,In_492,In_125);
and U272 (N_272,In_695,In_343);
or U273 (N_273,In_488,In_946);
nand U274 (N_274,In_406,In_463);
and U275 (N_275,In_258,In_596);
nor U276 (N_276,In_670,In_649);
nor U277 (N_277,In_103,In_939);
nor U278 (N_278,In_878,In_608);
or U279 (N_279,In_868,In_173);
nand U280 (N_280,In_275,In_612);
and U281 (N_281,In_716,In_439);
or U282 (N_282,In_207,In_405);
and U283 (N_283,In_992,In_680);
and U284 (N_284,In_3,In_894);
nor U285 (N_285,In_555,In_595);
and U286 (N_286,In_738,In_732);
nand U287 (N_287,In_679,In_10);
or U288 (N_288,In_423,In_436);
nor U289 (N_289,In_371,In_534);
xnor U290 (N_290,In_28,In_368);
nor U291 (N_291,In_585,In_415);
or U292 (N_292,In_628,In_437);
nor U293 (N_293,In_419,In_487);
or U294 (N_294,In_895,In_548);
or U295 (N_295,In_67,In_822);
and U296 (N_296,In_674,In_507);
nand U297 (N_297,In_884,In_626);
nor U298 (N_298,In_22,In_204);
and U299 (N_299,In_527,In_61);
or U300 (N_300,In_33,In_176);
nor U301 (N_301,In_930,In_47);
or U302 (N_302,In_744,In_675);
nand U303 (N_303,In_734,In_631);
and U304 (N_304,In_994,In_551);
nand U305 (N_305,In_342,In_913);
nand U306 (N_306,In_901,In_388);
or U307 (N_307,In_315,In_434);
nor U308 (N_308,In_206,In_216);
nand U309 (N_309,In_397,In_31);
nor U310 (N_310,In_929,In_880);
xnor U311 (N_311,In_413,In_62);
nor U312 (N_312,In_873,In_786);
nand U313 (N_313,In_162,In_119);
or U314 (N_314,In_844,In_15);
nand U315 (N_315,In_165,In_95);
nor U316 (N_316,In_174,In_964);
nand U317 (N_317,In_257,In_842);
or U318 (N_318,In_320,In_668);
nand U319 (N_319,In_689,In_792);
or U320 (N_320,In_879,In_621);
or U321 (N_321,In_523,In_262);
nand U322 (N_322,In_127,In_938);
nand U323 (N_323,In_906,In_661);
and U324 (N_324,In_243,In_836);
nor U325 (N_325,In_925,In_341);
nand U326 (N_326,In_933,In_370);
and U327 (N_327,In_709,In_99);
nand U328 (N_328,In_592,In_494);
nor U329 (N_329,In_897,In_493);
or U330 (N_330,In_849,In_502);
nand U331 (N_331,In_591,In_961);
and U332 (N_332,In_292,In_549);
nor U333 (N_333,In_851,In_73);
and U334 (N_334,In_118,In_333);
xnor U335 (N_335,In_916,In_541);
and U336 (N_336,In_75,In_859);
or U337 (N_337,In_870,In_256);
nand U338 (N_338,In_633,In_852);
xnor U339 (N_339,In_623,In_196);
and U340 (N_340,In_464,In_247);
and U341 (N_341,In_776,In_352);
nand U342 (N_342,In_637,In_411);
xnor U343 (N_343,In_890,In_104);
nor U344 (N_344,In_871,In_735);
nor U345 (N_345,In_360,In_907);
nand U346 (N_346,In_91,In_719);
nor U347 (N_347,In_745,In_949);
and U348 (N_348,In_345,In_910);
and U349 (N_349,In_228,In_578);
and U350 (N_350,In_958,In_139);
or U351 (N_351,In_349,In_948);
and U352 (N_352,In_944,In_959);
or U353 (N_353,In_455,In_50);
or U354 (N_354,In_651,In_252);
and U355 (N_355,In_774,In_305);
nor U356 (N_356,In_163,In_902);
nor U357 (N_357,In_730,In_156);
nor U358 (N_358,In_684,In_882);
nand U359 (N_359,In_641,In_727);
nand U360 (N_360,In_318,In_130);
xor U361 (N_361,In_809,In_509);
nand U362 (N_362,In_569,In_115);
nand U363 (N_363,In_601,In_211);
or U364 (N_364,In_145,In_496);
nor U365 (N_365,In_783,In_653);
or U366 (N_366,In_967,In_193);
and U367 (N_367,In_736,In_30);
nand U368 (N_368,In_618,In_382);
and U369 (N_369,In_768,In_903);
or U370 (N_370,In_990,In_90);
nor U371 (N_371,In_187,In_794);
or U372 (N_372,In_586,In_560);
or U373 (N_373,In_770,In_199);
xnor U374 (N_374,In_609,In_325);
nand U375 (N_375,In_151,In_681);
nor U376 (N_376,In_20,In_755);
and U377 (N_377,In_367,In_919);
xnor U378 (N_378,In_711,In_673);
nor U379 (N_379,In_834,In_729);
nand U380 (N_380,In_418,In_105);
xor U381 (N_381,In_760,In_576);
or U382 (N_382,In_703,In_571);
xnor U383 (N_383,In_639,In_510);
nand U384 (N_384,In_647,In_453);
nor U385 (N_385,In_479,In_129);
and U386 (N_386,In_444,In_797);
or U387 (N_387,In_798,In_166);
or U388 (N_388,In_904,In_657);
or U389 (N_389,In_553,In_121);
nand U390 (N_390,In_529,In_223);
nand U391 (N_391,In_164,In_518);
or U392 (N_392,In_922,In_702);
nor U393 (N_393,In_291,In_58);
nand U394 (N_394,In_332,In_380);
nor U395 (N_395,In_737,In_470);
nor U396 (N_396,In_440,In_587);
nor U397 (N_397,In_746,In_183);
nor U398 (N_398,In_269,In_763);
nor U399 (N_399,In_588,In_386);
and U400 (N_400,In_677,In_25);
nor U401 (N_401,In_276,In_824);
xnor U402 (N_402,In_54,In_301);
nor U403 (N_403,In_446,In_425);
nor U404 (N_404,In_23,In_385);
and U405 (N_405,In_282,In_280);
or U406 (N_406,In_468,In_421);
and U407 (N_407,In_659,In_227);
nand U408 (N_408,In_324,In_816);
or U409 (N_409,In_953,In_339);
nor U410 (N_410,In_181,In_678);
nand U411 (N_411,In_462,In_416);
or U412 (N_412,In_220,In_685);
nor U413 (N_413,In_331,In_602);
or U414 (N_414,In_538,In_611);
nand U415 (N_415,In_478,In_272);
and U416 (N_416,In_567,In_87);
or U417 (N_417,In_366,In_233);
xor U418 (N_418,In_987,In_723);
nand U419 (N_419,In_999,In_979);
or U420 (N_420,In_883,In_652);
nand U421 (N_421,In_40,In_399);
nor U422 (N_422,In_235,In_864);
nor U423 (N_423,In_552,In_748);
or U424 (N_424,In_899,In_565);
and U425 (N_425,In_169,In_892);
or U426 (N_426,In_610,In_106);
nand U427 (N_427,In_704,In_584);
or U428 (N_428,In_707,In_554);
nand U429 (N_429,In_210,In_288);
or U430 (N_430,In_447,In_885);
nor U431 (N_431,In_826,In_160);
or U432 (N_432,In_0,In_336);
nand U433 (N_433,In_53,In_51);
and U434 (N_434,In_579,In_259);
nand U435 (N_435,In_547,In_951);
or U436 (N_436,In_968,In_710);
and U437 (N_437,In_546,In_558);
or U438 (N_438,In_819,In_472);
and U439 (N_439,In_483,In_302);
or U440 (N_440,In_393,In_821);
nand U441 (N_441,In_70,In_750);
or U442 (N_442,In_64,In_840);
nor U443 (N_443,In_85,In_497);
nor U444 (N_444,In_598,In_287);
and U445 (N_445,In_245,In_208);
nor U446 (N_446,In_742,In_295);
xor U447 (N_447,In_963,In_392);
nor U448 (N_448,In_825,In_224);
nand U449 (N_449,In_956,In_543);
nand U450 (N_450,In_654,In_441);
or U451 (N_451,In_514,In_114);
and U452 (N_452,In_777,In_696);
or U453 (N_453,In_452,In_712);
and U454 (N_454,In_184,In_513);
and U455 (N_455,In_666,In_80);
or U456 (N_456,In_168,In_36);
nand U457 (N_457,In_267,In_209);
nand U458 (N_458,In_234,In_984);
or U459 (N_459,In_581,In_2);
nor U460 (N_460,In_123,In_379);
nand U461 (N_461,In_896,In_831);
or U462 (N_462,In_728,In_142);
nor U463 (N_463,In_747,In_66);
and U464 (N_464,In_733,In_550);
nor U465 (N_465,In_636,In_44);
nor U466 (N_466,In_334,In_945);
and U467 (N_467,In_279,In_271);
nor U468 (N_468,In_691,In_829);
nand U469 (N_469,In_92,In_8);
and U470 (N_470,In_221,In_832);
nand U471 (N_471,In_921,In_299);
xnor U472 (N_472,In_694,In_566);
and U473 (N_473,In_133,In_754);
nand U474 (N_474,In_795,In_260);
nand U475 (N_475,In_926,In_442);
or U476 (N_476,In_218,In_222);
nand U477 (N_477,In_42,In_936);
nor U478 (N_478,In_920,In_721);
nor U479 (N_479,In_136,In_662);
and U480 (N_480,In_311,In_856);
and U481 (N_481,In_526,In_128);
nor U482 (N_482,In_928,In_717);
or U483 (N_483,In_705,In_499);
and U484 (N_484,In_965,In_801);
nor U485 (N_485,In_660,In_789);
xor U486 (N_486,In_74,In_285);
nor U487 (N_487,In_313,In_182);
or U488 (N_488,In_688,In_443);
and U489 (N_489,In_402,In_347);
and U490 (N_490,In_148,In_561);
nand U491 (N_491,In_17,In_634);
and U492 (N_492,In_63,In_59);
nor U493 (N_493,In_298,In_424);
nand U494 (N_494,In_249,In_522);
nand U495 (N_495,In_764,In_417);
nor U496 (N_496,In_126,In_83);
nor U497 (N_497,In_980,In_905);
nand U498 (N_498,In_359,In_917);
nand U499 (N_499,In_363,In_327);
nor U500 (N_500,N_328,N_385);
or U501 (N_501,N_497,N_139);
and U502 (N_502,N_227,N_112);
and U503 (N_503,N_127,N_162);
nand U504 (N_504,N_248,N_95);
nand U505 (N_505,N_234,N_450);
nand U506 (N_506,N_366,N_246);
or U507 (N_507,N_51,N_260);
nor U508 (N_508,N_157,N_67);
nand U509 (N_509,N_77,N_347);
nand U510 (N_510,N_436,N_109);
or U511 (N_511,N_206,N_318);
nor U512 (N_512,N_439,N_478);
or U513 (N_513,N_462,N_185);
and U514 (N_514,N_9,N_28);
nand U515 (N_515,N_433,N_331);
nor U516 (N_516,N_335,N_396);
nor U517 (N_517,N_36,N_339);
or U518 (N_518,N_147,N_62);
nor U519 (N_519,N_167,N_447);
or U520 (N_520,N_455,N_132);
nor U521 (N_521,N_448,N_445);
and U522 (N_522,N_255,N_75);
xor U523 (N_523,N_459,N_39);
xnor U524 (N_524,N_86,N_499);
and U525 (N_525,N_294,N_374);
xnor U526 (N_526,N_250,N_437);
nor U527 (N_527,N_201,N_176);
nand U528 (N_528,N_498,N_473);
and U529 (N_529,N_186,N_317);
nand U530 (N_530,N_244,N_40);
and U531 (N_531,N_191,N_474);
nor U532 (N_532,N_333,N_57);
and U533 (N_533,N_113,N_119);
or U534 (N_534,N_222,N_355);
and U535 (N_535,N_104,N_211);
nand U536 (N_536,N_232,N_135);
and U537 (N_537,N_419,N_470);
or U538 (N_538,N_428,N_172);
nor U539 (N_539,N_426,N_143);
xnor U540 (N_540,N_168,N_133);
or U541 (N_541,N_44,N_171);
nand U542 (N_542,N_224,N_103);
and U543 (N_543,N_251,N_332);
xor U544 (N_544,N_137,N_3);
nand U545 (N_545,N_376,N_410);
xnor U546 (N_546,N_43,N_116);
or U547 (N_547,N_397,N_142);
nand U548 (N_548,N_321,N_226);
xor U549 (N_549,N_280,N_373);
or U550 (N_550,N_60,N_151);
nor U551 (N_551,N_306,N_277);
and U552 (N_552,N_496,N_472);
nor U553 (N_553,N_298,N_492);
and U554 (N_554,N_189,N_22);
nor U555 (N_555,N_285,N_356);
xor U556 (N_556,N_384,N_230);
and U557 (N_557,N_466,N_268);
xnor U558 (N_558,N_461,N_111);
xnor U559 (N_559,N_33,N_93);
nor U560 (N_560,N_270,N_435);
and U561 (N_561,N_399,N_365);
or U562 (N_562,N_272,N_73);
nor U563 (N_563,N_405,N_491);
nand U564 (N_564,N_130,N_330);
and U565 (N_565,N_346,N_30);
xor U566 (N_566,N_386,N_90);
xnor U567 (N_567,N_345,N_307);
nor U568 (N_568,N_489,N_182);
nor U569 (N_569,N_418,N_249);
and U570 (N_570,N_202,N_129);
or U571 (N_571,N_41,N_278);
nor U572 (N_572,N_449,N_344);
or U573 (N_573,N_241,N_324);
and U574 (N_574,N_273,N_266);
and U575 (N_575,N_23,N_262);
nand U576 (N_576,N_19,N_247);
xor U577 (N_577,N_149,N_281);
nand U578 (N_578,N_102,N_263);
nor U579 (N_579,N_74,N_422);
nand U580 (N_580,N_488,N_456);
nand U581 (N_581,N_326,N_444);
and U582 (N_582,N_32,N_21);
or U583 (N_583,N_291,N_415);
and U584 (N_584,N_391,N_493);
xor U585 (N_585,N_259,N_343);
xnor U586 (N_586,N_423,N_297);
nand U587 (N_587,N_400,N_175);
nand U588 (N_588,N_220,N_468);
or U589 (N_589,N_115,N_380);
nor U590 (N_590,N_97,N_388);
nand U591 (N_591,N_398,N_166);
or U592 (N_592,N_184,N_308);
nand U593 (N_593,N_315,N_245);
nor U594 (N_594,N_377,N_427);
and U595 (N_595,N_408,N_451);
nand U596 (N_596,N_215,N_200);
nand U597 (N_597,N_94,N_411);
nand U598 (N_598,N_17,N_100);
nand U599 (N_599,N_31,N_293);
nand U600 (N_600,N_204,N_138);
nand U601 (N_601,N_359,N_229);
or U602 (N_602,N_197,N_364);
or U603 (N_603,N_209,N_253);
or U604 (N_604,N_153,N_37);
nor U605 (N_605,N_301,N_216);
or U606 (N_606,N_425,N_59);
and U607 (N_607,N_218,N_208);
and U608 (N_608,N_309,N_35);
nand U609 (N_609,N_487,N_25);
or U610 (N_610,N_379,N_163);
or U611 (N_611,N_231,N_336);
xnor U612 (N_612,N_389,N_296);
nand U613 (N_613,N_349,N_124);
nand U614 (N_614,N_342,N_121);
nand U615 (N_615,N_261,N_403);
nor U616 (N_616,N_190,N_367);
or U617 (N_617,N_63,N_72);
nand U618 (N_618,N_453,N_50);
or U619 (N_619,N_18,N_322);
and U620 (N_620,N_158,N_414);
nand U621 (N_621,N_114,N_480);
and U622 (N_622,N_430,N_454);
or U623 (N_623,N_290,N_5);
and U624 (N_624,N_26,N_193);
nand U625 (N_625,N_310,N_432);
nand U626 (N_626,N_71,N_394);
and U627 (N_627,N_392,N_479);
nand U628 (N_628,N_465,N_126);
or U629 (N_629,N_238,N_416);
and U630 (N_630,N_150,N_165);
and U631 (N_631,N_164,N_368);
nand U632 (N_632,N_76,N_337);
nor U633 (N_633,N_288,N_213);
or U634 (N_634,N_484,N_174);
and U635 (N_635,N_48,N_282);
xnor U636 (N_636,N_99,N_458);
xor U637 (N_637,N_457,N_141);
nand U638 (N_638,N_117,N_148);
or U639 (N_639,N_159,N_122);
and U640 (N_640,N_107,N_11);
nor U641 (N_641,N_4,N_486);
and U642 (N_642,N_6,N_275);
or U643 (N_643,N_303,N_199);
xnor U644 (N_644,N_8,N_240);
or U645 (N_645,N_88,N_481);
nand U646 (N_646,N_312,N_181);
and U647 (N_647,N_128,N_390);
nor U648 (N_648,N_283,N_329);
nor U649 (N_649,N_54,N_58);
nor U650 (N_650,N_160,N_289);
nand U651 (N_651,N_271,N_482);
or U652 (N_652,N_110,N_125);
and U653 (N_653,N_357,N_34);
nor U654 (N_654,N_89,N_20);
or U655 (N_655,N_1,N_78);
nand U656 (N_656,N_69,N_53);
nand U657 (N_657,N_434,N_383);
and U658 (N_658,N_304,N_12);
xor U659 (N_659,N_188,N_313);
or U660 (N_660,N_210,N_257);
nor U661 (N_661,N_452,N_471);
and U662 (N_662,N_299,N_311);
or U663 (N_663,N_363,N_169);
nand U664 (N_664,N_108,N_120);
and U665 (N_665,N_440,N_348);
nand U666 (N_666,N_91,N_161);
or U667 (N_667,N_217,N_45);
and U668 (N_668,N_205,N_460);
xor U669 (N_669,N_327,N_287);
xnor U670 (N_670,N_196,N_406);
or U671 (N_671,N_409,N_446);
nand U672 (N_672,N_494,N_475);
nand U673 (N_673,N_354,N_340);
and U674 (N_674,N_56,N_323);
nand U675 (N_675,N_61,N_178);
or U676 (N_676,N_469,N_276);
nor U677 (N_677,N_362,N_361);
and U678 (N_678,N_105,N_334);
nand U679 (N_679,N_319,N_412);
nor U680 (N_680,N_2,N_146);
and U681 (N_681,N_269,N_341);
xor U682 (N_682,N_214,N_29);
nand U683 (N_683,N_80,N_85);
and U684 (N_684,N_52,N_420);
nor U685 (N_685,N_360,N_413);
and U686 (N_686,N_221,N_180);
nor U687 (N_687,N_81,N_477);
or U688 (N_688,N_207,N_314);
xor U689 (N_689,N_279,N_431);
nor U690 (N_690,N_14,N_223);
nand U691 (N_691,N_438,N_225);
nand U692 (N_692,N_254,N_401);
or U693 (N_693,N_92,N_84);
or U694 (N_694,N_123,N_64);
nor U695 (N_695,N_265,N_55);
nor U696 (N_696,N_325,N_68);
nor U697 (N_697,N_476,N_252);
nor U698 (N_698,N_101,N_286);
nor U699 (N_699,N_136,N_179);
nand U700 (N_700,N_353,N_70);
nand U701 (N_701,N_198,N_442);
nand U702 (N_702,N_375,N_350);
or U703 (N_703,N_131,N_13);
nor U704 (N_704,N_404,N_42);
nand U705 (N_705,N_236,N_228);
nor U706 (N_706,N_7,N_219);
or U707 (N_707,N_378,N_264);
or U708 (N_708,N_87,N_300);
nand U709 (N_709,N_382,N_235);
nor U710 (N_710,N_118,N_134);
and U711 (N_711,N_387,N_239);
nor U712 (N_712,N_352,N_242);
or U713 (N_713,N_395,N_402);
and U714 (N_714,N_83,N_46);
nand U715 (N_715,N_302,N_173);
or U716 (N_716,N_490,N_144);
nor U717 (N_717,N_417,N_407);
or U718 (N_718,N_195,N_82);
nor U719 (N_719,N_443,N_154);
xnor U720 (N_720,N_66,N_233);
nor U721 (N_721,N_295,N_429);
and U722 (N_722,N_38,N_421);
or U723 (N_723,N_424,N_47);
and U724 (N_724,N_381,N_258);
nor U725 (N_725,N_320,N_237);
nand U726 (N_726,N_483,N_292);
or U727 (N_727,N_256,N_152);
and U728 (N_728,N_183,N_393);
or U729 (N_729,N_371,N_351);
nor U730 (N_730,N_369,N_212);
nor U731 (N_731,N_24,N_305);
nand U732 (N_732,N_495,N_372);
and U733 (N_733,N_203,N_98);
nor U734 (N_734,N_338,N_441);
and U735 (N_735,N_106,N_316);
and U736 (N_736,N_0,N_485);
and U737 (N_737,N_156,N_284);
nor U738 (N_738,N_370,N_464);
nor U739 (N_739,N_358,N_243);
or U740 (N_740,N_170,N_177);
or U741 (N_741,N_140,N_16);
and U742 (N_742,N_463,N_79);
nor U743 (N_743,N_27,N_96);
or U744 (N_744,N_467,N_274);
or U745 (N_745,N_49,N_194);
or U746 (N_746,N_15,N_65);
xor U747 (N_747,N_145,N_155);
or U748 (N_748,N_267,N_187);
nand U749 (N_749,N_10,N_192);
nor U750 (N_750,N_12,N_113);
nand U751 (N_751,N_218,N_377);
and U752 (N_752,N_273,N_467);
and U753 (N_753,N_478,N_375);
nand U754 (N_754,N_67,N_235);
nand U755 (N_755,N_111,N_5);
xnor U756 (N_756,N_10,N_183);
nor U757 (N_757,N_282,N_176);
nand U758 (N_758,N_480,N_365);
xor U759 (N_759,N_414,N_324);
nand U760 (N_760,N_236,N_188);
or U761 (N_761,N_355,N_273);
nand U762 (N_762,N_129,N_43);
xnor U763 (N_763,N_335,N_205);
nor U764 (N_764,N_242,N_20);
xnor U765 (N_765,N_334,N_58);
nand U766 (N_766,N_29,N_229);
and U767 (N_767,N_301,N_7);
nor U768 (N_768,N_280,N_281);
nor U769 (N_769,N_487,N_237);
nor U770 (N_770,N_218,N_328);
nor U771 (N_771,N_280,N_188);
or U772 (N_772,N_101,N_246);
and U773 (N_773,N_477,N_474);
nor U774 (N_774,N_496,N_183);
or U775 (N_775,N_326,N_124);
or U776 (N_776,N_138,N_48);
nand U777 (N_777,N_460,N_281);
and U778 (N_778,N_476,N_64);
nand U779 (N_779,N_495,N_244);
and U780 (N_780,N_169,N_372);
or U781 (N_781,N_29,N_112);
nand U782 (N_782,N_457,N_93);
nor U783 (N_783,N_254,N_322);
and U784 (N_784,N_437,N_361);
and U785 (N_785,N_351,N_356);
and U786 (N_786,N_148,N_470);
xor U787 (N_787,N_305,N_481);
or U788 (N_788,N_185,N_411);
or U789 (N_789,N_43,N_484);
xnor U790 (N_790,N_441,N_152);
nand U791 (N_791,N_335,N_268);
nor U792 (N_792,N_149,N_159);
and U793 (N_793,N_396,N_88);
or U794 (N_794,N_362,N_35);
nand U795 (N_795,N_131,N_109);
or U796 (N_796,N_212,N_295);
and U797 (N_797,N_62,N_250);
or U798 (N_798,N_198,N_498);
nor U799 (N_799,N_250,N_58);
nor U800 (N_800,N_62,N_465);
nor U801 (N_801,N_429,N_442);
nor U802 (N_802,N_499,N_62);
and U803 (N_803,N_10,N_412);
and U804 (N_804,N_460,N_23);
or U805 (N_805,N_91,N_76);
and U806 (N_806,N_117,N_127);
nor U807 (N_807,N_456,N_202);
nor U808 (N_808,N_158,N_235);
nand U809 (N_809,N_136,N_214);
xor U810 (N_810,N_201,N_409);
nand U811 (N_811,N_300,N_438);
or U812 (N_812,N_398,N_224);
nand U813 (N_813,N_36,N_181);
nand U814 (N_814,N_168,N_60);
and U815 (N_815,N_485,N_122);
and U816 (N_816,N_207,N_201);
and U817 (N_817,N_233,N_287);
and U818 (N_818,N_408,N_259);
or U819 (N_819,N_214,N_388);
nor U820 (N_820,N_460,N_70);
nand U821 (N_821,N_419,N_325);
xor U822 (N_822,N_315,N_123);
or U823 (N_823,N_313,N_104);
and U824 (N_824,N_454,N_477);
nand U825 (N_825,N_203,N_177);
nor U826 (N_826,N_152,N_188);
and U827 (N_827,N_149,N_347);
nor U828 (N_828,N_25,N_0);
nand U829 (N_829,N_273,N_26);
xnor U830 (N_830,N_120,N_362);
nand U831 (N_831,N_375,N_113);
xor U832 (N_832,N_137,N_58);
nand U833 (N_833,N_454,N_108);
and U834 (N_834,N_94,N_408);
nand U835 (N_835,N_390,N_460);
and U836 (N_836,N_116,N_219);
and U837 (N_837,N_399,N_328);
nor U838 (N_838,N_369,N_440);
nor U839 (N_839,N_410,N_52);
nor U840 (N_840,N_22,N_42);
xnor U841 (N_841,N_397,N_402);
nand U842 (N_842,N_363,N_131);
nor U843 (N_843,N_36,N_286);
nor U844 (N_844,N_195,N_330);
nor U845 (N_845,N_78,N_462);
nor U846 (N_846,N_228,N_317);
nor U847 (N_847,N_279,N_17);
nor U848 (N_848,N_397,N_118);
nor U849 (N_849,N_19,N_277);
nor U850 (N_850,N_491,N_295);
nor U851 (N_851,N_212,N_348);
nand U852 (N_852,N_222,N_197);
nor U853 (N_853,N_231,N_158);
and U854 (N_854,N_22,N_410);
nand U855 (N_855,N_102,N_407);
nor U856 (N_856,N_482,N_27);
xnor U857 (N_857,N_411,N_299);
or U858 (N_858,N_468,N_88);
and U859 (N_859,N_398,N_279);
nor U860 (N_860,N_242,N_419);
nand U861 (N_861,N_106,N_141);
nand U862 (N_862,N_291,N_243);
nor U863 (N_863,N_186,N_39);
nand U864 (N_864,N_314,N_327);
xor U865 (N_865,N_311,N_486);
nand U866 (N_866,N_290,N_408);
nand U867 (N_867,N_341,N_464);
and U868 (N_868,N_355,N_63);
or U869 (N_869,N_318,N_418);
nand U870 (N_870,N_388,N_219);
xor U871 (N_871,N_353,N_130);
and U872 (N_872,N_78,N_82);
xnor U873 (N_873,N_289,N_341);
nor U874 (N_874,N_162,N_367);
or U875 (N_875,N_292,N_425);
or U876 (N_876,N_265,N_494);
and U877 (N_877,N_455,N_167);
nand U878 (N_878,N_386,N_387);
nor U879 (N_879,N_175,N_363);
nor U880 (N_880,N_163,N_4);
and U881 (N_881,N_328,N_142);
nor U882 (N_882,N_422,N_73);
nand U883 (N_883,N_477,N_129);
nand U884 (N_884,N_181,N_108);
xnor U885 (N_885,N_173,N_311);
nand U886 (N_886,N_452,N_169);
or U887 (N_887,N_321,N_327);
nand U888 (N_888,N_363,N_341);
or U889 (N_889,N_449,N_238);
and U890 (N_890,N_127,N_70);
nand U891 (N_891,N_174,N_342);
and U892 (N_892,N_198,N_234);
nand U893 (N_893,N_232,N_60);
nor U894 (N_894,N_104,N_183);
nand U895 (N_895,N_491,N_220);
and U896 (N_896,N_153,N_69);
or U897 (N_897,N_216,N_274);
and U898 (N_898,N_193,N_361);
nand U899 (N_899,N_66,N_137);
xnor U900 (N_900,N_138,N_438);
nand U901 (N_901,N_41,N_87);
nor U902 (N_902,N_317,N_483);
nand U903 (N_903,N_369,N_180);
and U904 (N_904,N_38,N_320);
nor U905 (N_905,N_286,N_71);
nor U906 (N_906,N_349,N_97);
nor U907 (N_907,N_21,N_98);
nor U908 (N_908,N_445,N_447);
or U909 (N_909,N_458,N_252);
or U910 (N_910,N_324,N_480);
nor U911 (N_911,N_317,N_101);
nor U912 (N_912,N_373,N_448);
nand U913 (N_913,N_494,N_169);
and U914 (N_914,N_418,N_86);
xor U915 (N_915,N_22,N_278);
and U916 (N_916,N_284,N_350);
or U917 (N_917,N_238,N_205);
or U918 (N_918,N_83,N_123);
or U919 (N_919,N_139,N_36);
nor U920 (N_920,N_255,N_443);
and U921 (N_921,N_342,N_347);
or U922 (N_922,N_472,N_298);
and U923 (N_923,N_356,N_209);
and U924 (N_924,N_408,N_407);
or U925 (N_925,N_332,N_306);
or U926 (N_926,N_24,N_159);
nor U927 (N_927,N_324,N_112);
nor U928 (N_928,N_357,N_7);
and U929 (N_929,N_105,N_286);
xor U930 (N_930,N_135,N_137);
or U931 (N_931,N_347,N_145);
or U932 (N_932,N_320,N_259);
and U933 (N_933,N_271,N_492);
nand U934 (N_934,N_94,N_99);
nand U935 (N_935,N_212,N_294);
nor U936 (N_936,N_400,N_150);
xor U937 (N_937,N_44,N_95);
or U938 (N_938,N_327,N_272);
nand U939 (N_939,N_85,N_423);
or U940 (N_940,N_120,N_375);
or U941 (N_941,N_189,N_153);
nand U942 (N_942,N_495,N_437);
or U943 (N_943,N_133,N_407);
and U944 (N_944,N_278,N_177);
and U945 (N_945,N_281,N_311);
nor U946 (N_946,N_475,N_227);
nand U947 (N_947,N_294,N_141);
and U948 (N_948,N_178,N_69);
or U949 (N_949,N_452,N_477);
nand U950 (N_950,N_420,N_74);
or U951 (N_951,N_229,N_486);
nand U952 (N_952,N_323,N_238);
nand U953 (N_953,N_24,N_119);
and U954 (N_954,N_484,N_5);
xor U955 (N_955,N_5,N_197);
and U956 (N_956,N_279,N_393);
nor U957 (N_957,N_392,N_28);
or U958 (N_958,N_319,N_160);
nand U959 (N_959,N_431,N_459);
or U960 (N_960,N_240,N_58);
nor U961 (N_961,N_279,N_289);
xor U962 (N_962,N_268,N_117);
xor U963 (N_963,N_303,N_481);
nor U964 (N_964,N_218,N_90);
nand U965 (N_965,N_383,N_263);
nor U966 (N_966,N_115,N_481);
or U967 (N_967,N_236,N_215);
nand U968 (N_968,N_267,N_159);
and U969 (N_969,N_476,N_454);
nand U970 (N_970,N_441,N_403);
or U971 (N_971,N_0,N_356);
nor U972 (N_972,N_157,N_471);
and U973 (N_973,N_48,N_358);
nor U974 (N_974,N_46,N_289);
xnor U975 (N_975,N_141,N_131);
nand U976 (N_976,N_6,N_178);
xor U977 (N_977,N_359,N_296);
or U978 (N_978,N_332,N_337);
nand U979 (N_979,N_235,N_136);
and U980 (N_980,N_10,N_14);
or U981 (N_981,N_134,N_246);
nor U982 (N_982,N_393,N_5);
or U983 (N_983,N_160,N_477);
nand U984 (N_984,N_431,N_96);
or U985 (N_985,N_140,N_486);
and U986 (N_986,N_98,N_263);
or U987 (N_987,N_238,N_331);
xnor U988 (N_988,N_195,N_96);
nor U989 (N_989,N_38,N_452);
or U990 (N_990,N_224,N_96);
and U991 (N_991,N_414,N_290);
xor U992 (N_992,N_394,N_470);
nand U993 (N_993,N_145,N_66);
or U994 (N_994,N_339,N_70);
xor U995 (N_995,N_446,N_400);
nand U996 (N_996,N_465,N_168);
or U997 (N_997,N_216,N_439);
nor U998 (N_998,N_118,N_279);
or U999 (N_999,N_440,N_144);
nand U1000 (N_1000,N_540,N_635);
or U1001 (N_1001,N_831,N_763);
or U1002 (N_1002,N_968,N_526);
nor U1003 (N_1003,N_743,N_620);
nor U1004 (N_1004,N_863,N_917);
nor U1005 (N_1005,N_536,N_695);
nand U1006 (N_1006,N_762,N_508);
xnor U1007 (N_1007,N_975,N_898);
or U1008 (N_1008,N_881,N_836);
and U1009 (N_1009,N_712,N_608);
nand U1010 (N_1010,N_846,N_929);
and U1011 (N_1011,N_710,N_668);
or U1012 (N_1012,N_781,N_703);
nor U1013 (N_1013,N_765,N_741);
or U1014 (N_1014,N_871,N_532);
and U1015 (N_1015,N_740,N_691);
xnor U1016 (N_1016,N_570,N_979);
and U1017 (N_1017,N_517,N_921);
nand U1018 (N_1018,N_764,N_788);
and U1019 (N_1019,N_679,N_773);
and U1020 (N_1020,N_617,N_708);
xor U1021 (N_1021,N_623,N_817);
nor U1022 (N_1022,N_546,N_868);
or U1023 (N_1023,N_520,N_660);
nand U1024 (N_1024,N_512,N_803);
xnor U1025 (N_1025,N_847,N_566);
and U1026 (N_1026,N_916,N_530);
nand U1027 (N_1027,N_638,N_656);
nand U1028 (N_1028,N_553,N_939);
nand U1029 (N_1029,N_932,N_991);
nand U1030 (N_1030,N_922,N_580);
xor U1031 (N_1031,N_816,N_509);
and U1032 (N_1032,N_924,N_682);
nand U1033 (N_1033,N_661,N_720);
nand U1034 (N_1034,N_876,N_902);
nor U1035 (N_1035,N_958,N_533);
or U1036 (N_1036,N_890,N_875);
nor U1037 (N_1037,N_562,N_505);
nand U1038 (N_1038,N_966,N_676);
nor U1039 (N_1039,N_577,N_967);
and U1040 (N_1040,N_605,N_930);
and U1041 (N_1041,N_907,N_733);
or U1042 (N_1042,N_986,N_769);
nor U1043 (N_1043,N_529,N_624);
nor U1044 (N_1044,N_995,N_571);
and U1045 (N_1045,N_514,N_531);
nor U1046 (N_1046,N_787,N_798);
nor U1047 (N_1047,N_644,N_856);
nand U1048 (N_1048,N_851,N_853);
nand U1049 (N_1049,N_511,N_633);
and U1050 (N_1050,N_686,N_515);
nor U1051 (N_1051,N_632,N_665);
nand U1052 (N_1052,N_651,N_611);
nor U1053 (N_1053,N_889,N_750);
or U1054 (N_1054,N_774,N_565);
and U1055 (N_1055,N_675,N_945);
or U1056 (N_1056,N_688,N_911);
nor U1057 (N_1057,N_602,N_835);
xnor U1058 (N_1058,N_622,N_724);
xnor U1059 (N_1059,N_523,N_884);
and U1060 (N_1060,N_826,N_642);
and U1061 (N_1061,N_908,N_513);
or U1062 (N_1062,N_866,N_783);
nand U1063 (N_1063,N_507,N_717);
xor U1064 (N_1064,N_669,N_699);
and U1065 (N_1065,N_951,N_581);
and U1066 (N_1066,N_680,N_522);
or U1067 (N_1067,N_504,N_645);
nand U1068 (N_1068,N_542,N_521);
or U1069 (N_1069,N_827,N_718);
nor U1070 (N_1070,N_959,N_525);
nor U1071 (N_1071,N_524,N_653);
xor U1072 (N_1072,N_678,N_906);
or U1073 (N_1073,N_709,N_796);
and U1074 (N_1074,N_814,N_641);
or U1075 (N_1075,N_585,N_888);
nor U1076 (N_1076,N_983,N_510);
nor U1077 (N_1077,N_934,N_528);
xnor U1078 (N_1078,N_631,N_684);
nand U1079 (N_1079,N_747,N_961);
nor U1080 (N_1080,N_812,N_857);
nand U1081 (N_1081,N_713,N_603);
and U1082 (N_1082,N_606,N_912);
nor U1083 (N_1083,N_715,N_616);
xnor U1084 (N_1084,N_830,N_595);
and U1085 (N_1085,N_649,N_841);
and U1086 (N_1086,N_655,N_793);
nor U1087 (N_1087,N_972,N_833);
nand U1088 (N_1088,N_599,N_809);
nand U1089 (N_1089,N_941,N_707);
nand U1090 (N_1090,N_770,N_701);
or U1091 (N_1091,N_759,N_555);
nor U1092 (N_1092,N_625,N_819);
nor U1093 (N_1093,N_636,N_516);
xor U1094 (N_1094,N_936,N_914);
nor U1095 (N_1095,N_801,N_752);
and U1096 (N_1096,N_706,N_643);
nor U1097 (N_1097,N_618,N_799);
nand U1098 (N_1098,N_903,N_737);
nand U1099 (N_1099,N_782,N_896);
and U1100 (N_1100,N_760,N_698);
nor U1101 (N_1101,N_594,N_662);
nand U1102 (N_1102,N_503,N_893);
nor U1103 (N_1103,N_877,N_865);
nor U1104 (N_1104,N_766,N_705);
and U1105 (N_1105,N_744,N_987);
nor U1106 (N_1106,N_811,N_904);
or U1107 (N_1107,N_742,N_858);
nor U1108 (N_1108,N_558,N_820);
xnor U1109 (N_1109,N_702,N_692);
or U1110 (N_1110,N_552,N_854);
and U1111 (N_1111,N_985,N_861);
nor U1112 (N_1112,N_685,N_956);
and U1113 (N_1113,N_776,N_704);
nor U1114 (N_1114,N_937,N_823);
nand U1115 (N_1115,N_746,N_767);
nor U1116 (N_1116,N_739,N_790);
or U1117 (N_1117,N_664,N_593);
nand U1118 (N_1118,N_813,N_810);
xnor U1119 (N_1119,N_614,N_728);
xnor U1120 (N_1120,N_549,N_758);
or U1121 (N_1121,N_550,N_980);
and U1122 (N_1122,N_895,N_990);
xor U1123 (N_1123,N_547,N_970);
or U1124 (N_1124,N_953,N_648);
or U1125 (N_1125,N_748,N_537);
and U1126 (N_1126,N_805,N_640);
xnor U1127 (N_1127,N_761,N_591);
nand U1128 (N_1128,N_829,N_832);
or U1129 (N_1129,N_650,N_940);
nand U1130 (N_1130,N_926,N_538);
or U1131 (N_1131,N_974,N_501);
xnor U1132 (N_1132,N_629,N_824);
nand U1133 (N_1133,N_971,N_527);
nor U1134 (N_1134,N_800,N_900);
nor U1135 (N_1135,N_757,N_697);
and U1136 (N_1136,N_943,N_613);
and U1137 (N_1137,N_657,N_949);
and U1138 (N_1138,N_780,N_574);
and U1139 (N_1139,N_828,N_545);
or U1140 (N_1140,N_789,N_541);
and U1141 (N_1141,N_573,N_543);
and U1142 (N_1142,N_879,N_778);
xnor U1143 (N_1143,N_915,N_753);
nor U1144 (N_1144,N_821,N_909);
or U1145 (N_1145,N_962,N_725);
or U1146 (N_1146,N_654,N_913);
nand U1147 (N_1147,N_882,N_860);
xor U1148 (N_1148,N_597,N_659);
or U1149 (N_1149,N_583,N_869);
nor U1150 (N_1150,N_897,N_696);
or U1151 (N_1151,N_804,N_872);
nand U1152 (N_1152,N_716,N_982);
nor U1153 (N_1153,N_840,N_590);
and U1154 (N_1154,N_600,N_878);
or U1155 (N_1155,N_977,N_518);
or U1156 (N_1156,N_992,N_815);
xor U1157 (N_1157,N_891,N_948);
xnor U1158 (N_1158,N_568,N_969);
and U1159 (N_1159,N_864,N_619);
or U1160 (N_1160,N_919,N_610);
nand U1161 (N_1161,N_579,N_838);
and U1162 (N_1162,N_771,N_681);
nor U1163 (N_1163,N_626,N_918);
nor U1164 (N_1164,N_554,N_870);
nor U1165 (N_1165,N_960,N_777);
nand U1166 (N_1166,N_749,N_519);
nor U1167 (N_1167,N_775,N_925);
or U1168 (N_1168,N_721,N_938);
and U1169 (N_1169,N_957,N_848);
or U1170 (N_1170,N_779,N_690);
and U1171 (N_1171,N_963,N_892);
or U1172 (N_1172,N_751,N_947);
or U1173 (N_1173,N_647,N_946);
or U1174 (N_1174,N_923,N_575);
nand U1175 (N_1175,N_792,N_673);
or U1176 (N_1176,N_736,N_576);
nor U1177 (N_1177,N_920,N_630);
or U1178 (N_1178,N_700,N_842);
and U1179 (N_1179,N_785,N_582);
and U1180 (N_1180,N_955,N_663);
nand U1181 (N_1181,N_551,N_535);
nand U1182 (N_1182,N_874,N_612);
nand U1183 (N_1183,N_500,N_671);
or U1184 (N_1184,N_734,N_901);
nor U1185 (N_1185,N_844,N_694);
and U1186 (N_1186,N_639,N_996);
or U1187 (N_1187,N_731,N_927);
nor U1188 (N_1188,N_534,N_997);
or U1189 (N_1189,N_586,N_797);
nand U1190 (N_1190,N_652,N_693);
or U1191 (N_1191,N_572,N_806);
xor U1192 (N_1192,N_818,N_672);
nor U1193 (N_1193,N_984,N_714);
nand U1194 (N_1194,N_674,N_588);
or U1195 (N_1195,N_850,N_578);
and U1196 (N_1196,N_589,N_502);
or U1197 (N_1197,N_998,N_506);
and U1198 (N_1198,N_999,N_628);
and U1199 (N_1199,N_564,N_935);
or U1200 (N_1200,N_719,N_729);
and U1201 (N_1201,N_592,N_730);
nor U1202 (N_1202,N_786,N_886);
nand U1203 (N_1203,N_784,N_822);
nand U1204 (N_1204,N_942,N_965);
or U1205 (N_1205,N_883,N_839);
xor U1206 (N_1206,N_726,N_768);
nor U1207 (N_1207,N_584,N_899);
and U1208 (N_1208,N_607,N_852);
or U1209 (N_1209,N_973,N_905);
and U1210 (N_1210,N_993,N_756);
xnor U1211 (N_1211,N_834,N_802);
and U1212 (N_1212,N_735,N_807);
xor U1213 (N_1213,N_738,N_976);
xor U1214 (N_1214,N_637,N_931);
nor U1215 (N_1215,N_539,N_873);
nand U1216 (N_1216,N_933,N_952);
nor U1217 (N_1217,N_557,N_754);
or U1218 (N_1218,N_964,N_677);
nand U1219 (N_1219,N_880,N_569);
and U1220 (N_1220,N_627,N_849);
or U1221 (N_1221,N_689,N_621);
nor U1222 (N_1222,N_544,N_825);
or U1223 (N_1223,N_587,N_604);
xor U1224 (N_1224,N_683,N_855);
nand U1225 (N_1225,N_596,N_843);
and U1226 (N_1226,N_609,N_887);
or U1227 (N_1227,N_772,N_556);
or U1228 (N_1228,N_615,N_687);
nor U1229 (N_1229,N_988,N_601);
nor U1230 (N_1230,N_646,N_561);
nand U1231 (N_1231,N_859,N_954);
or U1232 (N_1232,N_755,N_666);
nor U1233 (N_1233,N_794,N_791);
or U1234 (N_1234,N_745,N_723);
nor U1235 (N_1235,N_867,N_658);
or U1236 (N_1236,N_978,N_670);
nor U1237 (N_1237,N_808,N_567);
nand U1238 (N_1238,N_928,N_981);
nand U1239 (N_1239,N_837,N_667);
or U1240 (N_1240,N_598,N_950);
nand U1241 (N_1241,N_862,N_944);
or U1242 (N_1242,N_727,N_711);
nor U1243 (N_1243,N_894,N_795);
and U1244 (N_1244,N_634,N_563);
nor U1245 (N_1245,N_885,N_722);
nand U1246 (N_1246,N_994,N_845);
nand U1247 (N_1247,N_560,N_548);
or U1248 (N_1248,N_732,N_989);
nor U1249 (N_1249,N_559,N_910);
or U1250 (N_1250,N_779,N_933);
xor U1251 (N_1251,N_679,N_532);
nor U1252 (N_1252,N_600,N_665);
nor U1253 (N_1253,N_896,N_673);
nor U1254 (N_1254,N_964,N_841);
nor U1255 (N_1255,N_896,N_915);
nor U1256 (N_1256,N_966,N_635);
or U1257 (N_1257,N_632,N_775);
nand U1258 (N_1258,N_628,N_680);
or U1259 (N_1259,N_697,N_881);
nor U1260 (N_1260,N_887,N_955);
or U1261 (N_1261,N_755,N_650);
and U1262 (N_1262,N_598,N_571);
nor U1263 (N_1263,N_802,N_983);
or U1264 (N_1264,N_596,N_674);
nor U1265 (N_1265,N_655,N_811);
or U1266 (N_1266,N_586,N_750);
and U1267 (N_1267,N_510,N_618);
nor U1268 (N_1268,N_678,N_803);
or U1269 (N_1269,N_633,N_738);
and U1270 (N_1270,N_637,N_731);
or U1271 (N_1271,N_815,N_543);
or U1272 (N_1272,N_843,N_848);
nand U1273 (N_1273,N_897,N_963);
nand U1274 (N_1274,N_613,N_520);
nand U1275 (N_1275,N_700,N_557);
and U1276 (N_1276,N_506,N_620);
nor U1277 (N_1277,N_913,N_934);
nor U1278 (N_1278,N_654,N_714);
nand U1279 (N_1279,N_717,N_769);
nand U1280 (N_1280,N_721,N_635);
nand U1281 (N_1281,N_513,N_547);
nand U1282 (N_1282,N_938,N_672);
or U1283 (N_1283,N_860,N_522);
or U1284 (N_1284,N_781,N_607);
or U1285 (N_1285,N_631,N_960);
or U1286 (N_1286,N_539,N_604);
and U1287 (N_1287,N_903,N_842);
and U1288 (N_1288,N_559,N_506);
or U1289 (N_1289,N_751,N_861);
nand U1290 (N_1290,N_527,N_714);
xnor U1291 (N_1291,N_834,N_995);
xor U1292 (N_1292,N_630,N_841);
nand U1293 (N_1293,N_809,N_764);
and U1294 (N_1294,N_740,N_905);
or U1295 (N_1295,N_875,N_755);
or U1296 (N_1296,N_993,N_955);
or U1297 (N_1297,N_842,N_722);
nor U1298 (N_1298,N_515,N_865);
and U1299 (N_1299,N_600,N_618);
or U1300 (N_1300,N_939,N_589);
xor U1301 (N_1301,N_693,N_615);
or U1302 (N_1302,N_778,N_931);
or U1303 (N_1303,N_829,N_503);
or U1304 (N_1304,N_646,N_675);
or U1305 (N_1305,N_628,N_715);
nor U1306 (N_1306,N_828,N_723);
and U1307 (N_1307,N_610,N_753);
nand U1308 (N_1308,N_534,N_889);
nand U1309 (N_1309,N_844,N_995);
and U1310 (N_1310,N_848,N_891);
nand U1311 (N_1311,N_609,N_961);
nor U1312 (N_1312,N_901,N_626);
and U1313 (N_1313,N_505,N_759);
nor U1314 (N_1314,N_631,N_727);
xnor U1315 (N_1315,N_689,N_821);
or U1316 (N_1316,N_505,N_957);
or U1317 (N_1317,N_752,N_526);
nand U1318 (N_1318,N_778,N_648);
nand U1319 (N_1319,N_570,N_785);
nand U1320 (N_1320,N_904,N_639);
nor U1321 (N_1321,N_545,N_689);
and U1322 (N_1322,N_558,N_556);
or U1323 (N_1323,N_918,N_850);
and U1324 (N_1324,N_597,N_595);
xor U1325 (N_1325,N_638,N_814);
or U1326 (N_1326,N_991,N_752);
nor U1327 (N_1327,N_714,N_947);
nand U1328 (N_1328,N_866,N_679);
and U1329 (N_1329,N_823,N_908);
nand U1330 (N_1330,N_560,N_771);
and U1331 (N_1331,N_717,N_927);
nor U1332 (N_1332,N_870,N_562);
nor U1333 (N_1333,N_626,N_910);
nor U1334 (N_1334,N_674,N_694);
nor U1335 (N_1335,N_529,N_894);
and U1336 (N_1336,N_511,N_868);
nor U1337 (N_1337,N_525,N_801);
or U1338 (N_1338,N_936,N_532);
nand U1339 (N_1339,N_868,N_550);
or U1340 (N_1340,N_770,N_983);
or U1341 (N_1341,N_683,N_768);
nand U1342 (N_1342,N_585,N_672);
nor U1343 (N_1343,N_669,N_526);
nor U1344 (N_1344,N_616,N_627);
and U1345 (N_1345,N_530,N_521);
xor U1346 (N_1346,N_608,N_949);
and U1347 (N_1347,N_887,N_890);
nand U1348 (N_1348,N_857,N_829);
xor U1349 (N_1349,N_853,N_605);
and U1350 (N_1350,N_992,N_685);
or U1351 (N_1351,N_630,N_632);
nor U1352 (N_1352,N_506,N_845);
nand U1353 (N_1353,N_782,N_730);
nand U1354 (N_1354,N_956,N_923);
and U1355 (N_1355,N_917,N_670);
xnor U1356 (N_1356,N_845,N_663);
and U1357 (N_1357,N_878,N_883);
nor U1358 (N_1358,N_664,N_527);
nand U1359 (N_1359,N_722,N_990);
or U1360 (N_1360,N_811,N_990);
or U1361 (N_1361,N_858,N_969);
nor U1362 (N_1362,N_633,N_652);
nor U1363 (N_1363,N_838,N_731);
nand U1364 (N_1364,N_732,N_513);
nor U1365 (N_1365,N_882,N_729);
nor U1366 (N_1366,N_671,N_865);
nor U1367 (N_1367,N_603,N_717);
nand U1368 (N_1368,N_801,N_603);
or U1369 (N_1369,N_512,N_711);
and U1370 (N_1370,N_625,N_592);
and U1371 (N_1371,N_992,N_698);
or U1372 (N_1372,N_954,N_632);
nor U1373 (N_1373,N_863,N_526);
or U1374 (N_1374,N_710,N_705);
nand U1375 (N_1375,N_966,N_792);
nor U1376 (N_1376,N_969,N_903);
and U1377 (N_1377,N_636,N_613);
nand U1378 (N_1378,N_714,N_511);
or U1379 (N_1379,N_776,N_878);
and U1380 (N_1380,N_765,N_980);
nand U1381 (N_1381,N_791,N_568);
or U1382 (N_1382,N_566,N_763);
xnor U1383 (N_1383,N_901,N_754);
xnor U1384 (N_1384,N_596,N_500);
nand U1385 (N_1385,N_869,N_761);
nand U1386 (N_1386,N_689,N_627);
nor U1387 (N_1387,N_991,N_668);
nand U1388 (N_1388,N_866,N_621);
or U1389 (N_1389,N_673,N_697);
and U1390 (N_1390,N_843,N_890);
nand U1391 (N_1391,N_806,N_536);
and U1392 (N_1392,N_657,N_548);
nor U1393 (N_1393,N_733,N_502);
nor U1394 (N_1394,N_677,N_799);
nor U1395 (N_1395,N_515,N_772);
nand U1396 (N_1396,N_624,N_699);
or U1397 (N_1397,N_536,N_802);
or U1398 (N_1398,N_872,N_815);
nand U1399 (N_1399,N_875,N_689);
nand U1400 (N_1400,N_855,N_540);
nand U1401 (N_1401,N_868,N_841);
nor U1402 (N_1402,N_713,N_872);
and U1403 (N_1403,N_571,N_681);
and U1404 (N_1404,N_903,N_775);
and U1405 (N_1405,N_645,N_614);
and U1406 (N_1406,N_915,N_520);
and U1407 (N_1407,N_756,N_580);
nand U1408 (N_1408,N_739,N_768);
nand U1409 (N_1409,N_936,N_771);
or U1410 (N_1410,N_649,N_855);
nor U1411 (N_1411,N_711,N_783);
nor U1412 (N_1412,N_551,N_529);
or U1413 (N_1413,N_728,N_935);
or U1414 (N_1414,N_881,N_589);
nor U1415 (N_1415,N_725,N_547);
nand U1416 (N_1416,N_893,N_748);
nand U1417 (N_1417,N_854,N_950);
or U1418 (N_1418,N_703,N_677);
and U1419 (N_1419,N_915,N_937);
xor U1420 (N_1420,N_855,N_550);
nor U1421 (N_1421,N_583,N_929);
nand U1422 (N_1422,N_612,N_619);
or U1423 (N_1423,N_574,N_822);
nand U1424 (N_1424,N_661,N_745);
or U1425 (N_1425,N_747,N_582);
nor U1426 (N_1426,N_561,N_744);
nand U1427 (N_1427,N_649,N_506);
xnor U1428 (N_1428,N_606,N_643);
and U1429 (N_1429,N_720,N_786);
or U1430 (N_1430,N_576,N_844);
nor U1431 (N_1431,N_642,N_843);
nand U1432 (N_1432,N_921,N_607);
nor U1433 (N_1433,N_893,N_974);
nand U1434 (N_1434,N_797,N_987);
xor U1435 (N_1435,N_573,N_557);
or U1436 (N_1436,N_906,N_656);
nand U1437 (N_1437,N_661,N_531);
and U1438 (N_1438,N_797,N_750);
nand U1439 (N_1439,N_834,N_906);
xor U1440 (N_1440,N_963,N_720);
or U1441 (N_1441,N_941,N_971);
nand U1442 (N_1442,N_867,N_799);
or U1443 (N_1443,N_502,N_907);
nor U1444 (N_1444,N_874,N_616);
nand U1445 (N_1445,N_937,N_979);
and U1446 (N_1446,N_599,N_844);
nand U1447 (N_1447,N_549,N_909);
or U1448 (N_1448,N_547,N_720);
and U1449 (N_1449,N_773,N_637);
nand U1450 (N_1450,N_885,N_582);
or U1451 (N_1451,N_641,N_531);
xnor U1452 (N_1452,N_560,N_848);
nand U1453 (N_1453,N_974,N_920);
and U1454 (N_1454,N_815,N_600);
nor U1455 (N_1455,N_618,N_752);
and U1456 (N_1456,N_825,N_851);
or U1457 (N_1457,N_568,N_810);
nor U1458 (N_1458,N_983,N_724);
and U1459 (N_1459,N_724,N_985);
xor U1460 (N_1460,N_766,N_951);
xor U1461 (N_1461,N_966,N_623);
nand U1462 (N_1462,N_737,N_849);
or U1463 (N_1463,N_867,N_869);
nand U1464 (N_1464,N_775,N_697);
or U1465 (N_1465,N_797,N_788);
nor U1466 (N_1466,N_770,N_750);
or U1467 (N_1467,N_682,N_575);
xnor U1468 (N_1468,N_719,N_765);
nand U1469 (N_1469,N_505,N_688);
nand U1470 (N_1470,N_957,N_506);
or U1471 (N_1471,N_588,N_644);
and U1472 (N_1472,N_586,N_659);
nand U1473 (N_1473,N_620,N_733);
xor U1474 (N_1474,N_819,N_832);
nor U1475 (N_1475,N_946,N_676);
or U1476 (N_1476,N_587,N_822);
nor U1477 (N_1477,N_791,N_668);
xnor U1478 (N_1478,N_889,N_724);
or U1479 (N_1479,N_602,N_844);
or U1480 (N_1480,N_654,N_931);
nand U1481 (N_1481,N_922,N_873);
or U1482 (N_1482,N_879,N_860);
nor U1483 (N_1483,N_912,N_988);
or U1484 (N_1484,N_692,N_631);
xor U1485 (N_1485,N_803,N_916);
nand U1486 (N_1486,N_689,N_829);
or U1487 (N_1487,N_683,N_818);
nand U1488 (N_1488,N_656,N_755);
and U1489 (N_1489,N_676,N_803);
xnor U1490 (N_1490,N_838,N_583);
xnor U1491 (N_1491,N_904,N_980);
nand U1492 (N_1492,N_572,N_800);
or U1493 (N_1493,N_617,N_974);
nor U1494 (N_1494,N_671,N_627);
nor U1495 (N_1495,N_799,N_657);
or U1496 (N_1496,N_668,N_625);
and U1497 (N_1497,N_626,N_578);
and U1498 (N_1498,N_824,N_953);
nand U1499 (N_1499,N_642,N_897);
or U1500 (N_1500,N_1209,N_1175);
and U1501 (N_1501,N_1060,N_1169);
or U1502 (N_1502,N_1413,N_1365);
and U1503 (N_1503,N_1054,N_1383);
and U1504 (N_1504,N_1113,N_1447);
nand U1505 (N_1505,N_1286,N_1010);
nand U1506 (N_1506,N_1048,N_1475);
or U1507 (N_1507,N_1129,N_1180);
or U1508 (N_1508,N_1190,N_1137);
and U1509 (N_1509,N_1319,N_1377);
nand U1510 (N_1510,N_1170,N_1229);
xnor U1511 (N_1511,N_1236,N_1000);
or U1512 (N_1512,N_1403,N_1157);
nor U1513 (N_1513,N_1486,N_1003);
xor U1514 (N_1514,N_1158,N_1015);
and U1515 (N_1515,N_1358,N_1408);
nand U1516 (N_1516,N_1259,N_1075);
xnor U1517 (N_1517,N_1212,N_1004);
and U1518 (N_1518,N_1093,N_1380);
and U1519 (N_1519,N_1355,N_1109);
or U1520 (N_1520,N_1061,N_1201);
nor U1521 (N_1521,N_1441,N_1466);
nor U1522 (N_1522,N_1214,N_1440);
nand U1523 (N_1523,N_1059,N_1041);
nor U1524 (N_1524,N_1361,N_1146);
nor U1525 (N_1525,N_1472,N_1404);
nor U1526 (N_1526,N_1057,N_1386);
nand U1527 (N_1527,N_1350,N_1186);
and U1528 (N_1528,N_1068,N_1345);
nor U1529 (N_1529,N_1240,N_1025);
or U1530 (N_1530,N_1388,N_1040);
xnor U1531 (N_1531,N_1016,N_1461);
xnor U1532 (N_1532,N_1489,N_1179);
nand U1533 (N_1533,N_1399,N_1200);
nor U1534 (N_1534,N_1116,N_1250);
and U1535 (N_1535,N_1262,N_1073);
or U1536 (N_1536,N_1477,N_1215);
nor U1537 (N_1537,N_1246,N_1370);
or U1538 (N_1538,N_1375,N_1219);
nand U1539 (N_1539,N_1470,N_1457);
nor U1540 (N_1540,N_1352,N_1342);
or U1541 (N_1541,N_1474,N_1035);
and U1542 (N_1542,N_1287,N_1464);
nand U1543 (N_1543,N_1478,N_1136);
and U1544 (N_1544,N_1120,N_1174);
xnor U1545 (N_1545,N_1285,N_1424);
or U1546 (N_1546,N_1481,N_1418);
nand U1547 (N_1547,N_1013,N_1428);
and U1548 (N_1548,N_1275,N_1230);
nor U1549 (N_1549,N_1426,N_1260);
nor U1550 (N_1550,N_1042,N_1191);
or U1551 (N_1551,N_1276,N_1034);
nand U1552 (N_1552,N_1297,N_1427);
or U1553 (N_1553,N_1449,N_1458);
and U1554 (N_1554,N_1288,N_1298);
or U1555 (N_1555,N_1320,N_1098);
xor U1556 (N_1556,N_1419,N_1198);
nand U1557 (N_1557,N_1227,N_1266);
nor U1558 (N_1558,N_1391,N_1206);
nand U1559 (N_1559,N_1484,N_1197);
nor U1560 (N_1560,N_1001,N_1125);
or U1561 (N_1561,N_1008,N_1301);
and U1562 (N_1562,N_1291,N_1066);
xnor U1563 (N_1563,N_1397,N_1467);
or U1564 (N_1564,N_1224,N_1228);
nand U1565 (N_1565,N_1353,N_1226);
and U1566 (N_1566,N_1487,N_1141);
and U1567 (N_1567,N_1492,N_1398);
or U1568 (N_1568,N_1064,N_1092);
or U1569 (N_1569,N_1460,N_1119);
nand U1570 (N_1570,N_1142,N_1165);
and U1571 (N_1571,N_1071,N_1412);
and U1572 (N_1572,N_1485,N_1134);
nand U1573 (N_1573,N_1394,N_1382);
or U1574 (N_1574,N_1002,N_1251);
nor U1575 (N_1575,N_1346,N_1312);
nand U1576 (N_1576,N_1306,N_1210);
or U1577 (N_1577,N_1029,N_1452);
nand U1578 (N_1578,N_1363,N_1314);
and U1579 (N_1579,N_1095,N_1011);
nand U1580 (N_1580,N_1498,N_1339);
xnor U1581 (N_1581,N_1154,N_1017);
nor U1582 (N_1582,N_1147,N_1400);
or U1583 (N_1583,N_1300,N_1128);
or U1584 (N_1584,N_1321,N_1032);
nand U1585 (N_1585,N_1131,N_1362);
or U1586 (N_1586,N_1330,N_1133);
and U1587 (N_1587,N_1315,N_1148);
or U1588 (N_1588,N_1305,N_1244);
nand U1589 (N_1589,N_1205,N_1279);
or U1590 (N_1590,N_1089,N_1030);
or U1591 (N_1591,N_1065,N_1039);
nor U1592 (N_1592,N_1491,N_1181);
nand U1593 (N_1593,N_1406,N_1463);
and U1594 (N_1594,N_1122,N_1446);
nand U1595 (N_1595,N_1316,N_1199);
or U1596 (N_1596,N_1465,N_1036);
nor U1597 (N_1597,N_1414,N_1367);
and U1598 (N_1598,N_1033,N_1145);
nand U1599 (N_1599,N_1257,N_1031);
nor U1600 (N_1600,N_1220,N_1493);
or U1601 (N_1601,N_1332,N_1431);
and U1602 (N_1602,N_1234,N_1153);
nand U1603 (N_1603,N_1333,N_1409);
nor U1604 (N_1604,N_1348,N_1407);
or U1605 (N_1605,N_1074,N_1046);
nand U1606 (N_1606,N_1326,N_1435);
xnor U1607 (N_1607,N_1282,N_1241);
xnor U1608 (N_1608,N_1273,N_1423);
nand U1609 (N_1609,N_1469,N_1233);
nand U1610 (N_1610,N_1182,N_1410);
and U1611 (N_1611,N_1106,N_1294);
and U1612 (N_1612,N_1138,N_1052);
and U1613 (N_1613,N_1176,N_1225);
nand U1614 (N_1614,N_1083,N_1221);
or U1615 (N_1615,N_1497,N_1256);
and U1616 (N_1616,N_1480,N_1313);
or U1617 (N_1617,N_1390,N_1351);
nor U1618 (N_1618,N_1270,N_1012);
and U1619 (N_1619,N_1265,N_1347);
nand U1620 (N_1620,N_1028,N_1184);
nand U1621 (N_1621,N_1223,N_1368);
nand U1622 (N_1622,N_1045,N_1334);
xnor U1623 (N_1623,N_1299,N_1378);
nor U1624 (N_1624,N_1005,N_1438);
or U1625 (N_1625,N_1395,N_1108);
nand U1626 (N_1626,N_1268,N_1100);
nand U1627 (N_1627,N_1443,N_1047);
and U1628 (N_1628,N_1281,N_1082);
nor U1629 (N_1629,N_1055,N_1254);
nor U1630 (N_1630,N_1231,N_1448);
and U1631 (N_1631,N_1417,N_1335);
and U1632 (N_1632,N_1252,N_1295);
and U1633 (N_1633,N_1196,N_1278);
nand U1634 (N_1634,N_1471,N_1127);
nor U1635 (N_1635,N_1014,N_1248);
and U1636 (N_1636,N_1193,N_1022);
xor U1637 (N_1637,N_1387,N_1393);
and U1638 (N_1638,N_1405,N_1177);
or U1639 (N_1639,N_1238,N_1150);
or U1640 (N_1640,N_1097,N_1101);
nand U1641 (N_1641,N_1344,N_1139);
nand U1642 (N_1642,N_1499,N_1296);
and U1643 (N_1643,N_1364,N_1271);
or U1644 (N_1644,N_1038,N_1253);
and U1645 (N_1645,N_1118,N_1372);
nand U1646 (N_1646,N_1303,N_1077);
or U1647 (N_1647,N_1178,N_1021);
nand U1648 (N_1648,N_1324,N_1144);
nor U1649 (N_1649,N_1123,N_1433);
or U1650 (N_1650,N_1267,N_1293);
nor U1651 (N_1651,N_1356,N_1085);
xor U1652 (N_1652,N_1043,N_1149);
nand U1653 (N_1653,N_1289,N_1105);
nand U1654 (N_1654,N_1337,N_1135);
and U1655 (N_1655,N_1121,N_1483);
and U1656 (N_1656,N_1366,N_1401);
and U1657 (N_1657,N_1284,N_1421);
or U1658 (N_1658,N_1189,N_1072);
and U1659 (N_1659,N_1202,N_1292);
nand U1660 (N_1660,N_1094,N_1331);
and U1661 (N_1661,N_1102,N_1204);
nor U1662 (N_1662,N_1430,N_1090);
nor U1663 (N_1663,N_1099,N_1308);
nand U1664 (N_1664,N_1024,N_1392);
nand U1665 (N_1665,N_1218,N_1425);
nand U1666 (N_1666,N_1080,N_1389);
or U1667 (N_1667,N_1103,N_1341);
nor U1668 (N_1668,N_1451,N_1185);
or U1669 (N_1669,N_1213,N_1087);
nor U1670 (N_1670,N_1274,N_1084);
and U1671 (N_1671,N_1156,N_1217);
or U1672 (N_1672,N_1247,N_1336);
or U1673 (N_1673,N_1049,N_1479);
nand U1674 (N_1674,N_1162,N_1143);
nor U1675 (N_1675,N_1402,N_1462);
and U1676 (N_1676,N_1371,N_1056);
nand U1677 (N_1677,N_1115,N_1232);
nand U1678 (N_1678,N_1163,N_1450);
nand U1679 (N_1679,N_1058,N_1086);
or U1680 (N_1680,N_1338,N_1183);
nand U1681 (N_1681,N_1429,N_1290);
or U1682 (N_1682,N_1208,N_1468);
nand U1683 (N_1683,N_1456,N_1311);
or U1684 (N_1684,N_1126,N_1173);
nand U1685 (N_1685,N_1384,N_1019);
nand U1686 (N_1686,N_1051,N_1194);
or U1687 (N_1687,N_1327,N_1053);
or U1688 (N_1688,N_1155,N_1340);
nand U1689 (N_1689,N_1070,N_1396);
and U1690 (N_1690,N_1195,N_1369);
nand U1691 (N_1691,N_1473,N_1020);
nor U1692 (N_1692,N_1187,N_1455);
nand U1693 (N_1693,N_1318,N_1374);
and U1694 (N_1694,N_1111,N_1310);
and U1695 (N_1695,N_1302,N_1096);
and U1696 (N_1696,N_1317,N_1476);
and U1697 (N_1697,N_1420,N_1140);
nor U1698 (N_1698,N_1454,N_1280);
or U1699 (N_1699,N_1117,N_1006);
xnor U1700 (N_1700,N_1037,N_1415);
nand U1701 (N_1701,N_1063,N_1283);
and U1702 (N_1702,N_1385,N_1263);
and U1703 (N_1703,N_1027,N_1050);
nor U1704 (N_1704,N_1081,N_1411);
nand U1705 (N_1705,N_1130,N_1249);
and U1706 (N_1706,N_1151,N_1009);
or U1707 (N_1707,N_1264,N_1494);
nand U1708 (N_1708,N_1436,N_1329);
or U1709 (N_1709,N_1359,N_1132);
nor U1710 (N_1710,N_1437,N_1067);
nor U1711 (N_1711,N_1323,N_1349);
xnor U1712 (N_1712,N_1432,N_1459);
nor U1713 (N_1713,N_1360,N_1442);
or U1714 (N_1714,N_1107,N_1245);
or U1715 (N_1715,N_1490,N_1167);
or U1716 (N_1716,N_1239,N_1322);
and U1717 (N_1717,N_1207,N_1255);
nor U1718 (N_1718,N_1269,N_1243);
nor U1719 (N_1719,N_1216,N_1171);
and U1720 (N_1720,N_1357,N_1110);
or U1721 (N_1721,N_1168,N_1379);
and U1722 (N_1722,N_1272,N_1079);
or U1723 (N_1723,N_1088,N_1235);
nor U1724 (N_1724,N_1160,N_1166);
or U1725 (N_1725,N_1325,N_1309);
or U1726 (N_1726,N_1488,N_1172);
and U1727 (N_1727,N_1152,N_1078);
nand U1728 (N_1728,N_1482,N_1211);
nor U1729 (N_1729,N_1453,N_1496);
nand U1730 (N_1730,N_1277,N_1164);
and U1731 (N_1731,N_1495,N_1434);
nor U1732 (N_1732,N_1422,N_1076);
or U1733 (N_1733,N_1381,N_1328);
nand U1734 (N_1734,N_1124,N_1416);
nor U1735 (N_1735,N_1373,N_1159);
or U1736 (N_1736,N_1258,N_1343);
nand U1737 (N_1737,N_1188,N_1007);
xor U1738 (N_1738,N_1439,N_1192);
nor U1739 (N_1739,N_1112,N_1026);
xor U1740 (N_1740,N_1242,N_1091);
or U1741 (N_1741,N_1445,N_1161);
nor U1742 (N_1742,N_1104,N_1237);
nand U1743 (N_1743,N_1044,N_1023);
nand U1744 (N_1744,N_1018,N_1376);
nand U1745 (N_1745,N_1261,N_1222);
nor U1746 (N_1746,N_1114,N_1307);
or U1747 (N_1747,N_1444,N_1069);
and U1748 (N_1748,N_1354,N_1203);
nand U1749 (N_1749,N_1062,N_1304);
and U1750 (N_1750,N_1412,N_1009);
xor U1751 (N_1751,N_1136,N_1042);
and U1752 (N_1752,N_1489,N_1448);
and U1753 (N_1753,N_1442,N_1195);
nor U1754 (N_1754,N_1346,N_1215);
nor U1755 (N_1755,N_1235,N_1223);
nor U1756 (N_1756,N_1187,N_1051);
or U1757 (N_1757,N_1018,N_1189);
or U1758 (N_1758,N_1286,N_1098);
or U1759 (N_1759,N_1033,N_1412);
nand U1760 (N_1760,N_1280,N_1362);
nand U1761 (N_1761,N_1014,N_1432);
xnor U1762 (N_1762,N_1364,N_1470);
nand U1763 (N_1763,N_1007,N_1458);
and U1764 (N_1764,N_1436,N_1469);
or U1765 (N_1765,N_1101,N_1390);
and U1766 (N_1766,N_1453,N_1423);
xor U1767 (N_1767,N_1052,N_1174);
and U1768 (N_1768,N_1129,N_1085);
or U1769 (N_1769,N_1214,N_1259);
and U1770 (N_1770,N_1498,N_1045);
nand U1771 (N_1771,N_1272,N_1107);
and U1772 (N_1772,N_1416,N_1369);
or U1773 (N_1773,N_1213,N_1364);
nand U1774 (N_1774,N_1439,N_1126);
xnor U1775 (N_1775,N_1393,N_1312);
nor U1776 (N_1776,N_1192,N_1195);
and U1777 (N_1777,N_1360,N_1215);
xor U1778 (N_1778,N_1269,N_1279);
or U1779 (N_1779,N_1092,N_1193);
xnor U1780 (N_1780,N_1289,N_1465);
nand U1781 (N_1781,N_1162,N_1075);
and U1782 (N_1782,N_1279,N_1097);
nand U1783 (N_1783,N_1398,N_1439);
nor U1784 (N_1784,N_1181,N_1062);
or U1785 (N_1785,N_1242,N_1086);
nand U1786 (N_1786,N_1110,N_1039);
nor U1787 (N_1787,N_1144,N_1277);
and U1788 (N_1788,N_1096,N_1389);
nor U1789 (N_1789,N_1162,N_1076);
xor U1790 (N_1790,N_1412,N_1464);
or U1791 (N_1791,N_1160,N_1013);
and U1792 (N_1792,N_1340,N_1046);
nand U1793 (N_1793,N_1056,N_1197);
and U1794 (N_1794,N_1446,N_1197);
and U1795 (N_1795,N_1074,N_1020);
nand U1796 (N_1796,N_1216,N_1173);
xor U1797 (N_1797,N_1232,N_1165);
and U1798 (N_1798,N_1046,N_1075);
nor U1799 (N_1799,N_1258,N_1296);
and U1800 (N_1800,N_1451,N_1175);
and U1801 (N_1801,N_1462,N_1227);
and U1802 (N_1802,N_1438,N_1171);
xnor U1803 (N_1803,N_1368,N_1042);
nor U1804 (N_1804,N_1344,N_1282);
or U1805 (N_1805,N_1407,N_1233);
xnor U1806 (N_1806,N_1341,N_1061);
or U1807 (N_1807,N_1354,N_1189);
nand U1808 (N_1808,N_1279,N_1188);
or U1809 (N_1809,N_1496,N_1086);
nor U1810 (N_1810,N_1042,N_1376);
or U1811 (N_1811,N_1368,N_1288);
nor U1812 (N_1812,N_1025,N_1126);
nor U1813 (N_1813,N_1376,N_1109);
nand U1814 (N_1814,N_1435,N_1378);
nand U1815 (N_1815,N_1219,N_1028);
and U1816 (N_1816,N_1081,N_1045);
or U1817 (N_1817,N_1145,N_1195);
or U1818 (N_1818,N_1302,N_1472);
or U1819 (N_1819,N_1390,N_1347);
nand U1820 (N_1820,N_1328,N_1485);
nand U1821 (N_1821,N_1331,N_1281);
nor U1822 (N_1822,N_1177,N_1345);
or U1823 (N_1823,N_1268,N_1151);
nand U1824 (N_1824,N_1494,N_1326);
nor U1825 (N_1825,N_1498,N_1337);
nor U1826 (N_1826,N_1393,N_1271);
and U1827 (N_1827,N_1183,N_1264);
or U1828 (N_1828,N_1309,N_1426);
or U1829 (N_1829,N_1450,N_1286);
or U1830 (N_1830,N_1424,N_1284);
nor U1831 (N_1831,N_1448,N_1053);
nand U1832 (N_1832,N_1017,N_1049);
nand U1833 (N_1833,N_1449,N_1105);
and U1834 (N_1834,N_1292,N_1438);
or U1835 (N_1835,N_1415,N_1439);
nor U1836 (N_1836,N_1131,N_1449);
xor U1837 (N_1837,N_1174,N_1496);
nor U1838 (N_1838,N_1044,N_1112);
nor U1839 (N_1839,N_1058,N_1249);
nand U1840 (N_1840,N_1356,N_1018);
or U1841 (N_1841,N_1219,N_1328);
nand U1842 (N_1842,N_1185,N_1327);
or U1843 (N_1843,N_1479,N_1495);
and U1844 (N_1844,N_1248,N_1136);
or U1845 (N_1845,N_1345,N_1126);
nor U1846 (N_1846,N_1168,N_1103);
or U1847 (N_1847,N_1240,N_1398);
or U1848 (N_1848,N_1495,N_1469);
nor U1849 (N_1849,N_1118,N_1292);
nor U1850 (N_1850,N_1326,N_1138);
and U1851 (N_1851,N_1424,N_1472);
or U1852 (N_1852,N_1155,N_1188);
or U1853 (N_1853,N_1085,N_1155);
nand U1854 (N_1854,N_1338,N_1058);
and U1855 (N_1855,N_1438,N_1129);
and U1856 (N_1856,N_1416,N_1388);
nand U1857 (N_1857,N_1356,N_1076);
nor U1858 (N_1858,N_1271,N_1336);
and U1859 (N_1859,N_1066,N_1109);
nand U1860 (N_1860,N_1319,N_1181);
nor U1861 (N_1861,N_1150,N_1037);
nor U1862 (N_1862,N_1153,N_1292);
or U1863 (N_1863,N_1448,N_1108);
nand U1864 (N_1864,N_1416,N_1134);
or U1865 (N_1865,N_1305,N_1229);
nor U1866 (N_1866,N_1154,N_1249);
nor U1867 (N_1867,N_1104,N_1217);
or U1868 (N_1868,N_1351,N_1388);
or U1869 (N_1869,N_1460,N_1062);
and U1870 (N_1870,N_1152,N_1335);
nand U1871 (N_1871,N_1117,N_1362);
or U1872 (N_1872,N_1235,N_1155);
or U1873 (N_1873,N_1364,N_1405);
nor U1874 (N_1874,N_1496,N_1312);
nand U1875 (N_1875,N_1422,N_1062);
nand U1876 (N_1876,N_1160,N_1082);
or U1877 (N_1877,N_1491,N_1362);
xor U1878 (N_1878,N_1178,N_1060);
nor U1879 (N_1879,N_1029,N_1181);
nand U1880 (N_1880,N_1218,N_1325);
nor U1881 (N_1881,N_1173,N_1230);
and U1882 (N_1882,N_1405,N_1399);
nor U1883 (N_1883,N_1188,N_1457);
xnor U1884 (N_1884,N_1420,N_1123);
xor U1885 (N_1885,N_1334,N_1486);
nor U1886 (N_1886,N_1140,N_1234);
and U1887 (N_1887,N_1353,N_1465);
and U1888 (N_1888,N_1449,N_1098);
nor U1889 (N_1889,N_1323,N_1417);
nand U1890 (N_1890,N_1201,N_1222);
or U1891 (N_1891,N_1428,N_1390);
nor U1892 (N_1892,N_1485,N_1133);
nor U1893 (N_1893,N_1129,N_1012);
or U1894 (N_1894,N_1136,N_1398);
and U1895 (N_1895,N_1261,N_1472);
or U1896 (N_1896,N_1062,N_1244);
or U1897 (N_1897,N_1393,N_1115);
or U1898 (N_1898,N_1064,N_1159);
nor U1899 (N_1899,N_1422,N_1146);
nor U1900 (N_1900,N_1461,N_1384);
and U1901 (N_1901,N_1262,N_1292);
nand U1902 (N_1902,N_1453,N_1017);
nor U1903 (N_1903,N_1165,N_1311);
nor U1904 (N_1904,N_1179,N_1131);
nand U1905 (N_1905,N_1423,N_1185);
or U1906 (N_1906,N_1356,N_1460);
and U1907 (N_1907,N_1161,N_1374);
nor U1908 (N_1908,N_1348,N_1448);
nor U1909 (N_1909,N_1334,N_1254);
nor U1910 (N_1910,N_1196,N_1303);
and U1911 (N_1911,N_1006,N_1214);
or U1912 (N_1912,N_1111,N_1016);
xnor U1913 (N_1913,N_1161,N_1006);
nor U1914 (N_1914,N_1224,N_1249);
nand U1915 (N_1915,N_1082,N_1253);
nor U1916 (N_1916,N_1157,N_1066);
and U1917 (N_1917,N_1308,N_1023);
or U1918 (N_1918,N_1126,N_1013);
nor U1919 (N_1919,N_1266,N_1143);
nor U1920 (N_1920,N_1032,N_1023);
or U1921 (N_1921,N_1032,N_1027);
nor U1922 (N_1922,N_1489,N_1033);
nand U1923 (N_1923,N_1150,N_1323);
xnor U1924 (N_1924,N_1394,N_1475);
or U1925 (N_1925,N_1290,N_1333);
xnor U1926 (N_1926,N_1363,N_1164);
and U1927 (N_1927,N_1499,N_1102);
nor U1928 (N_1928,N_1263,N_1410);
xnor U1929 (N_1929,N_1279,N_1471);
and U1930 (N_1930,N_1431,N_1389);
nand U1931 (N_1931,N_1437,N_1056);
and U1932 (N_1932,N_1453,N_1177);
nand U1933 (N_1933,N_1180,N_1060);
nand U1934 (N_1934,N_1071,N_1391);
and U1935 (N_1935,N_1438,N_1210);
nor U1936 (N_1936,N_1305,N_1147);
nand U1937 (N_1937,N_1192,N_1079);
or U1938 (N_1938,N_1440,N_1248);
nor U1939 (N_1939,N_1080,N_1025);
nand U1940 (N_1940,N_1326,N_1226);
and U1941 (N_1941,N_1182,N_1302);
and U1942 (N_1942,N_1204,N_1161);
xnor U1943 (N_1943,N_1328,N_1119);
nor U1944 (N_1944,N_1014,N_1404);
or U1945 (N_1945,N_1270,N_1281);
xor U1946 (N_1946,N_1174,N_1365);
nor U1947 (N_1947,N_1240,N_1405);
and U1948 (N_1948,N_1264,N_1424);
or U1949 (N_1949,N_1366,N_1419);
nand U1950 (N_1950,N_1320,N_1430);
or U1951 (N_1951,N_1496,N_1002);
nand U1952 (N_1952,N_1267,N_1457);
nand U1953 (N_1953,N_1317,N_1163);
or U1954 (N_1954,N_1116,N_1109);
or U1955 (N_1955,N_1271,N_1409);
nand U1956 (N_1956,N_1090,N_1187);
nor U1957 (N_1957,N_1189,N_1431);
nand U1958 (N_1958,N_1246,N_1305);
and U1959 (N_1959,N_1096,N_1412);
and U1960 (N_1960,N_1346,N_1094);
xnor U1961 (N_1961,N_1239,N_1483);
or U1962 (N_1962,N_1428,N_1416);
or U1963 (N_1963,N_1223,N_1190);
xor U1964 (N_1964,N_1133,N_1499);
nand U1965 (N_1965,N_1315,N_1337);
or U1966 (N_1966,N_1348,N_1423);
nor U1967 (N_1967,N_1240,N_1251);
nand U1968 (N_1968,N_1358,N_1077);
nor U1969 (N_1969,N_1349,N_1450);
and U1970 (N_1970,N_1335,N_1324);
or U1971 (N_1971,N_1495,N_1476);
nor U1972 (N_1972,N_1234,N_1362);
and U1973 (N_1973,N_1112,N_1188);
nand U1974 (N_1974,N_1403,N_1103);
xor U1975 (N_1975,N_1098,N_1142);
nor U1976 (N_1976,N_1446,N_1318);
or U1977 (N_1977,N_1117,N_1454);
nor U1978 (N_1978,N_1190,N_1050);
and U1979 (N_1979,N_1348,N_1078);
nand U1980 (N_1980,N_1454,N_1341);
nand U1981 (N_1981,N_1274,N_1312);
and U1982 (N_1982,N_1222,N_1051);
nor U1983 (N_1983,N_1300,N_1427);
nand U1984 (N_1984,N_1277,N_1002);
nand U1985 (N_1985,N_1151,N_1156);
nor U1986 (N_1986,N_1230,N_1217);
nor U1987 (N_1987,N_1300,N_1198);
and U1988 (N_1988,N_1097,N_1460);
xnor U1989 (N_1989,N_1417,N_1218);
or U1990 (N_1990,N_1204,N_1141);
and U1991 (N_1991,N_1269,N_1316);
nor U1992 (N_1992,N_1372,N_1178);
or U1993 (N_1993,N_1072,N_1316);
and U1994 (N_1994,N_1171,N_1020);
and U1995 (N_1995,N_1129,N_1139);
or U1996 (N_1996,N_1142,N_1037);
nor U1997 (N_1997,N_1238,N_1246);
xnor U1998 (N_1998,N_1383,N_1467);
xor U1999 (N_1999,N_1334,N_1111);
nand U2000 (N_2000,N_1656,N_1670);
and U2001 (N_2001,N_1815,N_1558);
nand U2002 (N_2002,N_1706,N_1619);
nand U2003 (N_2003,N_1780,N_1796);
and U2004 (N_2004,N_1548,N_1809);
or U2005 (N_2005,N_1887,N_1657);
or U2006 (N_2006,N_1914,N_1766);
or U2007 (N_2007,N_1529,N_1873);
xnor U2008 (N_2008,N_1992,N_1562);
and U2009 (N_2009,N_1697,N_1842);
nor U2010 (N_2010,N_1909,N_1924);
nor U2011 (N_2011,N_1526,N_1935);
and U2012 (N_2012,N_1776,N_1812);
or U2013 (N_2013,N_1635,N_1816);
nor U2014 (N_2014,N_1690,N_1911);
nor U2015 (N_2015,N_1535,N_1857);
and U2016 (N_2016,N_1577,N_1718);
nor U2017 (N_2017,N_1856,N_1707);
or U2018 (N_2018,N_1549,N_1981);
or U2019 (N_2019,N_1721,N_1506);
xnor U2020 (N_2020,N_1557,N_1500);
nor U2021 (N_2021,N_1797,N_1917);
xor U2022 (N_2022,N_1987,N_1801);
nor U2023 (N_2023,N_1773,N_1973);
nor U2024 (N_2024,N_1689,N_1705);
nand U2025 (N_2025,N_1971,N_1692);
nor U2026 (N_2026,N_1531,N_1753);
nand U2027 (N_2027,N_1966,N_1946);
or U2028 (N_2028,N_1869,N_1700);
nor U2029 (N_2029,N_1573,N_1701);
and U2030 (N_2030,N_1872,N_1617);
nand U2031 (N_2031,N_1941,N_1505);
nor U2032 (N_2032,N_1612,N_1998);
or U2033 (N_2033,N_1953,N_1551);
and U2034 (N_2034,N_1746,N_1623);
or U2035 (N_2035,N_1546,N_1912);
xor U2036 (N_2036,N_1524,N_1595);
or U2037 (N_2037,N_1940,N_1640);
nand U2038 (N_2038,N_1686,N_1839);
or U2039 (N_2039,N_1850,N_1592);
nor U2040 (N_2040,N_1970,N_1982);
and U2041 (N_2041,N_1758,N_1583);
nor U2042 (N_2042,N_1566,N_1662);
or U2043 (N_2043,N_1702,N_1593);
or U2044 (N_2044,N_1737,N_1890);
and U2045 (N_2045,N_1667,N_1503);
or U2046 (N_2046,N_1810,N_1717);
nand U2047 (N_2047,N_1731,N_1674);
nand U2048 (N_2048,N_1969,N_1539);
or U2049 (N_2049,N_1808,N_1511);
and U2050 (N_2050,N_1794,N_1568);
nand U2051 (N_2051,N_1778,N_1598);
nor U2052 (N_2052,N_1615,N_1575);
nor U2053 (N_2053,N_1787,N_1921);
and U2054 (N_2054,N_1823,N_1680);
nand U2055 (N_2055,N_1691,N_1894);
or U2056 (N_2056,N_1938,N_1545);
and U2057 (N_2057,N_1906,N_1508);
and U2058 (N_2058,N_1734,N_1893);
and U2059 (N_2059,N_1846,N_1963);
nor U2060 (N_2060,N_1782,N_1587);
and U2061 (N_2061,N_1581,N_1789);
nor U2062 (N_2062,N_1603,N_1819);
and U2063 (N_2063,N_1723,N_1519);
or U2064 (N_2064,N_1552,N_1967);
nor U2065 (N_2065,N_1844,N_1870);
xor U2066 (N_2066,N_1915,N_1919);
or U2067 (N_2067,N_1621,N_1783);
or U2068 (N_2068,N_1620,N_1838);
nor U2069 (N_2069,N_1854,N_1806);
and U2070 (N_2070,N_1898,N_1507);
or U2071 (N_2071,N_1530,N_1678);
or U2072 (N_2072,N_1876,N_1534);
nand U2073 (N_2073,N_1565,N_1613);
and U2074 (N_2074,N_1832,N_1672);
and U2075 (N_2075,N_1540,N_1895);
or U2076 (N_2076,N_1588,N_1871);
nand U2077 (N_2077,N_1650,N_1708);
xor U2078 (N_2078,N_1892,N_1685);
nand U2079 (N_2079,N_1831,N_1528);
nor U2080 (N_2080,N_1936,N_1749);
and U2081 (N_2081,N_1750,N_1896);
or U2082 (N_2082,N_1543,N_1916);
nand U2083 (N_2083,N_1533,N_1561);
or U2084 (N_2084,N_1569,N_1885);
nand U2085 (N_2085,N_1851,N_1625);
nor U2086 (N_2086,N_1837,N_1790);
nor U2087 (N_2087,N_1563,N_1522);
and U2088 (N_2088,N_1805,N_1673);
and U2089 (N_2089,N_1772,N_1745);
or U2090 (N_2090,N_1618,N_1742);
and U2091 (N_2091,N_1814,N_1605);
xor U2092 (N_2092,N_1888,N_1743);
and U2093 (N_2093,N_1571,N_1997);
and U2094 (N_2094,N_1687,N_1875);
and U2095 (N_2095,N_1990,N_1658);
xor U2096 (N_2096,N_1983,N_1811);
or U2097 (N_2097,N_1822,N_1803);
nand U2098 (N_2098,N_1864,N_1785);
or U2099 (N_2099,N_1828,N_1570);
and U2100 (N_2100,N_1727,N_1740);
nand U2101 (N_2101,N_1611,N_1884);
or U2102 (N_2102,N_1863,N_1853);
nand U2103 (N_2103,N_1922,N_1675);
nor U2104 (N_2104,N_1859,N_1879);
and U2105 (N_2105,N_1891,N_1514);
and U2106 (N_2106,N_1653,N_1958);
or U2107 (N_2107,N_1800,N_1923);
or U2108 (N_2108,N_1616,N_1733);
xor U2109 (N_2109,N_1834,N_1537);
nor U2110 (N_2110,N_1732,N_1770);
nand U2111 (N_2111,N_1993,N_1724);
and U2112 (N_2112,N_1761,N_1920);
nor U2113 (N_2113,N_1984,N_1722);
and U2114 (N_2114,N_1688,N_1584);
and U2115 (N_2115,N_1676,N_1858);
and U2116 (N_2116,N_1594,N_1933);
and U2117 (N_2117,N_1974,N_1948);
or U2118 (N_2118,N_1843,N_1826);
or U2119 (N_2119,N_1677,N_1538);
and U2120 (N_2120,N_1682,N_1845);
and U2121 (N_2121,N_1760,N_1726);
nand U2122 (N_2122,N_1601,N_1523);
or U2123 (N_2123,N_1972,N_1755);
nor U2124 (N_2124,N_1719,N_1754);
nor U2125 (N_2125,N_1599,N_1713);
nor U2126 (N_2126,N_1880,N_1934);
xnor U2127 (N_2127,N_1883,N_1976);
nor U2128 (N_2128,N_1720,N_1631);
and U2129 (N_2129,N_1913,N_1665);
nand U2130 (N_2130,N_1937,N_1957);
or U2131 (N_2131,N_1881,N_1991);
nand U2132 (N_2132,N_1798,N_1986);
or U2133 (N_2133,N_1978,N_1532);
and U2134 (N_2134,N_1784,N_1696);
nand U2135 (N_2135,N_1738,N_1579);
nor U2136 (N_2136,N_1556,N_1627);
or U2137 (N_2137,N_1704,N_1602);
nor U2138 (N_2138,N_1596,N_1897);
or U2139 (N_2139,N_1628,N_1567);
nor U2140 (N_2140,N_1752,N_1554);
or U2141 (N_2141,N_1840,N_1517);
nor U2142 (N_2142,N_1693,N_1630);
and U2143 (N_2143,N_1867,N_1827);
nor U2144 (N_2144,N_1609,N_1835);
nor U2145 (N_2145,N_1736,N_1501);
or U2146 (N_2146,N_1756,N_1950);
nor U2147 (N_2147,N_1715,N_1759);
nor U2148 (N_2148,N_1975,N_1681);
nand U2149 (N_2149,N_1520,N_1502);
and U2150 (N_2150,N_1910,N_1779);
xnor U2151 (N_2151,N_1559,N_1899);
or U2152 (N_2152,N_1930,N_1716);
nand U2153 (N_2153,N_1550,N_1555);
nand U2154 (N_2154,N_1589,N_1791);
nor U2155 (N_2155,N_1542,N_1952);
and U2156 (N_2156,N_1652,N_1960);
and U2157 (N_2157,N_1764,N_1849);
nand U2158 (N_2158,N_1516,N_1882);
and U2159 (N_2159,N_1739,N_1626);
nand U2160 (N_2160,N_1638,N_1925);
nand U2161 (N_2161,N_1660,N_1943);
nand U2162 (N_2162,N_1886,N_1847);
nand U2163 (N_2163,N_1999,N_1632);
and U2164 (N_2164,N_1955,N_1641);
nor U2165 (N_2165,N_1661,N_1852);
and U2166 (N_2166,N_1829,N_1645);
xor U2167 (N_2167,N_1637,N_1679);
xnor U2168 (N_2168,N_1932,N_1703);
nor U2169 (N_2169,N_1907,N_1668);
and U2170 (N_2170,N_1931,N_1735);
and U2171 (N_2171,N_1515,N_1949);
and U2172 (N_2172,N_1860,N_1813);
xor U2173 (N_2173,N_1865,N_1698);
nor U2174 (N_2174,N_1709,N_1591);
xor U2175 (N_2175,N_1684,N_1807);
and U2176 (N_2176,N_1830,N_1954);
and U2177 (N_2177,N_1833,N_1655);
or U2178 (N_2178,N_1699,N_1564);
or U2179 (N_2179,N_1767,N_1965);
and U2180 (N_2180,N_1939,N_1547);
and U2181 (N_2181,N_1964,N_1989);
or U2182 (N_2182,N_1765,N_1824);
or U2183 (N_2183,N_1710,N_1714);
nand U2184 (N_2184,N_1771,N_1729);
nor U2185 (N_2185,N_1694,N_1862);
or U2186 (N_2186,N_1928,N_1580);
nor U2187 (N_2187,N_1929,N_1777);
nor U2188 (N_2188,N_1634,N_1763);
and U2189 (N_2189,N_1585,N_1942);
and U2190 (N_2190,N_1994,N_1586);
and U2191 (N_2191,N_1947,N_1544);
nor U2192 (N_2192,N_1995,N_1985);
xor U2193 (N_2193,N_1578,N_1600);
or U2194 (N_2194,N_1927,N_1874);
nor U2195 (N_2195,N_1817,N_1504);
nor U2196 (N_2196,N_1751,N_1642);
or U2197 (N_2197,N_1769,N_1848);
nand U2198 (N_2198,N_1741,N_1597);
or U2199 (N_2199,N_1802,N_1961);
or U2200 (N_2200,N_1792,N_1624);
nand U2201 (N_2201,N_1825,N_1945);
or U2202 (N_2202,N_1748,N_1518);
xnor U2203 (N_2203,N_1663,N_1683);
nand U2204 (N_2204,N_1622,N_1590);
nor U2205 (N_2205,N_1521,N_1644);
and U2206 (N_2206,N_1926,N_1944);
or U2207 (N_2207,N_1610,N_1855);
and U2208 (N_2208,N_1513,N_1861);
nand U2209 (N_2209,N_1744,N_1576);
and U2210 (N_2210,N_1560,N_1633);
xnor U2211 (N_2211,N_1608,N_1614);
nor U2212 (N_2212,N_1804,N_1977);
and U2213 (N_2213,N_1962,N_1541);
or U2214 (N_2214,N_1903,N_1725);
nand U2215 (N_2215,N_1536,N_1509);
or U2216 (N_2216,N_1889,N_1868);
and U2217 (N_2217,N_1979,N_1666);
nor U2218 (N_2218,N_1639,N_1553);
nor U2219 (N_2219,N_1664,N_1788);
or U2220 (N_2220,N_1510,N_1951);
xor U2221 (N_2221,N_1799,N_1900);
nor U2222 (N_2222,N_1786,N_1902);
xnor U2223 (N_2223,N_1757,N_1730);
or U2224 (N_2224,N_1712,N_1905);
or U2225 (N_2225,N_1768,N_1651);
nor U2226 (N_2226,N_1747,N_1908);
nand U2227 (N_2227,N_1582,N_1525);
nor U2228 (N_2228,N_1836,N_1866);
and U2229 (N_2229,N_1649,N_1629);
xnor U2230 (N_2230,N_1728,N_1968);
or U2231 (N_2231,N_1901,N_1820);
and U2232 (N_2232,N_1654,N_1527);
nor U2233 (N_2233,N_1878,N_1841);
nand U2234 (N_2234,N_1956,N_1659);
or U2235 (N_2235,N_1572,N_1643);
and U2236 (N_2236,N_1762,N_1604);
or U2237 (N_2237,N_1647,N_1980);
and U2238 (N_2238,N_1821,N_1695);
or U2239 (N_2239,N_1918,N_1636);
nor U2240 (N_2240,N_1818,N_1781);
xor U2241 (N_2241,N_1795,N_1648);
nor U2242 (N_2242,N_1512,N_1711);
and U2243 (N_2243,N_1646,N_1606);
or U2244 (N_2244,N_1574,N_1988);
or U2245 (N_2245,N_1671,N_1774);
xor U2246 (N_2246,N_1607,N_1996);
nor U2247 (N_2247,N_1669,N_1793);
nor U2248 (N_2248,N_1775,N_1959);
nand U2249 (N_2249,N_1877,N_1904);
nor U2250 (N_2250,N_1926,N_1521);
nand U2251 (N_2251,N_1655,N_1938);
nand U2252 (N_2252,N_1504,N_1731);
and U2253 (N_2253,N_1585,N_1853);
nand U2254 (N_2254,N_1636,N_1927);
nand U2255 (N_2255,N_1960,N_1836);
nand U2256 (N_2256,N_1509,N_1669);
and U2257 (N_2257,N_1536,N_1583);
or U2258 (N_2258,N_1776,N_1993);
or U2259 (N_2259,N_1715,N_1647);
nor U2260 (N_2260,N_1880,N_1951);
and U2261 (N_2261,N_1695,N_1781);
or U2262 (N_2262,N_1889,N_1703);
xor U2263 (N_2263,N_1730,N_1586);
or U2264 (N_2264,N_1777,N_1592);
and U2265 (N_2265,N_1794,N_1931);
or U2266 (N_2266,N_1611,N_1572);
nand U2267 (N_2267,N_1730,N_1598);
or U2268 (N_2268,N_1805,N_1598);
or U2269 (N_2269,N_1649,N_1634);
nand U2270 (N_2270,N_1519,N_1552);
or U2271 (N_2271,N_1943,N_1516);
nand U2272 (N_2272,N_1706,N_1705);
nand U2273 (N_2273,N_1961,N_1801);
nand U2274 (N_2274,N_1581,N_1615);
nor U2275 (N_2275,N_1653,N_1963);
nor U2276 (N_2276,N_1967,N_1994);
xnor U2277 (N_2277,N_1689,N_1735);
or U2278 (N_2278,N_1949,N_1915);
or U2279 (N_2279,N_1838,N_1573);
xnor U2280 (N_2280,N_1844,N_1530);
nor U2281 (N_2281,N_1954,N_1946);
or U2282 (N_2282,N_1855,N_1814);
nor U2283 (N_2283,N_1915,N_1674);
and U2284 (N_2284,N_1834,N_1611);
nor U2285 (N_2285,N_1573,N_1945);
nor U2286 (N_2286,N_1730,N_1932);
and U2287 (N_2287,N_1520,N_1542);
nand U2288 (N_2288,N_1696,N_1736);
and U2289 (N_2289,N_1631,N_1976);
nand U2290 (N_2290,N_1865,N_1513);
nor U2291 (N_2291,N_1747,N_1993);
or U2292 (N_2292,N_1990,N_1524);
xor U2293 (N_2293,N_1822,N_1873);
nor U2294 (N_2294,N_1582,N_1880);
or U2295 (N_2295,N_1976,N_1715);
or U2296 (N_2296,N_1915,N_1896);
nand U2297 (N_2297,N_1731,N_1801);
nand U2298 (N_2298,N_1615,N_1683);
or U2299 (N_2299,N_1730,N_1820);
xor U2300 (N_2300,N_1588,N_1820);
nor U2301 (N_2301,N_1729,N_1600);
and U2302 (N_2302,N_1961,N_1572);
or U2303 (N_2303,N_1738,N_1910);
nor U2304 (N_2304,N_1664,N_1909);
nor U2305 (N_2305,N_1850,N_1864);
or U2306 (N_2306,N_1691,N_1658);
or U2307 (N_2307,N_1573,N_1746);
or U2308 (N_2308,N_1753,N_1623);
and U2309 (N_2309,N_1970,N_1958);
and U2310 (N_2310,N_1854,N_1893);
nor U2311 (N_2311,N_1806,N_1769);
and U2312 (N_2312,N_1585,N_1678);
or U2313 (N_2313,N_1949,N_1811);
xnor U2314 (N_2314,N_1575,N_1580);
nor U2315 (N_2315,N_1656,N_1885);
nand U2316 (N_2316,N_1864,N_1722);
nand U2317 (N_2317,N_1900,N_1895);
nor U2318 (N_2318,N_1647,N_1877);
and U2319 (N_2319,N_1719,N_1808);
nand U2320 (N_2320,N_1721,N_1722);
nor U2321 (N_2321,N_1939,N_1979);
and U2322 (N_2322,N_1661,N_1859);
and U2323 (N_2323,N_1539,N_1529);
or U2324 (N_2324,N_1756,N_1519);
xor U2325 (N_2325,N_1591,N_1630);
nand U2326 (N_2326,N_1706,N_1697);
xor U2327 (N_2327,N_1551,N_1553);
nand U2328 (N_2328,N_1739,N_1871);
and U2329 (N_2329,N_1865,N_1510);
and U2330 (N_2330,N_1530,N_1536);
and U2331 (N_2331,N_1956,N_1904);
or U2332 (N_2332,N_1698,N_1872);
or U2333 (N_2333,N_1602,N_1702);
nand U2334 (N_2334,N_1656,N_1940);
nand U2335 (N_2335,N_1940,N_1755);
nor U2336 (N_2336,N_1832,N_1725);
or U2337 (N_2337,N_1935,N_1654);
xnor U2338 (N_2338,N_1936,N_1566);
or U2339 (N_2339,N_1674,N_1784);
nand U2340 (N_2340,N_1551,N_1763);
nor U2341 (N_2341,N_1509,N_1673);
and U2342 (N_2342,N_1985,N_1852);
nand U2343 (N_2343,N_1644,N_1511);
or U2344 (N_2344,N_1608,N_1587);
nor U2345 (N_2345,N_1691,N_1731);
nor U2346 (N_2346,N_1541,N_1753);
nor U2347 (N_2347,N_1825,N_1501);
and U2348 (N_2348,N_1892,N_1580);
and U2349 (N_2349,N_1758,N_1702);
nor U2350 (N_2350,N_1644,N_1703);
nand U2351 (N_2351,N_1821,N_1790);
nand U2352 (N_2352,N_1580,N_1644);
nand U2353 (N_2353,N_1673,N_1760);
nand U2354 (N_2354,N_1955,N_1913);
and U2355 (N_2355,N_1819,N_1977);
nand U2356 (N_2356,N_1746,N_1860);
nor U2357 (N_2357,N_1537,N_1533);
nor U2358 (N_2358,N_1576,N_1535);
or U2359 (N_2359,N_1789,N_1654);
nand U2360 (N_2360,N_1959,N_1789);
and U2361 (N_2361,N_1981,N_1743);
nor U2362 (N_2362,N_1559,N_1866);
and U2363 (N_2363,N_1887,N_1919);
nand U2364 (N_2364,N_1652,N_1991);
nor U2365 (N_2365,N_1832,N_1680);
nor U2366 (N_2366,N_1816,N_1819);
nand U2367 (N_2367,N_1929,N_1837);
nor U2368 (N_2368,N_1996,N_1876);
or U2369 (N_2369,N_1797,N_1541);
or U2370 (N_2370,N_1542,N_1514);
nor U2371 (N_2371,N_1777,N_1828);
nand U2372 (N_2372,N_1562,N_1789);
or U2373 (N_2373,N_1808,N_1730);
nand U2374 (N_2374,N_1970,N_1783);
xor U2375 (N_2375,N_1837,N_1781);
and U2376 (N_2376,N_1844,N_1952);
and U2377 (N_2377,N_1905,N_1990);
and U2378 (N_2378,N_1755,N_1862);
and U2379 (N_2379,N_1815,N_1911);
nor U2380 (N_2380,N_1629,N_1594);
nor U2381 (N_2381,N_1575,N_1898);
or U2382 (N_2382,N_1808,N_1967);
and U2383 (N_2383,N_1647,N_1566);
or U2384 (N_2384,N_1897,N_1985);
nand U2385 (N_2385,N_1634,N_1743);
xor U2386 (N_2386,N_1975,N_1830);
or U2387 (N_2387,N_1828,N_1510);
nor U2388 (N_2388,N_1833,N_1572);
or U2389 (N_2389,N_1684,N_1593);
nand U2390 (N_2390,N_1541,N_1512);
nor U2391 (N_2391,N_1882,N_1977);
and U2392 (N_2392,N_1711,N_1504);
xor U2393 (N_2393,N_1780,N_1799);
or U2394 (N_2394,N_1557,N_1934);
and U2395 (N_2395,N_1845,N_1532);
and U2396 (N_2396,N_1856,N_1584);
or U2397 (N_2397,N_1875,N_1615);
or U2398 (N_2398,N_1723,N_1705);
or U2399 (N_2399,N_1885,N_1560);
nand U2400 (N_2400,N_1966,N_1749);
and U2401 (N_2401,N_1884,N_1797);
nand U2402 (N_2402,N_1544,N_1774);
nand U2403 (N_2403,N_1558,N_1628);
or U2404 (N_2404,N_1656,N_1628);
xor U2405 (N_2405,N_1607,N_1712);
and U2406 (N_2406,N_1588,N_1710);
and U2407 (N_2407,N_1952,N_1560);
xnor U2408 (N_2408,N_1533,N_1570);
nor U2409 (N_2409,N_1770,N_1801);
or U2410 (N_2410,N_1713,N_1926);
and U2411 (N_2411,N_1645,N_1738);
nand U2412 (N_2412,N_1715,N_1728);
nand U2413 (N_2413,N_1684,N_1591);
xor U2414 (N_2414,N_1599,N_1993);
or U2415 (N_2415,N_1694,N_1970);
nor U2416 (N_2416,N_1979,N_1974);
nor U2417 (N_2417,N_1822,N_1568);
xor U2418 (N_2418,N_1799,N_1961);
and U2419 (N_2419,N_1750,N_1709);
nor U2420 (N_2420,N_1873,N_1800);
xor U2421 (N_2421,N_1606,N_1878);
or U2422 (N_2422,N_1728,N_1877);
nand U2423 (N_2423,N_1738,N_1946);
or U2424 (N_2424,N_1722,N_1887);
and U2425 (N_2425,N_1868,N_1528);
nor U2426 (N_2426,N_1537,N_1548);
nor U2427 (N_2427,N_1669,N_1801);
or U2428 (N_2428,N_1760,N_1846);
xor U2429 (N_2429,N_1733,N_1839);
nand U2430 (N_2430,N_1800,N_1850);
and U2431 (N_2431,N_1960,N_1553);
xnor U2432 (N_2432,N_1684,N_1895);
or U2433 (N_2433,N_1947,N_1604);
nor U2434 (N_2434,N_1703,N_1841);
nor U2435 (N_2435,N_1974,N_1583);
and U2436 (N_2436,N_1628,N_1970);
nor U2437 (N_2437,N_1566,N_1637);
and U2438 (N_2438,N_1873,N_1700);
nand U2439 (N_2439,N_1671,N_1718);
and U2440 (N_2440,N_1521,N_1971);
nand U2441 (N_2441,N_1769,N_1726);
or U2442 (N_2442,N_1783,N_1604);
nand U2443 (N_2443,N_1787,N_1923);
nor U2444 (N_2444,N_1971,N_1769);
and U2445 (N_2445,N_1777,N_1712);
nor U2446 (N_2446,N_1992,N_1919);
and U2447 (N_2447,N_1621,N_1863);
xnor U2448 (N_2448,N_1579,N_1610);
xnor U2449 (N_2449,N_1553,N_1732);
nand U2450 (N_2450,N_1641,N_1925);
and U2451 (N_2451,N_1525,N_1764);
and U2452 (N_2452,N_1633,N_1865);
nand U2453 (N_2453,N_1507,N_1709);
or U2454 (N_2454,N_1848,N_1863);
or U2455 (N_2455,N_1521,N_1561);
nor U2456 (N_2456,N_1646,N_1688);
or U2457 (N_2457,N_1515,N_1806);
nand U2458 (N_2458,N_1754,N_1687);
nor U2459 (N_2459,N_1855,N_1637);
xor U2460 (N_2460,N_1831,N_1653);
nor U2461 (N_2461,N_1625,N_1777);
or U2462 (N_2462,N_1928,N_1574);
nor U2463 (N_2463,N_1753,N_1822);
xor U2464 (N_2464,N_1557,N_1876);
and U2465 (N_2465,N_1700,N_1769);
and U2466 (N_2466,N_1559,N_1948);
and U2467 (N_2467,N_1608,N_1768);
or U2468 (N_2468,N_1777,N_1619);
nand U2469 (N_2469,N_1929,N_1903);
nand U2470 (N_2470,N_1660,N_1539);
or U2471 (N_2471,N_1837,N_1640);
nor U2472 (N_2472,N_1753,N_1528);
or U2473 (N_2473,N_1860,N_1950);
nand U2474 (N_2474,N_1608,N_1834);
and U2475 (N_2475,N_1726,N_1606);
nor U2476 (N_2476,N_1612,N_1982);
nor U2477 (N_2477,N_1969,N_1846);
and U2478 (N_2478,N_1549,N_1753);
or U2479 (N_2479,N_1535,N_1686);
nor U2480 (N_2480,N_1522,N_1718);
or U2481 (N_2481,N_1923,N_1824);
and U2482 (N_2482,N_1617,N_1534);
and U2483 (N_2483,N_1765,N_1522);
nand U2484 (N_2484,N_1600,N_1867);
or U2485 (N_2485,N_1725,N_1729);
and U2486 (N_2486,N_1886,N_1712);
or U2487 (N_2487,N_1849,N_1950);
nor U2488 (N_2488,N_1561,N_1893);
or U2489 (N_2489,N_1748,N_1902);
nand U2490 (N_2490,N_1889,N_1930);
or U2491 (N_2491,N_1611,N_1664);
nand U2492 (N_2492,N_1732,N_1793);
nor U2493 (N_2493,N_1817,N_1531);
nor U2494 (N_2494,N_1810,N_1660);
nand U2495 (N_2495,N_1743,N_1972);
and U2496 (N_2496,N_1944,N_1947);
and U2497 (N_2497,N_1601,N_1918);
or U2498 (N_2498,N_1554,N_1859);
and U2499 (N_2499,N_1749,N_1932);
nor U2500 (N_2500,N_2354,N_2467);
xnor U2501 (N_2501,N_2459,N_2012);
nor U2502 (N_2502,N_2396,N_2143);
xnor U2503 (N_2503,N_2443,N_2042);
nand U2504 (N_2504,N_2260,N_2233);
nand U2505 (N_2505,N_2375,N_2149);
nor U2506 (N_2506,N_2295,N_2245);
or U2507 (N_2507,N_2264,N_2325);
and U2508 (N_2508,N_2166,N_2452);
or U2509 (N_2509,N_2155,N_2040);
xor U2510 (N_2510,N_2446,N_2081);
nor U2511 (N_2511,N_2213,N_2301);
and U2512 (N_2512,N_2196,N_2019);
or U2513 (N_2513,N_2400,N_2358);
or U2514 (N_2514,N_2219,N_2072);
or U2515 (N_2515,N_2193,N_2460);
nand U2516 (N_2516,N_2335,N_2328);
xor U2517 (N_2517,N_2435,N_2076);
or U2518 (N_2518,N_2357,N_2331);
xor U2519 (N_2519,N_2444,N_2015);
nand U2520 (N_2520,N_2360,N_2432);
xor U2521 (N_2521,N_2231,N_2367);
nand U2522 (N_2522,N_2212,N_2159);
and U2523 (N_2523,N_2063,N_2027);
nand U2524 (N_2524,N_2437,N_2230);
nor U2525 (N_2525,N_2294,N_2383);
or U2526 (N_2526,N_2172,N_2109);
nor U2527 (N_2527,N_2261,N_2158);
and U2528 (N_2528,N_2322,N_2116);
or U2529 (N_2529,N_2393,N_2346);
nand U2530 (N_2530,N_2226,N_2255);
nand U2531 (N_2531,N_2201,N_2487);
nor U2532 (N_2532,N_2096,N_2471);
nor U2533 (N_2533,N_2408,N_2309);
nor U2534 (N_2534,N_2266,N_2180);
xor U2535 (N_2535,N_2385,N_2398);
or U2536 (N_2536,N_2221,N_2074);
or U2537 (N_2537,N_2314,N_2484);
and U2538 (N_2538,N_2362,N_2284);
nand U2539 (N_2539,N_2333,N_2110);
and U2540 (N_2540,N_2115,N_2227);
nor U2541 (N_2541,N_2183,N_2399);
nand U2542 (N_2542,N_2038,N_2177);
nand U2543 (N_2543,N_2218,N_2006);
nor U2544 (N_2544,N_2217,N_2268);
and U2545 (N_2545,N_2348,N_2239);
nor U2546 (N_2546,N_2472,N_2039);
xnor U2547 (N_2547,N_2355,N_2064);
xor U2548 (N_2548,N_2361,N_2428);
xor U2549 (N_2549,N_2496,N_2407);
nand U2550 (N_2550,N_2124,N_2028);
or U2551 (N_2551,N_2251,N_2389);
xor U2552 (N_2552,N_2178,N_2468);
nand U2553 (N_2553,N_2454,N_2495);
nor U2554 (N_2554,N_2161,N_2480);
or U2555 (N_2555,N_2136,N_2037);
nor U2556 (N_2556,N_2303,N_2121);
nor U2557 (N_2557,N_2341,N_2368);
nand U2558 (N_2558,N_2320,N_2469);
and U2559 (N_2559,N_2244,N_2272);
nor U2560 (N_2560,N_2413,N_2364);
nor U2561 (N_2561,N_2223,N_2225);
and U2562 (N_2562,N_2321,N_2098);
nor U2563 (N_2563,N_2319,N_2253);
xor U2564 (N_2564,N_2285,N_2162);
nand U2565 (N_2565,N_2047,N_2243);
and U2566 (N_2566,N_2440,N_2278);
nor U2567 (N_2567,N_2065,N_2448);
and U2568 (N_2568,N_2023,N_2008);
or U2569 (N_2569,N_2356,N_2482);
nor U2570 (N_2570,N_2486,N_2147);
or U2571 (N_2571,N_2492,N_2061);
nor U2572 (N_2572,N_2171,N_2237);
or U2573 (N_2573,N_2401,N_2347);
nand U2574 (N_2574,N_2186,N_2145);
nor U2575 (N_2575,N_2153,N_2169);
nor U2576 (N_2576,N_2418,N_2334);
xor U2577 (N_2577,N_2483,N_2010);
xnor U2578 (N_2578,N_2093,N_2494);
or U2579 (N_2579,N_2094,N_2007);
nor U2580 (N_2580,N_2215,N_2350);
nor U2581 (N_2581,N_2133,N_2105);
nor U2582 (N_2582,N_2447,N_2100);
nand U2583 (N_2583,N_2293,N_2099);
and U2584 (N_2584,N_2307,N_2412);
nand U2585 (N_2585,N_2417,N_2277);
or U2586 (N_2586,N_2323,N_2044);
or U2587 (N_2587,N_2438,N_2299);
or U2588 (N_2588,N_2129,N_2214);
and U2589 (N_2589,N_2411,N_2296);
nor U2590 (N_2590,N_2263,N_2493);
nand U2591 (N_2591,N_2033,N_2194);
nand U2592 (N_2592,N_2423,N_2250);
nand U2593 (N_2593,N_2372,N_2306);
or U2594 (N_2594,N_2324,N_2479);
nor U2595 (N_2595,N_2477,N_2387);
nand U2596 (N_2596,N_2031,N_2466);
nor U2597 (N_2597,N_2071,N_2127);
xor U2598 (N_2598,N_2123,N_2126);
xnor U2599 (N_2599,N_2157,N_2386);
nand U2600 (N_2600,N_2343,N_2210);
nor U2601 (N_2601,N_2415,N_2282);
nand U2602 (N_2602,N_2252,N_2025);
nor U2603 (N_2603,N_2187,N_2113);
nand U2604 (N_2604,N_2165,N_2017);
nand U2605 (N_2605,N_2232,N_2198);
xnor U2606 (N_2606,N_2035,N_2315);
xnor U2607 (N_2607,N_2142,N_2489);
and U2608 (N_2608,N_2088,N_2046);
or U2609 (N_2609,N_2290,N_2283);
nor U2610 (N_2610,N_2340,N_2405);
and U2611 (N_2611,N_2337,N_2330);
and U2612 (N_2612,N_2391,N_2406);
and U2613 (N_2613,N_2429,N_2059);
or U2614 (N_2614,N_2490,N_2144);
or U2615 (N_2615,N_2185,N_2478);
nor U2616 (N_2616,N_2404,N_2339);
or U2617 (N_2617,N_2045,N_2270);
or U2618 (N_2618,N_2199,N_2114);
and U2619 (N_2619,N_2052,N_2271);
or U2620 (N_2620,N_2050,N_2485);
nor U2621 (N_2621,N_2181,N_2422);
nand U2622 (N_2622,N_2461,N_2376);
nor U2623 (N_2623,N_2238,N_2104);
and U2624 (N_2624,N_2138,N_2475);
xnor U2625 (N_2625,N_2032,N_2465);
nor U2626 (N_2626,N_2421,N_2281);
nand U2627 (N_2627,N_2190,N_2414);
and U2628 (N_2628,N_2055,N_2207);
nor U2629 (N_2629,N_2004,N_2388);
nor U2630 (N_2630,N_2235,N_2327);
or U2631 (N_2631,N_2326,N_2370);
and U2632 (N_2632,N_2229,N_2305);
and U2633 (N_2633,N_2451,N_2135);
nand U2634 (N_2634,N_2195,N_2431);
xor U2635 (N_2635,N_2345,N_2286);
xor U2636 (N_2636,N_2242,N_2156);
and U2637 (N_2637,N_2426,N_2003);
or U2638 (N_2638,N_2392,N_2338);
and U2639 (N_2639,N_2020,N_2304);
nor U2640 (N_2640,N_2211,N_2202);
xor U2641 (N_2641,N_2259,N_2204);
or U2642 (N_2642,N_2349,N_2410);
or U2643 (N_2643,N_2164,N_2043);
or U2644 (N_2644,N_2409,N_2462);
or U2645 (N_2645,N_2382,N_2085);
nand U2646 (N_2646,N_2456,N_2236);
and U2647 (N_2647,N_2103,N_2051);
nor U2648 (N_2648,N_2311,N_2359);
nor U2649 (N_2649,N_2170,N_2097);
nor U2650 (N_2650,N_2464,N_2298);
nor U2651 (N_2651,N_2441,N_2473);
nor U2652 (N_2652,N_2234,N_2089);
and U2653 (N_2653,N_2075,N_2139);
and U2654 (N_2654,N_2248,N_2101);
and U2655 (N_2655,N_2371,N_2146);
nor U2656 (N_2656,N_2336,N_2292);
or U2657 (N_2657,N_2112,N_2106);
or U2658 (N_2658,N_2182,N_2216);
nor U2659 (N_2659,N_2070,N_2256);
or U2660 (N_2660,N_2208,N_2080);
nor U2661 (N_2661,N_2403,N_2427);
or U2662 (N_2662,N_2318,N_2189);
nand U2663 (N_2663,N_2108,N_2381);
or U2664 (N_2664,N_2273,N_2068);
nor U2665 (N_2665,N_2002,N_2488);
nand U2666 (N_2666,N_2117,N_2384);
or U2667 (N_2667,N_2022,N_2481);
and U2668 (N_2668,N_2470,N_2317);
nor U2669 (N_2669,N_2424,N_2005);
or U2670 (N_2670,N_2176,N_2167);
nand U2671 (N_2671,N_2086,N_2206);
or U2672 (N_2672,N_2018,N_2352);
xor U2673 (N_2673,N_2257,N_2134);
nor U2674 (N_2674,N_2455,N_2302);
nand U2675 (N_2675,N_2291,N_2378);
nand U2676 (N_2676,N_2366,N_2353);
nand U2677 (N_2677,N_2119,N_2095);
or U2678 (N_2678,N_2390,N_2016);
nand U2679 (N_2679,N_2363,N_2374);
nand U2680 (N_2680,N_2154,N_2150);
xnor U2681 (N_2681,N_2030,N_2091);
and U2682 (N_2682,N_2151,N_2184);
and U2683 (N_2683,N_2377,N_2056);
and U2684 (N_2684,N_2083,N_2344);
nor U2685 (N_2685,N_2011,N_2498);
nor U2686 (N_2686,N_2394,N_2024);
or U2687 (N_2687,N_2474,N_2262);
nor U2688 (N_2688,N_2200,N_2137);
nor U2689 (N_2689,N_2308,N_2453);
nor U2690 (N_2690,N_2141,N_2192);
or U2691 (N_2691,N_2087,N_2258);
nor U2692 (N_2692,N_2001,N_2160);
and U2693 (N_2693,N_2249,N_2049);
nor U2694 (N_2694,N_2092,N_2082);
or U2695 (N_2695,N_2275,N_2289);
xor U2696 (N_2696,N_2048,N_2224);
and U2697 (N_2697,N_2310,N_2279);
nand U2698 (N_2698,N_2036,N_2420);
or U2699 (N_2699,N_2365,N_2220);
or U2700 (N_2700,N_2497,N_2491);
or U2701 (N_2701,N_2179,N_2434);
nor U2702 (N_2702,N_2118,N_2274);
and U2703 (N_2703,N_2288,N_2297);
or U2704 (N_2704,N_2128,N_2457);
nand U2705 (N_2705,N_2203,N_2058);
or U2706 (N_2706,N_2077,N_2152);
nand U2707 (N_2707,N_2130,N_2276);
or U2708 (N_2708,N_2369,N_2313);
nor U2709 (N_2709,N_2342,N_2163);
or U2710 (N_2710,N_2188,N_2060);
or U2711 (N_2711,N_2168,N_2332);
and U2712 (N_2712,N_2107,N_2174);
and U2713 (N_2713,N_2079,N_2034);
and U2714 (N_2714,N_2402,N_2111);
or U2715 (N_2715,N_2029,N_2312);
nand U2716 (N_2716,N_2449,N_2222);
nor U2717 (N_2717,N_2247,N_2067);
or U2718 (N_2718,N_2439,N_2265);
or U2719 (N_2719,N_2000,N_2009);
or U2720 (N_2720,N_2054,N_2078);
nor U2721 (N_2721,N_2090,N_2241);
or U2722 (N_2722,N_2026,N_2351);
or U2723 (N_2723,N_2267,N_2269);
and U2724 (N_2724,N_2175,N_2102);
nand U2725 (N_2725,N_2120,N_2316);
and U2726 (N_2726,N_2122,N_2013);
nand U2727 (N_2727,N_2425,N_2476);
nor U2728 (N_2728,N_2073,N_2132);
nor U2729 (N_2729,N_2373,N_2066);
or U2730 (N_2730,N_2433,N_2021);
and U2731 (N_2731,N_2300,N_2499);
or U2732 (N_2732,N_2062,N_2458);
or U2733 (N_2733,N_2380,N_2395);
nand U2734 (N_2734,N_2084,N_2379);
nor U2735 (N_2735,N_2430,N_2041);
nand U2736 (N_2736,N_2053,N_2280);
or U2737 (N_2737,N_2140,N_2463);
nor U2738 (N_2738,N_2197,N_2436);
nand U2739 (N_2739,N_2014,N_2329);
nor U2740 (N_2740,N_2450,N_2131);
or U2741 (N_2741,N_2191,N_2069);
and U2742 (N_2742,N_2397,N_2246);
and U2743 (N_2743,N_2209,N_2254);
and U2744 (N_2744,N_2057,N_2173);
nor U2745 (N_2745,N_2442,N_2240);
nor U2746 (N_2746,N_2419,N_2228);
nand U2747 (N_2747,N_2205,N_2287);
nor U2748 (N_2748,N_2125,N_2445);
or U2749 (N_2749,N_2416,N_2148);
nor U2750 (N_2750,N_2332,N_2157);
xnor U2751 (N_2751,N_2102,N_2142);
and U2752 (N_2752,N_2079,N_2319);
and U2753 (N_2753,N_2207,N_2040);
or U2754 (N_2754,N_2248,N_2298);
nand U2755 (N_2755,N_2334,N_2205);
and U2756 (N_2756,N_2308,N_2484);
nor U2757 (N_2757,N_2448,N_2278);
nor U2758 (N_2758,N_2153,N_2441);
or U2759 (N_2759,N_2316,N_2257);
or U2760 (N_2760,N_2389,N_2483);
nand U2761 (N_2761,N_2186,N_2313);
nor U2762 (N_2762,N_2467,N_2264);
and U2763 (N_2763,N_2398,N_2176);
and U2764 (N_2764,N_2082,N_2203);
or U2765 (N_2765,N_2342,N_2048);
or U2766 (N_2766,N_2277,N_2088);
nand U2767 (N_2767,N_2283,N_2093);
or U2768 (N_2768,N_2455,N_2346);
nor U2769 (N_2769,N_2056,N_2165);
xnor U2770 (N_2770,N_2007,N_2470);
and U2771 (N_2771,N_2137,N_2378);
nand U2772 (N_2772,N_2447,N_2034);
or U2773 (N_2773,N_2315,N_2233);
nand U2774 (N_2774,N_2054,N_2297);
or U2775 (N_2775,N_2406,N_2173);
nand U2776 (N_2776,N_2265,N_2078);
or U2777 (N_2777,N_2318,N_2365);
and U2778 (N_2778,N_2105,N_2056);
nor U2779 (N_2779,N_2013,N_2356);
nand U2780 (N_2780,N_2215,N_2366);
nor U2781 (N_2781,N_2465,N_2431);
or U2782 (N_2782,N_2262,N_2087);
nand U2783 (N_2783,N_2159,N_2006);
and U2784 (N_2784,N_2372,N_2029);
nor U2785 (N_2785,N_2376,N_2184);
nand U2786 (N_2786,N_2028,N_2174);
nand U2787 (N_2787,N_2081,N_2101);
xnor U2788 (N_2788,N_2273,N_2026);
nand U2789 (N_2789,N_2378,N_2359);
or U2790 (N_2790,N_2148,N_2381);
or U2791 (N_2791,N_2288,N_2444);
nand U2792 (N_2792,N_2385,N_2458);
and U2793 (N_2793,N_2141,N_2332);
and U2794 (N_2794,N_2316,N_2402);
or U2795 (N_2795,N_2034,N_2284);
nand U2796 (N_2796,N_2133,N_2307);
or U2797 (N_2797,N_2106,N_2088);
nand U2798 (N_2798,N_2424,N_2190);
nor U2799 (N_2799,N_2344,N_2452);
or U2800 (N_2800,N_2179,N_2203);
xnor U2801 (N_2801,N_2409,N_2303);
and U2802 (N_2802,N_2489,N_2327);
or U2803 (N_2803,N_2232,N_2449);
or U2804 (N_2804,N_2432,N_2301);
or U2805 (N_2805,N_2345,N_2090);
or U2806 (N_2806,N_2057,N_2443);
nand U2807 (N_2807,N_2466,N_2270);
nor U2808 (N_2808,N_2259,N_2361);
nand U2809 (N_2809,N_2351,N_2402);
nor U2810 (N_2810,N_2223,N_2455);
nor U2811 (N_2811,N_2341,N_2404);
xnor U2812 (N_2812,N_2292,N_2463);
and U2813 (N_2813,N_2477,N_2122);
nor U2814 (N_2814,N_2087,N_2193);
and U2815 (N_2815,N_2262,N_2060);
nand U2816 (N_2816,N_2318,N_2120);
xor U2817 (N_2817,N_2342,N_2379);
and U2818 (N_2818,N_2332,N_2114);
or U2819 (N_2819,N_2475,N_2301);
xor U2820 (N_2820,N_2043,N_2266);
nand U2821 (N_2821,N_2250,N_2013);
or U2822 (N_2822,N_2421,N_2278);
nand U2823 (N_2823,N_2228,N_2176);
xnor U2824 (N_2824,N_2371,N_2225);
or U2825 (N_2825,N_2377,N_2393);
nand U2826 (N_2826,N_2268,N_2168);
or U2827 (N_2827,N_2489,N_2027);
or U2828 (N_2828,N_2343,N_2054);
nand U2829 (N_2829,N_2082,N_2074);
and U2830 (N_2830,N_2354,N_2377);
nand U2831 (N_2831,N_2110,N_2055);
xor U2832 (N_2832,N_2265,N_2131);
nor U2833 (N_2833,N_2328,N_2319);
nor U2834 (N_2834,N_2349,N_2301);
nor U2835 (N_2835,N_2211,N_2140);
nand U2836 (N_2836,N_2286,N_2089);
nand U2837 (N_2837,N_2176,N_2464);
nor U2838 (N_2838,N_2003,N_2436);
xor U2839 (N_2839,N_2415,N_2189);
nand U2840 (N_2840,N_2315,N_2041);
xor U2841 (N_2841,N_2477,N_2456);
or U2842 (N_2842,N_2457,N_2024);
or U2843 (N_2843,N_2202,N_2174);
nand U2844 (N_2844,N_2373,N_2315);
and U2845 (N_2845,N_2166,N_2444);
or U2846 (N_2846,N_2480,N_2278);
xor U2847 (N_2847,N_2308,N_2298);
and U2848 (N_2848,N_2372,N_2245);
and U2849 (N_2849,N_2476,N_2201);
nor U2850 (N_2850,N_2107,N_2447);
nor U2851 (N_2851,N_2244,N_2308);
nand U2852 (N_2852,N_2282,N_2216);
or U2853 (N_2853,N_2419,N_2408);
and U2854 (N_2854,N_2059,N_2467);
nor U2855 (N_2855,N_2212,N_2039);
and U2856 (N_2856,N_2462,N_2395);
nand U2857 (N_2857,N_2135,N_2213);
and U2858 (N_2858,N_2081,N_2408);
and U2859 (N_2859,N_2387,N_2096);
nand U2860 (N_2860,N_2108,N_2143);
nor U2861 (N_2861,N_2124,N_2072);
and U2862 (N_2862,N_2220,N_2232);
xnor U2863 (N_2863,N_2074,N_2243);
nor U2864 (N_2864,N_2471,N_2469);
nor U2865 (N_2865,N_2011,N_2140);
nand U2866 (N_2866,N_2458,N_2396);
xnor U2867 (N_2867,N_2129,N_2208);
and U2868 (N_2868,N_2368,N_2434);
or U2869 (N_2869,N_2054,N_2088);
nor U2870 (N_2870,N_2406,N_2286);
nor U2871 (N_2871,N_2029,N_2068);
nor U2872 (N_2872,N_2409,N_2249);
nor U2873 (N_2873,N_2445,N_2468);
xnor U2874 (N_2874,N_2114,N_2422);
xor U2875 (N_2875,N_2033,N_2191);
or U2876 (N_2876,N_2259,N_2293);
nor U2877 (N_2877,N_2096,N_2020);
and U2878 (N_2878,N_2423,N_2384);
nor U2879 (N_2879,N_2023,N_2211);
nand U2880 (N_2880,N_2355,N_2474);
nor U2881 (N_2881,N_2486,N_2065);
nor U2882 (N_2882,N_2119,N_2251);
nor U2883 (N_2883,N_2096,N_2073);
or U2884 (N_2884,N_2312,N_2147);
nor U2885 (N_2885,N_2124,N_2468);
and U2886 (N_2886,N_2201,N_2078);
xnor U2887 (N_2887,N_2182,N_2386);
nand U2888 (N_2888,N_2156,N_2259);
nor U2889 (N_2889,N_2058,N_2463);
nor U2890 (N_2890,N_2044,N_2065);
xor U2891 (N_2891,N_2203,N_2266);
xnor U2892 (N_2892,N_2041,N_2400);
nand U2893 (N_2893,N_2147,N_2479);
and U2894 (N_2894,N_2316,N_2239);
and U2895 (N_2895,N_2268,N_2183);
nor U2896 (N_2896,N_2432,N_2048);
nand U2897 (N_2897,N_2031,N_2242);
or U2898 (N_2898,N_2218,N_2458);
nand U2899 (N_2899,N_2349,N_2251);
nand U2900 (N_2900,N_2051,N_2168);
and U2901 (N_2901,N_2073,N_2285);
nand U2902 (N_2902,N_2098,N_2382);
or U2903 (N_2903,N_2028,N_2293);
and U2904 (N_2904,N_2037,N_2152);
nand U2905 (N_2905,N_2144,N_2150);
and U2906 (N_2906,N_2075,N_2071);
or U2907 (N_2907,N_2258,N_2131);
nor U2908 (N_2908,N_2095,N_2429);
and U2909 (N_2909,N_2357,N_2310);
nand U2910 (N_2910,N_2440,N_2279);
and U2911 (N_2911,N_2450,N_2142);
and U2912 (N_2912,N_2177,N_2248);
and U2913 (N_2913,N_2183,N_2069);
nand U2914 (N_2914,N_2119,N_2489);
nand U2915 (N_2915,N_2335,N_2475);
nand U2916 (N_2916,N_2176,N_2098);
nor U2917 (N_2917,N_2285,N_2143);
or U2918 (N_2918,N_2499,N_2137);
nor U2919 (N_2919,N_2234,N_2235);
or U2920 (N_2920,N_2491,N_2347);
or U2921 (N_2921,N_2291,N_2362);
and U2922 (N_2922,N_2344,N_2332);
nand U2923 (N_2923,N_2084,N_2470);
xnor U2924 (N_2924,N_2489,N_2339);
nand U2925 (N_2925,N_2100,N_2183);
and U2926 (N_2926,N_2268,N_2372);
or U2927 (N_2927,N_2462,N_2365);
nor U2928 (N_2928,N_2113,N_2229);
nor U2929 (N_2929,N_2433,N_2461);
nor U2930 (N_2930,N_2401,N_2446);
and U2931 (N_2931,N_2029,N_2479);
and U2932 (N_2932,N_2023,N_2253);
and U2933 (N_2933,N_2104,N_2355);
or U2934 (N_2934,N_2337,N_2322);
or U2935 (N_2935,N_2209,N_2384);
nand U2936 (N_2936,N_2249,N_2210);
nor U2937 (N_2937,N_2321,N_2323);
or U2938 (N_2938,N_2397,N_2191);
xnor U2939 (N_2939,N_2009,N_2028);
or U2940 (N_2940,N_2324,N_2227);
or U2941 (N_2941,N_2163,N_2449);
and U2942 (N_2942,N_2415,N_2134);
nand U2943 (N_2943,N_2240,N_2293);
or U2944 (N_2944,N_2041,N_2342);
nor U2945 (N_2945,N_2164,N_2256);
nand U2946 (N_2946,N_2302,N_2280);
xnor U2947 (N_2947,N_2104,N_2163);
and U2948 (N_2948,N_2056,N_2128);
nor U2949 (N_2949,N_2023,N_2475);
nor U2950 (N_2950,N_2434,N_2349);
and U2951 (N_2951,N_2149,N_2431);
nor U2952 (N_2952,N_2041,N_2062);
nor U2953 (N_2953,N_2358,N_2141);
or U2954 (N_2954,N_2216,N_2199);
xnor U2955 (N_2955,N_2403,N_2480);
and U2956 (N_2956,N_2373,N_2388);
nor U2957 (N_2957,N_2409,N_2225);
nor U2958 (N_2958,N_2087,N_2283);
and U2959 (N_2959,N_2438,N_2361);
nor U2960 (N_2960,N_2207,N_2396);
and U2961 (N_2961,N_2288,N_2324);
nand U2962 (N_2962,N_2393,N_2418);
nand U2963 (N_2963,N_2368,N_2207);
nor U2964 (N_2964,N_2436,N_2351);
xor U2965 (N_2965,N_2171,N_2374);
nor U2966 (N_2966,N_2279,N_2220);
nand U2967 (N_2967,N_2148,N_2179);
nand U2968 (N_2968,N_2267,N_2089);
nand U2969 (N_2969,N_2095,N_2416);
and U2970 (N_2970,N_2412,N_2402);
and U2971 (N_2971,N_2426,N_2311);
and U2972 (N_2972,N_2439,N_2351);
and U2973 (N_2973,N_2065,N_2032);
or U2974 (N_2974,N_2039,N_2294);
or U2975 (N_2975,N_2023,N_2442);
nor U2976 (N_2976,N_2123,N_2352);
or U2977 (N_2977,N_2346,N_2039);
nand U2978 (N_2978,N_2063,N_2354);
nand U2979 (N_2979,N_2179,N_2402);
and U2980 (N_2980,N_2456,N_2280);
nor U2981 (N_2981,N_2233,N_2327);
nor U2982 (N_2982,N_2314,N_2239);
and U2983 (N_2983,N_2459,N_2471);
and U2984 (N_2984,N_2204,N_2095);
nand U2985 (N_2985,N_2174,N_2463);
nor U2986 (N_2986,N_2164,N_2435);
or U2987 (N_2987,N_2296,N_2434);
xnor U2988 (N_2988,N_2462,N_2011);
or U2989 (N_2989,N_2008,N_2149);
nand U2990 (N_2990,N_2347,N_2053);
or U2991 (N_2991,N_2168,N_2220);
or U2992 (N_2992,N_2090,N_2190);
nor U2993 (N_2993,N_2362,N_2118);
nand U2994 (N_2994,N_2090,N_2139);
and U2995 (N_2995,N_2493,N_2108);
nor U2996 (N_2996,N_2319,N_2234);
xor U2997 (N_2997,N_2002,N_2221);
nor U2998 (N_2998,N_2332,N_2266);
or U2999 (N_2999,N_2236,N_2415);
and U3000 (N_3000,N_2564,N_2632);
nand U3001 (N_3001,N_2706,N_2927);
nor U3002 (N_3002,N_2704,N_2579);
nor U3003 (N_3003,N_2533,N_2872);
or U3004 (N_3004,N_2532,N_2740);
and U3005 (N_3005,N_2785,N_2646);
or U3006 (N_3006,N_2589,N_2879);
or U3007 (N_3007,N_2655,N_2771);
nand U3008 (N_3008,N_2814,N_2778);
nand U3009 (N_3009,N_2698,N_2701);
nor U3010 (N_3010,N_2866,N_2898);
nand U3011 (N_3011,N_2587,N_2851);
and U3012 (N_3012,N_2958,N_2604);
or U3013 (N_3013,N_2614,N_2743);
nor U3014 (N_3014,N_2984,N_2877);
nand U3015 (N_3015,N_2858,N_2748);
nand U3016 (N_3016,N_2934,N_2810);
and U3017 (N_3017,N_2702,N_2730);
or U3018 (N_3018,N_2721,N_2765);
or U3019 (N_3019,N_2691,N_2925);
nand U3020 (N_3020,N_2912,N_2825);
nor U3021 (N_3021,N_2525,N_2878);
or U3022 (N_3022,N_2648,N_2507);
or U3023 (N_3023,N_2959,N_2857);
xor U3024 (N_3024,N_2513,N_2869);
xnor U3025 (N_3025,N_2907,N_2895);
or U3026 (N_3026,N_2913,N_2852);
or U3027 (N_3027,N_2804,N_2742);
nor U3028 (N_3028,N_2696,N_2952);
or U3029 (N_3029,N_2617,N_2954);
nor U3030 (N_3030,N_2900,N_2733);
nor U3031 (N_3031,N_2839,N_2893);
nand U3032 (N_3032,N_2968,N_2591);
nand U3033 (N_3033,N_2574,N_2874);
or U3034 (N_3034,N_2552,N_2654);
xnor U3035 (N_3035,N_2961,N_2974);
and U3036 (N_3036,N_2556,N_2642);
and U3037 (N_3037,N_2714,N_2571);
nor U3038 (N_3038,N_2658,N_2528);
or U3039 (N_3039,N_2668,N_2670);
and U3040 (N_3040,N_2559,N_2826);
or U3041 (N_3041,N_2685,N_2786);
nor U3042 (N_3042,N_2752,N_2787);
or U3043 (N_3043,N_2505,N_2745);
and U3044 (N_3044,N_2833,N_2626);
and U3045 (N_3045,N_2982,N_2883);
nor U3046 (N_3046,N_2988,N_2682);
nand U3047 (N_3047,N_2817,N_2942);
and U3048 (N_3048,N_2590,N_2502);
xnor U3049 (N_3049,N_2763,N_2815);
and U3050 (N_3050,N_2803,N_2845);
nand U3051 (N_3051,N_2792,N_2791);
nand U3052 (N_3052,N_2676,N_2754);
and U3053 (N_3053,N_2534,N_2977);
and U3054 (N_3054,N_2797,N_2636);
or U3055 (N_3055,N_2768,N_2660);
and U3056 (N_3056,N_2821,N_2688);
nand U3057 (N_3057,N_2638,N_2910);
and U3058 (N_3058,N_2728,N_2541);
nand U3059 (N_3059,N_2635,N_2863);
xor U3060 (N_3060,N_2920,N_2527);
and U3061 (N_3061,N_2715,N_2592);
or U3062 (N_3062,N_2609,N_2530);
or U3063 (N_3063,N_2819,N_2630);
or U3064 (N_3064,N_2669,N_2756);
nand U3065 (N_3065,N_2949,N_2567);
nand U3066 (N_3066,N_2653,N_2948);
and U3067 (N_3067,N_2856,N_2849);
xor U3068 (N_3068,N_2842,N_2508);
and U3069 (N_3069,N_2601,N_2649);
or U3070 (N_3070,N_2569,N_2985);
nand U3071 (N_3071,N_2549,N_2906);
nand U3072 (N_3072,N_2725,N_2724);
and U3073 (N_3073,N_2750,N_2511);
nand U3074 (N_3074,N_2562,N_2599);
nor U3075 (N_3075,N_2773,N_2554);
or U3076 (N_3076,N_2557,N_2572);
nor U3077 (N_3077,N_2551,N_2506);
xor U3078 (N_3078,N_2894,N_2995);
nor U3079 (N_3079,N_2627,N_2739);
xor U3080 (N_3080,N_2620,N_2521);
nor U3081 (N_3081,N_2844,N_2924);
nand U3082 (N_3082,N_2686,N_2841);
xor U3083 (N_3083,N_2998,N_2713);
nor U3084 (N_3084,N_2707,N_2994);
xnor U3085 (N_3085,N_2529,N_2767);
xnor U3086 (N_3086,N_2608,N_2890);
or U3087 (N_3087,N_2840,N_2902);
xor U3088 (N_3088,N_2602,N_2595);
and U3089 (N_3089,N_2624,N_2770);
and U3090 (N_3090,N_2918,N_2618);
and U3091 (N_3091,N_2662,N_2736);
xnor U3092 (N_3092,N_2885,N_2899);
and U3093 (N_3093,N_2990,N_2711);
or U3094 (N_3094,N_2975,N_2518);
nor U3095 (N_3095,N_2989,N_2776);
nor U3096 (N_3096,N_2594,N_2846);
nand U3097 (N_3097,N_2999,N_2577);
xor U3098 (N_3098,N_2809,N_2903);
and U3099 (N_3099,N_2689,N_2760);
or U3100 (N_3100,N_2876,N_2573);
or U3101 (N_3101,N_2798,N_2970);
nand U3102 (N_3102,N_2789,N_2867);
or U3103 (N_3103,N_2848,N_2645);
nor U3104 (N_3104,N_2526,N_2873);
xnor U3105 (N_3105,N_2586,N_2880);
nor U3106 (N_3106,N_2517,N_2565);
and U3107 (N_3107,N_2794,N_2811);
nand U3108 (N_3108,N_2500,N_2911);
and U3109 (N_3109,N_2629,N_2853);
nor U3110 (N_3110,N_2611,N_2619);
and U3111 (N_3111,N_2650,N_2523);
nor U3112 (N_3112,N_2991,N_2746);
nand U3113 (N_3113,N_2687,N_2621);
nor U3114 (N_3114,N_2788,N_2566);
nand U3115 (N_3115,N_2932,N_2663);
nor U3116 (N_3116,N_2580,N_2610);
and U3117 (N_3117,N_2919,N_2545);
nor U3118 (N_3118,N_2824,N_2836);
nor U3119 (N_3119,N_2922,N_2537);
xnor U3120 (N_3120,N_2812,N_2993);
nor U3121 (N_3121,N_2539,N_2855);
or U3122 (N_3122,N_2757,N_2967);
and U3123 (N_3123,N_2940,N_2973);
and U3124 (N_3124,N_2928,N_2795);
nand U3125 (N_3125,N_2625,N_2875);
and U3126 (N_3126,N_2909,N_2700);
and U3127 (N_3127,N_2941,N_2615);
xnor U3128 (N_3128,N_2931,N_2892);
or U3129 (N_3129,N_2923,N_2901);
xor U3130 (N_3130,N_2695,N_2504);
nor U3131 (N_3131,N_2865,N_2980);
nand U3132 (N_3132,N_2677,N_2543);
and U3133 (N_3133,N_2584,N_2963);
or U3134 (N_3134,N_2732,N_2829);
nor U3135 (N_3135,N_2777,N_2503);
xnor U3136 (N_3136,N_2753,N_2678);
nand U3137 (N_3137,N_2761,N_2807);
and U3138 (N_3138,N_2956,N_2850);
or U3139 (N_3139,N_2960,N_2697);
and U3140 (N_3140,N_2806,N_2664);
and U3141 (N_3141,N_2652,N_2986);
or U3142 (N_3142,N_2926,N_2884);
nor U3143 (N_3143,N_2515,N_2782);
or U3144 (N_3144,N_2593,N_2957);
nor U3145 (N_3145,N_2764,N_2690);
nor U3146 (N_3146,N_2780,N_2738);
and U3147 (N_3147,N_2886,N_2675);
or U3148 (N_3148,N_2553,N_2955);
nand U3149 (N_3149,N_2981,N_2633);
xor U3150 (N_3150,N_2783,N_2860);
or U3151 (N_3151,N_2870,N_2978);
or U3152 (N_3152,N_2943,N_2656);
or U3153 (N_3153,N_2800,N_2935);
or U3154 (N_3154,N_2813,N_2613);
nand U3155 (N_3155,N_2607,N_2827);
or U3156 (N_3156,N_2921,N_2692);
nand U3157 (N_3157,N_2801,N_2510);
and U3158 (N_3158,N_2908,N_2712);
nor U3159 (N_3159,N_2847,N_2772);
nand U3160 (N_3160,N_2519,N_2759);
nand U3161 (N_3161,N_2637,N_2904);
nor U3162 (N_3162,N_2734,N_2583);
or U3163 (N_3163,N_2622,N_2679);
nor U3164 (N_3164,N_2996,N_2570);
nor U3165 (N_3165,N_2843,N_2735);
xnor U3166 (N_3166,N_2634,N_2945);
or U3167 (N_3167,N_2936,N_2501);
and U3168 (N_3168,N_2699,N_2747);
nor U3169 (N_3169,N_2681,N_2784);
nor U3170 (N_3170,N_2522,N_2540);
nand U3171 (N_3171,N_2775,N_2793);
nand U3172 (N_3172,N_2603,N_2914);
and U3173 (N_3173,N_2966,N_2969);
nand U3174 (N_3174,N_2758,N_2558);
or U3175 (N_3175,N_2640,N_2716);
nor U3176 (N_3176,N_2972,N_2520);
nand U3177 (N_3177,N_2983,N_2944);
nor U3178 (N_3178,N_2965,N_2717);
nand U3179 (N_3179,N_2805,N_2727);
nor U3180 (N_3180,N_2644,N_2612);
or U3181 (N_3181,N_2799,N_2672);
nand U3182 (N_3182,N_2744,N_2871);
nand U3183 (N_3183,N_2762,N_2751);
or U3184 (N_3184,N_2830,N_2544);
and U3185 (N_3185,N_2888,N_2661);
nand U3186 (N_3186,N_2524,N_2823);
and U3187 (N_3187,N_2997,N_2937);
nand U3188 (N_3188,N_2719,N_2693);
and U3189 (N_3189,N_2828,N_2684);
or U3190 (N_3190,N_2673,N_2889);
and U3191 (N_3191,N_2731,N_2838);
nor U3192 (N_3192,N_2561,N_2651);
and U3193 (N_3193,N_2516,N_2512);
or U3194 (N_3194,N_2887,N_2818);
or U3195 (N_3195,N_2915,N_2837);
or U3196 (N_3196,N_2623,N_2546);
and U3197 (N_3197,N_2709,N_2929);
nand U3198 (N_3198,N_2581,N_2816);
nor U3199 (N_3199,N_2971,N_2683);
or U3200 (N_3200,N_2962,N_2694);
xor U3201 (N_3201,N_2930,N_2596);
nand U3202 (N_3202,N_2665,N_2769);
or U3203 (N_3203,N_2862,N_2514);
nor U3204 (N_3204,N_2868,N_2864);
or U3205 (N_3205,N_2779,N_2835);
or U3206 (N_3206,N_2951,N_2938);
xor U3207 (N_3207,N_2859,N_2939);
or U3208 (N_3208,N_2953,N_2796);
nand U3209 (N_3209,N_2703,N_2891);
nor U3210 (N_3210,N_2832,N_2737);
nand U3211 (N_3211,N_2597,N_2536);
or U3212 (N_3212,N_2588,N_2905);
and U3213 (N_3213,N_2950,N_2987);
and U3214 (N_3214,N_2979,N_2535);
nor U3215 (N_3215,N_2741,N_2560);
nor U3216 (N_3216,N_2834,N_2946);
nand U3217 (N_3217,N_2710,N_2643);
xnor U3218 (N_3218,N_2947,N_2820);
and U3219 (N_3219,N_2933,N_2831);
and U3220 (N_3220,N_2585,N_2726);
and U3221 (N_3221,N_2749,N_2578);
and U3222 (N_3222,N_2657,N_2550);
nor U3223 (N_3223,N_2666,N_2755);
xor U3224 (N_3224,N_2854,N_2671);
and U3225 (N_3225,N_2917,N_2722);
nor U3226 (N_3226,N_2606,N_2729);
nand U3227 (N_3227,N_2639,N_2509);
and U3228 (N_3228,N_2659,N_2531);
and U3229 (N_3229,N_2674,N_2774);
nor U3230 (N_3230,N_2616,N_2822);
and U3231 (N_3231,N_2897,N_2600);
or U3232 (N_3232,N_2882,N_2542);
or U3233 (N_3233,N_2802,N_2568);
and U3234 (N_3234,N_2628,N_2766);
nor U3235 (N_3235,N_2631,N_2720);
or U3236 (N_3236,N_2548,N_2861);
and U3237 (N_3237,N_2916,N_2598);
nand U3238 (N_3238,N_2563,N_2575);
nor U3239 (N_3239,N_2667,N_2881);
nand U3240 (N_3240,N_2605,N_2708);
nor U3241 (N_3241,N_2705,N_2547);
xor U3242 (N_3242,N_2896,N_2555);
nand U3243 (N_3243,N_2582,N_2976);
nor U3244 (N_3244,N_2718,N_2576);
nor U3245 (N_3245,N_2538,N_2647);
or U3246 (N_3246,N_2808,N_2992);
or U3247 (N_3247,N_2723,N_2964);
xor U3248 (N_3248,N_2781,N_2790);
nand U3249 (N_3249,N_2680,N_2641);
nand U3250 (N_3250,N_2714,N_2646);
or U3251 (N_3251,N_2994,N_2634);
nand U3252 (N_3252,N_2883,N_2607);
or U3253 (N_3253,N_2560,N_2808);
nor U3254 (N_3254,N_2903,N_2741);
and U3255 (N_3255,N_2895,N_2796);
and U3256 (N_3256,N_2857,N_2894);
and U3257 (N_3257,N_2656,N_2559);
and U3258 (N_3258,N_2852,N_2740);
nand U3259 (N_3259,N_2834,N_2907);
nor U3260 (N_3260,N_2573,N_2740);
nand U3261 (N_3261,N_2717,N_2560);
and U3262 (N_3262,N_2695,N_2548);
and U3263 (N_3263,N_2966,N_2849);
or U3264 (N_3264,N_2672,N_2509);
nor U3265 (N_3265,N_2694,N_2569);
xor U3266 (N_3266,N_2831,N_2967);
and U3267 (N_3267,N_2788,N_2906);
or U3268 (N_3268,N_2548,N_2565);
and U3269 (N_3269,N_2599,N_2865);
nor U3270 (N_3270,N_2829,N_2736);
and U3271 (N_3271,N_2903,N_2607);
nand U3272 (N_3272,N_2560,N_2712);
or U3273 (N_3273,N_2519,N_2843);
or U3274 (N_3274,N_2819,N_2712);
nand U3275 (N_3275,N_2650,N_2937);
xor U3276 (N_3276,N_2527,N_2540);
and U3277 (N_3277,N_2528,N_2836);
nor U3278 (N_3278,N_2795,N_2505);
nand U3279 (N_3279,N_2774,N_2804);
and U3280 (N_3280,N_2588,N_2814);
nor U3281 (N_3281,N_2613,N_2721);
nor U3282 (N_3282,N_2951,N_2663);
nor U3283 (N_3283,N_2617,N_2509);
nand U3284 (N_3284,N_2863,N_2607);
and U3285 (N_3285,N_2878,N_2734);
nand U3286 (N_3286,N_2683,N_2650);
nor U3287 (N_3287,N_2857,N_2662);
nand U3288 (N_3288,N_2836,N_2749);
and U3289 (N_3289,N_2975,N_2783);
and U3290 (N_3290,N_2936,N_2941);
or U3291 (N_3291,N_2740,N_2689);
nor U3292 (N_3292,N_2819,N_2617);
or U3293 (N_3293,N_2911,N_2906);
nor U3294 (N_3294,N_2792,N_2601);
or U3295 (N_3295,N_2576,N_2971);
nor U3296 (N_3296,N_2526,N_2960);
or U3297 (N_3297,N_2508,N_2757);
or U3298 (N_3298,N_2700,N_2678);
nor U3299 (N_3299,N_2770,N_2573);
or U3300 (N_3300,N_2710,N_2635);
or U3301 (N_3301,N_2696,N_2852);
nor U3302 (N_3302,N_2831,N_2888);
and U3303 (N_3303,N_2930,N_2544);
nand U3304 (N_3304,N_2804,N_2981);
nor U3305 (N_3305,N_2970,N_2987);
and U3306 (N_3306,N_2929,N_2827);
and U3307 (N_3307,N_2857,N_2766);
xnor U3308 (N_3308,N_2604,N_2880);
nor U3309 (N_3309,N_2923,N_2940);
or U3310 (N_3310,N_2545,N_2566);
nand U3311 (N_3311,N_2941,N_2639);
and U3312 (N_3312,N_2654,N_2780);
nand U3313 (N_3313,N_2616,N_2854);
and U3314 (N_3314,N_2644,N_2590);
nand U3315 (N_3315,N_2758,N_2723);
nand U3316 (N_3316,N_2757,N_2619);
nand U3317 (N_3317,N_2517,N_2889);
nor U3318 (N_3318,N_2783,N_2822);
xor U3319 (N_3319,N_2708,N_2948);
and U3320 (N_3320,N_2762,N_2781);
nand U3321 (N_3321,N_2989,N_2962);
and U3322 (N_3322,N_2784,N_2765);
and U3323 (N_3323,N_2546,N_2960);
nand U3324 (N_3324,N_2709,N_2512);
or U3325 (N_3325,N_2808,N_2580);
and U3326 (N_3326,N_2619,N_2813);
and U3327 (N_3327,N_2740,N_2759);
nand U3328 (N_3328,N_2639,N_2883);
nand U3329 (N_3329,N_2621,N_2534);
nor U3330 (N_3330,N_2681,N_2684);
xor U3331 (N_3331,N_2741,N_2841);
and U3332 (N_3332,N_2836,N_2530);
nor U3333 (N_3333,N_2981,N_2596);
or U3334 (N_3334,N_2892,N_2651);
nand U3335 (N_3335,N_2671,N_2935);
and U3336 (N_3336,N_2930,N_2834);
nand U3337 (N_3337,N_2666,N_2858);
nor U3338 (N_3338,N_2782,N_2956);
and U3339 (N_3339,N_2553,N_2506);
nand U3340 (N_3340,N_2765,N_2600);
nor U3341 (N_3341,N_2543,N_2933);
xor U3342 (N_3342,N_2644,N_2684);
and U3343 (N_3343,N_2515,N_2679);
xor U3344 (N_3344,N_2801,N_2858);
or U3345 (N_3345,N_2937,N_2691);
nor U3346 (N_3346,N_2775,N_2719);
and U3347 (N_3347,N_2896,N_2919);
and U3348 (N_3348,N_2766,N_2639);
or U3349 (N_3349,N_2504,N_2904);
xor U3350 (N_3350,N_2868,N_2597);
nand U3351 (N_3351,N_2815,N_2692);
and U3352 (N_3352,N_2596,N_2650);
and U3353 (N_3353,N_2708,N_2976);
and U3354 (N_3354,N_2699,N_2653);
and U3355 (N_3355,N_2658,N_2814);
and U3356 (N_3356,N_2646,N_2842);
or U3357 (N_3357,N_2635,N_2542);
nand U3358 (N_3358,N_2714,N_2802);
nand U3359 (N_3359,N_2798,N_2552);
or U3360 (N_3360,N_2852,N_2866);
or U3361 (N_3361,N_2967,N_2694);
or U3362 (N_3362,N_2896,N_2562);
nor U3363 (N_3363,N_2507,N_2805);
and U3364 (N_3364,N_2927,N_2985);
nor U3365 (N_3365,N_2552,N_2924);
xor U3366 (N_3366,N_2504,N_2545);
or U3367 (N_3367,N_2709,N_2809);
nand U3368 (N_3368,N_2705,N_2793);
nor U3369 (N_3369,N_2673,N_2875);
nand U3370 (N_3370,N_2598,N_2867);
nor U3371 (N_3371,N_2699,N_2986);
nor U3372 (N_3372,N_2675,N_2914);
or U3373 (N_3373,N_2911,N_2556);
and U3374 (N_3374,N_2594,N_2604);
nand U3375 (N_3375,N_2830,N_2604);
nand U3376 (N_3376,N_2968,N_2610);
nor U3377 (N_3377,N_2926,N_2579);
nand U3378 (N_3378,N_2787,N_2556);
xnor U3379 (N_3379,N_2860,N_2720);
and U3380 (N_3380,N_2972,N_2521);
and U3381 (N_3381,N_2692,N_2505);
nand U3382 (N_3382,N_2927,N_2561);
or U3383 (N_3383,N_2643,N_2704);
nand U3384 (N_3384,N_2969,N_2586);
nor U3385 (N_3385,N_2722,N_2746);
or U3386 (N_3386,N_2964,N_2855);
nand U3387 (N_3387,N_2563,N_2601);
nor U3388 (N_3388,N_2600,N_2810);
nand U3389 (N_3389,N_2851,N_2528);
nor U3390 (N_3390,N_2961,N_2916);
and U3391 (N_3391,N_2665,N_2680);
nand U3392 (N_3392,N_2562,N_2686);
nor U3393 (N_3393,N_2763,N_2616);
and U3394 (N_3394,N_2523,N_2892);
nand U3395 (N_3395,N_2641,N_2638);
or U3396 (N_3396,N_2946,N_2867);
and U3397 (N_3397,N_2937,N_2704);
or U3398 (N_3398,N_2814,N_2809);
or U3399 (N_3399,N_2671,N_2568);
xnor U3400 (N_3400,N_2679,N_2635);
or U3401 (N_3401,N_2641,N_2556);
xnor U3402 (N_3402,N_2865,N_2637);
nand U3403 (N_3403,N_2746,N_2796);
and U3404 (N_3404,N_2737,N_2988);
nor U3405 (N_3405,N_2575,N_2887);
and U3406 (N_3406,N_2883,N_2878);
nand U3407 (N_3407,N_2569,N_2918);
nor U3408 (N_3408,N_2639,N_2947);
and U3409 (N_3409,N_2575,N_2932);
nand U3410 (N_3410,N_2770,N_2781);
or U3411 (N_3411,N_2981,N_2934);
or U3412 (N_3412,N_2546,N_2680);
xor U3413 (N_3413,N_2670,N_2800);
xnor U3414 (N_3414,N_2773,N_2795);
xor U3415 (N_3415,N_2600,N_2860);
or U3416 (N_3416,N_2710,N_2878);
or U3417 (N_3417,N_2952,N_2700);
nor U3418 (N_3418,N_2683,N_2531);
and U3419 (N_3419,N_2673,N_2992);
or U3420 (N_3420,N_2503,N_2785);
nor U3421 (N_3421,N_2670,N_2762);
or U3422 (N_3422,N_2740,N_2571);
nand U3423 (N_3423,N_2704,N_2502);
nand U3424 (N_3424,N_2774,N_2688);
and U3425 (N_3425,N_2626,N_2928);
nor U3426 (N_3426,N_2953,N_2616);
or U3427 (N_3427,N_2588,N_2893);
nor U3428 (N_3428,N_2772,N_2897);
nor U3429 (N_3429,N_2899,N_2767);
and U3430 (N_3430,N_2758,N_2975);
nor U3431 (N_3431,N_2603,N_2965);
nor U3432 (N_3432,N_2715,N_2750);
and U3433 (N_3433,N_2930,N_2572);
nor U3434 (N_3434,N_2922,N_2562);
xor U3435 (N_3435,N_2993,N_2642);
nor U3436 (N_3436,N_2833,N_2963);
nand U3437 (N_3437,N_2899,N_2869);
or U3438 (N_3438,N_2821,N_2700);
or U3439 (N_3439,N_2867,N_2559);
and U3440 (N_3440,N_2850,N_2535);
nand U3441 (N_3441,N_2861,N_2694);
or U3442 (N_3442,N_2876,N_2833);
and U3443 (N_3443,N_2613,N_2652);
xor U3444 (N_3444,N_2893,N_2628);
or U3445 (N_3445,N_2832,N_2934);
nor U3446 (N_3446,N_2685,N_2735);
nor U3447 (N_3447,N_2650,N_2983);
or U3448 (N_3448,N_2561,N_2853);
and U3449 (N_3449,N_2951,N_2958);
or U3450 (N_3450,N_2983,N_2917);
and U3451 (N_3451,N_2694,N_2516);
nor U3452 (N_3452,N_2705,N_2807);
and U3453 (N_3453,N_2617,N_2672);
and U3454 (N_3454,N_2761,N_2600);
or U3455 (N_3455,N_2976,N_2845);
or U3456 (N_3456,N_2920,N_2902);
and U3457 (N_3457,N_2612,N_2771);
and U3458 (N_3458,N_2975,N_2668);
and U3459 (N_3459,N_2611,N_2975);
and U3460 (N_3460,N_2508,N_2642);
nand U3461 (N_3461,N_2787,N_2510);
nand U3462 (N_3462,N_2940,N_2882);
and U3463 (N_3463,N_2821,N_2751);
xor U3464 (N_3464,N_2898,N_2733);
nor U3465 (N_3465,N_2572,N_2609);
nor U3466 (N_3466,N_2762,N_2977);
nand U3467 (N_3467,N_2866,N_2976);
and U3468 (N_3468,N_2819,N_2930);
or U3469 (N_3469,N_2604,N_2762);
nor U3470 (N_3470,N_2857,N_2970);
nor U3471 (N_3471,N_2735,N_2741);
and U3472 (N_3472,N_2638,N_2659);
and U3473 (N_3473,N_2950,N_2564);
nor U3474 (N_3474,N_2744,N_2510);
nor U3475 (N_3475,N_2507,N_2727);
nand U3476 (N_3476,N_2807,N_2995);
nand U3477 (N_3477,N_2660,N_2902);
or U3478 (N_3478,N_2541,N_2824);
and U3479 (N_3479,N_2987,N_2724);
or U3480 (N_3480,N_2509,N_2671);
xor U3481 (N_3481,N_2732,N_2748);
or U3482 (N_3482,N_2697,N_2820);
and U3483 (N_3483,N_2787,N_2915);
or U3484 (N_3484,N_2638,N_2972);
or U3485 (N_3485,N_2684,N_2732);
nand U3486 (N_3486,N_2654,N_2793);
nor U3487 (N_3487,N_2753,N_2563);
nand U3488 (N_3488,N_2911,N_2843);
nor U3489 (N_3489,N_2619,N_2975);
and U3490 (N_3490,N_2968,N_2550);
nand U3491 (N_3491,N_2922,N_2823);
or U3492 (N_3492,N_2574,N_2624);
nor U3493 (N_3493,N_2500,N_2795);
nor U3494 (N_3494,N_2723,N_2912);
nand U3495 (N_3495,N_2874,N_2525);
or U3496 (N_3496,N_2690,N_2753);
and U3497 (N_3497,N_2646,N_2799);
or U3498 (N_3498,N_2891,N_2953);
nor U3499 (N_3499,N_2860,N_2853);
nand U3500 (N_3500,N_3387,N_3448);
and U3501 (N_3501,N_3488,N_3281);
nand U3502 (N_3502,N_3408,N_3370);
or U3503 (N_3503,N_3157,N_3143);
and U3504 (N_3504,N_3252,N_3349);
nor U3505 (N_3505,N_3374,N_3068);
or U3506 (N_3506,N_3376,N_3158);
or U3507 (N_3507,N_3210,N_3415);
nor U3508 (N_3508,N_3156,N_3194);
or U3509 (N_3509,N_3226,N_3219);
or U3510 (N_3510,N_3424,N_3207);
or U3511 (N_3511,N_3003,N_3411);
or U3512 (N_3512,N_3109,N_3309);
nor U3513 (N_3513,N_3327,N_3437);
nand U3514 (N_3514,N_3190,N_3315);
and U3515 (N_3515,N_3301,N_3269);
nand U3516 (N_3516,N_3254,N_3005);
nor U3517 (N_3517,N_3289,N_3319);
nand U3518 (N_3518,N_3340,N_3064);
and U3519 (N_3519,N_3114,N_3388);
and U3520 (N_3520,N_3482,N_3014);
xor U3521 (N_3521,N_3168,N_3443);
or U3522 (N_3522,N_3329,N_3086);
or U3523 (N_3523,N_3429,N_3077);
xor U3524 (N_3524,N_3067,N_3293);
nand U3525 (N_3525,N_3091,N_3242);
xnor U3526 (N_3526,N_3140,N_3222);
or U3527 (N_3527,N_3233,N_3307);
or U3528 (N_3528,N_3008,N_3166);
and U3529 (N_3529,N_3181,N_3031);
nor U3530 (N_3530,N_3476,N_3095);
nor U3531 (N_3531,N_3137,N_3006);
or U3532 (N_3532,N_3028,N_3154);
xor U3533 (N_3533,N_3467,N_3398);
or U3534 (N_3534,N_3416,N_3348);
or U3535 (N_3535,N_3170,N_3243);
or U3536 (N_3536,N_3292,N_3193);
nand U3537 (N_3537,N_3453,N_3481);
or U3538 (N_3538,N_3343,N_3283);
nand U3539 (N_3539,N_3299,N_3359);
nand U3540 (N_3540,N_3103,N_3162);
xnor U3541 (N_3541,N_3291,N_3149);
and U3542 (N_3542,N_3044,N_3232);
or U3543 (N_3543,N_3320,N_3350);
nand U3544 (N_3544,N_3393,N_3366);
xor U3545 (N_3545,N_3490,N_3208);
nor U3546 (N_3546,N_3225,N_3088);
nand U3547 (N_3547,N_3294,N_3395);
xnor U3548 (N_3548,N_3120,N_3155);
and U3549 (N_3549,N_3465,N_3177);
nor U3550 (N_3550,N_3023,N_3065);
nand U3551 (N_3551,N_3211,N_3438);
nand U3552 (N_3552,N_3262,N_3128);
or U3553 (N_3553,N_3385,N_3256);
or U3554 (N_3554,N_3336,N_3427);
and U3555 (N_3555,N_3297,N_3331);
nor U3556 (N_3556,N_3464,N_3425);
nand U3557 (N_3557,N_3392,N_3375);
nand U3558 (N_3558,N_3039,N_3097);
xnor U3559 (N_3559,N_3380,N_3072);
and U3560 (N_3560,N_3037,N_3337);
nand U3561 (N_3561,N_3275,N_3197);
and U3562 (N_3562,N_3125,N_3246);
nor U3563 (N_3563,N_3217,N_3280);
and U3564 (N_3564,N_3442,N_3368);
xnor U3565 (N_3565,N_3163,N_3200);
or U3566 (N_3566,N_3123,N_3248);
nor U3567 (N_3567,N_3347,N_3494);
nor U3568 (N_3568,N_3061,N_3078);
or U3569 (N_3569,N_3394,N_3019);
nand U3570 (N_3570,N_3363,N_3334);
and U3571 (N_3571,N_3002,N_3377);
nand U3572 (N_3572,N_3477,N_3321);
or U3573 (N_3573,N_3027,N_3201);
nor U3574 (N_3574,N_3209,N_3391);
or U3575 (N_3575,N_3169,N_3053);
and U3576 (N_3576,N_3130,N_3179);
or U3577 (N_3577,N_3167,N_3263);
nor U3578 (N_3578,N_3051,N_3129);
and U3579 (N_3579,N_3213,N_3253);
nor U3580 (N_3580,N_3025,N_3258);
nand U3581 (N_3581,N_3076,N_3290);
nand U3582 (N_3582,N_3412,N_3303);
nand U3583 (N_3583,N_3241,N_3127);
and U3584 (N_3584,N_3326,N_3100);
or U3585 (N_3585,N_3378,N_3332);
nand U3586 (N_3586,N_3029,N_3308);
nor U3587 (N_3587,N_3196,N_3265);
nand U3588 (N_3588,N_3409,N_3428);
and U3589 (N_3589,N_3202,N_3038);
and U3590 (N_3590,N_3312,N_3117);
nand U3591 (N_3591,N_3447,N_3055);
nand U3592 (N_3592,N_3112,N_3236);
and U3593 (N_3593,N_3013,N_3228);
nand U3594 (N_3594,N_3151,N_3054);
nor U3595 (N_3595,N_3043,N_3485);
xnor U3596 (N_3596,N_3282,N_3144);
nand U3597 (N_3597,N_3383,N_3105);
nand U3598 (N_3598,N_3180,N_3462);
and U3599 (N_3599,N_3188,N_3354);
and U3600 (N_3600,N_3135,N_3066);
and U3601 (N_3601,N_3238,N_3115);
or U3602 (N_3602,N_3082,N_3139);
nor U3603 (N_3603,N_3259,N_3199);
and U3604 (N_3604,N_3034,N_3497);
or U3605 (N_3605,N_3257,N_3325);
or U3606 (N_3606,N_3161,N_3471);
nand U3607 (N_3607,N_3063,N_3274);
nor U3608 (N_3608,N_3345,N_3410);
or U3609 (N_3609,N_3119,N_3470);
nand U3610 (N_3610,N_3272,N_3205);
and U3611 (N_3611,N_3267,N_3404);
nand U3612 (N_3612,N_3369,N_3405);
nor U3613 (N_3613,N_3356,N_3328);
nor U3614 (N_3614,N_3324,N_3413);
nor U3615 (N_3615,N_3224,N_3052);
and U3616 (N_3616,N_3148,N_3486);
nand U3617 (N_3617,N_3367,N_3449);
xor U3618 (N_3618,N_3342,N_3472);
nand U3619 (N_3619,N_3284,N_3096);
or U3620 (N_3620,N_3033,N_3358);
and U3621 (N_3621,N_3142,N_3365);
or U3622 (N_3622,N_3473,N_3421);
and U3623 (N_3623,N_3397,N_3386);
and U3624 (N_3624,N_3191,N_3346);
xor U3625 (N_3625,N_3314,N_3451);
and U3626 (N_3626,N_3070,N_3244);
nand U3627 (N_3627,N_3396,N_3040);
xnor U3628 (N_3628,N_3004,N_3174);
or U3629 (N_3629,N_3175,N_3011);
and U3630 (N_3630,N_3302,N_3110);
and U3631 (N_3631,N_3480,N_3098);
or U3632 (N_3632,N_3474,N_3015);
or U3633 (N_3633,N_3300,N_3460);
and U3634 (N_3634,N_3104,N_3007);
or U3635 (N_3635,N_3059,N_3164);
nor U3636 (N_3636,N_3439,N_3152);
or U3637 (N_3637,N_3344,N_3434);
or U3638 (N_3638,N_3456,N_3311);
and U3639 (N_3639,N_3400,N_3231);
nor U3640 (N_3640,N_3261,N_3230);
xnor U3641 (N_3641,N_3371,N_3126);
xor U3642 (N_3642,N_3009,N_3381);
xor U3643 (N_3643,N_3138,N_3172);
nor U3644 (N_3644,N_3183,N_3499);
nor U3645 (N_3645,N_3189,N_3288);
nor U3646 (N_3646,N_3136,N_3455);
nor U3647 (N_3647,N_3215,N_3074);
nand U3648 (N_3648,N_3178,N_3237);
or U3649 (N_3649,N_3333,N_3229);
nor U3650 (N_3650,N_3479,N_3160);
nand U3651 (N_3651,N_3466,N_3195);
or U3652 (N_3652,N_3277,N_3216);
or U3653 (N_3653,N_3498,N_3446);
xor U3654 (N_3654,N_3106,N_3270);
or U3655 (N_3655,N_3220,N_3094);
nand U3656 (N_3656,N_3018,N_3032);
or U3657 (N_3657,N_3218,N_3185);
nor U3658 (N_3658,N_3056,N_3322);
nor U3659 (N_3659,N_3026,N_3173);
nor U3660 (N_3660,N_3171,N_3122);
nor U3661 (N_3661,N_3108,N_3399);
or U3662 (N_3662,N_3085,N_3390);
or U3663 (N_3663,N_3468,N_3022);
and U3664 (N_3664,N_3030,N_3251);
nand U3665 (N_3665,N_3012,N_3245);
xnor U3666 (N_3666,N_3050,N_3478);
or U3667 (N_3667,N_3436,N_3124);
nand U3668 (N_3668,N_3083,N_3084);
nand U3669 (N_3669,N_3045,N_3389);
or U3670 (N_3670,N_3121,N_3310);
and U3671 (N_3671,N_3240,N_3483);
and U3672 (N_3672,N_3454,N_3420);
nand U3673 (N_3673,N_3418,N_3227);
or U3674 (N_3674,N_3384,N_3223);
nor U3675 (N_3675,N_3047,N_3147);
nand U3676 (N_3676,N_3278,N_3081);
nand U3677 (N_3677,N_3010,N_3042);
or U3678 (N_3678,N_3339,N_3020);
or U3679 (N_3679,N_3492,N_3071);
and U3680 (N_3680,N_3234,N_3295);
or U3681 (N_3681,N_3276,N_3035);
nand U3682 (N_3682,N_3133,N_3250);
or U3683 (N_3683,N_3484,N_3024);
and U3684 (N_3684,N_3461,N_3419);
nand U3685 (N_3685,N_3036,N_3092);
xor U3686 (N_3686,N_3255,N_3260);
or U3687 (N_3687,N_3355,N_3192);
and U3688 (N_3688,N_3159,N_3401);
nand U3689 (N_3689,N_3316,N_3184);
nor U3690 (N_3690,N_3134,N_3041);
and U3691 (N_3691,N_3382,N_3430);
or U3692 (N_3692,N_3351,N_3417);
nand U3693 (N_3693,N_3432,N_3279);
and U3694 (N_3694,N_3318,N_3221);
nor U3695 (N_3695,N_3239,N_3206);
nor U3696 (N_3696,N_3450,N_3493);
and U3697 (N_3697,N_3285,N_3017);
and U3698 (N_3698,N_3264,N_3075);
nand U3699 (N_3699,N_3452,N_3153);
or U3700 (N_3700,N_3132,N_3330);
or U3701 (N_3701,N_3102,N_3145);
nor U3702 (N_3702,N_3048,N_3150);
nand U3703 (N_3703,N_3489,N_3203);
xnor U3704 (N_3704,N_3089,N_3093);
and U3705 (N_3705,N_3165,N_3214);
nand U3706 (N_3706,N_3204,N_3440);
or U3707 (N_3707,N_3235,N_3414);
nand U3708 (N_3708,N_3458,N_3445);
or U3709 (N_3709,N_3286,N_3423);
and U3710 (N_3710,N_3090,N_3113);
nor U3711 (N_3711,N_3116,N_3335);
or U3712 (N_3712,N_3062,N_3058);
or U3713 (N_3713,N_3463,N_3305);
or U3714 (N_3714,N_3357,N_3457);
xor U3715 (N_3715,N_3426,N_3372);
xor U3716 (N_3716,N_3362,N_3176);
nor U3717 (N_3717,N_3057,N_3273);
xnor U3718 (N_3718,N_3271,N_3001);
nor U3719 (N_3719,N_3249,N_3079);
nor U3720 (N_3720,N_3373,N_3435);
nor U3721 (N_3721,N_3495,N_3268);
nor U3722 (N_3722,N_3198,N_3403);
nor U3723 (N_3723,N_3496,N_3016);
xnor U3724 (N_3724,N_3101,N_3073);
and U3725 (N_3725,N_3379,N_3049);
nor U3726 (N_3726,N_3422,N_3131);
or U3727 (N_3727,N_3187,N_3266);
or U3728 (N_3728,N_3360,N_3469);
nand U3729 (N_3729,N_3361,N_3287);
xnor U3730 (N_3730,N_3021,N_3146);
and U3731 (N_3731,N_3406,N_3364);
nand U3732 (N_3732,N_3099,N_3298);
and U3733 (N_3733,N_3402,N_3069);
or U3734 (N_3734,N_3087,N_3182);
and U3735 (N_3735,N_3296,N_3000);
and U3736 (N_3736,N_3475,N_3459);
and U3737 (N_3737,N_3352,N_3111);
nor U3738 (N_3738,N_3431,N_3487);
xnor U3739 (N_3739,N_3212,N_3313);
xor U3740 (N_3740,N_3304,N_3433);
and U3741 (N_3741,N_3141,N_3338);
or U3742 (N_3742,N_3317,N_3341);
nor U3743 (N_3743,N_3444,N_3323);
nand U3744 (N_3744,N_3046,N_3491);
and U3745 (N_3745,N_3353,N_3247);
and U3746 (N_3746,N_3060,N_3306);
and U3747 (N_3747,N_3080,N_3107);
and U3748 (N_3748,N_3441,N_3186);
or U3749 (N_3749,N_3118,N_3407);
or U3750 (N_3750,N_3394,N_3436);
or U3751 (N_3751,N_3282,N_3329);
and U3752 (N_3752,N_3065,N_3405);
nand U3753 (N_3753,N_3221,N_3084);
nand U3754 (N_3754,N_3351,N_3060);
nand U3755 (N_3755,N_3122,N_3128);
and U3756 (N_3756,N_3101,N_3297);
nor U3757 (N_3757,N_3380,N_3253);
or U3758 (N_3758,N_3218,N_3365);
xnor U3759 (N_3759,N_3343,N_3485);
and U3760 (N_3760,N_3285,N_3398);
and U3761 (N_3761,N_3105,N_3397);
nor U3762 (N_3762,N_3482,N_3228);
and U3763 (N_3763,N_3290,N_3135);
nor U3764 (N_3764,N_3487,N_3490);
nor U3765 (N_3765,N_3479,N_3376);
nor U3766 (N_3766,N_3091,N_3477);
nor U3767 (N_3767,N_3331,N_3084);
and U3768 (N_3768,N_3285,N_3433);
or U3769 (N_3769,N_3253,N_3196);
nand U3770 (N_3770,N_3467,N_3144);
or U3771 (N_3771,N_3449,N_3123);
nand U3772 (N_3772,N_3324,N_3355);
nor U3773 (N_3773,N_3058,N_3076);
or U3774 (N_3774,N_3453,N_3141);
or U3775 (N_3775,N_3488,N_3106);
nor U3776 (N_3776,N_3033,N_3163);
nand U3777 (N_3777,N_3111,N_3222);
xnor U3778 (N_3778,N_3496,N_3467);
and U3779 (N_3779,N_3449,N_3296);
and U3780 (N_3780,N_3298,N_3482);
or U3781 (N_3781,N_3425,N_3432);
nand U3782 (N_3782,N_3303,N_3268);
or U3783 (N_3783,N_3106,N_3443);
or U3784 (N_3784,N_3440,N_3257);
or U3785 (N_3785,N_3490,N_3067);
and U3786 (N_3786,N_3398,N_3244);
and U3787 (N_3787,N_3177,N_3188);
or U3788 (N_3788,N_3079,N_3179);
and U3789 (N_3789,N_3458,N_3495);
and U3790 (N_3790,N_3252,N_3061);
or U3791 (N_3791,N_3076,N_3185);
or U3792 (N_3792,N_3040,N_3345);
and U3793 (N_3793,N_3444,N_3326);
or U3794 (N_3794,N_3387,N_3165);
or U3795 (N_3795,N_3150,N_3217);
and U3796 (N_3796,N_3448,N_3319);
xor U3797 (N_3797,N_3446,N_3499);
nand U3798 (N_3798,N_3298,N_3376);
or U3799 (N_3799,N_3196,N_3151);
and U3800 (N_3800,N_3351,N_3183);
nor U3801 (N_3801,N_3459,N_3186);
xnor U3802 (N_3802,N_3268,N_3025);
and U3803 (N_3803,N_3278,N_3005);
and U3804 (N_3804,N_3328,N_3320);
or U3805 (N_3805,N_3488,N_3450);
nand U3806 (N_3806,N_3216,N_3212);
nor U3807 (N_3807,N_3471,N_3304);
nand U3808 (N_3808,N_3046,N_3186);
or U3809 (N_3809,N_3034,N_3381);
nand U3810 (N_3810,N_3027,N_3380);
nor U3811 (N_3811,N_3004,N_3309);
or U3812 (N_3812,N_3339,N_3171);
and U3813 (N_3813,N_3026,N_3267);
nor U3814 (N_3814,N_3029,N_3403);
and U3815 (N_3815,N_3337,N_3057);
xnor U3816 (N_3816,N_3204,N_3493);
or U3817 (N_3817,N_3420,N_3252);
and U3818 (N_3818,N_3333,N_3245);
xnor U3819 (N_3819,N_3141,N_3494);
nor U3820 (N_3820,N_3186,N_3409);
and U3821 (N_3821,N_3296,N_3148);
or U3822 (N_3822,N_3005,N_3262);
nand U3823 (N_3823,N_3186,N_3114);
nor U3824 (N_3824,N_3067,N_3190);
nand U3825 (N_3825,N_3176,N_3300);
nor U3826 (N_3826,N_3079,N_3034);
and U3827 (N_3827,N_3403,N_3425);
nor U3828 (N_3828,N_3365,N_3292);
and U3829 (N_3829,N_3350,N_3042);
or U3830 (N_3830,N_3166,N_3139);
and U3831 (N_3831,N_3026,N_3076);
and U3832 (N_3832,N_3358,N_3143);
nand U3833 (N_3833,N_3151,N_3195);
nor U3834 (N_3834,N_3085,N_3018);
or U3835 (N_3835,N_3397,N_3216);
nand U3836 (N_3836,N_3394,N_3367);
or U3837 (N_3837,N_3084,N_3482);
or U3838 (N_3838,N_3060,N_3323);
or U3839 (N_3839,N_3455,N_3246);
nor U3840 (N_3840,N_3484,N_3079);
nor U3841 (N_3841,N_3012,N_3193);
or U3842 (N_3842,N_3347,N_3310);
or U3843 (N_3843,N_3232,N_3296);
or U3844 (N_3844,N_3074,N_3493);
xnor U3845 (N_3845,N_3018,N_3102);
xor U3846 (N_3846,N_3062,N_3260);
and U3847 (N_3847,N_3018,N_3461);
nand U3848 (N_3848,N_3255,N_3437);
nand U3849 (N_3849,N_3453,N_3386);
or U3850 (N_3850,N_3408,N_3280);
or U3851 (N_3851,N_3108,N_3401);
nor U3852 (N_3852,N_3235,N_3055);
and U3853 (N_3853,N_3223,N_3013);
nor U3854 (N_3854,N_3410,N_3006);
and U3855 (N_3855,N_3356,N_3185);
or U3856 (N_3856,N_3374,N_3437);
and U3857 (N_3857,N_3131,N_3148);
xor U3858 (N_3858,N_3458,N_3220);
nor U3859 (N_3859,N_3161,N_3364);
nor U3860 (N_3860,N_3435,N_3404);
or U3861 (N_3861,N_3351,N_3109);
or U3862 (N_3862,N_3149,N_3418);
nor U3863 (N_3863,N_3323,N_3278);
or U3864 (N_3864,N_3438,N_3012);
nand U3865 (N_3865,N_3148,N_3491);
nor U3866 (N_3866,N_3273,N_3211);
nor U3867 (N_3867,N_3467,N_3393);
nor U3868 (N_3868,N_3060,N_3097);
and U3869 (N_3869,N_3282,N_3302);
nand U3870 (N_3870,N_3387,N_3096);
nor U3871 (N_3871,N_3000,N_3399);
or U3872 (N_3872,N_3496,N_3478);
and U3873 (N_3873,N_3199,N_3347);
xnor U3874 (N_3874,N_3116,N_3454);
and U3875 (N_3875,N_3138,N_3490);
xor U3876 (N_3876,N_3139,N_3228);
or U3877 (N_3877,N_3363,N_3003);
xnor U3878 (N_3878,N_3398,N_3135);
xor U3879 (N_3879,N_3217,N_3368);
nand U3880 (N_3880,N_3468,N_3140);
nand U3881 (N_3881,N_3266,N_3131);
xor U3882 (N_3882,N_3293,N_3137);
or U3883 (N_3883,N_3041,N_3393);
nand U3884 (N_3884,N_3449,N_3117);
and U3885 (N_3885,N_3210,N_3499);
and U3886 (N_3886,N_3219,N_3437);
nand U3887 (N_3887,N_3022,N_3443);
nor U3888 (N_3888,N_3497,N_3174);
nand U3889 (N_3889,N_3487,N_3219);
nand U3890 (N_3890,N_3221,N_3472);
nand U3891 (N_3891,N_3136,N_3225);
xor U3892 (N_3892,N_3044,N_3159);
nor U3893 (N_3893,N_3419,N_3170);
or U3894 (N_3894,N_3171,N_3389);
or U3895 (N_3895,N_3318,N_3470);
or U3896 (N_3896,N_3300,N_3114);
nor U3897 (N_3897,N_3194,N_3056);
nor U3898 (N_3898,N_3179,N_3013);
and U3899 (N_3899,N_3001,N_3026);
nor U3900 (N_3900,N_3421,N_3007);
nand U3901 (N_3901,N_3112,N_3329);
or U3902 (N_3902,N_3063,N_3064);
xor U3903 (N_3903,N_3078,N_3433);
nor U3904 (N_3904,N_3456,N_3420);
nor U3905 (N_3905,N_3239,N_3238);
and U3906 (N_3906,N_3125,N_3027);
xor U3907 (N_3907,N_3192,N_3188);
and U3908 (N_3908,N_3065,N_3283);
nand U3909 (N_3909,N_3324,N_3165);
xor U3910 (N_3910,N_3015,N_3350);
and U3911 (N_3911,N_3212,N_3310);
and U3912 (N_3912,N_3104,N_3166);
or U3913 (N_3913,N_3308,N_3497);
nor U3914 (N_3914,N_3494,N_3435);
or U3915 (N_3915,N_3203,N_3191);
nand U3916 (N_3916,N_3361,N_3118);
nor U3917 (N_3917,N_3185,N_3328);
nor U3918 (N_3918,N_3394,N_3067);
or U3919 (N_3919,N_3128,N_3115);
nor U3920 (N_3920,N_3097,N_3130);
nor U3921 (N_3921,N_3339,N_3025);
nand U3922 (N_3922,N_3067,N_3135);
nand U3923 (N_3923,N_3472,N_3353);
and U3924 (N_3924,N_3393,N_3485);
xnor U3925 (N_3925,N_3351,N_3345);
or U3926 (N_3926,N_3488,N_3100);
and U3927 (N_3927,N_3259,N_3072);
nor U3928 (N_3928,N_3180,N_3465);
and U3929 (N_3929,N_3347,N_3200);
and U3930 (N_3930,N_3045,N_3242);
or U3931 (N_3931,N_3308,N_3368);
nand U3932 (N_3932,N_3314,N_3297);
nor U3933 (N_3933,N_3088,N_3074);
nand U3934 (N_3934,N_3240,N_3276);
or U3935 (N_3935,N_3068,N_3007);
xnor U3936 (N_3936,N_3233,N_3212);
nor U3937 (N_3937,N_3057,N_3139);
xnor U3938 (N_3938,N_3041,N_3204);
nor U3939 (N_3939,N_3350,N_3329);
or U3940 (N_3940,N_3045,N_3008);
and U3941 (N_3941,N_3062,N_3348);
and U3942 (N_3942,N_3173,N_3035);
or U3943 (N_3943,N_3082,N_3486);
or U3944 (N_3944,N_3387,N_3223);
or U3945 (N_3945,N_3249,N_3040);
nor U3946 (N_3946,N_3291,N_3267);
nand U3947 (N_3947,N_3271,N_3268);
or U3948 (N_3948,N_3087,N_3481);
nand U3949 (N_3949,N_3481,N_3050);
xnor U3950 (N_3950,N_3196,N_3254);
or U3951 (N_3951,N_3070,N_3077);
nand U3952 (N_3952,N_3032,N_3083);
or U3953 (N_3953,N_3114,N_3269);
nand U3954 (N_3954,N_3044,N_3091);
or U3955 (N_3955,N_3422,N_3216);
or U3956 (N_3956,N_3271,N_3090);
xnor U3957 (N_3957,N_3486,N_3015);
nor U3958 (N_3958,N_3315,N_3276);
xor U3959 (N_3959,N_3198,N_3279);
xor U3960 (N_3960,N_3136,N_3325);
nand U3961 (N_3961,N_3404,N_3161);
nand U3962 (N_3962,N_3463,N_3116);
and U3963 (N_3963,N_3375,N_3057);
nand U3964 (N_3964,N_3396,N_3086);
xor U3965 (N_3965,N_3324,N_3054);
nor U3966 (N_3966,N_3252,N_3309);
or U3967 (N_3967,N_3001,N_3012);
nand U3968 (N_3968,N_3270,N_3180);
nand U3969 (N_3969,N_3143,N_3353);
xor U3970 (N_3970,N_3163,N_3468);
nor U3971 (N_3971,N_3139,N_3397);
nand U3972 (N_3972,N_3154,N_3066);
and U3973 (N_3973,N_3192,N_3420);
and U3974 (N_3974,N_3299,N_3065);
and U3975 (N_3975,N_3265,N_3317);
xnor U3976 (N_3976,N_3203,N_3014);
xor U3977 (N_3977,N_3240,N_3031);
nand U3978 (N_3978,N_3460,N_3411);
nand U3979 (N_3979,N_3471,N_3148);
nor U3980 (N_3980,N_3406,N_3132);
nand U3981 (N_3981,N_3340,N_3084);
and U3982 (N_3982,N_3444,N_3165);
and U3983 (N_3983,N_3230,N_3140);
nor U3984 (N_3984,N_3180,N_3182);
or U3985 (N_3985,N_3123,N_3028);
or U3986 (N_3986,N_3011,N_3350);
nand U3987 (N_3987,N_3295,N_3206);
xnor U3988 (N_3988,N_3174,N_3295);
xnor U3989 (N_3989,N_3148,N_3285);
and U3990 (N_3990,N_3460,N_3359);
nor U3991 (N_3991,N_3494,N_3073);
and U3992 (N_3992,N_3461,N_3350);
nor U3993 (N_3993,N_3202,N_3237);
and U3994 (N_3994,N_3103,N_3109);
nor U3995 (N_3995,N_3149,N_3355);
or U3996 (N_3996,N_3223,N_3378);
nor U3997 (N_3997,N_3425,N_3244);
nor U3998 (N_3998,N_3364,N_3240);
or U3999 (N_3999,N_3035,N_3107);
or U4000 (N_4000,N_3978,N_3522);
nand U4001 (N_4001,N_3715,N_3951);
nand U4002 (N_4002,N_3628,N_3799);
or U4003 (N_4003,N_3863,N_3829);
and U4004 (N_4004,N_3935,N_3776);
nor U4005 (N_4005,N_3549,N_3985);
or U4006 (N_4006,N_3762,N_3945);
and U4007 (N_4007,N_3584,N_3828);
nor U4008 (N_4008,N_3564,N_3916);
or U4009 (N_4009,N_3646,N_3929);
or U4010 (N_4010,N_3906,N_3663);
or U4011 (N_4011,N_3565,N_3666);
nor U4012 (N_4012,N_3813,N_3831);
xnor U4013 (N_4013,N_3835,N_3639);
or U4014 (N_4014,N_3939,N_3669);
nand U4015 (N_4015,N_3533,N_3980);
or U4016 (N_4016,N_3636,N_3735);
and U4017 (N_4017,N_3538,N_3970);
and U4018 (N_4018,N_3789,N_3977);
xor U4019 (N_4019,N_3548,N_3782);
or U4020 (N_4020,N_3972,N_3708);
and U4021 (N_4021,N_3519,N_3790);
and U4022 (N_4022,N_3902,N_3784);
nor U4023 (N_4023,N_3817,N_3756);
xor U4024 (N_4024,N_3734,N_3897);
and U4025 (N_4025,N_3974,N_3919);
nor U4026 (N_4026,N_3687,N_3883);
nand U4027 (N_4027,N_3909,N_3960);
nand U4028 (N_4028,N_3913,N_3516);
or U4029 (N_4029,N_3573,N_3948);
or U4030 (N_4030,N_3562,N_3764);
and U4031 (N_4031,N_3637,N_3848);
nor U4032 (N_4032,N_3768,N_3606);
or U4033 (N_4033,N_3921,N_3791);
and U4034 (N_4034,N_3924,N_3745);
or U4035 (N_4035,N_3633,N_3733);
nand U4036 (N_4036,N_3988,N_3650);
nand U4037 (N_4037,N_3803,N_3661);
or U4038 (N_4038,N_3975,N_3622);
and U4039 (N_4039,N_3686,N_3870);
or U4040 (N_4040,N_3868,N_3800);
nor U4041 (N_4041,N_3504,N_3994);
or U4042 (N_4042,N_3627,N_3895);
nor U4043 (N_4043,N_3918,N_3904);
nor U4044 (N_4044,N_3809,N_3967);
and U4045 (N_4045,N_3954,N_3613);
nand U4046 (N_4046,N_3859,N_3728);
and U4047 (N_4047,N_3957,N_3552);
nor U4048 (N_4048,N_3551,N_3662);
or U4049 (N_4049,N_3585,N_3737);
xnor U4050 (N_4050,N_3648,N_3617);
and U4051 (N_4051,N_3757,N_3944);
nor U4052 (N_4052,N_3556,N_3647);
nor U4053 (N_4053,N_3840,N_3629);
nor U4054 (N_4054,N_3683,N_3788);
or U4055 (N_4055,N_3827,N_3881);
nor U4056 (N_4056,N_3591,N_3610);
nor U4057 (N_4057,N_3999,N_3910);
nor U4058 (N_4058,N_3882,N_3580);
and U4059 (N_4059,N_3676,N_3819);
nand U4060 (N_4060,N_3814,N_3792);
xnor U4061 (N_4061,N_3727,N_3947);
nand U4062 (N_4062,N_3583,N_3760);
nor U4063 (N_4063,N_3587,N_3596);
or U4064 (N_4064,N_3574,N_3664);
nor U4065 (N_4065,N_3680,N_3582);
or U4066 (N_4066,N_3971,N_3701);
or U4067 (N_4067,N_3810,N_3915);
xor U4068 (N_4068,N_3566,N_3763);
nand U4069 (N_4069,N_3656,N_3511);
nor U4070 (N_4070,N_3842,N_3779);
nor U4071 (N_4071,N_3898,N_3815);
nor U4072 (N_4072,N_3801,N_3794);
nand U4073 (N_4073,N_3624,N_3884);
or U4074 (N_4074,N_3570,N_3940);
or U4075 (N_4075,N_3642,N_3861);
or U4076 (N_4076,N_3612,N_3682);
and U4077 (N_4077,N_3597,N_3665);
and U4078 (N_4078,N_3890,N_3532);
xor U4079 (N_4079,N_3787,N_3524);
nor U4080 (N_4080,N_3502,N_3774);
or U4081 (N_4081,N_3990,N_3846);
or U4082 (N_4082,N_3654,N_3812);
or U4083 (N_4083,N_3555,N_3705);
or U4084 (N_4084,N_3693,N_3702);
nand U4085 (N_4085,N_3604,N_3885);
or U4086 (N_4086,N_3722,N_3630);
nor U4087 (N_4087,N_3738,N_3933);
nor U4088 (N_4088,N_3865,N_3816);
nand U4089 (N_4089,N_3507,N_3963);
nand U4090 (N_4090,N_3931,N_3891);
nor U4091 (N_4091,N_3755,N_3928);
nand U4092 (N_4092,N_3917,N_3547);
nor U4093 (N_4093,N_3867,N_3672);
nor U4094 (N_4094,N_3786,N_3880);
and U4095 (N_4095,N_3725,N_3806);
and U4096 (N_4096,N_3690,N_3601);
and U4097 (N_4097,N_3771,N_3905);
nor U4098 (N_4098,N_3938,N_3927);
or U4099 (N_4099,N_3560,N_3930);
or U4100 (N_4100,N_3608,N_3506);
or U4101 (N_4101,N_3925,N_3856);
nand U4102 (N_4102,N_3703,N_3991);
nand U4103 (N_4103,N_3589,N_3546);
and U4104 (N_4104,N_3864,N_3710);
nand U4105 (N_4105,N_3989,N_3839);
or U4106 (N_4106,N_3862,N_3694);
nor U4107 (N_4107,N_3770,N_3577);
nand U4108 (N_4108,N_3785,N_3855);
nor U4109 (N_4109,N_3979,N_3652);
and U4110 (N_4110,N_3553,N_3833);
or U4111 (N_4111,N_3718,N_3926);
and U4112 (N_4112,N_3568,N_3778);
or U4113 (N_4113,N_3563,N_3805);
nor U4114 (N_4114,N_3509,N_3998);
nand U4115 (N_4115,N_3501,N_3525);
nor U4116 (N_4116,N_3670,N_3607);
xnor U4117 (N_4117,N_3623,N_3539);
nor U4118 (N_4118,N_3808,N_3667);
nor U4119 (N_4119,N_3802,N_3640);
and U4120 (N_4120,N_3559,N_3598);
or U4121 (N_4121,N_3530,N_3550);
nand U4122 (N_4122,N_3730,N_3781);
nand U4123 (N_4123,N_3542,N_3679);
nand U4124 (N_4124,N_3558,N_3973);
nand U4125 (N_4125,N_3886,N_3888);
and U4126 (N_4126,N_3632,N_3937);
nand U4127 (N_4127,N_3594,N_3941);
and U4128 (N_4128,N_3586,N_3903);
nand U4129 (N_4129,N_3922,N_3520);
and U4130 (N_4130,N_3887,N_3993);
and U4131 (N_4131,N_3876,N_3961);
nor U4132 (N_4132,N_3657,N_3969);
or U4133 (N_4133,N_3739,N_3866);
and U4134 (N_4134,N_3626,N_3521);
or U4135 (N_4135,N_3712,N_3692);
nand U4136 (N_4136,N_3619,N_3673);
nand U4137 (N_4137,N_3943,N_3982);
and U4138 (N_4138,N_3995,N_3912);
nand U4139 (N_4139,N_3615,N_3820);
and U4140 (N_4140,N_3668,N_3860);
or U4141 (N_4141,N_3536,N_3753);
and U4142 (N_4142,N_3696,N_3685);
xor U4143 (N_4143,N_3523,N_3513);
and U4144 (N_4144,N_3602,N_3614);
xnor U4145 (N_4145,N_3968,N_3750);
nor U4146 (N_4146,N_3849,N_3505);
nand U4147 (N_4147,N_3625,N_3748);
nor U4148 (N_4148,N_3798,N_3581);
nor U4149 (N_4149,N_3503,N_3716);
nor U4150 (N_4150,N_3878,N_3908);
or U4151 (N_4151,N_3643,N_3605);
xnor U4152 (N_4152,N_3644,N_3832);
or U4153 (N_4153,N_3987,N_3877);
nor U4154 (N_4154,N_3854,N_3953);
nand U4155 (N_4155,N_3588,N_3823);
and U4156 (N_4156,N_3783,N_3869);
xnor U4157 (N_4157,N_3958,N_3746);
nand U4158 (N_4158,N_3804,N_3510);
nand U4159 (N_4159,N_3658,N_3966);
nand U4160 (N_4160,N_3620,N_3599);
nand U4161 (N_4161,N_3649,N_3894);
and U4162 (N_4162,N_3952,N_3834);
nor U4163 (N_4163,N_3811,N_3700);
xor U4164 (N_4164,N_3731,N_3675);
nand U4165 (N_4165,N_3659,N_3514);
nand U4166 (N_4166,N_3660,N_3777);
xor U4167 (N_4167,N_3871,N_3752);
xor U4168 (N_4168,N_3914,N_3576);
or U4169 (N_4169,N_3653,N_3706);
and U4170 (N_4170,N_3618,N_3853);
nor U4171 (N_4171,N_3508,N_3932);
and U4172 (N_4172,N_3709,N_3765);
or U4173 (N_4173,N_3751,N_3537);
nor U4174 (N_4174,N_3590,N_3651);
nor U4175 (N_4175,N_3850,N_3535);
xor U4176 (N_4176,N_3826,N_3681);
nand U4177 (N_4177,N_3892,N_3603);
nand U4178 (N_4178,N_3796,N_3841);
or U4179 (N_4179,N_3851,N_3795);
and U4180 (N_4180,N_3571,N_3529);
nand U4181 (N_4181,N_3674,N_3852);
or U4182 (N_4182,N_3836,N_3689);
or U4183 (N_4183,N_3911,N_3517);
and U4184 (N_4184,N_3699,N_3554);
and U4185 (N_4185,N_3698,N_3754);
nand U4186 (N_4186,N_3996,N_3950);
nand U4187 (N_4187,N_3893,N_3749);
or U4188 (N_4188,N_3825,N_3830);
and U4189 (N_4189,N_3515,N_3879);
and U4190 (N_4190,N_3724,N_3512);
or U4191 (N_4191,N_3736,N_3743);
or U4192 (N_4192,N_3534,N_3645);
nor U4193 (N_4193,N_3714,N_3688);
nand U4194 (N_4194,N_3723,N_3824);
or U4195 (N_4195,N_3616,N_3976);
xor U4196 (N_4196,N_3634,N_3992);
or U4197 (N_4197,N_3780,N_3747);
xor U4198 (N_4198,N_3697,N_3874);
or U4199 (N_4199,N_3997,N_3964);
nor U4200 (N_4200,N_3729,N_3838);
or U4201 (N_4201,N_3631,N_3741);
nor U4202 (N_4202,N_3569,N_3845);
or U4203 (N_4203,N_3773,N_3704);
nor U4204 (N_4204,N_3593,N_3769);
or U4205 (N_4205,N_3531,N_3678);
xnor U4206 (N_4206,N_3557,N_3942);
or U4207 (N_4207,N_3844,N_3872);
or U4208 (N_4208,N_3843,N_3740);
and U4209 (N_4209,N_3920,N_3684);
xor U4210 (N_4210,N_3873,N_3986);
nand U4211 (N_4211,N_3720,N_3578);
nor U4212 (N_4212,N_3595,N_3600);
xor U4213 (N_4213,N_3821,N_3767);
nand U4214 (N_4214,N_3719,N_3732);
and U4215 (N_4215,N_3934,N_3857);
nand U4216 (N_4216,N_3543,N_3711);
or U4217 (N_4217,N_3956,N_3959);
and U4218 (N_4218,N_3858,N_3772);
or U4219 (N_4219,N_3707,N_3567);
nand U4220 (N_4220,N_3655,N_3984);
nor U4221 (N_4221,N_3946,N_3526);
or U4222 (N_4222,N_3758,N_3561);
nand U4223 (N_4223,N_3775,N_3899);
xnor U4224 (N_4224,N_3575,N_3572);
and U4225 (N_4225,N_3923,N_3896);
xor U4226 (N_4226,N_3592,N_3540);
and U4227 (N_4227,N_3900,N_3742);
nor U4228 (N_4228,N_3907,N_3875);
nand U4229 (N_4229,N_3981,N_3744);
or U4230 (N_4230,N_3713,N_3949);
nor U4231 (N_4231,N_3677,N_3635);
or U4232 (N_4232,N_3936,N_3641);
nand U4233 (N_4233,N_3609,N_3717);
and U4234 (N_4234,N_3889,N_3544);
and U4235 (N_4235,N_3847,N_3962);
nor U4236 (N_4236,N_3695,N_3621);
nor U4237 (N_4237,N_3638,N_3691);
or U4238 (N_4238,N_3837,N_3759);
xnor U4239 (N_4239,N_3766,N_3761);
nor U4240 (N_4240,N_3671,N_3528);
and U4241 (N_4241,N_3965,N_3983);
or U4242 (N_4242,N_3545,N_3797);
or U4243 (N_4243,N_3527,N_3955);
and U4244 (N_4244,N_3726,N_3611);
or U4245 (N_4245,N_3901,N_3818);
and U4246 (N_4246,N_3500,N_3541);
or U4247 (N_4247,N_3822,N_3793);
nor U4248 (N_4248,N_3579,N_3518);
nand U4249 (N_4249,N_3721,N_3807);
nor U4250 (N_4250,N_3776,N_3934);
or U4251 (N_4251,N_3880,N_3848);
or U4252 (N_4252,N_3956,N_3939);
or U4253 (N_4253,N_3511,N_3749);
nand U4254 (N_4254,N_3693,N_3524);
nor U4255 (N_4255,N_3813,N_3595);
and U4256 (N_4256,N_3938,N_3736);
nand U4257 (N_4257,N_3548,N_3720);
and U4258 (N_4258,N_3843,N_3604);
nor U4259 (N_4259,N_3715,N_3719);
and U4260 (N_4260,N_3758,N_3510);
and U4261 (N_4261,N_3788,N_3764);
and U4262 (N_4262,N_3829,N_3504);
or U4263 (N_4263,N_3546,N_3913);
nand U4264 (N_4264,N_3608,N_3693);
and U4265 (N_4265,N_3738,N_3670);
nand U4266 (N_4266,N_3884,N_3613);
nor U4267 (N_4267,N_3527,N_3923);
and U4268 (N_4268,N_3588,N_3602);
nand U4269 (N_4269,N_3951,N_3629);
nor U4270 (N_4270,N_3988,N_3922);
nor U4271 (N_4271,N_3738,N_3775);
and U4272 (N_4272,N_3558,N_3561);
nand U4273 (N_4273,N_3626,N_3660);
xnor U4274 (N_4274,N_3548,N_3944);
and U4275 (N_4275,N_3930,N_3618);
nand U4276 (N_4276,N_3526,N_3864);
xnor U4277 (N_4277,N_3710,N_3813);
nand U4278 (N_4278,N_3769,N_3527);
and U4279 (N_4279,N_3555,N_3690);
xnor U4280 (N_4280,N_3787,N_3564);
nand U4281 (N_4281,N_3633,N_3634);
or U4282 (N_4282,N_3601,N_3925);
nor U4283 (N_4283,N_3635,N_3579);
and U4284 (N_4284,N_3986,N_3671);
and U4285 (N_4285,N_3663,N_3787);
or U4286 (N_4286,N_3695,N_3880);
or U4287 (N_4287,N_3883,N_3991);
xnor U4288 (N_4288,N_3728,N_3795);
nor U4289 (N_4289,N_3501,N_3957);
nand U4290 (N_4290,N_3815,N_3740);
nor U4291 (N_4291,N_3956,N_3691);
and U4292 (N_4292,N_3648,N_3900);
and U4293 (N_4293,N_3692,N_3604);
and U4294 (N_4294,N_3923,N_3515);
or U4295 (N_4295,N_3570,N_3622);
or U4296 (N_4296,N_3637,N_3799);
nand U4297 (N_4297,N_3642,N_3794);
nor U4298 (N_4298,N_3624,N_3792);
or U4299 (N_4299,N_3541,N_3658);
xnor U4300 (N_4300,N_3806,N_3865);
or U4301 (N_4301,N_3914,N_3706);
and U4302 (N_4302,N_3879,N_3630);
xor U4303 (N_4303,N_3706,N_3726);
and U4304 (N_4304,N_3530,N_3672);
or U4305 (N_4305,N_3891,N_3539);
and U4306 (N_4306,N_3512,N_3840);
or U4307 (N_4307,N_3711,N_3947);
nor U4308 (N_4308,N_3520,N_3667);
nor U4309 (N_4309,N_3945,N_3904);
and U4310 (N_4310,N_3699,N_3536);
or U4311 (N_4311,N_3863,N_3531);
nand U4312 (N_4312,N_3594,N_3917);
nor U4313 (N_4313,N_3750,N_3839);
nor U4314 (N_4314,N_3824,N_3558);
nor U4315 (N_4315,N_3919,N_3915);
and U4316 (N_4316,N_3995,N_3589);
or U4317 (N_4317,N_3558,N_3669);
nand U4318 (N_4318,N_3513,N_3762);
nor U4319 (N_4319,N_3869,N_3972);
and U4320 (N_4320,N_3910,N_3751);
or U4321 (N_4321,N_3647,N_3870);
xnor U4322 (N_4322,N_3979,N_3943);
and U4323 (N_4323,N_3691,N_3757);
nor U4324 (N_4324,N_3761,N_3782);
nor U4325 (N_4325,N_3709,N_3968);
and U4326 (N_4326,N_3529,N_3720);
or U4327 (N_4327,N_3536,N_3887);
nand U4328 (N_4328,N_3787,N_3837);
or U4329 (N_4329,N_3921,N_3938);
or U4330 (N_4330,N_3882,N_3726);
nand U4331 (N_4331,N_3668,N_3980);
or U4332 (N_4332,N_3504,N_3741);
or U4333 (N_4333,N_3610,N_3585);
or U4334 (N_4334,N_3987,N_3978);
or U4335 (N_4335,N_3661,N_3526);
xor U4336 (N_4336,N_3564,N_3660);
and U4337 (N_4337,N_3653,N_3780);
nand U4338 (N_4338,N_3686,N_3911);
and U4339 (N_4339,N_3647,N_3826);
nand U4340 (N_4340,N_3979,N_3782);
nand U4341 (N_4341,N_3662,N_3703);
and U4342 (N_4342,N_3653,N_3589);
or U4343 (N_4343,N_3675,N_3565);
nor U4344 (N_4344,N_3506,N_3871);
and U4345 (N_4345,N_3978,N_3857);
or U4346 (N_4346,N_3846,N_3849);
or U4347 (N_4347,N_3856,N_3638);
or U4348 (N_4348,N_3581,N_3977);
or U4349 (N_4349,N_3567,N_3889);
and U4350 (N_4350,N_3527,N_3571);
or U4351 (N_4351,N_3587,N_3883);
nor U4352 (N_4352,N_3839,N_3970);
nor U4353 (N_4353,N_3889,N_3734);
and U4354 (N_4354,N_3794,N_3554);
nor U4355 (N_4355,N_3577,N_3677);
and U4356 (N_4356,N_3750,N_3931);
nor U4357 (N_4357,N_3901,N_3694);
xor U4358 (N_4358,N_3777,N_3768);
or U4359 (N_4359,N_3951,N_3511);
and U4360 (N_4360,N_3535,N_3774);
or U4361 (N_4361,N_3680,N_3684);
or U4362 (N_4362,N_3848,N_3668);
nand U4363 (N_4363,N_3568,N_3745);
or U4364 (N_4364,N_3504,N_3681);
and U4365 (N_4365,N_3681,N_3890);
or U4366 (N_4366,N_3970,N_3571);
nand U4367 (N_4367,N_3616,N_3579);
and U4368 (N_4368,N_3953,N_3694);
or U4369 (N_4369,N_3764,N_3679);
or U4370 (N_4370,N_3725,N_3828);
nand U4371 (N_4371,N_3992,N_3555);
or U4372 (N_4372,N_3877,N_3849);
xor U4373 (N_4373,N_3862,N_3872);
nor U4374 (N_4374,N_3774,N_3669);
or U4375 (N_4375,N_3743,N_3932);
and U4376 (N_4376,N_3584,N_3672);
nor U4377 (N_4377,N_3904,N_3982);
nor U4378 (N_4378,N_3774,N_3650);
nand U4379 (N_4379,N_3821,N_3886);
nor U4380 (N_4380,N_3554,N_3560);
xnor U4381 (N_4381,N_3894,N_3799);
nor U4382 (N_4382,N_3600,N_3517);
and U4383 (N_4383,N_3703,N_3912);
nand U4384 (N_4384,N_3621,N_3737);
xor U4385 (N_4385,N_3815,N_3667);
nand U4386 (N_4386,N_3854,N_3828);
nor U4387 (N_4387,N_3665,N_3760);
nand U4388 (N_4388,N_3630,N_3616);
nor U4389 (N_4389,N_3525,N_3900);
and U4390 (N_4390,N_3742,N_3670);
or U4391 (N_4391,N_3503,N_3840);
nand U4392 (N_4392,N_3548,N_3730);
nor U4393 (N_4393,N_3808,N_3787);
nor U4394 (N_4394,N_3938,N_3937);
nor U4395 (N_4395,N_3863,N_3936);
and U4396 (N_4396,N_3853,N_3691);
nor U4397 (N_4397,N_3814,N_3741);
xnor U4398 (N_4398,N_3714,N_3501);
nand U4399 (N_4399,N_3824,N_3607);
nand U4400 (N_4400,N_3785,N_3860);
nand U4401 (N_4401,N_3866,N_3960);
or U4402 (N_4402,N_3766,N_3631);
nor U4403 (N_4403,N_3733,N_3790);
and U4404 (N_4404,N_3912,N_3746);
nand U4405 (N_4405,N_3581,N_3897);
nand U4406 (N_4406,N_3611,N_3548);
or U4407 (N_4407,N_3711,N_3591);
or U4408 (N_4408,N_3801,N_3581);
or U4409 (N_4409,N_3930,N_3980);
and U4410 (N_4410,N_3951,N_3568);
nor U4411 (N_4411,N_3948,N_3807);
or U4412 (N_4412,N_3750,N_3614);
or U4413 (N_4413,N_3981,N_3970);
or U4414 (N_4414,N_3661,N_3688);
nand U4415 (N_4415,N_3618,N_3660);
or U4416 (N_4416,N_3557,N_3771);
nor U4417 (N_4417,N_3583,N_3828);
or U4418 (N_4418,N_3999,N_3503);
nand U4419 (N_4419,N_3911,N_3745);
and U4420 (N_4420,N_3826,N_3921);
xnor U4421 (N_4421,N_3585,N_3575);
nor U4422 (N_4422,N_3625,N_3716);
and U4423 (N_4423,N_3931,N_3966);
and U4424 (N_4424,N_3633,N_3614);
nor U4425 (N_4425,N_3520,N_3664);
or U4426 (N_4426,N_3697,N_3655);
nor U4427 (N_4427,N_3790,N_3757);
and U4428 (N_4428,N_3933,N_3590);
or U4429 (N_4429,N_3607,N_3880);
or U4430 (N_4430,N_3722,N_3963);
and U4431 (N_4431,N_3780,N_3758);
or U4432 (N_4432,N_3829,N_3601);
and U4433 (N_4433,N_3686,N_3954);
or U4434 (N_4434,N_3751,N_3982);
nand U4435 (N_4435,N_3614,N_3884);
or U4436 (N_4436,N_3643,N_3967);
or U4437 (N_4437,N_3604,N_3681);
nor U4438 (N_4438,N_3865,N_3968);
nor U4439 (N_4439,N_3726,N_3999);
xnor U4440 (N_4440,N_3519,N_3711);
nor U4441 (N_4441,N_3791,N_3666);
nand U4442 (N_4442,N_3944,N_3824);
and U4443 (N_4443,N_3914,N_3837);
and U4444 (N_4444,N_3806,N_3978);
nor U4445 (N_4445,N_3722,N_3691);
and U4446 (N_4446,N_3510,N_3548);
nand U4447 (N_4447,N_3750,N_3546);
nand U4448 (N_4448,N_3865,N_3758);
nand U4449 (N_4449,N_3661,N_3524);
nand U4450 (N_4450,N_3519,N_3621);
or U4451 (N_4451,N_3622,N_3884);
and U4452 (N_4452,N_3788,N_3821);
and U4453 (N_4453,N_3565,N_3837);
nand U4454 (N_4454,N_3818,N_3592);
xor U4455 (N_4455,N_3517,N_3664);
nor U4456 (N_4456,N_3597,N_3930);
nor U4457 (N_4457,N_3795,N_3706);
nand U4458 (N_4458,N_3848,N_3529);
and U4459 (N_4459,N_3639,N_3728);
nand U4460 (N_4460,N_3507,N_3526);
and U4461 (N_4461,N_3504,N_3891);
xnor U4462 (N_4462,N_3931,N_3651);
nand U4463 (N_4463,N_3661,N_3670);
or U4464 (N_4464,N_3776,N_3896);
and U4465 (N_4465,N_3507,N_3773);
nor U4466 (N_4466,N_3912,N_3532);
xor U4467 (N_4467,N_3518,N_3918);
nand U4468 (N_4468,N_3555,N_3585);
nor U4469 (N_4469,N_3523,N_3643);
or U4470 (N_4470,N_3954,N_3620);
or U4471 (N_4471,N_3904,N_3753);
xor U4472 (N_4472,N_3748,N_3829);
nor U4473 (N_4473,N_3563,N_3726);
or U4474 (N_4474,N_3502,N_3948);
nand U4475 (N_4475,N_3527,N_3737);
xor U4476 (N_4476,N_3836,N_3927);
nor U4477 (N_4477,N_3607,N_3621);
nor U4478 (N_4478,N_3668,N_3647);
and U4479 (N_4479,N_3825,N_3876);
nor U4480 (N_4480,N_3656,N_3851);
and U4481 (N_4481,N_3917,N_3891);
nand U4482 (N_4482,N_3993,N_3538);
nor U4483 (N_4483,N_3519,N_3560);
or U4484 (N_4484,N_3954,N_3787);
and U4485 (N_4485,N_3751,N_3876);
and U4486 (N_4486,N_3715,N_3552);
nor U4487 (N_4487,N_3608,N_3750);
nor U4488 (N_4488,N_3709,N_3663);
nand U4489 (N_4489,N_3722,N_3869);
nand U4490 (N_4490,N_3764,N_3648);
xor U4491 (N_4491,N_3876,N_3507);
or U4492 (N_4492,N_3921,N_3548);
or U4493 (N_4493,N_3643,N_3889);
xor U4494 (N_4494,N_3700,N_3627);
nor U4495 (N_4495,N_3574,N_3642);
or U4496 (N_4496,N_3877,N_3581);
xor U4497 (N_4497,N_3562,N_3650);
nor U4498 (N_4498,N_3874,N_3914);
or U4499 (N_4499,N_3812,N_3604);
and U4500 (N_4500,N_4056,N_4080);
nor U4501 (N_4501,N_4187,N_4250);
nand U4502 (N_4502,N_4165,N_4248);
and U4503 (N_4503,N_4284,N_4263);
nand U4504 (N_4504,N_4271,N_4355);
or U4505 (N_4505,N_4148,N_4132);
nand U4506 (N_4506,N_4314,N_4329);
nor U4507 (N_4507,N_4398,N_4053);
nor U4508 (N_4508,N_4048,N_4036);
or U4509 (N_4509,N_4328,N_4473);
nand U4510 (N_4510,N_4443,N_4421);
and U4511 (N_4511,N_4188,N_4228);
or U4512 (N_4512,N_4315,N_4466);
nand U4513 (N_4513,N_4190,N_4456);
or U4514 (N_4514,N_4418,N_4462);
and U4515 (N_4515,N_4390,N_4335);
or U4516 (N_4516,N_4130,N_4268);
or U4517 (N_4517,N_4078,N_4186);
xor U4518 (N_4518,N_4363,N_4380);
or U4519 (N_4519,N_4256,N_4361);
nor U4520 (N_4520,N_4150,N_4246);
or U4521 (N_4521,N_4478,N_4157);
or U4522 (N_4522,N_4205,N_4341);
nor U4523 (N_4523,N_4270,N_4230);
nor U4524 (N_4524,N_4326,N_4229);
xor U4525 (N_4525,N_4495,N_4136);
and U4526 (N_4526,N_4274,N_4345);
nand U4527 (N_4527,N_4338,N_4392);
nor U4528 (N_4528,N_4389,N_4360);
xnor U4529 (N_4529,N_4425,N_4038);
nor U4530 (N_4530,N_4379,N_4451);
nor U4531 (N_4531,N_4318,N_4342);
nand U4532 (N_4532,N_4202,N_4484);
nor U4533 (N_4533,N_4181,N_4195);
and U4534 (N_4534,N_4383,N_4377);
nand U4535 (N_4535,N_4498,N_4412);
nor U4536 (N_4536,N_4305,N_4135);
and U4537 (N_4537,N_4481,N_4381);
or U4538 (N_4538,N_4204,N_4405);
or U4539 (N_4539,N_4233,N_4175);
nor U4540 (N_4540,N_4309,N_4403);
and U4541 (N_4541,N_4156,N_4127);
or U4542 (N_4542,N_4023,N_4450);
nor U4543 (N_4543,N_4082,N_4168);
and U4544 (N_4544,N_4171,N_4468);
and U4545 (N_4545,N_4051,N_4073);
and U4546 (N_4546,N_4200,N_4416);
nand U4547 (N_4547,N_4084,N_4428);
xor U4548 (N_4548,N_4308,N_4296);
nand U4549 (N_4549,N_4417,N_4359);
nor U4550 (N_4550,N_4266,N_4126);
or U4551 (N_4551,N_4217,N_4034);
and U4552 (N_4552,N_4365,N_4141);
xnor U4553 (N_4553,N_4475,N_4069);
nand U4554 (N_4554,N_4460,N_4358);
and U4555 (N_4555,N_4112,N_4139);
nor U4556 (N_4556,N_4254,N_4159);
nand U4557 (N_4557,N_4154,N_4120);
or U4558 (N_4558,N_4201,N_4144);
nand U4559 (N_4559,N_4430,N_4324);
and U4560 (N_4560,N_4004,N_4226);
nand U4561 (N_4561,N_4114,N_4104);
and U4562 (N_4562,N_4407,N_4123);
or U4563 (N_4563,N_4457,N_4325);
xor U4564 (N_4564,N_4350,N_4477);
nand U4565 (N_4565,N_4424,N_4353);
or U4566 (N_4566,N_4062,N_4232);
nand U4567 (N_4567,N_4406,N_4452);
nand U4568 (N_4568,N_4098,N_4367);
nand U4569 (N_4569,N_4423,N_4373);
nand U4570 (N_4570,N_4280,N_4420);
and U4571 (N_4571,N_4458,N_4221);
and U4572 (N_4572,N_4153,N_4486);
and U4573 (N_4573,N_4317,N_4343);
nor U4574 (N_4574,N_4009,N_4033);
and U4575 (N_4575,N_4439,N_4362);
nand U4576 (N_4576,N_4485,N_4149);
nand U4577 (N_4577,N_4162,N_4267);
and U4578 (N_4578,N_4238,N_4313);
xnor U4579 (N_4579,N_4102,N_4010);
and U4580 (N_4580,N_4447,N_4099);
nor U4581 (N_4581,N_4283,N_4075);
and U4582 (N_4582,N_4087,N_4470);
and U4583 (N_4583,N_4286,N_4349);
or U4584 (N_4584,N_4101,N_4320);
xor U4585 (N_4585,N_4368,N_4241);
nand U4586 (N_4586,N_4096,N_4259);
nand U4587 (N_4587,N_4088,N_4289);
nand U4588 (N_4588,N_4411,N_4081);
or U4589 (N_4589,N_4322,N_4278);
nand U4590 (N_4590,N_4223,N_4437);
or U4591 (N_4591,N_4442,N_4323);
or U4592 (N_4592,N_4446,N_4196);
nor U4593 (N_4593,N_4108,N_4086);
and U4594 (N_4594,N_4163,N_4001);
and U4595 (N_4595,N_4167,N_4191);
and U4596 (N_4596,N_4354,N_4334);
and U4597 (N_4597,N_4454,N_4337);
nand U4598 (N_4598,N_4453,N_4306);
or U4599 (N_4599,N_4094,N_4044);
nor U4600 (N_4600,N_4237,N_4109);
xnor U4601 (N_4601,N_4319,N_4193);
nor U4602 (N_4602,N_4291,N_4106);
and U4603 (N_4603,N_4269,N_4002);
and U4604 (N_4604,N_4093,N_4275);
and U4605 (N_4605,N_4170,N_4216);
nand U4606 (N_4606,N_4046,N_4068);
and U4607 (N_4607,N_4340,N_4000);
nand U4608 (N_4608,N_4474,N_4077);
or U4609 (N_4609,N_4448,N_4281);
nor U4610 (N_4610,N_4372,N_4143);
nand U4611 (N_4611,N_4387,N_4017);
or U4612 (N_4612,N_4436,N_4006);
nand U4613 (N_4613,N_4219,N_4067);
or U4614 (N_4614,N_4161,N_4197);
or U4615 (N_4615,N_4152,N_4321);
or U4616 (N_4616,N_4332,N_4185);
and U4617 (N_4617,N_4066,N_4176);
nand U4618 (N_4618,N_4116,N_4255);
xor U4619 (N_4619,N_4210,N_4307);
nor U4620 (N_4620,N_4333,N_4414);
nand U4621 (N_4621,N_4287,N_4465);
xnor U4622 (N_4622,N_4261,N_4007);
or U4623 (N_4623,N_4169,N_4083);
and U4624 (N_4624,N_4312,N_4276);
nand U4625 (N_4625,N_4364,N_4397);
and U4626 (N_4626,N_4199,N_4218);
and U4627 (N_4627,N_4282,N_4013);
nand U4628 (N_4628,N_4074,N_4045);
xnor U4629 (N_4629,N_4297,N_4131);
nor U4630 (N_4630,N_4018,N_4061);
or U4631 (N_4631,N_4455,N_4145);
or U4632 (N_4632,N_4396,N_4124);
nand U4633 (N_4633,N_4408,N_4103);
xor U4634 (N_4634,N_4395,N_4265);
or U4635 (N_4635,N_4253,N_4234);
or U4636 (N_4636,N_4180,N_4203);
or U4637 (N_4637,N_4370,N_4240);
or U4638 (N_4638,N_4304,N_4371);
nor U4639 (N_4639,N_4311,N_4140);
nand U4640 (N_4640,N_4129,N_4060);
nor U4641 (N_4641,N_4290,N_4251);
and U4642 (N_4642,N_4438,N_4435);
nor U4643 (N_4643,N_4085,N_4483);
nand U4644 (N_4644,N_4327,N_4294);
or U4645 (N_4645,N_4121,N_4277);
or U4646 (N_4646,N_4347,N_4258);
nor U4647 (N_4647,N_4015,N_4493);
nand U4648 (N_4648,N_4142,N_4206);
or U4649 (N_4649,N_4182,N_4419);
xnor U4650 (N_4650,N_4260,N_4118);
nor U4651 (N_4651,N_4344,N_4492);
and U4652 (N_4652,N_4050,N_4295);
nor U4653 (N_4653,N_4415,N_4441);
nor U4654 (N_4654,N_4279,N_4490);
and U4655 (N_4655,N_4429,N_4166);
xnor U4656 (N_4656,N_4298,N_4264);
and U4657 (N_4657,N_4054,N_4330);
and U4658 (N_4658,N_4352,N_4225);
nor U4659 (N_4659,N_4422,N_4339);
nor U4660 (N_4660,N_4198,N_4461);
nand U4661 (N_4661,N_4027,N_4164);
nand U4662 (N_4662,N_4331,N_4024);
nor U4663 (N_4663,N_4310,N_4160);
nor U4664 (N_4664,N_4463,N_4091);
nand U4665 (N_4665,N_4026,N_4480);
nand U4666 (N_4666,N_4348,N_4028);
and U4667 (N_4667,N_4346,N_4158);
and U4668 (N_4668,N_4400,N_4394);
or U4669 (N_4669,N_4244,N_4172);
xor U4670 (N_4670,N_4496,N_4440);
nand U4671 (N_4671,N_4300,N_4385);
xor U4672 (N_4672,N_4467,N_4211);
or U4673 (N_4673,N_4243,N_4155);
nand U4674 (N_4674,N_4316,N_4137);
or U4675 (N_4675,N_4292,N_4090);
nand U4676 (N_4676,N_4374,N_4151);
nor U4677 (N_4677,N_4183,N_4378);
nand U4678 (N_4678,N_4014,N_4031);
nand U4679 (N_4679,N_4147,N_4499);
and U4680 (N_4680,N_4071,N_4449);
or U4681 (N_4681,N_4035,N_4366);
nor U4682 (N_4682,N_4356,N_4097);
xor U4683 (N_4683,N_4043,N_4011);
and U4684 (N_4684,N_4065,N_4111);
xor U4685 (N_4685,N_4273,N_4138);
xor U4686 (N_4686,N_4236,N_4491);
and U4687 (N_4687,N_4174,N_4189);
nor U4688 (N_4688,N_4494,N_4427);
nand U4689 (N_4689,N_4016,N_4012);
nand U4690 (N_4690,N_4376,N_4469);
and U4691 (N_4691,N_4113,N_4459);
xor U4692 (N_4692,N_4299,N_4285);
or U4693 (N_4693,N_4433,N_4122);
nand U4694 (N_4694,N_4386,N_4262);
nand U4695 (N_4695,N_4092,N_4245);
or U4696 (N_4696,N_4030,N_4444);
and U4697 (N_4697,N_4057,N_4063);
or U4698 (N_4698,N_4215,N_4041);
nor U4699 (N_4699,N_4076,N_4487);
nor U4700 (N_4700,N_4375,N_4357);
nor U4701 (N_4701,N_4242,N_4489);
nor U4702 (N_4702,N_4293,N_4224);
nand U4703 (N_4703,N_4212,N_4302);
nand U4704 (N_4704,N_4184,N_4039);
or U4705 (N_4705,N_4404,N_4472);
nand U4706 (N_4706,N_4208,N_4471);
xnor U4707 (N_4707,N_4052,N_4005);
and U4708 (N_4708,N_4047,N_4133);
or U4709 (N_4709,N_4476,N_4058);
nand U4710 (N_4710,N_4008,N_4072);
and U4711 (N_4711,N_4432,N_4105);
nor U4712 (N_4712,N_4445,N_4207);
nand U4713 (N_4713,N_4059,N_4431);
or U4714 (N_4714,N_4095,N_4235);
and U4715 (N_4715,N_4301,N_4369);
and U4716 (N_4716,N_4021,N_4049);
or U4717 (N_4717,N_4192,N_4464);
xnor U4718 (N_4718,N_4288,N_4179);
or U4719 (N_4719,N_4037,N_4107);
nand U4720 (N_4720,N_4336,N_4214);
or U4721 (N_4721,N_4064,N_4388);
nor U4722 (N_4722,N_4222,N_4413);
nor U4723 (N_4723,N_4134,N_4257);
or U4724 (N_4724,N_4488,N_4384);
nor U4725 (N_4725,N_4402,N_4220);
nand U4726 (N_4726,N_4019,N_4177);
or U4727 (N_4727,N_4040,N_4194);
or U4728 (N_4728,N_4089,N_4213);
or U4729 (N_4729,N_4125,N_4231);
nand U4730 (N_4730,N_4032,N_4003);
nand U4731 (N_4731,N_4247,N_4110);
and U4732 (N_4732,N_4128,N_4173);
nand U4733 (N_4733,N_4401,N_4482);
or U4734 (N_4734,N_4391,N_4029);
xnor U4735 (N_4735,N_4351,N_4249);
and U4736 (N_4736,N_4410,N_4022);
and U4737 (N_4737,N_4115,N_4272);
nor U4738 (N_4738,N_4252,N_4227);
nand U4739 (N_4739,N_4178,N_4146);
and U4740 (N_4740,N_4025,N_4399);
xor U4741 (N_4741,N_4434,N_4479);
or U4742 (N_4742,N_4209,N_4426);
xnor U4743 (N_4743,N_4409,N_4393);
nor U4744 (N_4744,N_4079,N_4100);
nor U4745 (N_4745,N_4070,N_4119);
and U4746 (N_4746,N_4055,N_4042);
or U4747 (N_4747,N_4020,N_4303);
nand U4748 (N_4748,N_4117,N_4239);
nor U4749 (N_4749,N_4382,N_4497);
and U4750 (N_4750,N_4364,N_4002);
and U4751 (N_4751,N_4053,N_4104);
xor U4752 (N_4752,N_4028,N_4018);
nand U4753 (N_4753,N_4291,N_4393);
or U4754 (N_4754,N_4488,N_4190);
and U4755 (N_4755,N_4051,N_4002);
and U4756 (N_4756,N_4351,N_4037);
and U4757 (N_4757,N_4264,N_4089);
nand U4758 (N_4758,N_4332,N_4158);
nand U4759 (N_4759,N_4497,N_4203);
nand U4760 (N_4760,N_4028,N_4341);
nor U4761 (N_4761,N_4473,N_4102);
nor U4762 (N_4762,N_4462,N_4444);
or U4763 (N_4763,N_4281,N_4074);
nor U4764 (N_4764,N_4160,N_4191);
or U4765 (N_4765,N_4271,N_4000);
or U4766 (N_4766,N_4436,N_4184);
or U4767 (N_4767,N_4026,N_4483);
nand U4768 (N_4768,N_4194,N_4057);
and U4769 (N_4769,N_4115,N_4107);
xor U4770 (N_4770,N_4170,N_4139);
nand U4771 (N_4771,N_4429,N_4045);
xnor U4772 (N_4772,N_4469,N_4159);
nor U4773 (N_4773,N_4437,N_4421);
nor U4774 (N_4774,N_4189,N_4344);
nand U4775 (N_4775,N_4177,N_4425);
and U4776 (N_4776,N_4341,N_4244);
xnor U4777 (N_4777,N_4263,N_4433);
nand U4778 (N_4778,N_4444,N_4177);
nand U4779 (N_4779,N_4390,N_4030);
and U4780 (N_4780,N_4381,N_4009);
nor U4781 (N_4781,N_4454,N_4152);
or U4782 (N_4782,N_4367,N_4036);
nand U4783 (N_4783,N_4034,N_4173);
nand U4784 (N_4784,N_4329,N_4438);
or U4785 (N_4785,N_4198,N_4209);
nor U4786 (N_4786,N_4288,N_4091);
nor U4787 (N_4787,N_4376,N_4061);
nand U4788 (N_4788,N_4394,N_4234);
xnor U4789 (N_4789,N_4026,N_4448);
nor U4790 (N_4790,N_4321,N_4347);
and U4791 (N_4791,N_4251,N_4205);
and U4792 (N_4792,N_4177,N_4012);
and U4793 (N_4793,N_4338,N_4275);
nand U4794 (N_4794,N_4056,N_4071);
nor U4795 (N_4795,N_4163,N_4330);
or U4796 (N_4796,N_4456,N_4009);
and U4797 (N_4797,N_4431,N_4193);
xor U4798 (N_4798,N_4101,N_4212);
nor U4799 (N_4799,N_4387,N_4220);
xor U4800 (N_4800,N_4457,N_4372);
or U4801 (N_4801,N_4004,N_4386);
nand U4802 (N_4802,N_4400,N_4180);
nand U4803 (N_4803,N_4322,N_4248);
and U4804 (N_4804,N_4398,N_4006);
nor U4805 (N_4805,N_4107,N_4340);
nor U4806 (N_4806,N_4447,N_4074);
nor U4807 (N_4807,N_4134,N_4438);
nand U4808 (N_4808,N_4120,N_4173);
nand U4809 (N_4809,N_4301,N_4144);
nand U4810 (N_4810,N_4123,N_4129);
nor U4811 (N_4811,N_4198,N_4238);
or U4812 (N_4812,N_4131,N_4389);
and U4813 (N_4813,N_4273,N_4375);
nor U4814 (N_4814,N_4344,N_4075);
nor U4815 (N_4815,N_4434,N_4230);
xor U4816 (N_4816,N_4427,N_4120);
or U4817 (N_4817,N_4048,N_4073);
and U4818 (N_4818,N_4039,N_4151);
nand U4819 (N_4819,N_4317,N_4146);
nand U4820 (N_4820,N_4246,N_4082);
and U4821 (N_4821,N_4464,N_4367);
nand U4822 (N_4822,N_4315,N_4141);
and U4823 (N_4823,N_4025,N_4462);
nor U4824 (N_4824,N_4353,N_4241);
nor U4825 (N_4825,N_4359,N_4379);
nand U4826 (N_4826,N_4046,N_4014);
and U4827 (N_4827,N_4124,N_4479);
nor U4828 (N_4828,N_4299,N_4436);
xor U4829 (N_4829,N_4244,N_4456);
and U4830 (N_4830,N_4013,N_4104);
and U4831 (N_4831,N_4384,N_4252);
or U4832 (N_4832,N_4471,N_4282);
nand U4833 (N_4833,N_4103,N_4141);
or U4834 (N_4834,N_4091,N_4280);
or U4835 (N_4835,N_4263,N_4166);
nor U4836 (N_4836,N_4194,N_4324);
or U4837 (N_4837,N_4084,N_4062);
and U4838 (N_4838,N_4167,N_4031);
or U4839 (N_4839,N_4293,N_4314);
and U4840 (N_4840,N_4207,N_4384);
and U4841 (N_4841,N_4253,N_4173);
or U4842 (N_4842,N_4117,N_4328);
nand U4843 (N_4843,N_4321,N_4437);
and U4844 (N_4844,N_4424,N_4023);
nand U4845 (N_4845,N_4397,N_4085);
and U4846 (N_4846,N_4452,N_4255);
or U4847 (N_4847,N_4496,N_4494);
and U4848 (N_4848,N_4329,N_4463);
nor U4849 (N_4849,N_4222,N_4032);
and U4850 (N_4850,N_4337,N_4215);
and U4851 (N_4851,N_4312,N_4457);
nor U4852 (N_4852,N_4295,N_4131);
nor U4853 (N_4853,N_4279,N_4437);
or U4854 (N_4854,N_4090,N_4337);
and U4855 (N_4855,N_4207,N_4065);
nand U4856 (N_4856,N_4265,N_4125);
or U4857 (N_4857,N_4049,N_4008);
and U4858 (N_4858,N_4343,N_4177);
nor U4859 (N_4859,N_4374,N_4450);
or U4860 (N_4860,N_4221,N_4096);
and U4861 (N_4861,N_4206,N_4108);
and U4862 (N_4862,N_4299,N_4094);
or U4863 (N_4863,N_4412,N_4425);
or U4864 (N_4864,N_4247,N_4147);
or U4865 (N_4865,N_4470,N_4095);
xor U4866 (N_4866,N_4088,N_4262);
nand U4867 (N_4867,N_4177,N_4046);
nor U4868 (N_4868,N_4018,N_4400);
and U4869 (N_4869,N_4310,N_4062);
and U4870 (N_4870,N_4353,N_4249);
and U4871 (N_4871,N_4043,N_4345);
nand U4872 (N_4872,N_4278,N_4093);
or U4873 (N_4873,N_4246,N_4162);
and U4874 (N_4874,N_4302,N_4303);
nand U4875 (N_4875,N_4048,N_4458);
nand U4876 (N_4876,N_4105,N_4006);
nand U4877 (N_4877,N_4280,N_4309);
nor U4878 (N_4878,N_4478,N_4319);
and U4879 (N_4879,N_4251,N_4442);
and U4880 (N_4880,N_4369,N_4437);
or U4881 (N_4881,N_4341,N_4209);
nor U4882 (N_4882,N_4369,N_4076);
nand U4883 (N_4883,N_4465,N_4003);
nor U4884 (N_4884,N_4347,N_4170);
or U4885 (N_4885,N_4334,N_4350);
and U4886 (N_4886,N_4450,N_4425);
xor U4887 (N_4887,N_4393,N_4262);
or U4888 (N_4888,N_4453,N_4305);
nor U4889 (N_4889,N_4139,N_4424);
nand U4890 (N_4890,N_4318,N_4306);
nand U4891 (N_4891,N_4101,N_4300);
and U4892 (N_4892,N_4011,N_4168);
nand U4893 (N_4893,N_4236,N_4259);
nand U4894 (N_4894,N_4475,N_4038);
nand U4895 (N_4895,N_4030,N_4014);
and U4896 (N_4896,N_4247,N_4285);
or U4897 (N_4897,N_4288,N_4152);
nor U4898 (N_4898,N_4376,N_4054);
and U4899 (N_4899,N_4399,N_4335);
nor U4900 (N_4900,N_4455,N_4407);
nand U4901 (N_4901,N_4268,N_4061);
and U4902 (N_4902,N_4304,N_4353);
nor U4903 (N_4903,N_4336,N_4480);
nand U4904 (N_4904,N_4371,N_4441);
nand U4905 (N_4905,N_4299,N_4414);
nand U4906 (N_4906,N_4112,N_4359);
and U4907 (N_4907,N_4115,N_4407);
xor U4908 (N_4908,N_4052,N_4193);
xor U4909 (N_4909,N_4208,N_4233);
nand U4910 (N_4910,N_4057,N_4493);
xnor U4911 (N_4911,N_4121,N_4000);
nand U4912 (N_4912,N_4313,N_4364);
and U4913 (N_4913,N_4138,N_4236);
and U4914 (N_4914,N_4011,N_4248);
nand U4915 (N_4915,N_4201,N_4284);
nand U4916 (N_4916,N_4160,N_4040);
xnor U4917 (N_4917,N_4269,N_4104);
or U4918 (N_4918,N_4303,N_4015);
and U4919 (N_4919,N_4257,N_4139);
and U4920 (N_4920,N_4390,N_4274);
or U4921 (N_4921,N_4258,N_4100);
nand U4922 (N_4922,N_4491,N_4285);
nor U4923 (N_4923,N_4468,N_4084);
nand U4924 (N_4924,N_4137,N_4213);
nand U4925 (N_4925,N_4339,N_4107);
and U4926 (N_4926,N_4417,N_4280);
nor U4927 (N_4927,N_4377,N_4233);
nor U4928 (N_4928,N_4351,N_4462);
nor U4929 (N_4929,N_4289,N_4388);
or U4930 (N_4930,N_4322,N_4122);
and U4931 (N_4931,N_4154,N_4334);
nor U4932 (N_4932,N_4104,N_4025);
or U4933 (N_4933,N_4422,N_4055);
nor U4934 (N_4934,N_4139,N_4284);
and U4935 (N_4935,N_4483,N_4059);
or U4936 (N_4936,N_4311,N_4491);
nand U4937 (N_4937,N_4294,N_4259);
nor U4938 (N_4938,N_4222,N_4138);
nor U4939 (N_4939,N_4309,N_4341);
and U4940 (N_4940,N_4341,N_4427);
or U4941 (N_4941,N_4442,N_4385);
and U4942 (N_4942,N_4460,N_4021);
nand U4943 (N_4943,N_4064,N_4407);
and U4944 (N_4944,N_4101,N_4172);
nor U4945 (N_4945,N_4341,N_4248);
or U4946 (N_4946,N_4227,N_4407);
and U4947 (N_4947,N_4066,N_4324);
nor U4948 (N_4948,N_4103,N_4428);
and U4949 (N_4949,N_4421,N_4388);
or U4950 (N_4950,N_4358,N_4308);
nand U4951 (N_4951,N_4217,N_4297);
nand U4952 (N_4952,N_4166,N_4027);
nand U4953 (N_4953,N_4094,N_4375);
nor U4954 (N_4954,N_4270,N_4338);
and U4955 (N_4955,N_4030,N_4294);
and U4956 (N_4956,N_4073,N_4109);
nand U4957 (N_4957,N_4370,N_4266);
nor U4958 (N_4958,N_4014,N_4357);
or U4959 (N_4959,N_4344,N_4232);
nand U4960 (N_4960,N_4201,N_4185);
nand U4961 (N_4961,N_4394,N_4450);
nor U4962 (N_4962,N_4455,N_4345);
or U4963 (N_4963,N_4308,N_4306);
nand U4964 (N_4964,N_4290,N_4221);
nor U4965 (N_4965,N_4105,N_4391);
nand U4966 (N_4966,N_4044,N_4032);
and U4967 (N_4967,N_4247,N_4004);
nand U4968 (N_4968,N_4184,N_4438);
nor U4969 (N_4969,N_4414,N_4436);
nor U4970 (N_4970,N_4423,N_4481);
and U4971 (N_4971,N_4481,N_4147);
nand U4972 (N_4972,N_4401,N_4060);
nand U4973 (N_4973,N_4312,N_4319);
xor U4974 (N_4974,N_4018,N_4166);
or U4975 (N_4975,N_4006,N_4273);
xor U4976 (N_4976,N_4297,N_4117);
nor U4977 (N_4977,N_4031,N_4159);
nor U4978 (N_4978,N_4225,N_4210);
or U4979 (N_4979,N_4126,N_4054);
and U4980 (N_4980,N_4415,N_4034);
nor U4981 (N_4981,N_4292,N_4278);
nand U4982 (N_4982,N_4122,N_4146);
nor U4983 (N_4983,N_4001,N_4057);
and U4984 (N_4984,N_4482,N_4219);
or U4985 (N_4985,N_4021,N_4106);
nand U4986 (N_4986,N_4208,N_4271);
nand U4987 (N_4987,N_4306,N_4096);
nor U4988 (N_4988,N_4379,N_4073);
nor U4989 (N_4989,N_4038,N_4248);
nand U4990 (N_4990,N_4040,N_4191);
nand U4991 (N_4991,N_4094,N_4205);
nor U4992 (N_4992,N_4168,N_4149);
nand U4993 (N_4993,N_4490,N_4207);
nand U4994 (N_4994,N_4105,N_4390);
and U4995 (N_4995,N_4334,N_4320);
or U4996 (N_4996,N_4283,N_4416);
and U4997 (N_4997,N_4208,N_4225);
and U4998 (N_4998,N_4017,N_4355);
and U4999 (N_4999,N_4317,N_4498);
nor U5000 (N_5000,N_4585,N_4849);
or U5001 (N_5001,N_4761,N_4663);
nand U5002 (N_5002,N_4624,N_4878);
and U5003 (N_5003,N_4809,N_4760);
xor U5004 (N_5004,N_4548,N_4994);
nand U5005 (N_5005,N_4867,N_4512);
nor U5006 (N_5006,N_4529,N_4909);
and U5007 (N_5007,N_4749,N_4623);
or U5008 (N_5008,N_4908,N_4816);
xnor U5009 (N_5009,N_4708,N_4590);
or U5010 (N_5010,N_4626,N_4521);
nand U5011 (N_5011,N_4975,N_4934);
nand U5012 (N_5012,N_4921,N_4891);
and U5013 (N_5013,N_4596,N_4756);
xor U5014 (N_5014,N_4656,N_4610);
nor U5015 (N_5015,N_4841,N_4915);
nand U5016 (N_5016,N_4592,N_4635);
or U5017 (N_5017,N_4573,N_4851);
nor U5018 (N_5018,N_4976,N_4781);
nand U5019 (N_5019,N_4959,N_4574);
xnor U5020 (N_5020,N_4614,N_4740);
and U5021 (N_5021,N_4981,N_4914);
and U5022 (N_5022,N_4741,N_4715);
nor U5023 (N_5023,N_4861,N_4834);
xor U5024 (N_5024,N_4580,N_4515);
xnor U5025 (N_5025,N_4848,N_4765);
or U5026 (N_5026,N_4714,N_4992);
or U5027 (N_5027,N_4968,N_4964);
nand U5028 (N_5028,N_4846,N_4583);
or U5029 (N_5029,N_4905,N_4742);
and U5030 (N_5030,N_4775,N_4784);
nand U5031 (N_5031,N_4653,N_4864);
or U5032 (N_5032,N_4997,N_4786);
and U5033 (N_5033,N_4900,N_4758);
or U5034 (N_5034,N_4526,N_4817);
and U5035 (N_5035,N_4931,N_4895);
or U5036 (N_5036,N_4984,N_4776);
and U5037 (N_5037,N_4979,N_4570);
and U5038 (N_5038,N_4683,N_4510);
and U5039 (N_5039,N_4854,N_4906);
nand U5040 (N_5040,N_4743,N_4812);
xor U5041 (N_5041,N_4607,N_4866);
xor U5042 (N_5042,N_4597,N_4824);
nor U5043 (N_5043,N_4606,N_4554);
and U5044 (N_5044,N_4733,N_4511);
and U5045 (N_5045,N_4990,N_4813);
and U5046 (N_5046,N_4528,N_4807);
or U5047 (N_5047,N_4978,N_4995);
nor U5048 (N_5048,N_4581,N_4639);
nand U5049 (N_5049,N_4871,N_4886);
or U5050 (N_5050,N_4540,N_4734);
xor U5051 (N_5051,N_4998,N_4702);
xnor U5052 (N_5052,N_4821,N_4564);
nor U5053 (N_5053,N_4599,N_4501);
or U5054 (N_5054,N_4919,N_4601);
and U5055 (N_5055,N_4869,N_4575);
nor U5056 (N_5056,N_4710,N_4693);
or U5057 (N_5057,N_4790,N_4520);
or U5058 (N_5058,N_4612,N_4666);
or U5059 (N_5059,N_4603,N_4772);
and U5060 (N_5060,N_4704,N_4634);
nor U5061 (N_5061,N_4883,N_4739);
or U5062 (N_5062,N_4945,N_4896);
or U5063 (N_5063,N_4766,N_4525);
or U5064 (N_5064,N_4796,N_4774);
or U5065 (N_5065,N_4565,N_4602);
and U5066 (N_5066,N_4753,N_4778);
nand U5067 (N_5067,N_4899,N_4865);
or U5068 (N_5068,N_4729,N_4609);
or U5069 (N_5069,N_4569,N_4792);
nor U5070 (N_5070,N_4587,N_4750);
or U5071 (N_5071,N_4991,N_4800);
nand U5072 (N_5072,N_4698,N_4611);
nor U5073 (N_5073,N_4810,N_4682);
nand U5074 (N_5074,N_4688,N_4549);
nor U5075 (N_5075,N_4628,N_4955);
and U5076 (N_5076,N_4657,N_4543);
and U5077 (N_5077,N_4694,N_4855);
nand U5078 (N_5078,N_4860,N_4880);
xor U5079 (N_5079,N_4811,N_4620);
or U5080 (N_5080,N_4689,N_4672);
xnor U5081 (N_5081,N_4820,N_4745);
nor U5082 (N_5082,N_4873,N_4922);
nor U5083 (N_5083,N_4884,N_4941);
and U5084 (N_5084,N_4731,N_4705);
and U5085 (N_5085,N_4932,N_4889);
and U5086 (N_5086,N_4948,N_4930);
or U5087 (N_5087,N_4957,N_4629);
nor U5088 (N_5088,N_4696,N_4722);
nor U5089 (N_5089,N_4579,N_4627);
and U5090 (N_5090,N_4982,N_4777);
or U5091 (N_5091,N_4615,N_4863);
nor U5092 (N_5092,N_4842,N_4539);
nand U5093 (N_5093,N_4736,N_4535);
nand U5094 (N_5094,N_4576,N_4716);
or U5095 (N_5095,N_4591,N_4928);
nor U5096 (N_5096,N_4522,N_4799);
and U5097 (N_5097,N_4578,N_4844);
and U5098 (N_5098,N_4801,N_4853);
xor U5099 (N_5099,N_4500,N_4542);
or U5100 (N_5100,N_4856,N_4648);
nand U5101 (N_5101,N_4970,N_4559);
nor U5102 (N_5102,N_4951,N_4996);
or U5103 (N_5103,N_4943,N_4637);
nand U5104 (N_5104,N_4840,N_4700);
xor U5105 (N_5105,N_4887,N_4684);
or U5106 (N_5106,N_4641,N_4665);
and U5107 (N_5107,N_4724,N_4795);
nand U5108 (N_5108,N_4897,N_4885);
and U5109 (N_5109,N_4757,N_4678);
or U5110 (N_5110,N_4551,N_4594);
and U5111 (N_5111,N_4797,N_4712);
and U5112 (N_5112,N_4836,N_4662);
and U5113 (N_5113,N_4654,N_4960);
and U5114 (N_5114,N_4793,N_4507);
nor U5115 (N_5115,N_4751,N_4822);
and U5116 (N_5116,N_4874,N_4649);
or U5117 (N_5117,N_4808,N_4767);
and U5118 (N_5118,N_4532,N_4787);
nor U5119 (N_5119,N_4933,N_4912);
and U5120 (N_5120,N_4725,N_4534);
nand U5121 (N_5121,N_4805,N_4942);
and U5122 (N_5122,N_4514,N_4862);
xor U5123 (N_5123,N_4572,N_4680);
and U5124 (N_5124,N_4843,N_4789);
nor U5125 (N_5125,N_4685,N_4831);
nand U5126 (N_5126,N_4927,N_4798);
nor U5127 (N_5127,N_4898,N_4769);
and U5128 (N_5128,N_4727,N_4903);
nand U5129 (N_5129,N_4910,N_4988);
and U5130 (N_5130,N_4770,N_4971);
and U5131 (N_5131,N_4806,N_4699);
and U5132 (N_5132,N_4818,N_4938);
nand U5133 (N_5133,N_4829,N_4621);
nand U5134 (N_5134,N_4558,N_4726);
xnor U5135 (N_5135,N_4827,N_4561);
or U5136 (N_5136,N_4950,N_4691);
nand U5137 (N_5137,N_4819,N_4783);
and U5138 (N_5138,N_4901,N_4717);
nand U5139 (N_5139,N_4850,N_4815);
nand U5140 (N_5140,N_4589,N_4646);
or U5141 (N_5141,N_4566,N_4703);
nand U5142 (N_5142,N_4872,N_4967);
and U5143 (N_5143,N_4645,N_4547);
or U5144 (N_5144,N_4926,N_4509);
or U5145 (N_5145,N_4764,N_4987);
or U5146 (N_5146,N_4524,N_4814);
xor U5147 (N_5147,N_4923,N_4674);
xor U5148 (N_5148,N_4593,N_4643);
nor U5149 (N_5149,N_4826,N_4692);
or U5150 (N_5150,N_4917,N_4782);
nor U5151 (N_5151,N_4954,N_4632);
or U5152 (N_5152,N_4527,N_4986);
nor U5153 (N_5153,N_4892,N_4619);
and U5154 (N_5154,N_4837,N_4730);
or U5155 (N_5155,N_4661,N_4961);
nor U5156 (N_5156,N_4802,N_4916);
or U5157 (N_5157,N_4616,N_4879);
nand U5158 (N_5158,N_4768,N_4659);
or U5159 (N_5159,N_4613,N_4541);
nor U5160 (N_5160,N_4845,N_4625);
and U5161 (N_5161,N_4630,N_4956);
nand U5162 (N_5162,N_4728,N_4748);
nand U5163 (N_5163,N_4870,N_4642);
or U5164 (N_5164,N_4553,N_4852);
nand U5165 (N_5165,N_4546,N_4631);
nor U5166 (N_5166,N_4838,N_4833);
xor U5167 (N_5167,N_4924,N_4664);
and U5168 (N_5168,N_4538,N_4735);
nand U5169 (N_5169,N_4754,N_4977);
nand U5170 (N_5170,N_4857,N_4859);
or U5171 (N_5171,N_4571,N_4771);
nor U5172 (N_5172,N_4647,N_4894);
and U5173 (N_5173,N_4505,N_4686);
nand U5174 (N_5174,N_4697,N_4962);
or U5175 (N_5175,N_4746,N_4839);
and U5176 (N_5176,N_4972,N_4747);
nor U5177 (N_5177,N_4737,N_4562);
nand U5178 (N_5178,N_4660,N_4669);
or U5179 (N_5179,N_4973,N_4552);
nor U5180 (N_5180,N_4881,N_4709);
nand U5181 (N_5181,N_4673,N_4517);
nand U5182 (N_5182,N_4598,N_4963);
nand U5183 (N_5183,N_4633,N_4832);
or U5184 (N_5184,N_4763,N_4701);
xnor U5185 (N_5185,N_4902,N_4536);
and U5186 (N_5186,N_4999,N_4513);
nor U5187 (N_5187,N_4965,N_4882);
xor U5188 (N_5188,N_4516,N_4877);
nand U5189 (N_5189,N_4706,N_4503);
xor U5190 (N_5190,N_4600,N_4586);
or U5191 (N_5191,N_4738,N_4533);
or U5192 (N_5192,N_4582,N_4711);
and U5193 (N_5193,N_4944,N_4780);
nor U5194 (N_5194,N_4779,N_4893);
and U5195 (N_5195,N_4502,N_4622);
nand U5196 (N_5196,N_4605,N_4707);
and U5197 (N_5197,N_4545,N_4675);
nand U5198 (N_5198,N_4584,N_4828);
and U5199 (N_5199,N_4560,N_4537);
nand U5200 (N_5200,N_4953,N_4555);
and U5201 (N_5201,N_4925,N_4695);
nand U5202 (N_5202,N_4556,N_4875);
and U5203 (N_5203,N_4658,N_4618);
nor U5204 (N_5204,N_4937,N_4785);
and U5205 (N_5205,N_4929,N_4550);
or U5206 (N_5206,N_4762,N_4519);
and U5207 (N_5207,N_4651,N_4723);
or U5208 (N_5208,N_4752,N_4989);
nand U5209 (N_5209,N_4687,N_4506);
nand U5210 (N_5210,N_4794,N_4876);
xor U5211 (N_5211,N_4835,N_4668);
or U5212 (N_5212,N_4980,N_4679);
xor U5213 (N_5213,N_4544,N_4907);
or U5214 (N_5214,N_4888,N_4531);
xor U5215 (N_5215,N_4718,N_4577);
nor U5216 (N_5216,N_4567,N_4719);
or U5217 (N_5217,N_4640,N_4523);
nor U5218 (N_5218,N_4935,N_4825);
and U5219 (N_5219,N_4670,N_4868);
xnor U5220 (N_5220,N_4791,N_4676);
or U5221 (N_5221,N_4755,N_4913);
and U5222 (N_5222,N_4847,N_4721);
nor U5223 (N_5223,N_4650,N_4563);
and U5224 (N_5224,N_4974,N_4604);
xnor U5225 (N_5225,N_4823,N_4947);
and U5226 (N_5226,N_4690,N_4918);
xor U5227 (N_5227,N_4904,N_4504);
or U5228 (N_5228,N_4671,N_4744);
nand U5229 (N_5229,N_4557,N_4940);
nand U5230 (N_5230,N_4608,N_4952);
and U5231 (N_5231,N_4949,N_4969);
or U5232 (N_5232,N_4568,N_4652);
and U5233 (N_5233,N_4636,N_4830);
and U5234 (N_5234,N_4518,N_4936);
nand U5235 (N_5235,N_4773,N_4788);
xor U5236 (N_5236,N_4911,N_4804);
nand U5237 (N_5237,N_4713,N_4588);
or U5238 (N_5238,N_4890,N_4966);
nor U5239 (N_5239,N_4638,N_4681);
nand U5240 (N_5240,N_4983,N_4858);
xor U5241 (N_5241,N_4958,N_4939);
nand U5242 (N_5242,N_4920,N_4732);
or U5243 (N_5243,N_4803,N_4667);
xnor U5244 (N_5244,N_4617,N_4595);
or U5245 (N_5245,N_4946,N_4530);
nand U5246 (N_5246,N_4985,N_4644);
and U5247 (N_5247,N_4677,N_4720);
nor U5248 (N_5248,N_4508,N_4759);
nand U5249 (N_5249,N_4993,N_4655);
nand U5250 (N_5250,N_4708,N_4599);
nand U5251 (N_5251,N_4707,N_4690);
or U5252 (N_5252,N_4928,N_4594);
nor U5253 (N_5253,N_4598,N_4697);
xor U5254 (N_5254,N_4801,N_4704);
or U5255 (N_5255,N_4756,N_4766);
and U5256 (N_5256,N_4690,N_4855);
or U5257 (N_5257,N_4703,N_4949);
xor U5258 (N_5258,N_4796,N_4770);
or U5259 (N_5259,N_4886,N_4587);
or U5260 (N_5260,N_4648,N_4986);
or U5261 (N_5261,N_4748,N_4679);
xor U5262 (N_5262,N_4593,N_4539);
nand U5263 (N_5263,N_4906,N_4782);
nor U5264 (N_5264,N_4737,N_4802);
xor U5265 (N_5265,N_4767,N_4570);
nor U5266 (N_5266,N_4621,N_4872);
and U5267 (N_5267,N_4834,N_4557);
nor U5268 (N_5268,N_4911,N_4638);
nand U5269 (N_5269,N_4616,N_4913);
nor U5270 (N_5270,N_4566,N_4927);
nor U5271 (N_5271,N_4836,N_4544);
or U5272 (N_5272,N_4535,N_4801);
nor U5273 (N_5273,N_4563,N_4583);
nand U5274 (N_5274,N_4587,N_4665);
nand U5275 (N_5275,N_4969,N_4611);
nand U5276 (N_5276,N_4520,N_4932);
nand U5277 (N_5277,N_4538,N_4646);
nand U5278 (N_5278,N_4994,N_4906);
xor U5279 (N_5279,N_4842,N_4777);
nand U5280 (N_5280,N_4692,N_4931);
and U5281 (N_5281,N_4939,N_4870);
or U5282 (N_5282,N_4579,N_4830);
or U5283 (N_5283,N_4524,N_4697);
and U5284 (N_5284,N_4836,N_4649);
nand U5285 (N_5285,N_4576,N_4634);
or U5286 (N_5286,N_4668,N_4691);
nor U5287 (N_5287,N_4950,N_4662);
nand U5288 (N_5288,N_4614,N_4698);
nand U5289 (N_5289,N_4692,N_4970);
and U5290 (N_5290,N_4568,N_4793);
nand U5291 (N_5291,N_4967,N_4779);
nor U5292 (N_5292,N_4627,N_4586);
and U5293 (N_5293,N_4548,N_4684);
or U5294 (N_5294,N_4880,N_4711);
nor U5295 (N_5295,N_4557,N_4563);
and U5296 (N_5296,N_4790,N_4634);
xnor U5297 (N_5297,N_4917,N_4683);
nor U5298 (N_5298,N_4756,N_4956);
or U5299 (N_5299,N_4931,N_4806);
nand U5300 (N_5300,N_4781,N_4605);
nor U5301 (N_5301,N_4508,N_4670);
and U5302 (N_5302,N_4726,N_4552);
nor U5303 (N_5303,N_4715,N_4736);
and U5304 (N_5304,N_4979,N_4567);
nor U5305 (N_5305,N_4711,N_4527);
and U5306 (N_5306,N_4786,N_4735);
xnor U5307 (N_5307,N_4724,N_4963);
nand U5308 (N_5308,N_4840,N_4858);
or U5309 (N_5309,N_4628,N_4507);
or U5310 (N_5310,N_4586,N_4801);
and U5311 (N_5311,N_4676,N_4764);
nor U5312 (N_5312,N_4782,N_4589);
or U5313 (N_5313,N_4874,N_4766);
nand U5314 (N_5314,N_4611,N_4960);
xnor U5315 (N_5315,N_4952,N_4684);
and U5316 (N_5316,N_4871,N_4640);
and U5317 (N_5317,N_4917,N_4738);
nor U5318 (N_5318,N_4747,N_4507);
or U5319 (N_5319,N_4825,N_4861);
xor U5320 (N_5320,N_4677,N_4843);
and U5321 (N_5321,N_4769,N_4831);
or U5322 (N_5322,N_4723,N_4926);
nor U5323 (N_5323,N_4853,N_4834);
nor U5324 (N_5324,N_4808,N_4526);
or U5325 (N_5325,N_4602,N_4807);
or U5326 (N_5326,N_4849,N_4897);
and U5327 (N_5327,N_4796,N_4810);
nor U5328 (N_5328,N_4604,N_4529);
nand U5329 (N_5329,N_4838,N_4700);
nand U5330 (N_5330,N_4565,N_4670);
or U5331 (N_5331,N_4660,N_4666);
nor U5332 (N_5332,N_4728,N_4714);
nor U5333 (N_5333,N_4923,N_4700);
or U5334 (N_5334,N_4790,N_4555);
or U5335 (N_5335,N_4586,N_4712);
and U5336 (N_5336,N_4869,N_4883);
or U5337 (N_5337,N_4798,N_4893);
or U5338 (N_5338,N_4766,N_4585);
xor U5339 (N_5339,N_4708,N_4739);
and U5340 (N_5340,N_4558,N_4751);
nor U5341 (N_5341,N_4541,N_4887);
xor U5342 (N_5342,N_4811,N_4977);
and U5343 (N_5343,N_4722,N_4920);
nand U5344 (N_5344,N_4699,N_4758);
nor U5345 (N_5345,N_4931,N_4855);
nand U5346 (N_5346,N_4932,N_4610);
and U5347 (N_5347,N_4894,N_4677);
and U5348 (N_5348,N_4603,N_4695);
or U5349 (N_5349,N_4768,N_4995);
and U5350 (N_5350,N_4761,N_4790);
nand U5351 (N_5351,N_4853,N_4540);
nand U5352 (N_5352,N_4941,N_4617);
or U5353 (N_5353,N_4887,N_4972);
nor U5354 (N_5354,N_4772,N_4591);
nand U5355 (N_5355,N_4523,N_4871);
nor U5356 (N_5356,N_4603,N_4842);
xnor U5357 (N_5357,N_4534,N_4598);
and U5358 (N_5358,N_4614,N_4833);
and U5359 (N_5359,N_4516,N_4638);
or U5360 (N_5360,N_4903,N_4851);
or U5361 (N_5361,N_4781,N_4506);
or U5362 (N_5362,N_4619,N_4779);
xnor U5363 (N_5363,N_4932,N_4716);
xnor U5364 (N_5364,N_4704,N_4979);
nor U5365 (N_5365,N_4931,N_4767);
xor U5366 (N_5366,N_4662,N_4722);
or U5367 (N_5367,N_4550,N_4851);
and U5368 (N_5368,N_4509,N_4663);
nor U5369 (N_5369,N_4705,N_4548);
or U5370 (N_5370,N_4531,N_4647);
nand U5371 (N_5371,N_4978,N_4500);
nor U5372 (N_5372,N_4756,N_4989);
nor U5373 (N_5373,N_4927,N_4583);
and U5374 (N_5374,N_4757,N_4877);
nor U5375 (N_5375,N_4851,N_4845);
nand U5376 (N_5376,N_4828,N_4602);
or U5377 (N_5377,N_4620,N_4851);
or U5378 (N_5378,N_4767,N_4956);
or U5379 (N_5379,N_4902,N_4561);
or U5380 (N_5380,N_4986,N_4643);
nand U5381 (N_5381,N_4937,N_4885);
nand U5382 (N_5382,N_4585,N_4926);
nand U5383 (N_5383,N_4745,N_4922);
xor U5384 (N_5384,N_4873,N_4563);
nor U5385 (N_5385,N_4578,N_4660);
or U5386 (N_5386,N_4891,N_4557);
and U5387 (N_5387,N_4624,N_4756);
nand U5388 (N_5388,N_4633,N_4669);
nor U5389 (N_5389,N_4960,N_4776);
nand U5390 (N_5390,N_4898,N_4529);
nand U5391 (N_5391,N_4526,N_4993);
xnor U5392 (N_5392,N_4863,N_4698);
and U5393 (N_5393,N_4937,N_4577);
nand U5394 (N_5394,N_4506,N_4841);
and U5395 (N_5395,N_4822,N_4674);
xor U5396 (N_5396,N_4737,N_4805);
and U5397 (N_5397,N_4931,N_4780);
and U5398 (N_5398,N_4718,N_4836);
nor U5399 (N_5399,N_4535,N_4536);
xor U5400 (N_5400,N_4685,N_4861);
nand U5401 (N_5401,N_4559,N_4603);
nor U5402 (N_5402,N_4689,N_4567);
nand U5403 (N_5403,N_4968,N_4887);
and U5404 (N_5404,N_4957,N_4551);
nand U5405 (N_5405,N_4886,N_4849);
and U5406 (N_5406,N_4540,N_4822);
nand U5407 (N_5407,N_4854,N_4836);
and U5408 (N_5408,N_4597,N_4839);
nand U5409 (N_5409,N_4626,N_4656);
or U5410 (N_5410,N_4712,N_4637);
and U5411 (N_5411,N_4549,N_4992);
or U5412 (N_5412,N_4704,N_4838);
xnor U5413 (N_5413,N_4605,N_4586);
nand U5414 (N_5414,N_4806,N_4602);
nor U5415 (N_5415,N_4671,N_4523);
nor U5416 (N_5416,N_4858,N_4853);
nand U5417 (N_5417,N_4605,N_4802);
nor U5418 (N_5418,N_4663,N_4949);
nand U5419 (N_5419,N_4748,N_4960);
nand U5420 (N_5420,N_4824,N_4706);
nor U5421 (N_5421,N_4618,N_4570);
or U5422 (N_5422,N_4666,N_4973);
and U5423 (N_5423,N_4684,N_4580);
xor U5424 (N_5424,N_4835,N_4640);
and U5425 (N_5425,N_4787,N_4938);
nand U5426 (N_5426,N_4542,N_4756);
nand U5427 (N_5427,N_4914,N_4720);
or U5428 (N_5428,N_4581,N_4708);
nor U5429 (N_5429,N_4795,N_4558);
or U5430 (N_5430,N_4998,N_4576);
nand U5431 (N_5431,N_4612,N_4797);
nand U5432 (N_5432,N_4653,N_4960);
and U5433 (N_5433,N_4547,N_4628);
or U5434 (N_5434,N_4938,N_4891);
nor U5435 (N_5435,N_4544,N_4809);
or U5436 (N_5436,N_4926,N_4749);
nand U5437 (N_5437,N_4839,N_4667);
nand U5438 (N_5438,N_4912,N_4683);
nand U5439 (N_5439,N_4696,N_4733);
nor U5440 (N_5440,N_4579,N_4687);
xnor U5441 (N_5441,N_4919,N_4930);
nand U5442 (N_5442,N_4854,N_4686);
and U5443 (N_5443,N_4868,N_4930);
nor U5444 (N_5444,N_4501,N_4855);
or U5445 (N_5445,N_4884,N_4683);
nor U5446 (N_5446,N_4748,N_4894);
nor U5447 (N_5447,N_4704,N_4985);
xnor U5448 (N_5448,N_4850,N_4776);
nand U5449 (N_5449,N_4754,N_4641);
nor U5450 (N_5450,N_4606,N_4551);
xnor U5451 (N_5451,N_4743,N_4912);
xor U5452 (N_5452,N_4712,N_4980);
nor U5453 (N_5453,N_4651,N_4986);
nor U5454 (N_5454,N_4518,N_4657);
and U5455 (N_5455,N_4638,N_4566);
and U5456 (N_5456,N_4699,N_4744);
nor U5457 (N_5457,N_4594,N_4744);
and U5458 (N_5458,N_4731,N_4923);
or U5459 (N_5459,N_4681,N_4752);
nor U5460 (N_5460,N_4982,N_4927);
nand U5461 (N_5461,N_4577,N_4693);
nand U5462 (N_5462,N_4800,N_4996);
or U5463 (N_5463,N_4692,N_4890);
nand U5464 (N_5464,N_4826,N_4870);
xor U5465 (N_5465,N_4813,N_4672);
or U5466 (N_5466,N_4546,N_4842);
or U5467 (N_5467,N_4721,N_4517);
nor U5468 (N_5468,N_4521,N_4818);
nor U5469 (N_5469,N_4579,N_4714);
or U5470 (N_5470,N_4571,N_4615);
and U5471 (N_5471,N_4853,N_4992);
or U5472 (N_5472,N_4963,N_4642);
nand U5473 (N_5473,N_4739,N_4596);
xor U5474 (N_5474,N_4807,N_4647);
or U5475 (N_5475,N_4561,N_4567);
nor U5476 (N_5476,N_4617,N_4613);
or U5477 (N_5477,N_4966,N_4797);
xnor U5478 (N_5478,N_4659,N_4650);
or U5479 (N_5479,N_4988,N_4992);
nand U5480 (N_5480,N_4725,N_4988);
or U5481 (N_5481,N_4804,N_4573);
nand U5482 (N_5482,N_4768,N_4806);
xnor U5483 (N_5483,N_4626,N_4794);
nor U5484 (N_5484,N_4590,N_4939);
and U5485 (N_5485,N_4607,N_4531);
or U5486 (N_5486,N_4798,N_4636);
nand U5487 (N_5487,N_4769,N_4906);
nand U5488 (N_5488,N_4563,N_4966);
xnor U5489 (N_5489,N_4906,N_4718);
and U5490 (N_5490,N_4731,N_4832);
or U5491 (N_5491,N_4978,N_4829);
or U5492 (N_5492,N_4510,N_4546);
nor U5493 (N_5493,N_4569,N_4522);
and U5494 (N_5494,N_4869,N_4800);
nor U5495 (N_5495,N_4525,N_4906);
and U5496 (N_5496,N_4905,N_4638);
nand U5497 (N_5497,N_4950,N_4508);
and U5498 (N_5498,N_4863,N_4665);
or U5499 (N_5499,N_4813,N_4833);
nor U5500 (N_5500,N_5113,N_5396);
or U5501 (N_5501,N_5102,N_5017);
nand U5502 (N_5502,N_5150,N_5246);
nor U5503 (N_5503,N_5047,N_5477);
nor U5504 (N_5504,N_5373,N_5060);
nand U5505 (N_5505,N_5189,N_5272);
and U5506 (N_5506,N_5316,N_5206);
and U5507 (N_5507,N_5357,N_5331);
and U5508 (N_5508,N_5273,N_5442);
and U5509 (N_5509,N_5302,N_5268);
nor U5510 (N_5510,N_5185,N_5480);
nand U5511 (N_5511,N_5235,N_5204);
nand U5512 (N_5512,N_5391,N_5203);
nand U5513 (N_5513,N_5300,N_5455);
nand U5514 (N_5514,N_5147,N_5319);
and U5515 (N_5515,N_5158,N_5079);
nand U5516 (N_5516,N_5106,N_5036);
nand U5517 (N_5517,N_5080,N_5146);
or U5518 (N_5518,N_5436,N_5467);
and U5519 (N_5519,N_5062,N_5001);
or U5520 (N_5520,N_5037,N_5205);
nand U5521 (N_5521,N_5303,N_5194);
nand U5522 (N_5522,N_5159,N_5252);
nor U5523 (N_5523,N_5026,N_5210);
and U5524 (N_5524,N_5100,N_5489);
nand U5525 (N_5525,N_5438,N_5264);
nor U5526 (N_5526,N_5231,N_5177);
and U5527 (N_5527,N_5108,N_5021);
nand U5528 (N_5528,N_5307,N_5253);
xnor U5529 (N_5529,N_5462,N_5071);
nor U5530 (N_5530,N_5109,N_5151);
nand U5531 (N_5531,N_5383,N_5228);
xor U5532 (N_5532,N_5408,N_5077);
or U5533 (N_5533,N_5173,N_5139);
nand U5534 (N_5534,N_5003,N_5294);
or U5535 (N_5535,N_5039,N_5207);
nand U5536 (N_5536,N_5019,N_5333);
nor U5537 (N_5537,N_5095,N_5117);
and U5538 (N_5538,N_5061,N_5058);
nor U5539 (N_5539,N_5221,N_5445);
and U5540 (N_5540,N_5220,N_5188);
or U5541 (N_5541,N_5486,N_5362);
or U5542 (N_5542,N_5367,N_5082);
nand U5543 (N_5543,N_5352,N_5224);
nor U5544 (N_5544,N_5353,N_5441);
nand U5545 (N_5545,N_5305,N_5422);
nand U5546 (N_5546,N_5327,N_5284);
and U5547 (N_5547,N_5468,N_5306);
nand U5548 (N_5548,N_5007,N_5174);
nor U5549 (N_5549,N_5238,N_5363);
xnor U5550 (N_5550,N_5010,N_5359);
and U5551 (N_5551,N_5072,N_5286);
and U5552 (N_5552,N_5122,N_5129);
nand U5553 (N_5553,N_5440,N_5290);
and U5554 (N_5554,N_5370,N_5354);
and U5555 (N_5555,N_5218,N_5481);
nor U5556 (N_5556,N_5141,N_5490);
and U5557 (N_5557,N_5499,N_5075);
nor U5558 (N_5558,N_5463,N_5176);
nand U5559 (N_5559,N_5089,N_5378);
nor U5560 (N_5560,N_5012,N_5155);
nor U5561 (N_5561,N_5073,N_5393);
and U5562 (N_5562,N_5308,N_5078);
nor U5563 (N_5563,N_5092,N_5435);
or U5564 (N_5564,N_5488,N_5278);
nand U5565 (N_5565,N_5227,N_5245);
nand U5566 (N_5566,N_5450,N_5121);
nand U5567 (N_5567,N_5143,N_5156);
nor U5568 (N_5568,N_5426,N_5215);
nand U5569 (N_5569,N_5195,N_5293);
nand U5570 (N_5570,N_5279,N_5377);
and U5571 (N_5571,N_5397,N_5417);
nand U5572 (N_5572,N_5454,N_5386);
or U5573 (N_5573,N_5269,N_5291);
or U5574 (N_5574,N_5076,N_5222);
or U5575 (N_5575,N_5097,N_5361);
nand U5576 (N_5576,N_5444,N_5223);
xor U5577 (N_5577,N_5289,N_5356);
nand U5578 (N_5578,N_5285,N_5029);
nor U5579 (N_5579,N_5309,N_5042);
and U5580 (N_5580,N_5119,N_5365);
nor U5581 (N_5581,N_5270,N_5255);
xnor U5582 (N_5582,N_5250,N_5416);
and U5583 (N_5583,N_5111,N_5484);
and U5584 (N_5584,N_5498,N_5107);
nor U5585 (N_5585,N_5430,N_5038);
nor U5586 (N_5586,N_5199,N_5474);
nand U5587 (N_5587,N_5027,N_5494);
nor U5588 (N_5588,N_5427,N_5398);
or U5589 (N_5589,N_5483,N_5461);
nor U5590 (N_5590,N_5138,N_5413);
or U5591 (N_5591,N_5243,N_5153);
and U5592 (N_5592,N_5265,N_5201);
or U5593 (N_5593,N_5094,N_5035);
or U5594 (N_5594,N_5380,N_5162);
nor U5595 (N_5595,N_5142,N_5382);
nor U5596 (N_5596,N_5219,N_5496);
nand U5597 (N_5597,N_5288,N_5181);
or U5598 (N_5598,N_5394,N_5161);
nand U5599 (N_5599,N_5103,N_5345);
or U5600 (N_5600,N_5297,N_5315);
xor U5601 (N_5601,N_5475,N_5387);
xor U5602 (N_5602,N_5453,N_5091);
nor U5603 (N_5603,N_5028,N_5433);
xor U5604 (N_5604,N_5419,N_5310);
and U5605 (N_5605,N_5464,N_5392);
nor U5606 (N_5606,N_5301,N_5013);
nor U5607 (N_5607,N_5005,N_5263);
nand U5608 (N_5608,N_5325,N_5170);
nor U5609 (N_5609,N_5041,N_5184);
or U5610 (N_5610,N_5020,N_5443);
or U5611 (N_5611,N_5131,N_5083);
or U5612 (N_5612,N_5348,N_5134);
or U5613 (N_5613,N_5266,N_5217);
or U5614 (N_5614,N_5198,N_5186);
nand U5615 (N_5615,N_5154,N_5414);
nor U5616 (N_5616,N_5262,N_5030);
or U5617 (N_5617,N_5163,N_5469);
nor U5618 (N_5618,N_5145,N_5298);
nand U5619 (N_5619,N_5208,N_5130);
nand U5620 (N_5620,N_5209,N_5407);
nand U5621 (N_5621,N_5355,N_5456);
and U5622 (N_5622,N_5418,N_5261);
or U5623 (N_5623,N_5420,N_5105);
nand U5624 (N_5624,N_5381,N_5025);
nand U5625 (N_5625,N_5011,N_5063);
xor U5626 (N_5626,N_5379,N_5335);
nand U5627 (N_5627,N_5428,N_5226);
or U5628 (N_5628,N_5135,N_5330);
nand U5629 (N_5629,N_5312,N_5487);
nor U5630 (N_5630,N_5406,N_5295);
or U5631 (N_5631,N_5339,N_5049);
and U5632 (N_5632,N_5110,N_5347);
nand U5633 (N_5633,N_5329,N_5104);
nand U5634 (N_5634,N_5304,N_5179);
or U5635 (N_5635,N_5299,N_5178);
and U5636 (N_5636,N_5409,N_5167);
and U5637 (N_5637,N_5459,N_5234);
xor U5638 (N_5638,N_5470,N_5127);
and U5639 (N_5639,N_5086,N_5016);
or U5640 (N_5640,N_5180,N_5314);
and U5641 (N_5641,N_5410,N_5317);
xor U5642 (N_5642,N_5473,N_5472);
and U5643 (N_5643,N_5341,N_5343);
nor U5644 (N_5644,N_5040,N_5115);
or U5645 (N_5645,N_5225,N_5344);
nor U5646 (N_5646,N_5258,N_5249);
nand U5647 (N_5647,N_5485,N_5326);
or U5648 (N_5648,N_5283,N_5057);
nand U5649 (N_5649,N_5251,N_5175);
xnor U5650 (N_5650,N_5338,N_5059);
nand U5651 (N_5651,N_5006,N_5112);
and U5652 (N_5652,N_5402,N_5123);
xor U5653 (N_5653,N_5048,N_5101);
nor U5654 (N_5654,N_5451,N_5066);
nand U5655 (N_5655,N_5014,N_5081);
or U5656 (N_5656,N_5050,N_5247);
and U5657 (N_5657,N_5087,N_5191);
nor U5658 (N_5658,N_5320,N_5133);
nor U5659 (N_5659,N_5004,N_5033);
nand U5660 (N_5660,N_5390,N_5334);
and U5661 (N_5661,N_5476,N_5403);
or U5662 (N_5662,N_5324,N_5183);
nor U5663 (N_5663,N_5099,N_5271);
xnor U5664 (N_5664,N_5360,N_5052);
or U5665 (N_5665,N_5148,N_5169);
and U5666 (N_5666,N_5212,N_5412);
or U5667 (N_5667,N_5478,N_5248);
and U5668 (N_5668,N_5065,N_5034);
nor U5669 (N_5669,N_5349,N_5157);
nand U5670 (N_5670,N_5068,N_5144);
nand U5671 (N_5671,N_5482,N_5351);
xnor U5672 (N_5672,N_5172,N_5200);
nand U5673 (N_5673,N_5492,N_5152);
nor U5674 (N_5674,N_5374,N_5260);
xnor U5675 (N_5675,N_5008,N_5281);
nand U5676 (N_5676,N_5193,N_5311);
nand U5677 (N_5677,N_5276,N_5192);
nor U5678 (N_5678,N_5056,N_5375);
or U5679 (N_5679,N_5090,N_5015);
and U5680 (N_5680,N_5332,N_5166);
and U5681 (N_5681,N_5321,N_5256);
nor U5682 (N_5682,N_5031,N_5211);
and U5683 (N_5683,N_5069,N_5275);
nor U5684 (N_5684,N_5364,N_5282);
and U5685 (N_5685,N_5448,N_5216);
nand U5686 (N_5686,N_5471,N_5244);
nor U5687 (N_5687,N_5126,N_5096);
nand U5688 (N_5688,N_5128,N_5053);
xor U5689 (N_5689,N_5239,N_5267);
nor U5690 (N_5690,N_5160,N_5322);
nand U5691 (N_5691,N_5368,N_5371);
or U5692 (N_5692,N_5495,N_5366);
and U5693 (N_5693,N_5214,N_5399);
xor U5694 (N_5694,N_5024,N_5350);
or U5695 (N_5695,N_5296,N_5241);
and U5696 (N_5696,N_5044,N_5164);
and U5697 (N_5697,N_5369,N_5337);
xnor U5698 (N_5698,N_5457,N_5116);
or U5699 (N_5699,N_5280,N_5385);
nor U5700 (N_5700,N_5340,N_5196);
nand U5701 (N_5701,N_5423,N_5400);
nand U5702 (N_5702,N_5318,N_5232);
nor U5703 (N_5703,N_5055,N_5452);
and U5704 (N_5704,N_5067,N_5018);
and U5705 (N_5705,N_5197,N_5054);
nand U5706 (N_5706,N_5460,N_5032);
and U5707 (N_5707,N_5389,N_5046);
or U5708 (N_5708,N_5132,N_5045);
or U5709 (N_5709,N_5165,N_5292);
nand U5710 (N_5710,N_5240,N_5358);
xor U5711 (N_5711,N_5439,N_5051);
nor U5712 (N_5712,N_5257,N_5388);
or U5713 (N_5713,N_5136,N_5230);
nand U5714 (N_5714,N_5085,N_5213);
or U5715 (N_5715,N_5202,N_5395);
and U5716 (N_5716,N_5254,N_5168);
nand U5717 (N_5717,N_5446,N_5434);
nand U5718 (N_5718,N_5415,N_5404);
and U5719 (N_5719,N_5229,N_5120);
or U5720 (N_5720,N_5064,N_5466);
or U5721 (N_5721,N_5497,N_5182);
nor U5722 (N_5722,N_5491,N_5432);
nor U5723 (N_5723,N_5043,N_5421);
and U5724 (N_5724,N_5447,N_5287);
nand U5725 (N_5725,N_5259,N_5323);
or U5726 (N_5726,N_5088,N_5171);
nor U5727 (N_5727,N_5405,N_5242);
nor U5728 (N_5728,N_5124,N_5233);
or U5729 (N_5729,N_5098,N_5401);
nor U5730 (N_5730,N_5424,N_5342);
and U5731 (N_5731,N_5236,N_5000);
xor U5732 (N_5732,N_5190,N_5237);
nand U5733 (N_5733,N_5277,N_5140);
nand U5734 (N_5734,N_5137,N_5479);
and U5735 (N_5735,N_5084,N_5009);
or U5736 (N_5736,N_5313,N_5429);
nor U5737 (N_5737,N_5437,N_5411);
and U5738 (N_5738,N_5431,N_5425);
nor U5739 (N_5739,N_5274,N_5002);
nor U5740 (N_5740,N_5118,N_5384);
or U5741 (N_5741,N_5114,N_5376);
xor U5742 (N_5742,N_5336,N_5328);
nand U5743 (N_5743,N_5187,N_5465);
and U5744 (N_5744,N_5074,N_5093);
nand U5745 (N_5745,N_5372,N_5023);
or U5746 (N_5746,N_5070,N_5458);
or U5747 (N_5747,N_5493,N_5125);
and U5748 (N_5748,N_5149,N_5022);
nor U5749 (N_5749,N_5346,N_5449);
nand U5750 (N_5750,N_5291,N_5188);
nor U5751 (N_5751,N_5079,N_5128);
nor U5752 (N_5752,N_5278,N_5398);
nand U5753 (N_5753,N_5497,N_5468);
xnor U5754 (N_5754,N_5121,N_5362);
or U5755 (N_5755,N_5310,N_5411);
nand U5756 (N_5756,N_5191,N_5231);
and U5757 (N_5757,N_5386,N_5446);
xnor U5758 (N_5758,N_5424,N_5402);
or U5759 (N_5759,N_5476,N_5020);
nor U5760 (N_5760,N_5485,N_5172);
nand U5761 (N_5761,N_5279,N_5327);
or U5762 (N_5762,N_5070,N_5447);
nand U5763 (N_5763,N_5446,N_5075);
or U5764 (N_5764,N_5401,N_5034);
and U5765 (N_5765,N_5122,N_5486);
and U5766 (N_5766,N_5098,N_5226);
nand U5767 (N_5767,N_5204,N_5272);
nor U5768 (N_5768,N_5328,N_5446);
nor U5769 (N_5769,N_5308,N_5454);
nor U5770 (N_5770,N_5110,N_5330);
or U5771 (N_5771,N_5337,N_5380);
nand U5772 (N_5772,N_5387,N_5487);
or U5773 (N_5773,N_5259,N_5397);
and U5774 (N_5774,N_5023,N_5190);
and U5775 (N_5775,N_5118,N_5494);
nand U5776 (N_5776,N_5396,N_5417);
or U5777 (N_5777,N_5311,N_5320);
nand U5778 (N_5778,N_5189,N_5034);
and U5779 (N_5779,N_5320,N_5273);
or U5780 (N_5780,N_5351,N_5432);
nor U5781 (N_5781,N_5127,N_5003);
nor U5782 (N_5782,N_5206,N_5411);
or U5783 (N_5783,N_5376,N_5435);
xnor U5784 (N_5784,N_5154,N_5455);
nor U5785 (N_5785,N_5170,N_5098);
or U5786 (N_5786,N_5007,N_5496);
and U5787 (N_5787,N_5069,N_5182);
nand U5788 (N_5788,N_5119,N_5490);
nand U5789 (N_5789,N_5299,N_5129);
nand U5790 (N_5790,N_5030,N_5287);
nand U5791 (N_5791,N_5074,N_5328);
nor U5792 (N_5792,N_5487,N_5441);
or U5793 (N_5793,N_5332,N_5050);
or U5794 (N_5794,N_5108,N_5346);
and U5795 (N_5795,N_5099,N_5132);
nand U5796 (N_5796,N_5316,N_5262);
or U5797 (N_5797,N_5413,N_5453);
or U5798 (N_5798,N_5287,N_5162);
nand U5799 (N_5799,N_5234,N_5126);
nand U5800 (N_5800,N_5190,N_5241);
nor U5801 (N_5801,N_5083,N_5154);
or U5802 (N_5802,N_5062,N_5049);
or U5803 (N_5803,N_5262,N_5474);
nor U5804 (N_5804,N_5245,N_5294);
nand U5805 (N_5805,N_5499,N_5447);
or U5806 (N_5806,N_5301,N_5201);
nor U5807 (N_5807,N_5320,N_5376);
nor U5808 (N_5808,N_5354,N_5114);
or U5809 (N_5809,N_5342,N_5068);
nand U5810 (N_5810,N_5411,N_5114);
or U5811 (N_5811,N_5069,N_5304);
nor U5812 (N_5812,N_5413,N_5458);
or U5813 (N_5813,N_5277,N_5349);
or U5814 (N_5814,N_5059,N_5479);
nor U5815 (N_5815,N_5243,N_5028);
nand U5816 (N_5816,N_5231,N_5433);
nand U5817 (N_5817,N_5476,N_5374);
nor U5818 (N_5818,N_5331,N_5093);
nor U5819 (N_5819,N_5200,N_5335);
or U5820 (N_5820,N_5001,N_5363);
or U5821 (N_5821,N_5101,N_5438);
nand U5822 (N_5822,N_5145,N_5261);
or U5823 (N_5823,N_5351,N_5069);
and U5824 (N_5824,N_5432,N_5264);
and U5825 (N_5825,N_5185,N_5390);
and U5826 (N_5826,N_5279,N_5023);
xnor U5827 (N_5827,N_5439,N_5101);
and U5828 (N_5828,N_5209,N_5106);
nand U5829 (N_5829,N_5227,N_5287);
nand U5830 (N_5830,N_5177,N_5141);
xnor U5831 (N_5831,N_5167,N_5359);
xnor U5832 (N_5832,N_5114,N_5283);
or U5833 (N_5833,N_5086,N_5161);
nor U5834 (N_5834,N_5391,N_5149);
nor U5835 (N_5835,N_5122,N_5473);
nor U5836 (N_5836,N_5199,N_5088);
nor U5837 (N_5837,N_5407,N_5127);
nand U5838 (N_5838,N_5150,N_5232);
and U5839 (N_5839,N_5366,N_5124);
or U5840 (N_5840,N_5070,N_5332);
nor U5841 (N_5841,N_5146,N_5179);
or U5842 (N_5842,N_5188,N_5021);
nand U5843 (N_5843,N_5037,N_5478);
and U5844 (N_5844,N_5342,N_5372);
or U5845 (N_5845,N_5021,N_5178);
nand U5846 (N_5846,N_5312,N_5253);
and U5847 (N_5847,N_5317,N_5173);
and U5848 (N_5848,N_5358,N_5029);
or U5849 (N_5849,N_5049,N_5259);
nor U5850 (N_5850,N_5457,N_5058);
nor U5851 (N_5851,N_5032,N_5479);
nand U5852 (N_5852,N_5480,N_5343);
nand U5853 (N_5853,N_5162,N_5374);
and U5854 (N_5854,N_5355,N_5037);
nor U5855 (N_5855,N_5423,N_5436);
and U5856 (N_5856,N_5358,N_5156);
nor U5857 (N_5857,N_5458,N_5304);
xor U5858 (N_5858,N_5064,N_5191);
xor U5859 (N_5859,N_5134,N_5030);
xor U5860 (N_5860,N_5309,N_5279);
or U5861 (N_5861,N_5297,N_5314);
or U5862 (N_5862,N_5213,N_5495);
nand U5863 (N_5863,N_5456,N_5176);
and U5864 (N_5864,N_5085,N_5108);
nand U5865 (N_5865,N_5272,N_5443);
or U5866 (N_5866,N_5425,N_5037);
or U5867 (N_5867,N_5216,N_5100);
nand U5868 (N_5868,N_5085,N_5178);
and U5869 (N_5869,N_5166,N_5252);
and U5870 (N_5870,N_5002,N_5196);
nand U5871 (N_5871,N_5355,N_5349);
nand U5872 (N_5872,N_5132,N_5194);
xnor U5873 (N_5873,N_5258,N_5016);
or U5874 (N_5874,N_5156,N_5385);
nand U5875 (N_5875,N_5313,N_5448);
and U5876 (N_5876,N_5419,N_5255);
xor U5877 (N_5877,N_5408,N_5264);
nor U5878 (N_5878,N_5346,N_5414);
and U5879 (N_5879,N_5139,N_5230);
nand U5880 (N_5880,N_5120,N_5485);
or U5881 (N_5881,N_5328,N_5269);
nor U5882 (N_5882,N_5293,N_5424);
nor U5883 (N_5883,N_5392,N_5287);
and U5884 (N_5884,N_5002,N_5197);
xor U5885 (N_5885,N_5234,N_5200);
nor U5886 (N_5886,N_5178,N_5262);
nor U5887 (N_5887,N_5354,N_5364);
or U5888 (N_5888,N_5328,N_5118);
nand U5889 (N_5889,N_5256,N_5175);
nor U5890 (N_5890,N_5043,N_5006);
and U5891 (N_5891,N_5089,N_5009);
nand U5892 (N_5892,N_5387,N_5287);
and U5893 (N_5893,N_5375,N_5285);
nor U5894 (N_5894,N_5481,N_5056);
and U5895 (N_5895,N_5137,N_5076);
xor U5896 (N_5896,N_5258,N_5452);
nor U5897 (N_5897,N_5205,N_5039);
and U5898 (N_5898,N_5224,N_5137);
nor U5899 (N_5899,N_5142,N_5179);
and U5900 (N_5900,N_5222,N_5145);
or U5901 (N_5901,N_5221,N_5147);
nand U5902 (N_5902,N_5195,N_5411);
and U5903 (N_5903,N_5318,N_5368);
nand U5904 (N_5904,N_5094,N_5058);
nand U5905 (N_5905,N_5186,N_5130);
nand U5906 (N_5906,N_5292,N_5258);
nor U5907 (N_5907,N_5356,N_5455);
xnor U5908 (N_5908,N_5386,N_5228);
nand U5909 (N_5909,N_5287,N_5420);
nor U5910 (N_5910,N_5264,N_5342);
and U5911 (N_5911,N_5179,N_5150);
or U5912 (N_5912,N_5263,N_5278);
or U5913 (N_5913,N_5494,N_5171);
nand U5914 (N_5914,N_5292,N_5231);
or U5915 (N_5915,N_5378,N_5498);
xor U5916 (N_5916,N_5376,N_5036);
nand U5917 (N_5917,N_5338,N_5182);
or U5918 (N_5918,N_5162,N_5171);
nand U5919 (N_5919,N_5107,N_5325);
and U5920 (N_5920,N_5241,N_5311);
and U5921 (N_5921,N_5082,N_5127);
and U5922 (N_5922,N_5312,N_5034);
nor U5923 (N_5923,N_5107,N_5088);
and U5924 (N_5924,N_5255,N_5116);
nand U5925 (N_5925,N_5475,N_5332);
nor U5926 (N_5926,N_5315,N_5425);
and U5927 (N_5927,N_5303,N_5288);
nand U5928 (N_5928,N_5111,N_5396);
and U5929 (N_5929,N_5284,N_5497);
xor U5930 (N_5930,N_5129,N_5118);
or U5931 (N_5931,N_5353,N_5240);
nor U5932 (N_5932,N_5072,N_5192);
nand U5933 (N_5933,N_5354,N_5162);
or U5934 (N_5934,N_5343,N_5302);
or U5935 (N_5935,N_5304,N_5077);
nand U5936 (N_5936,N_5423,N_5147);
nand U5937 (N_5937,N_5144,N_5069);
nand U5938 (N_5938,N_5040,N_5349);
or U5939 (N_5939,N_5470,N_5303);
or U5940 (N_5940,N_5495,N_5055);
and U5941 (N_5941,N_5244,N_5497);
nand U5942 (N_5942,N_5344,N_5008);
or U5943 (N_5943,N_5221,N_5462);
nor U5944 (N_5944,N_5248,N_5042);
nor U5945 (N_5945,N_5172,N_5183);
or U5946 (N_5946,N_5346,N_5441);
nand U5947 (N_5947,N_5277,N_5402);
nand U5948 (N_5948,N_5352,N_5036);
or U5949 (N_5949,N_5087,N_5486);
nand U5950 (N_5950,N_5265,N_5175);
xor U5951 (N_5951,N_5058,N_5085);
xor U5952 (N_5952,N_5047,N_5288);
and U5953 (N_5953,N_5110,N_5054);
nor U5954 (N_5954,N_5476,N_5155);
and U5955 (N_5955,N_5466,N_5431);
nand U5956 (N_5956,N_5482,N_5431);
and U5957 (N_5957,N_5095,N_5409);
or U5958 (N_5958,N_5066,N_5275);
or U5959 (N_5959,N_5378,N_5067);
nor U5960 (N_5960,N_5180,N_5395);
nor U5961 (N_5961,N_5130,N_5122);
nand U5962 (N_5962,N_5284,N_5176);
nor U5963 (N_5963,N_5477,N_5053);
and U5964 (N_5964,N_5103,N_5109);
nand U5965 (N_5965,N_5424,N_5305);
nor U5966 (N_5966,N_5243,N_5116);
or U5967 (N_5967,N_5376,N_5079);
nor U5968 (N_5968,N_5227,N_5005);
nand U5969 (N_5969,N_5337,N_5007);
and U5970 (N_5970,N_5068,N_5313);
nand U5971 (N_5971,N_5457,N_5234);
nand U5972 (N_5972,N_5444,N_5499);
xnor U5973 (N_5973,N_5165,N_5334);
and U5974 (N_5974,N_5091,N_5270);
nor U5975 (N_5975,N_5088,N_5308);
nor U5976 (N_5976,N_5375,N_5119);
nand U5977 (N_5977,N_5135,N_5393);
nand U5978 (N_5978,N_5203,N_5262);
nor U5979 (N_5979,N_5392,N_5333);
nand U5980 (N_5980,N_5094,N_5297);
or U5981 (N_5981,N_5352,N_5391);
nor U5982 (N_5982,N_5230,N_5337);
nor U5983 (N_5983,N_5013,N_5136);
nand U5984 (N_5984,N_5086,N_5499);
and U5985 (N_5985,N_5282,N_5187);
and U5986 (N_5986,N_5407,N_5220);
and U5987 (N_5987,N_5406,N_5388);
or U5988 (N_5988,N_5141,N_5409);
and U5989 (N_5989,N_5400,N_5011);
nand U5990 (N_5990,N_5367,N_5029);
and U5991 (N_5991,N_5159,N_5314);
xor U5992 (N_5992,N_5285,N_5371);
nor U5993 (N_5993,N_5471,N_5071);
or U5994 (N_5994,N_5342,N_5044);
nor U5995 (N_5995,N_5219,N_5494);
and U5996 (N_5996,N_5197,N_5233);
xor U5997 (N_5997,N_5058,N_5081);
nor U5998 (N_5998,N_5166,N_5304);
nand U5999 (N_5999,N_5153,N_5247);
and U6000 (N_6000,N_5932,N_5754);
xor U6001 (N_6001,N_5680,N_5855);
nand U6002 (N_6002,N_5878,N_5779);
and U6003 (N_6003,N_5781,N_5573);
or U6004 (N_6004,N_5609,N_5674);
or U6005 (N_6005,N_5615,N_5876);
and U6006 (N_6006,N_5873,N_5831);
and U6007 (N_6007,N_5999,N_5505);
and U6008 (N_6008,N_5975,N_5552);
or U6009 (N_6009,N_5849,N_5942);
nand U6010 (N_6010,N_5550,N_5738);
nor U6011 (N_6011,N_5933,N_5830);
nand U6012 (N_6012,N_5623,N_5811);
nand U6013 (N_6013,N_5983,N_5663);
nand U6014 (N_6014,N_5950,N_5970);
or U6015 (N_6015,N_5760,N_5574);
nand U6016 (N_6016,N_5561,N_5636);
or U6017 (N_6017,N_5582,N_5778);
or U6018 (N_6018,N_5732,N_5884);
or U6019 (N_6019,N_5536,N_5971);
or U6020 (N_6020,N_5828,N_5515);
xnor U6021 (N_6021,N_5722,N_5958);
nand U6022 (N_6022,N_5572,N_5587);
nand U6023 (N_6023,N_5799,N_5549);
nor U6024 (N_6024,N_5929,N_5939);
and U6025 (N_6025,N_5522,N_5954);
and U6026 (N_6026,N_5686,N_5729);
and U6027 (N_6027,N_5621,N_5585);
nand U6028 (N_6028,N_5665,N_5710);
and U6029 (N_6029,N_5687,N_5912);
and U6030 (N_6030,N_5743,N_5907);
or U6031 (N_6031,N_5734,N_5789);
or U6032 (N_6032,N_5945,N_5642);
nor U6033 (N_6033,N_5920,N_5557);
nand U6034 (N_6034,N_5879,N_5616);
nor U6035 (N_6035,N_5769,N_5540);
nand U6036 (N_6036,N_5617,N_5500);
nor U6037 (N_6037,N_5541,N_5510);
or U6038 (N_6038,N_5521,N_5916);
or U6039 (N_6039,N_5957,N_5834);
or U6040 (N_6040,N_5785,N_5562);
and U6041 (N_6041,N_5986,N_5968);
or U6042 (N_6042,N_5701,N_5964);
nor U6043 (N_6043,N_5997,N_5787);
nor U6044 (N_6044,N_5886,N_5918);
nand U6045 (N_6045,N_5625,N_5668);
nor U6046 (N_6046,N_5944,N_5535);
or U6047 (N_6047,N_5948,N_5527);
nand U6048 (N_6048,N_5813,N_5824);
nand U6049 (N_6049,N_5809,N_5543);
nor U6050 (N_6050,N_5571,N_5883);
and U6051 (N_6051,N_5832,N_5606);
nand U6052 (N_6052,N_5766,N_5837);
nor U6053 (N_6053,N_5534,N_5901);
nor U6054 (N_6054,N_5633,N_5653);
or U6055 (N_6055,N_5919,N_5504);
and U6056 (N_6056,N_5586,N_5961);
nand U6057 (N_6057,N_5807,N_5648);
xor U6058 (N_6058,N_5869,N_5608);
nand U6059 (N_6059,N_5871,N_5896);
nand U6060 (N_6060,N_5672,N_5993);
nand U6061 (N_6061,N_5851,N_5863);
nand U6062 (N_6062,N_5555,N_5897);
nand U6063 (N_6063,N_5657,N_5815);
nor U6064 (N_6064,N_5723,N_5563);
and U6065 (N_6065,N_5707,N_5940);
nand U6066 (N_6066,N_5755,N_5514);
nor U6067 (N_6067,N_5539,N_5800);
nor U6068 (N_6068,N_5548,N_5516);
and U6069 (N_6069,N_5823,N_5730);
or U6070 (N_6070,N_5767,N_5731);
nor U6071 (N_6071,N_5782,N_5531);
and U6072 (N_6072,N_5894,N_5793);
and U6073 (N_6073,N_5796,N_5567);
nand U6074 (N_6074,N_5761,N_5614);
nand U6075 (N_6075,N_5565,N_5853);
nor U6076 (N_6076,N_5757,N_5895);
nand U6077 (N_6077,N_5553,N_5861);
nand U6078 (N_6078,N_5801,N_5607);
nand U6079 (N_6079,N_5599,N_5752);
nand U6080 (N_6080,N_5590,N_5704);
nand U6081 (N_6081,N_5844,N_5794);
or U6082 (N_6082,N_5699,N_5905);
and U6083 (N_6083,N_5620,N_5913);
and U6084 (N_6084,N_5671,N_5915);
nor U6085 (N_6085,N_5847,N_5751);
xnor U6086 (N_6086,N_5872,N_5717);
or U6087 (N_6087,N_5745,N_5601);
and U6088 (N_6088,N_5917,N_5598);
or U6089 (N_6089,N_5776,N_5888);
and U6090 (N_6090,N_5772,N_5693);
nand U6091 (N_6091,N_5914,N_5736);
nand U6092 (N_6092,N_5508,N_5770);
and U6093 (N_6093,N_5949,N_5864);
and U6094 (N_6094,N_5798,N_5695);
xor U6095 (N_6095,N_5644,N_5637);
xnor U6096 (N_6096,N_5524,N_5804);
or U6097 (N_6097,N_5670,N_5597);
nor U6098 (N_6098,N_5712,N_5688);
and U6099 (N_6099,N_5908,N_5960);
and U6100 (N_6100,N_5835,N_5619);
and U6101 (N_6101,N_5882,N_5887);
and U6102 (N_6102,N_5788,N_5783);
and U6103 (N_6103,N_5852,N_5934);
nand U6104 (N_6104,N_5867,N_5556);
and U6105 (N_6105,N_5705,N_5771);
or U6106 (N_6106,N_5881,N_5507);
and U6107 (N_6107,N_5649,N_5880);
and U6108 (N_6108,N_5578,N_5825);
or U6109 (N_6109,N_5792,N_5622);
nor U6110 (N_6110,N_5820,N_5669);
nor U6111 (N_6111,N_5904,N_5709);
and U6112 (N_6112,N_5951,N_5660);
nand U6113 (N_6113,N_5545,N_5513);
nand U6114 (N_6114,N_5860,N_5546);
nand U6115 (N_6115,N_5646,N_5697);
nand U6116 (N_6116,N_5509,N_5972);
or U6117 (N_6117,N_5927,N_5923);
xor U6118 (N_6118,N_5523,N_5865);
nor U6119 (N_6119,N_5877,N_5626);
nand U6120 (N_6120,N_5511,N_5750);
or U6121 (N_6121,N_5805,N_5909);
and U6122 (N_6122,N_5826,N_5978);
and U6123 (N_6123,N_5737,N_5856);
xor U6124 (N_6124,N_5937,N_5791);
and U6125 (N_6125,N_5612,N_5976);
or U6126 (N_6126,N_5594,N_5526);
and U6127 (N_6127,N_5708,N_5875);
and U6128 (N_6128,N_5533,N_5581);
and U6129 (N_6129,N_5786,N_5506);
or U6130 (N_6130,N_5739,N_5726);
and U6131 (N_6131,N_5827,N_5874);
nor U6132 (N_6132,N_5711,N_5603);
or U6133 (N_6133,N_5822,N_5850);
or U6134 (N_6134,N_5512,N_5977);
nor U6135 (N_6135,N_5746,N_5664);
or U6136 (N_6136,N_5678,N_5931);
nor U6137 (N_6137,N_5890,N_5655);
or U6138 (N_6138,N_5613,N_5839);
and U6139 (N_6139,N_5763,N_5967);
nand U6140 (N_6140,N_5652,N_5638);
nor U6141 (N_6141,N_5673,N_5683);
or U6142 (N_6142,N_5728,N_5990);
nor U6143 (N_6143,N_5952,N_5889);
nor U6144 (N_6144,N_5714,N_5542);
nand U6145 (N_6145,N_5816,N_5593);
and U6146 (N_6146,N_5906,N_5554);
nor U6147 (N_6147,N_5747,N_5803);
and U6148 (N_6148,N_5628,N_5995);
xnor U6149 (N_6149,N_5857,N_5899);
or U6150 (N_6150,N_5530,N_5632);
or U6151 (N_6151,N_5602,N_5575);
nand U6152 (N_6152,N_5965,N_5690);
and U6153 (N_6153,N_5532,N_5579);
nor U6154 (N_6154,N_5596,N_5935);
nor U6155 (N_6155,N_5706,N_5987);
nand U6156 (N_6156,N_5818,N_5519);
nor U6157 (N_6157,N_5740,N_5624);
nor U6158 (N_6158,N_5592,N_5963);
or U6159 (N_6159,N_5900,N_5696);
and U6160 (N_6160,N_5955,N_5893);
and U6161 (N_6161,N_5682,N_5790);
or U6162 (N_6162,N_5777,N_5806);
and U6163 (N_6163,N_5762,N_5947);
and U6164 (N_6164,N_5992,N_5833);
or U6165 (N_6165,N_5996,N_5930);
nand U6166 (N_6166,N_5661,N_5694);
xor U6167 (N_6167,N_5784,N_5639);
and U6168 (N_6168,N_5892,N_5946);
xor U6169 (N_6169,N_5774,N_5858);
and U6170 (N_6170,N_5538,N_5610);
or U6171 (N_6171,N_5640,N_5570);
xor U6172 (N_6172,N_5654,N_5566);
nor U6173 (N_6173,N_5645,N_5765);
nand U6174 (N_6174,N_5698,N_5716);
nand U6175 (N_6175,N_5662,N_5584);
or U6176 (N_6176,N_5583,N_5600);
or U6177 (N_6177,N_5501,N_5719);
and U6178 (N_6178,N_5848,N_5910);
or U6179 (N_6179,N_5922,N_5721);
and U6180 (N_6180,N_5692,N_5854);
nor U6181 (N_6181,N_5689,N_5588);
nand U6182 (N_6182,N_5862,N_5604);
nand U6183 (N_6183,N_5868,N_5560);
nor U6184 (N_6184,N_5795,N_5650);
nor U6185 (N_6185,N_5502,N_5666);
or U6186 (N_6186,N_5921,N_5568);
or U6187 (N_6187,N_5715,N_5768);
nand U6188 (N_6188,N_5595,N_5685);
and U6189 (N_6189,N_5870,N_5677);
or U6190 (N_6190,N_5753,N_5810);
nand U6191 (N_6191,N_5924,N_5559);
nor U6192 (N_6192,N_5814,N_5713);
and U6193 (N_6193,N_5979,N_5956);
nor U6194 (N_6194,N_5675,N_5656);
and U6195 (N_6195,N_5982,N_5741);
or U6196 (N_6196,N_5758,N_5981);
and U6197 (N_6197,N_5756,N_5551);
nand U6198 (N_6198,N_5647,N_5627);
or U6199 (N_6199,N_5643,N_5891);
or U6200 (N_6200,N_5759,N_5681);
nor U6201 (N_6201,N_5898,N_5938);
or U6202 (N_6202,N_5984,N_5577);
and U6203 (N_6203,N_5727,N_5589);
and U6204 (N_6204,N_5724,N_5611);
or U6205 (N_6205,N_5773,N_5775);
or U6206 (N_6206,N_5840,N_5700);
nand U6207 (N_6207,N_5989,N_5634);
nor U6208 (N_6208,N_5842,N_5928);
or U6209 (N_6209,N_5936,N_5841);
xnor U6210 (N_6210,N_5576,N_5529);
or U6211 (N_6211,N_5911,N_5866);
or U6212 (N_6212,N_5985,N_5651);
xor U6213 (N_6213,N_5558,N_5829);
and U6214 (N_6214,N_5926,N_5659);
and U6215 (N_6215,N_5503,N_5903);
nor U6216 (N_6216,N_5973,N_5537);
nand U6217 (N_6217,N_5802,N_5517);
and U6218 (N_6218,N_5974,N_5518);
nand U6219 (N_6219,N_5630,N_5812);
and U6220 (N_6220,N_5941,N_5943);
or U6221 (N_6221,N_5635,N_5591);
nand U6222 (N_6222,N_5658,N_5528);
or U6223 (N_6223,N_5618,N_5838);
xor U6224 (N_6224,N_5764,N_5845);
nor U6225 (N_6225,N_5547,N_5821);
and U6226 (N_6226,N_5885,N_5544);
or U6227 (N_6227,N_5749,N_5720);
nand U6228 (N_6228,N_5525,N_5748);
or U6229 (N_6229,N_5564,N_5962);
nor U6230 (N_6230,N_5797,N_5702);
and U6231 (N_6231,N_5925,N_5843);
and U6232 (N_6232,N_5580,N_5605);
or U6233 (N_6233,N_5998,N_5953);
or U6234 (N_6234,N_5846,N_5808);
nand U6235 (N_6235,N_5691,N_5641);
xnor U6236 (N_6236,N_5819,N_5817);
nand U6237 (N_6237,N_5991,N_5859);
and U6238 (N_6238,N_5744,N_5703);
nor U6239 (N_6239,N_5836,N_5780);
nand U6240 (N_6240,N_5735,N_5569);
or U6241 (N_6241,N_5631,N_5742);
nor U6242 (N_6242,N_5684,N_5718);
nor U6243 (N_6243,N_5520,N_5902);
xor U6244 (N_6244,N_5969,N_5629);
xor U6245 (N_6245,N_5679,N_5733);
and U6246 (N_6246,N_5994,N_5959);
and U6247 (N_6247,N_5966,N_5988);
xor U6248 (N_6248,N_5725,N_5667);
nand U6249 (N_6249,N_5980,N_5676);
or U6250 (N_6250,N_5618,N_5887);
nand U6251 (N_6251,N_5669,N_5734);
or U6252 (N_6252,N_5649,N_5953);
and U6253 (N_6253,N_5975,N_5665);
nor U6254 (N_6254,N_5876,N_5727);
nor U6255 (N_6255,N_5838,N_5769);
nand U6256 (N_6256,N_5666,N_5556);
or U6257 (N_6257,N_5584,N_5586);
nor U6258 (N_6258,N_5725,N_5555);
nand U6259 (N_6259,N_5662,N_5955);
nand U6260 (N_6260,N_5926,N_5783);
or U6261 (N_6261,N_5618,N_5596);
nand U6262 (N_6262,N_5514,N_5987);
xor U6263 (N_6263,N_5702,N_5735);
nand U6264 (N_6264,N_5950,N_5513);
or U6265 (N_6265,N_5772,N_5978);
nor U6266 (N_6266,N_5703,N_5982);
or U6267 (N_6267,N_5855,N_5533);
and U6268 (N_6268,N_5972,N_5981);
or U6269 (N_6269,N_5531,N_5845);
and U6270 (N_6270,N_5723,N_5616);
and U6271 (N_6271,N_5893,N_5695);
nand U6272 (N_6272,N_5682,N_5948);
or U6273 (N_6273,N_5567,N_5757);
and U6274 (N_6274,N_5963,N_5897);
nor U6275 (N_6275,N_5763,N_5736);
and U6276 (N_6276,N_5795,N_5660);
nor U6277 (N_6277,N_5672,N_5955);
nand U6278 (N_6278,N_5829,N_5932);
nor U6279 (N_6279,N_5598,N_5966);
xor U6280 (N_6280,N_5942,N_5670);
nand U6281 (N_6281,N_5636,N_5907);
nor U6282 (N_6282,N_5725,N_5818);
nor U6283 (N_6283,N_5738,N_5592);
nor U6284 (N_6284,N_5797,N_5925);
nand U6285 (N_6285,N_5992,N_5789);
or U6286 (N_6286,N_5561,N_5547);
and U6287 (N_6287,N_5677,N_5672);
or U6288 (N_6288,N_5951,N_5619);
nand U6289 (N_6289,N_5743,N_5697);
xnor U6290 (N_6290,N_5898,N_5517);
xor U6291 (N_6291,N_5657,N_5904);
and U6292 (N_6292,N_5984,N_5728);
and U6293 (N_6293,N_5974,N_5692);
nor U6294 (N_6294,N_5980,N_5894);
and U6295 (N_6295,N_5547,N_5707);
nor U6296 (N_6296,N_5932,N_5535);
or U6297 (N_6297,N_5868,N_5620);
nor U6298 (N_6298,N_5894,N_5891);
nor U6299 (N_6299,N_5712,N_5707);
nand U6300 (N_6300,N_5967,N_5658);
nor U6301 (N_6301,N_5887,N_5753);
nor U6302 (N_6302,N_5615,N_5854);
nand U6303 (N_6303,N_5979,N_5761);
nor U6304 (N_6304,N_5705,N_5902);
and U6305 (N_6305,N_5690,N_5696);
nand U6306 (N_6306,N_5836,N_5797);
nand U6307 (N_6307,N_5576,N_5660);
and U6308 (N_6308,N_5658,N_5698);
and U6309 (N_6309,N_5706,N_5712);
nand U6310 (N_6310,N_5585,N_5530);
nand U6311 (N_6311,N_5542,N_5807);
or U6312 (N_6312,N_5809,N_5939);
nand U6313 (N_6313,N_5789,N_5630);
and U6314 (N_6314,N_5806,N_5680);
nor U6315 (N_6315,N_5502,N_5817);
or U6316 (N_6316,N_5543,N_5629);
or U6317 (N_6317,N_5957,N_5852);
or U6318 (N_6318,N_5525,N_5860);
nand U6319 (N_6319,N_5998,N_5518);
and U6320 (N_6320,N_5977,N_5681);
nor U6321 (N_6321,N_5576,N_5920);
and U6322 (N_6322,N_5543,N_5854);
or U6323 (N_6323,N_5553,N_5820);
xnor U6324 (N_6324,N_5819,N_5788);
nor U6325 (N_6325,N_5775,N_5820);
xnor U6326 (N_6326,N_5522,N_5702);
nor U6327 (N_6327,N_5919,N_5534);
nor U6328 (N_6328,N_5542,N_5680);
nand U6329 (N_6329,N_5885,N_5980);
nand U6330 (N_6330,N_5855,N_5742);
and U6331 (N_6331,N_5872,N_5760);
or U6332 (N_6332,N_5906,N_5739);
nor U6333 (N_6333,N_5696,N_5761);
or U6334 (N_6334,N_5908,N_5708);
and U6335 (N_6335,N_5960,N_5941);
and U6336 (N_6336,N_5637,N_5664);
and U6337 (N_6337,N_5611,N_5766);
or U6338 (N_6338,N_5582,N_5911);
nor U6339 (N_6339,N_5820,N_5827);
and U6340 (N_6340,N_5618,N_5831);
nor U6341 (N_6341,N_5611,N_5506);
xnor U6342 (N_6342,N_5770,N_5806);
or U6343 (N_6343,N_5829,N_5514);
and U6344 (N_6344,N_5841,N_5989);
and U6345 (N_6345,N_5975,N_5553);
or U6346 (N_6346,N_5582,N_5810);
xnor U6347 (N_6347,N_5633,N_5741);
nor U6348 (N_6348,N_5501,N_5626);
and U6349 (N_6349,N_5585,N_5934);
or U6350 (N_6350,N_5688,N_5950);
xnor U6351 (N_6351,N_5779,N_5826);
nand U6352 (N_6352,N_5702,N_5563);
or U6353 (N_6353,N_5969,N_5971);
and U6354 (N_6354,N_5523,N_5968);
nor U6355 (N_6355,N_5981,N_5725);
and U6356 (N_6356,N_5753,N_5554);
nand U6357 (N_6357,N_5736,N_5871);
nor U6358 (N_6358,N_5677,N_5882);
nor U6359 (N_6359,N_5507,N_5863);
nand U6360 (N_6360,N_5675,N_5650);
or U6361 (N_6361,N_5848,N_5884);
or U6362 (N_6362,N_5626,N_5947);
or U6363 (N_6363,N_5623,N_5686);
or U6364 (N_6364,N_5679,N_5622);
nor U6365 (N_6365,N_5820,N_5720);
and U6366 (N_6366,N_5646,N_5651);
nand U6367 (N_6367,N_5992,N_5794);
nor U6368 (N_6368,N_5898,N_5937);
or U6369 (N_6369,N_5706,N_5789);
nor U6370 (N_6370,N_5929,N_5570);
and U6371 (N_6371,N_5518,N_5997);
and U6372 (N_6372,N_5921,N_5595);
nor U6373 (N_6373,N_5808,N_5837);
and U6374 (N_6374,N_5773,N_5628);
or U6375 (N_6375,N_5912,N_5914);
xor U6376 (N_6376,N_5846,N_5792);
nor U6377 (N_6377,N_5923,N_5806);
nor U6378 (N_6378,N_5966,N_5780);
nand U6379 (N_6379,N_5975,N_5593);
nand U6380 (N_6380,N_5928,N_5665);
nand U6381 (N_6381,N_5601,N_5629);
and U6382 (N_6382,N_5764,N_5880);
and U6383 (N_6383,N_5699,N_5867);
and U6384 (N_6384,N_5836,N_5867);
or U6385 (N_6385,N_5739,N_5541);
nand U6386 (N_6386,N_5554,N_5739);
and U6387 (N_6387,N_5588,N_5876);
nand U6388 (N_6388,N_5596,N_5611);
and U6389 (N_6389,N_5629,N_5696);
xor U6390 (N_6390,N_5891,N_5713);
nor U6391 (N_6391,N_5700,N_5829);
and U6392 (N_6392,N_5842,N_5583);
nor U6393 (N_6393,N_5940,N_5753);
or U6394 (N_6394,N_5675,N_5895);
nand U6395 (N_6395,N_5595,N_5855);
or U6396 (N_6396,N_5629,N_5952);
nand U6397 (N_6397,N_5774,N_5505);
or U6398 (N_6398,N_5564,N_5931);
nor U6399 (N_6399,N_5961,N_5826);
nand U6400 (N_6400,N_5624,N_5667);
or U6401 (N_6401,N_5909,N_5681);
nor U6402 (N_6402,N_5534,N_5793);
nand U6403 (N_6403,N_5794,N_5994);
or U6404 (N_6404,N_5532,N_5747);
and U6405 (N_6405,N_5930,N_5691);
nor U6406 (N_6406,N_5540,N_5991);
or U6407 (N_6407,N_5531,N_5521);
and U6408 (N_6408,N_5660,N_5913);
or U6409 (N_6409,N_5569,N_5537);
xor U6410 (N_6410,N_5509,N_5643);
and U6411 (N_6411,N_5888,N_5825);
nor U6412 (N_6412,N_5869,N_5900);
and U6413 (N_6413,N_5797,N_5844);
and U6414 (N_6414,N_5771,N_5897);
nand U6415 (N_6415,N_5613,N_5995);
nor U6416 (N_6416,N_5895,N_5970);
nor U6417 (N_6417,N_5703,N_5952);
or U6418 (N_6418,N_5889,N_5714);
and U6419 (N_6419,N_5626,N_5500);
or U6420 (N_6420,N_5643,N_5793);
nand U6421 (N_6421,N_5519,N_5875);
and U6422 (N_6422,N_5618,N_5998);
nor U6423 (N_6423,N_5523,N_5906);
and U6424 (N_6424,N_5956,N_5771);
nand U6425 (N_6425,N_5638,N_5943);
and U6426 (N_6426,N_5512,N_5921);
nor U6427 (N_6427,N_5668,N_5718);
and U6428 (N_6428,N_5678,N_5590);
and U6429 (N_6429,N_5657,N_5586);
and U6430 (N_6430,N_5988,N_5620);
nor U6431 (N_6431,N_5762,N_5615);
or U6432 (N_6432,N_5660,N_5762);
or U6433 (N_6433,N_5685,N_5647);
nor U6434 (N_6434,N_5912,N_5507);
and U6435 (N_6435,N_5939,N_5673);
or U6436 (N_6436,N_5740,N_5627);
nor U6437 (N_6437,N_5776,N_5577);
xor U6438 (N_6438,N_5831,N_5564);
nand U6439 (N_6439,N_5996,N_5809);
or U6440 (N_6440,N_5633,N_5983);
xor U6441 (N_6441,N_5884,N_5549);
xor U6442 (N_6442,N_5877,N_5955);
or U6443 (N_6443,N_5593,N_5624);
xor U6444 (N_6444,N_5641,N_5708);
nand U6445 (N_6445,N_5847,N_5673);
and U6446 (N_6446,N_5974,N_5641);
or U6447 (N_6447,N_5983,N_5771);
nand U6448 (N_6448,N_5773,N_5834);
or U6449 (N_6449,N_5907,N_5689);
or U6450 (N_6450,N_5676,N_5530);
and U6451 (N_6451,N_5901,N_5844);
or U6452 (N_6452,N_5608,N_5704);
or U6453 (N_6453,N_5950,N_5728);
nand U6454 (N_6454,N_5937,N_5774);
or U6455 (N_6455,N_5510,N_5864);
nor U6456 (N_6456,N_5506,N_5719);
nor U6457 (N_6457,N_5510,N_5686);
nor U6458 (N_6458,N_5812,N_5862);
nor U6459 (N_6459,N_5928,N_5752);
nor U6460 (N_6460,N_5761,N_5573);
nor U6461 (N_6461,N_5923,N_5942);
nand U6462 (N_6462,N_5616,N_5762);
and U6463 (N_6463,N_5509,N_5507);
and U6464 (N_6464,N_5955,N_5728);
nand U6465 (N_6465,N_5513,N_5915);
and U6466 (N_6466,N_5836,N_5566);
nor U6467 (N_6467,N_5982,N_5668);
nand U6468 (N_6468,N_5860,N_5631);
xor U6469 (N_6469,N_5923,N_5895);
nor U6470 (N_6470,N_5829,N_5845);
or U6471 (N_6471,N_5803,N_5726);
nand U6472 (N_6472,N_5944,N_5854);
or U6473 (N_6473,N_5698,N_5865);
nor U6474 (N_6474,N_5566,N_5716);
and U6475 (N_6475,N_5948,N_5700);
nand U6476 (N_6476,N_5704,N_5719);
nor U6477 (N_6477,N_5588,N_5728);
or U6478 (N_6478,N_5667,N_5933);
or U6479 (N_6479,N_5646,N_5912);
and U6480 (N_6480,N_5620,N_5824);
nand U6481 (N_6481,N_5675,N_5509);
or U6482 (N_6482,N_5500,N_5812);
or U6483 (N_6483,N_5730,N_5819);
and U6484 (N_6484,N_5947,N_5957);
nor U6485 (N_6485,N_5925,N_5719);
nor U6486 (N_6486,N_5690,N_5882);
and U6487 (N_6487,N_5506,N_5519);
or U6488 (N_6488,N_5840,N_5911);
xnor U6489 (N_6489,N_5815,N_5650);
nand U6490 (N_6490,N_5990,N_5906);
nand U6491 (N_6491,N_5929,N_5968);
and U6492 (N_6492,N_5774,N_5811);
and U6493 (N_6493,N_5530,N_5699);
nand U6494 (N_6494,N_5601,N_5795);
nor U6495 (N_6495,N_5799,N_5771);
nor U6496 (N_6496,N_5996,N_5830);
or U6497 (N_6497,N_5580,N_5600);
nor U6498 (N_6498,N_5882,N_5819);
and U6499 (N_6499,N_5755,N_5645);
or U6500 (N_6500,N_6497,N_6327);
and U6501 (N_6501,N_6000,N_6390);
nand U6502 (N_6502,N_6323,N_6269);
nor U6503 (N_6503,N_6300,N_6185);
nand U6504 (N_6504,N_6002,N_6080);
or U6505 (N_6505,N_6156,N_6238);
xor U6506 (N_6506,N_6141,N_6160);
nor U6507 (N_6507,N_6279,N_6313);
nand U6508 (N_6508,N_6006,N_6482);
nor U6509 (N_6509,N_6486,N_6363);
xnor U6510 (N_6510,N_6399,N_6217);
or U6511 (N_6511,N_6081,N_6395);
or U6512 (N_6512,N_6388,N_6094);
and U6513 (N_6513,N_6176,N_6367);
nor U6514 (N_6514,N_6396,N_6254);
and U6515 (N_6515,N_6010,N_6472);
nand U6516 (N_6516,N_6284,N_6349);
nand U6517 (N_6517,N_6423,N_6484);
xor U6518 (N_6518,N_6461,N_6274);
nor U6519 (N_6519,N_6030,N_6403);
nor U6520 (N_6520,N_6223,N_6014);
and U6521 (N_6521,N_6364,N_6085);
or U6522 (N_6522,N_6192,N_6197);
and U6523 (N_6523,N_6249,N_6177);
or U6524 (N_6524,N_6152,N_6454);
or U6525 (N_6525,N_6400,N_6431);
xor U6526 (N_6526,N_6491,N_6060);
nor U6527 (N_6527,N_6154,N_6077);
or U6528 (N_6528,N_6414,N_6195);
and U6529 (N_6529,N_6048,N_6096);
nand U6530 (N_6530,N_6161,N_6107);
or U6531 (N_6531,N_6070,N_6270);
and U6532 (N_6532,N_6487,N_6035);
nand U6533 (N_6533,N_6353,N_6265);
or U6534 (N_6534,N_6459,N_6375);
and U6535 (N_6535,N_6047,N_6319);
nand U6536 (N_6536,N_6291,N_6130);
nand U6537 (N_6537,N_6456,N_6286);
nor U6538 (N_6538,N_6278,N_6432);
nand U6539 (N_6539,N_6490,N_6138);
xor U6540 (N_6540,N_6241,N_6343);
nand U6541 (N_6541,N_6451,N_6131);
nand U6542 (N_6542,N_6452,N_6493);
nand U6543 (N_6543,N_6440,N_6088);
nand U6544 (N_6544,N_6236,N_6429);
or U6545 (N_6545,N_6023,N_6168);
or U6546 (N_6546,N_6372,N_6253);
or U6547 (N_6547,N_6449,N_6143);
and U6548 (N_6548,N_6317,N_6106);
nor U6549 (N_6549,N_6234,N_6444);
xnor U6550 (N_6550,N_6303,N_6113);
or U6551 (N_6551,N_6032,N_6090);
or U6552 (N_6552,N_6204,N_6275);
or U6553 (N_6553,N_6439,N_6139);
nor U6554 (N_6554,N_6295,N_6341);
and U6555 (N_6555,N_6261,N_6338);
xor U6556 (N_6556,N_6342,N_6436);
xor U6557 (N_6557,N_6147,N_6412);
nand U6558 (N_6558,N_6332,N_6049);
nor U6559 (N_6559,N_6103,N_6114);
nand U6560 (N_6560,N_6268,N_6345);
or U6561 (N_6561,N_6126,N_6215);
nand U6562 (N_6562,N_6335,N_6038);
or U6563 (N_6563,N_6173,N_6229);
and U6564 (N_6564,N_6251,N_6026);
or U6565 (N_6565,N_6473,N_6155);
or U6566 (N_6566,N_6157,N_6446);
and U6567 (N_6567,N_6329,N_6489);
nand U6568 (N_6568,N_6151,N_6443);
and U6569 (N_6569,N_6174,N_6166);
or U6570 (N_6570,N_6434,N_6101);
nand U6571 (N_6571,N_6153,N_6257);
or U6572 (N_6572,N_6277,N_6182);
nor U6573 (N_6573,N_6383,N_6015);
and U6574 (N_6574,N_6149,N_6306);
xnor U6575 (N_6575,N_6496,N_6029);
nand U6576 (N_6576,N_6424,N_6333);
and U6577 (N_6577,N_6072,N_6056);
nor U6578 (N_6578,N_6016,N_6425);
nor U6579 (N_6579,N_6453,N_6296);
nor U6580 (N_6580,N_6078,N_6122);
and U6581 (N_6581,N_6068,N_6172);
nor U6582 (N_6582,N_6137,N_6039);
or U6583 (N_6583,N_6045,N_6393);
and U6584 (N_6584,N_6361,N_6104);
or U6585 (N_6585,N_6178,N_6227);
and U6586 (N_6586,N_6162,N_6075);
nand U6587 (N_6587,N_6376,N_6159);
nand U6588 (N_6588,N_6328,N_6212);
or U6589 (N_6589,N_6012,N_6356);
nand U6590 (N_6590,N_6124,N_6437);
and U6591 (N_6591,N_6301,N_6109);
and U6592 (N_6592,N_6209,N_6442);
and U6593 (N_6593,N_6475,N_6460);
xnor U6594 (N_6594,N_6410,N_6211);
nand U6595 (N_6595,N_6381,N_6214);
nor U6596 (N_6596,N_6044,N_6441);
or U6597 (N_6597,N_6213,N_6042);
xor U6598 (N_6598,N_6339,N_6447);
nand U6599 (N_6599,N_6171,N_6387);
or U6600 (N_6600,N_6190,N_6478);
xor U6601 (N_6601,N_6320,N_6315);
or U6602 (N_6602,N_6189,N_6310);
nor U6603 (N_6603,N_6005,N_6028);
nand U6604 (N_6604,N_6224,N_6272);
nor U6605 (N_6605,N_6256,N_6470);
nor U6606 (N_6606,N_6054,N_6466);
or U6607 (N_6607,N_6200,N_6148);
or U6608 (N_6608,N_6464,N_6357);
nor U6609 (N_6609,N_6202,N_6108);
or U6610 (N_6610,N_6417,N_6179);
and U6611 (N_6611,N_6231,N_6293);
xnor U6612 (N_6612,N_6102,N_6145);
or U6613 (N_6613,N_6260,N_6302);
nor U6614 (N_6614,N_6298,N_6312);
and U6615 (N_6615,N_6405,N_6471);
nor U6616 (N_6616,N_6205,N_6347);
or U6617 (N_6617,N_6289,N_6061);
or U6618 (N_6618,N_6379,N_6389);
and U6619 (N_6619,N_6468,N_6422);
xor U6620 (N_6620,N_6116,N_6309);
or U6621 (N_6621,N_6017,N_6409);
nand U6622 (N_6622,N_6326,N_6184);
xnor U6623 (N_6623,N_6067,N_6201);
nor U6624 (N_6624,N_6084,N_6355);
nand U6625 (N_6625,N_6052,N_6426);
and U6626 (N_6626,N_6411,N_6243);
and U6627 (N_6627,N_6034,N_6239);
nand U6628 (N_6628,N_6262,N_6210);
or U6629 (N_6629,N_6398,N_6290);
nor U6630 (N_6630,N_6354,N_6105);
and U6631 (N_6631,N_6255,N_6371);
nand U6632 (N_6632,N_6311,N_6421);
nand U6633 (N_6633,N_6391,N_6180);
or U6634 (N_6634,N_6370,N_6271);
and U6635 (N_6635,N_6198,N_6001);
or U6636 (N_6636,N_6024,N_6233);
or U6637 (N_6637,N_6183,N_6066);
and U6638 (N_6638,N_6469,N_6420);
and U6639 (N_6639,N_6465,N_6494);
nor U6640 (N_6640,N_6165,N_6071);
and U6641 (N_6641,N_6076,N_6267);
or U6642 (N_6642,N_6093,N_6083);
xor U6643 (N_6643,N_6118,N_6053);
nand U6644 (N_6644,N_6033,N_6366);
xnor U6645 (N_6645,N_6373,N_6404);
nand U6646 (N_6646,N_6397,N_6134);
and U6647 (N_6647,N_6266,N_6158);
nand U6648 (N_6648,N_6402,N_6074);
nor U6649 (N_6649,N_6350,N_6430);
or U6650 (N_6650,N_6287,N_6457);
nor U6651 (N_6651,N_6352,N_6428);
nand U6652 (N_6652,N_6294,N_6374);
nand U6653 (N_6653,N_6462,N_6377);
xor U6654 (N_6654,N_6282,N_6021);
and U6655 (N_6655,N_6069,N_6082);
or U6656 (N_6656,N_6163,N_6401);
xnor U6657 (N_6657,N_6463,N_6427);
xor U6658 (N_6658,N_6040,N_6055);
nand U6659 (N_6659,N_6481,N_6100);
and U6660 (N_6660,N_6140,N_6142);
xnor U6661 (N_6661,N_6110,N_6089);
or U6662 (N_6662,N_6226,N_6499);
or U6663 (N_6663,N_6351,N_6498);
nor U6664 (N_6664,N_6119,N_6288);
or U6665 (N_6665,N_6416,N_6285);
and U6666 (N_6666,N_6479,N_6230);
nand U6667 (N_6667,N_6264,N_6276);
or U6668 (N_6668,N_6187,N_6120);
xnor U6669 (N_6669,N_6435,N_6087);
nor U6670 (N_6670,N_6348,N_6136);
and U6671 (N_6671,N_6369,N_6208);
nand U6672 (N_6672,N_6181,N_6123);
or U6673 (N_6673,N_6170,N_6216);
nor U6674 (N_6674,N_6359,N_6025);
or U6675 (N_6675,N_6413,N_6018);
or U6676 (N_6676,N_6477,N_6408);
or U6677 (N_6677,N_6304,N_6144);
nor U6678 (N_6678,N_6036,N_6091);
nand U6679 (N_6679,N_6228,N_6220);
and U6680 (N_6680,N_6191,N_6219);
nand U6681 (N_6681,N_6007,N_6199);
xor U6682 (N_6682,N_6150,N_6186);
nand U6683 (N_6683,N_6382,N_6225);
nor U6684 (N_6684,N_6135,N_6283);
nand U6685 (N_6685,N_6368,N_6237);
nor U6686 (N_6686,N_6059,N_6063);
nor U6687 (N_6687,N_6065,N_6246);
nand U6688 (N_6688,N_6194,N_6248);
nor U6689 (N_6689,N_6020,N_6308);
and U6690 (N_6690,N_6188,N_6128);
nor U6691 (N_6691,N_6314,N_6222);
or U6692 (N_6692,N_6167,N_6344);
nand U6693 (N_6693,N_6346,N_6146);
nand U6694 (N_6694,N_6221,N_6206);
and U6695 (N_6695,N_6235,N_6384);
xor U6696 (N_6696,N_6242,N_6438);
or U6697 (N_6697,N_6406,N_6419);
or U6698 (N_6698,N_6316,N_6095);
nand U6699 (N_6699,N_6232,N_6331);
nor U6700 (N_6700,N_6307,N_6098);
and U6701 (N_6701,N_6008,N_6474);
or U6702 (N_6702,N_6340,N_6051);
nor U6703 (N_6703,N_6132,N_6019);
or U6704 (N_6704,N_6245,N_6380);
or U6705 (N_6705,N_6495,N_6488);
nand U6706 (N_6706,N_6252,N_6013);
nor U6707 (N_6707,N_6458,N_6196);
or U6708 (N_6708,N_6111,N_6292);
or U6709 (N_6709,N_6322,N_6455);
and U6710 (N_6710,N_6492,N_6485);
xnor U6711 (N_6711,N_6041,N_6450);
nand U6712 (N_6712,N_6448,N_6378);
nor U6713 (N_6713,N_6133,N_6043);
nor U6714 (N_6714,N_6004,N_6297);
nand U6715 (N_6715,N_6476,N_6392);
nor U6716 (N_6716,N_6031,N_6099);
nor U6717 (N_6717,N_6097,N_6263);
or U6718 (N_6718,N_6480,N_6092);
nand U6719 (N_6719,N_6325,N_6299);
nand U6720 (N_6720,N_6250,N_6305);
nand U6721 (N_6721,N_6321,N_6445);
xnor U6722 (N_6722,N_6218,N_6467);
nand U6723 (N_6723,N_6244,N_6280);
or U6724 (N_6724,N_6324,N_6079);
and U6725 (N_6725,N_6037,N_6117);
and U6726 (N_6726,N_6062,N_6362);
nand U6727 (N_6727,N_6073,N_6330);
and U6728 (N_6728,N_6164,N_6009);
nor U6729 (N_6729,N_6046,N_6318);
nand U6730 (N_6730,N_6121,N_6281);
nand U6731 (N_6731,N_6386,N_6358);
and U6732 (N_6732,N_6129,N_6112);
and U6733 (N_6733,N_6193,N_6259);
nor U6734 (N_6734,N_6337,N_6125);
or U6735 (N_6735,N_6240,N_6336);
nand U6736 (N_6736,N_6334,N_6365);
or U6737 (N_6737,N_6011,N_6433);
xor U6738 (N_6738,N_6115,N_6022);
or U6739 (N_6739,N_6175,N_6247);
and U6740 (N_6740,N_6203,N_6127);
nor U6741 (N_6741,N_6050,N_6086);
or U6742 (N_6742,N_6418,N_6057);
nand U6743 (N_6743,N_6407,N_6385);
nand U6744 (N_6744,N_6415,N_6483);
nor U6745 (N_6745,N_6360,N_6058);
nor U6746 (N_6746,N_6027,N_6064);
or U6747 (N_6747,N_6394,N_6273);
xnor U6748 (N_6748,N_6258,N_6169);
and U6749 (N_6749,N_6003,N_6207);
and U6750 (N_6750,N_6147,N_6437);
nor U6751 (N_6751,N_6089,N_6395);
or U6752 (N_6752,N_6019,N_6271);
or U6753 (N_6753,N_6102,N_6299);
nand U6754 (N_6754,N_6043,N_6137);
nand U6755 (N_6755,N_6429,N_6228);
or U6756 (N_6756,N_6296,N_6145);
nor U6757 (N_6757,N_6346,N_6149);
nor U6758 (N_6758,N_6033,N_6462);
xor U6759 (N_6759,N_6207,N_6200);
or U6760 (N_6760,N_6223,N_6350);
nor U6761 (N_6761,N_6497,N_6379);
nand U6762 (N_6762,N_6450,N_6377);
nand U6763 (N_6763,N_6347,N_6408);
nand U6764 (N_6764,N_6204,N_6242);
nor U6765 (N_6765,N_6100,N_6343);
and U6766 (N_6766,N_6257,N_6020);
nor U6767 (N_6767,N_6126,N_6414);
and U6768 (N_6768,N_6491,N_6227);
or U6769 (N_6769,N_6480,N_6200);
and U6770 (N_6770,N_6257,N_6243);
and U6771 (N_6771,N_6152,N_6444);
xor U6772 (N_6772,N_6067,N_6414);
or U6773 (N_6773,N_6104,N_6316);
and U6774 (N_6774,N_6382,N_6147);
xor U6775 (N_6775,N_6419,N_6263);
and U6776 (N_6776,N_6332,N_6269);
or U6777 (N_6777,N_6470,N_6184);
nor U6778 (N_6778,N_6486,N_6480);
nand U6779 (N_6779,N_6175,N_6451);
and U6780 (N_6780,N_6214,N_6276);
and U6781 (N_6781,N_6019,N_6014);
nor U6782 (N_6782,N_6481,N_6096);
xnor U6783 (N_6783,N_6473,N_6154);
or U6784 (N_6784,N_6447,N_6317);
nor U6785 (N_6785,N_6320,N_6069);
nor U6786 (N_6786,N_6131,N_6281);
or U6787 (N_6787,N_6121,N_6026);
and U6788 (N_6788,N_6299,N_6132);
and U6789 (N_6789,N_6157,N_6123);
and U6790 (N_6790,N_6026,N_6359);
nand U6791 (N_6791,N_6114,N_6347);
or U6792 (N_6792,N_6160,N_6469);
and U6793 (N_6793,N_6299,N_6316);
xor U6794 (N_6794,N_6040,N_6231);
xnor U6795 (N_6795,N_6445,N_6305);
nand U6796 (N_6796,N_6422,N_6231);
xor U6797 (N_6797,N_6043,N_6020);
nand U6798 (N_6798,N_6495,N_6286);
xnor U6799 (N_6799,N_6386,N_6078);
nand U6800 (N_6800,N_6018,N_6458);
nor U6801 (N_6801,N_6194,N_6237);
xnor U6802 (N_6802,N_6277,N_6484);
or U6803 (N_6803,N_6117,N_6084);
and U6804 (N_6804,N_6322,N_6443);
nor U6805 (N_6805,N_6341,N_6423);
nand U6806 (N_6806,N_6104,N_6017);
and U6807 (N_6807,N_6428,N_6020);
nand U6808 (N_6808,N_6344,N_6281);
nand U6809 (N_6809,N_6378,N_6210);
or U6810 (N_6810,N_6056,N_6196);
or U6811 (N_6811,N_6073,N_6466);
nor U6812 (N_6812,N_6159,N_6243);
xnor U6813 (N_6813,N_6426,N_6363);
and U6814 (N_6814,N_6039,N_6466);
nor U6815 (N_6815,N_6019,N_6433);
nor U6816 (N_6816,N_6488,N_6362);
or U6817 (N_6817,N_6169,N_6450);
nand U6818 (N_6818,N_6367,N_6470);
nand U6819 (N_6819,N_6359,N_6443);
nand U6820 (N_6820,N_6463,N_6032);
or U6821 (N_6821,N_6414,N_6253);
nor U6822 (N_6822,N_6333,N_6290);
nand U6823 (N_6823,N_6048,N_6238);
nor U6824 (N_6824,N_6423,N_6057);
and U6825 (N_6825,N_6048,N_6188);
and U6826 (N_6826,N_6121,N_6108);
nor U6827 (N_6827,N_6283,N_6266);
nand U6828 (N_6828,N_6069,N_6188);
nor U6829 (N_6829,N_6445,N_6013);
nand U6830 (N_6830,N_6490,N_6304);
nand U6831 (N_6831,N_6287,N_6054);
or U6832 (N_6832,N_6064,N_6446);
nand U6833 (N_6833,N_6009,N_6207);
nand U6834 (N_6834,N_6322,N_6109);
nor U6835 (N_6835,N_6388,N_6060);
or U6836 (N_6836,N_6080,N_6318);
xor U6837 (N_6837,N_6388,N_6225);
nor U6838 (N_6838,N_6189,N_6373);
nor U6839 (N_6839,N_6224,N_6156);
xnor U6840 (N_6840,N_6096,N_6329);
and U6841 (N_6841,N_6159,N_6457);
nor U6842 (N_6842,N_6256,N_6104);
nor U6843 (N_6843,N_6278,N_6126);
and U6844 (N_6844,N_6484,N_6435);
xnor U6845 (N_6845,N_6003,N_6148);
or U6846 (N_6846,N_6071,N_6181);
nand U6847 (N_6847,N_6133,N_6129);
nand U6848 (N_6848,N_6235,N_6298);
nand U6849 (N_6849,N_6028,N_6171);
nand U6850 (N_6850,N_6370,N_6299);
or U6851 (N_6851,N_6047,N_6387);
and U6852 (N_6852,N_6104,N_6285);
and U6853 (N_6853,N_6258,N_6238);
xor U6854 (N_6854,N_6095,N_6122);
nor U6855 (N_6855,N_6029,N_6100);
or U6856 (N_6856,N_6467,N_6365);
nor U6857 (N_6857,N_6259,N_6042);
and U6858 (N_6858,N_6221,N_6385);
nand U6859 (N_6859,N_6492,N_6126);
and U6860 (N_6860,N_6108,N_6352);
nand U6861 (N_6861,N_6440,N_6277);
and U6862 (N_6862,N_6414,N_6375);
nor U6863 (N_6863,N_6370,N_6221);
nand U6864 (N_6864,N_6246,N_6359);
and U6865 (N_6865,N_6195,N_6132);
nand U6866 (N_6866,N_6313,N_6345);
and U6867 (N_6867,N_6209,N_6233);
xnor U6868 (N_6868,N_6435,N_6187);
nand U6869 (N_6869,N_6056,N_6452);
nand U6870 (N_6870,N_6334,N_6425);
xnor U6871 (N_6871,N_6358,N_6223);
nor U6872 (N_6872,N_6277,N_6488);
nor U6873 (N_6873,N_6356,N_6011);
or U6874 (N_6874,N_6227,N_6087);
nand U6875 (N_6875,N_6057,N_6102);
or U6876 (N_6876,N_6394,N_6097);
or U6877 (N_6877,N_6492,N_6312);
or U6878 (N_6878,N_6275,N_6008);
nand U6879 (N_6879,N_6414,N_6355);
nand U6880 (N_6880,N_6335,N_6128);
and U6881 (N_6881,N_6308,N_6298);
and U6882 (N_6882,N_6040,N_6266);
nand U6883 (N_6883,N_6215,N_6101);
and U6884 (N_6884,N_6323,N_6217);
nand U6885 (N_6885,N_6040,N_6076);
xor U6886 (N_6886,N_6048,N_6208);
nand U6887 (N_6887,N_6170,N_6352);
nand U6888 (N_6888,N_6313,N_6416);
xor U6889 (N_6889,N_6362,N_6178);
or U6890 (N_6890,N_6285,N_6346);
or U6891 (N_6891,N_6296,N_6442);
or U6892 (N_6892,N_6423,N_6249);
nand U6893 (N_6893,N_6368,N_6476);
nor U6894 (N_6894,N_6201,N_6479);
xnor U6895 (N_6895,N_6391,N_6412);
nand U6896 (N_6896,N_6288,N_6295);
or U6897 (N_6897,N_6057,N_6278);
or U6898 (N_6898,N_6109,N_6190);
and U6899 (N_6899,N_6269,N_6260);
or U6900 (N_6900,N_6264,N_6058);
and U6901 (N_6901,N_6499,N_6353);
and U6902 (N_6902,N_6205,N_6079);
or U6903 (N_6903,N_6233,N_6184);
nand U6904 (N_6904,N_6334,N_6187);
nand U6905 (N_6905,N_6233,N_6030);
nor U6906 (N_6906,N_6002,N_6042);
nor U6907 (N_6907,N_6177,N_6489);
nand U6908 (N_6908,N_6165,N_6249);
nand U6909 (N_6909,N_6428,N_6230);
nor U6910 (N_6910,N_6249,N_6267);
or U6911 (N_6911,N_6129,N_6423);
xnor U6912 (N_6912,N_6406,N_6281);
or U6913 (N_6913,N_6162,N_6088);
nor U6914 (N_6914,N_6028,N_6376);
and U6915 (N_6915,N_6015,N_6311);
nor U6916 (N_6916,N_6397,N_6362);
and U6917 (N_6917,N_6142,N_6297);
and U6918 (N_6918,N_6425,N_6406);
or U6919 (N_6919,N_6013,N_6107);
xor U6920 (N_6920,N_6459,N_6480);
or U6921 (N_6921,N_6236,N_6311);
xor U6922 (N_6922,N_6389,N_6003);
nor U6923 (N_6923,N_6403,N_6475);
xor U6924 (N_6924,N_6294,N_6495);
nand U6925 (N_6925,N_6450,N_6370);
or U6926 (N_6926,N_6316,N_6396);
and U6927 (N_6927,N_6422,N_6411);
and U6928 (N_6928,N_6335,N_6389);
xor U6929 (N_6929,N_6368,N_6271);
nand U6930 (N_6930,N_6031,N_6111);
or U6931 (N_6931,N_6275,N_6373);
or U6932 (N_6932,N_6451,N_6234);
or U6933 (N_6933,N_6321,N_6376);
nand U6934 (N_6934,N_6244,N_6041);
and U6935 (N_6935,N_6287,N_6337);
nor U6936 (N_6936,N_6204,N_6123);
nand U6937 (N_6937,N_6131,N_6490);
nor U6938 (N_6938,N_6484,N_6444);
nor U6939 (N_6939,N_6246,N_6085);
and U6940 (N_6940,N_6303,N_6292);
nor U6941 (N_6941,N_6354,N_6043);
and U6942 (N_6942,N_6123,N_6011);
and U6943 (N_6943,N_6147,N_6320);
nor U6944 (N_6944,N_6031,N_6291);
or U6945 (N_6945,N_6150,N_6452);
nand U6946 (N_6946,N_6331,N_6269);
nor U6947 (N_6947,N_6015,N_6013);
nand U6948 (N_6948,N_6124,N_6451);
and U6949 (N_6949,N_6331,N_6192);
nand U6950 (N_6950,N_6290,N_6356);
and U6951 (N_6951,N_6428,N_6204);
or U6952 (N_6952,N_6426,N_6180);
or U6953 (N_6953,N_6404,N_6014);
nand U6954 (N_6954,N_6077,N_6048);
or U6955 (N_6955,N_6010,N_6365);
xnor U6956 (N_6956,N_6158,N_6374);
or U6957 (N_6957,N_6393,N_6009);
or U6958 (N_6958,N_6391,N_6419);
and U6959 (N_6959,N_6103,N_6112);
nor U6960 (N_6960,N_6184,N_6064);
and U6961 (N_6961,N_6016,N_6133);
or U6962 (N_6962,N_6310,N_6285);
or U6963 (N_6963,N_6100,N_6211);
or U6964 (N_6964,N_6235,N_6243);
xor U6965 (N_6965,N_6365,N_6300);
or U6966 (N_6966,N_6004,N_6232);
or U6967 (N_6967,N_6435,N_6047);
and U6968 (N_6968,N_6265,N_6471);
or U6969 (N_6969,N_6467,N_6318);
nand U6970 (N_6970,N_6353,N_6345);
nand U6971 (N_6971,N_6288,N_6237);
and U6972 (N_6972,N_6324,N_6200);
nand U6973 (N_6973,N_6418,N_6028);
and U6974 (N_6974,N_6325,N_6261);
or U6975 (N_6975,N_6480,N_6118);
nor U6976 (N_6976,N_6156,N_6057);
or U6977 (N_6977,N_6252,N_6054);
nor U6978 (N_6978,N_6251,N_6346);
or U6979 (N_6979,N_6276,N_6312);
nand U6980 (N_6980,N_6240,N_6045);
or U6981 (N_6981,N_6116,N_6482);
and U6982 (N_6982,N_6272,N_6172);
nor U6983 (N_6983,N_6425,N_6391);
nand U6984 (N_6984,N_6340,N_6324);
xor U6985 (N_6985,N_6159,N_6484);
nor U6986 (N_6986,N_6022,N_6263);
nor U6987 (N_6987,N_6031,N_6176);
or U6988 (N_6988,N_6266,N_6386);
and U6989 (N_6989,N_6409,N_6073);
or U6990 (N_6990,N_6236,N_6133);
and U6991 (N_6991,N_6094,N_6259);
nand U6992 (N_6992,N_6365,N_6247);
nand U6993 (N_6993,N_6240,N_6082);
and U6994 (N_6994,N_6413,N_6039);
or U6995 (N_6995,N_6319,N_6160);
nor U6996 (N_6996,N_6293,N_6376);
xor U6997 (N_6997,N_6206,N_6192);
nor U6998 (N_6998,N_6205,N_6029);
nand U6999 (N_6999,N_6374,N_6469);
and U7000 (N_7000,N_6666,N_6676);
and U7001 (N_7001,N_6521,N_6974);
or U7002 (N_7002,N_6683,N_6819);
and U7003 (N_7003,N_6868,N_6716);
and U7004 (N_7004,N_6873,N_6708);
nand U7005 (N_7005,N_6580,N_6553);
xor U7006 (N_7006,N_6620,N_6972);
nor U7007 (N_7007,N_6679,N_6769);
or U7008 (N_7008,N_6557,N_6951);
nor U7009 (N_7009,N_6513,N_6907);
nor U7010 (N_7010,N_6969,N_6647);
and U7011 (N_7011,N_6793,N_6639);
nand U7012 (N_7012,N_6859,N_6688);
xnor U7013 (N_7013,N_6977,N_6667);
and U7014 (N_7014,N_6815,N_6837);
nor U7015 (N_7015,N_6656,N_6644);
and U7016 (N_7016,N_6905,N_6777);
xor U7017 (N_7017,N_6735,N_6697);
nor U7018 (N_7018,N_6502,N_6635);
nor U7019 (N_7019,N_6511,N_6600);
nor U7020 (N_7020,N_6918,N_6773);
xor U7021 (N_7021,N_6887,N_6929);
and U7022 (N_7022,N_6914,N_6806);
nand U7023 (N_7023,N_6698,N_6678);
xor U7024 (N_7024,N_6570,N_6724);
and U7025 (N_7025,N_6573,N_6725);
xor U7026 (N_7026,N_6751,N_6663);
nand U7027 (N_7027,N_6942,N_6799);
xor U7028 (N_7028,N_6541,N_6804);
and U7029 (N_7029,N_6925,N_6935);
or U7030 (N_7030,N_6991,N_6601);
or U7031 (N_7031,N_6911,N_6847);
or U7032 (N_7032,N_6934,N_6944);
and U7033 (N_7033,N_6693,N_6810);
or U7034 (N_7034,N_6870,N_6596);
xnor U7035 (N_7035,N_6861,N_6715);
nand U7036 (N_7036,N_6850,N_6864);
or U7037 (N_7037,N_6558,N_6758);
nor U7038 (N_7038,N_6984,N_6955);
nor U7039 (N_7039,N_6783,N_6665);
nand U7040 (N_7040,N_6782,N_6875);
and U7041 (N_7041,N_6794,N_6652);
nor U7042 (N_7042,N_6808,N_6909);
nand U7043 (N_7043,N_6771,N_6625);
nor U7044 (N_7044,N_6996,N_6768);
and U7045 (N_7045,N_6894,N_6638);
or U7046 (N_7046,N_6571,N_6577);
and U7047 (N_7047,N_6956,N_6877);
nand U7048 (N_7048,N_6726,N_6568);
nor U7049 (N_7049,N_6714,N_6817);
nor U7050 (N_7050,N_6843,N_6787);
or U7051 (N_7051,N_6841,N_6752);
nand U7052 (N_7052,N_6637,N_6921);
or U7053 (N_7053,N_6954,N_6985);
and U7054 (N_7054,N_6976,N_6582);
nand U7055 (N_7055,N_6805,N_6655);
or U7056 (N_7056,N_6785,N_6889);
or U7057 (N_7057,N_6871,N_6506);
and U7058 (N_7058,N_6610,N_6757);
nand U7059 (N_7059,N_6775,N_6917);
and U7060 (N_7060,N_6973,N_6534);
or U7061 (N_7061,N_6630,N_6755);
nor U7062 (N_7062,N_6618,N_6611);
nor U7063 (N_7063,N_6992,N_6556);
and U7064 (N_7064,N_6705,N_6807);
and U7065 (N_7065,N_6500,N_6711);
nor U7066 (N_7066,N_6723,N_6613);
or U7067 (N_7067,N_6649,N_6776);
nor U7068 (N_7068,N_6988,N_6765);
nand U7069 (N_7069,N_6950,N_6626);
or U7070 (N_7070,N_6772,N_6525);
and U7071 (N_7071,N_6707,N_6795);
and U7072 (N_7072,N_6827,N_6659);
nor U7073 (N_7073,N_6884,N_6961);
nand U7074 (N_7074,N_6614,N_6890);
or U7075 (N_7075,N_6750,N_6970);
xnor U7076 (N_7076,N_6981,N_6798);
nor U7077 (N_7077,N_6510,N_6661);
or U7078 (N_7078,N_6651,N_6615);
and U7079 (N_7079,N_6619,N_6780);
nand U7080 (N_7080,N_6763,N_6906);
nor U7081 (N_7081,N_6801,N_6575);
and U7082 (N_7082,N_6704,N_6701);
nor U7083 (N_7083,N_6535,N_6504);
and U7084 (N_7084,N_6590,N_6749);
nand U7085 (N_7085,N_6941,N_6860);
and U7086 (N_7086,N_6999,N_6857);
nor U7087 (N_7087,N_6529,N_6733);
and U7088 (N_7088,N_6963,N_6813);
and U7089 (N_7089,N_6778,N_6531);
xor U7090 (N_7090,N_6928,N_6910);
nor U7091 (N_7091,N_6943,N_6975);
nor U7092 (N_7092,N_6717,N_6824);
nand U7093 (N_7093,N_6881,N_6930);
and U7094 (N_7094,N_6731,N_6902);
or U7095 (N_7095,N_6931,N_6933);
nor U7096 (N_7096,N_6703,N_6628);
or U7097 (N_7097,N_6826,N_6527);
nand U7098 (N_7098,N_6567,N_6998);
nor U7099 (N_7099,N_6560,N_6669);
nand U7100 (N_7100,N_6713,N_6672);
nor U7101 (N_7101,N_6603,N_6836);
nor U7102 (N_7102,N_6722,N_6839);
nand U7103 (N_7103,N_6712,N_6702);
and U7104 (N_7104,N_6642,N_6846);
nand U7105 (N_7105,N_6770,N_6737);
and U7106 (N_7106,N_6788,N_6899);
or U7107 (N_7107,N_6888,N_6501);
and U7108 (N_7108,N_6822,N_6640);
or U7109 (N_7109,N_6736,N_6605);
and U7110 (N_7110,N_6938,N_6866);
nor U7111 (N_7111,N_6767,N_6515);
and U7112 (N_7112,N_6754,N_6650);
nor U7113 (N_7113,N_6882,N_6878);
xnor U7114 (N_7114,N_6689,N_6551);
or U7115 (N_7115,N_6690,N_6842);
or U7116 (N_7116,N_6654,N_6953);
nor U7117 (N_7117,N_6588,N_6893);
nor U7118 (N_7118,N_6790,N_6591);
and U7119 (N_7119,N_6563,N_6585);
and U7120 (N_7120,N_6609,N_6592);
or U7121 (N_7121,N_6595,N_6677);
nor U7122 (N_7122,N_6812,N_6830);
nor U7123 (N_7123,N_6604,N_6616);
nand U7124 (N_7124,N_6766,N_6645);
nor U7125 (N_7125,N_6668,N_6743);
or U7126 (N_7126,N_6990,N_6569);
nand U7127 (N_7127,N_6718,N_6634);
and U7128 (N_7128,N_6948,N_6900);
nor U7129 (N_7129,N_6648,N_6700);
and U7130 (N_7130,N_6526,N_6838);
and U7131 (N_7131,N_6781,N_6680);
or U7132 (N_7132,N_6895,N_6566);
or U7133 (N_7133,N_6612,N_6550);
nand U7134 (N_7134,N_6811,N_6710);
and U7135 (N_7135,N_6823,N_6641);
or U7136 (N_7136,N_6989,N_6740);
xnor U7137 (N_7137,N_6623,N_6892);
or U7138 (N_7138,N_6599,N_6548);
nand U7139 (N_7139,N_6853,N_6832);
xnor U7140 (N_7140,N_6920,N_6682);
and U7141 (N_7141,N_6997,N_6624);
or U7142 (N_7142,N_6865,N_6512);
or U7143 (N_7143,N_6919,N_6959);
nand U7144 (N_7144,N_6851,N_6574);
and U7145 (N_7145,N_6968,N_6741);
nand U7146 (N_7146,N_6524,N_6980);
or U7147 (N_7147,N_6995,N_6744);
nand U7148 (N_7148,N_6940,N_6987);
and U7149 (N_7149,N_6730,N_6589);
nand U7150 (N_7150,N_6924,N_6786);
and U7151 (N_7151,N_6897,N_6802);
nand U7152 (N_7152,N_6622,N_6664);
or U7153 (N_7153,N_6728,N_6848);
xnor U7154 (N_7154,N_6945,N_6994);
and U7155 (N_7155,N_6721,N_6519);
or U7156 (N_7156,N_6518,N_6932);
nand U7157 (N_7157,N_6631,N_6507);
nand U7158 (N_7158,N_6742,N_6581);
or U7159 (N_7159,N_6694,N_6530);
nand U7160 (N_7160,N_6686,N_6957);
or U7161 (N_7161,N_6632,N_6863);
and U7162 (N_7162,N_6692,N_6901);
xor U7163 (N_7163,N_6579,N_6818);
or U7164 (N_7164,N_6936,N_6503);
or U7165 (N_7165,N_6979,N_6761);
nand U7166 (N_7166,N_6947,N_6774);
and U7167 (N_7167,N_6709,N_6898);
and U7168 (N_7168,N_6546,N_6727);
or U7169 (N_7169,N_6593,N_6699);
and U7170 (N_7170,N_6797,N_6674);
or U7171 (N_7171,N_6879,N_6662);
nor U7172 (N_7172,N_6520,N_6965);
nand U7173 (N_7173,N_6695,N_6578);
or U7174 (N_7174,N_6671,N_6814);
nand U7175 (N_7175,N_6880,N_6594);
nand U7176 (N_7176,N_6544,N_6937);
nand U7177 (N_7177,N_6739,N_6952);
nand U7178 (N_7178,N_6572,N_6633);
nand U7179 (N_7179,N_6886,N_6653);
or U7180 (N_7180,N_6966,N_6779);
nand U7181 (N_7181,N_6516,N_6913);
xor U7182 (N_7182,N_6791,N_6816);
and U7183 (N_7183,N_6833,N_6675);
or U7184 (N_7184,N_6636,N_6927);
nor U7185 (N_7185,N_6896,N_6753);
and U7186 (N_7186,N_6658,N_6684);
nand U7187 (N_7187,N_6762,N_6554);
and U7188 (N_7188,N_6908,N_6982);
and U7189 (N_7189,N_6706,N_6584);
nand U7190 (N_7190,N_6845,N_6852);
and U7191 (N_7191,N_6685,N_6903);
or U7192 (N_7192,N_6809,N_6834);
nor U7193 (N_7193,N_6883,N_6746);
and U7194 (N_7194,N_6681,N_6756);
or U7195 (N_7195,N_6643,N_6967);
nand U7196 (N_7196,N_6646,N_6922);
or U7197 (N_7197,N_6803,N_6508);
xor U7198 (N_7198,N_6586,N_6583);
and U7199 (N_7199,N_6876,N_6912);
or U7200 (N_7200,N_6732,N_6738);
xnor U7201 (N_7201,N_6627,N_6617);
nor U7202 (N_7202,N_6960,N_6598);
nor U7203 (N_7203,N_6854,N_6862);
nand U7204 (N_7204,N_6673,N_6559);
nand U7205 (N_7205,N_6719,N_6720);
nand U7206 (N_7206,N_6829,N_6687);
nand U7207 (N_7207,N_6607,N_6986);
nor U7208 (N_7208,N_6536,N_6562);
nor U7209 (N_7209,N_6792,N_6858);
nor U7210 (N_7210,N_6835,N_6691);
and U7211 (N_7211,N_6542,N_6840);
or U7212 (N_7212,N_6891,N_6856);
nor U7213 (N_7213,N_6747,N_6971);
and U7214 (N_7214,N_6885,N_6545);
nor U7215 (N_7215,N_6825,N_6514);
nor U7216 (N_7216,N_6796,N_6855);
or U7217 (N_7217,N_6820,N_6555);
or U7218 (N_7218,N_6962,N_6949);
nor U7219 (N_7219,N_6946,N_6734);
and U7220 (N_7220,N_6547,N_6745);
or U7221 (N_7221,N_6533,N_6764);
xnor U7222 (N_7222,N_6505,N_6759);
or U7223 (N_7223,N_6602,N_6849);
and U7224 (N_7224,N_6509,N_6964);
nor U7225 (N_7225,N_6789,N_6760);
and U7226 (N_7226,N_6748,N_6537);
nor U7227 (N_7227,N_6587,N_6844);
or U7228 (N_7228,N_6552,N_6978);
nor U7229 (N_7229,N_6784,N_6821);
nand U7230 (N_7230,N_6597,N_6915);
nand U7231 (N_7231,N_6540,N_6621);
nor U7232 (N_7232,N_6869,N_6670);
nand U7233 (N_7233,N_6872,N_6993);
nand U7234 (N_7234,N_6729,N_6528);
nand U7235 (N_7235,N_6958,N_6874);
and U7236 (N_7236,N_6926,N_6983);
nor U7237 (N_7237,N_6543,N_6660);
nand U7238 (N_7238,N_6522,N_6608);
and U7239 (N_7239,N_6904,N_6576);
and U7240 (N_7240,N_6564,N_6696);
nor U7241 (N_7241,N_6561,N_6916);
nor U7242 (N_7242,N_6538,N_6800);
xor U7243 (N_7243,N_6828,N_6629);
and U7244 (N_7244,N_6539,N_6549);
or U7245 (N_7245,N_6565,N_6939);
xnor U7246 (N_7246,N_6606,N_6657);
nand U7247 (N_7247,N_6867,N_6532);
nor U7248 (N_7248,N_6831,N_6517);
xor U7249 (N_7249,N_6523,N_6923);
and U7250 (N_7250,N_6560,N_6751);
nor U7251 (N_7251,N_6855,N_6748);
or U7252 (N_7252,N_6838,N_6943);
nand U7253 (N_7253,N_6766,N_6937);
or U7254 (N_7254,N_6863,N_6667);
or U7255 (N_7255,N_6990,N_6884);
or U7256 (N_7256,N_6952,N_6893);
nand U7257 (N_7257,N_6963,N_6953);
nand U7258 (N_7258,N_6765,N_6956);
or U7259 (N_7259,N_6531,N_6873);
and U7260 (N_7260,N_6640,N_6860);
xnor U7261 (N_7261,N_6705,N_6797);
and U7262 (N_7262,N_6674,N_6911);
nand U7263 (N_7263,N_6892,N_6799);
and U7264 (N_7264,N_6800,N_6747);
and U7265 (N_7265,N_6916,N_6922);
and U7266 (N_7266,N_6654,N_6731);
or U7267 (N_7267,N_6776,N_6757);
nor U7268 (N_7268,N_6880,N_6578);
nor U7269 (N_7269,N_6800,N_6861);
and U7270 (N_7270,N_6740,N_6899);
nor U7271 (N_7271,N_6865,N_6809);
and U7272 (N_7272,N_6673,N_6935);
or U7273 (N_7273,N_6732,N_6670);
xnor U7274 (N_7274,N_6879,N_6726);
nand U7275 (N_7275,N_6907,N_6592);
nor U7276 (N_7276,N_6654,N_6544);
nor U7277 (N_7277,N_6505,N_6646);
and U7278 (N_7278,N_6882,N_6810);
nor U7279 (N_7279,N_6520,N_6977);
and U7280 (N_7280,N_6667,N_6594);
nand U7281 (N_7281,N_6710,N_6558);
xnor U7282 (N_7282,N_6804,N_6858);
nor U7283 (N_7283,N_6798,N_6939);
nand U7284 (N_7284,N_6682,N_6718);
or U7285 (N_7285,N_6856,N_6987);
nor U7286 (N_7286,N_6663,N_6946);
nand U7287 (N_7287,N_6843,N_6976);
and U7288 (N_7288,N_6590,N_6846);
and U7289 (N_7289,N_6884,N_6970);
nor U7290 (N_7290,N_6521,N_6517);
and U7291 (N_7291,N_6654,N_6843);
and U7292 (N_7292,N_6695,N_6551);
nand U7293 (N_7293,N_6623,N_6585);
nor U7294 (N_7294,N_6900,N_6895);
nand U7295 (N_7295,N_6937,N_6684);
nand U7296 (N_7296,N_6880,N_6617);
nor U7297 (N_7297,N_6862,N_6974);
nor U7298 (N_7298,N_6964,N_6995);
or U7299 (N_7299,N_6704,N_6714);
and U7300 (N_7300,N_6648,N_6802);
nor U7301 (N_7301,N_6898,N_6931);
nor U7302 (N_7302,N_6601,N_6560);
nand U7303 (N_7303,N_6922,N_6628);
nor U7304 (N_7304,N_6850,N_6799);
nor U7305 (N_7305,N_6746,N_6945);
nand U7306 (N_7306,N_6727,N_6998);
or U7307 (N_7307,N_6763,N_6869);
nand U7308 (N_7308,N_6735,N_6874);
and U7309 (N_7309,N_6949,N_6710);
xnor U7310 (N_7310,N_6833,N_6679);
nor U7311 (N_7311,N_6714,N_6870);
or U7312 (N_7312,N_6619,N_6997);
xor U7313 (N_7313,N_6543,N_6985);
and U7314 (N_7314,N_6970,N_6856);
and U7315 (N_7315,N_6685,N_6855);
or U7316 (N_7316,N_6831,N_6923);
nand U7317 (N_7317,N_6807,N_6522);
nand U7318 (N_7318,N_6590,N_6508);
and U7319 (N_7319,N_6818,N_6749);
and U7320 (N_7320,N_6904,N_6866);
or U7321 (N_7321,N_6782,N_6736);
and U7322 (N_7322,N_6624,N_6991);
or U7323 (N_7323,N_6668,N_6874);
and U7324 (N_7324,N_6867,N_6626);
or U7325 (N_7325,N_6545,N_6659);
or U7326 (N_7326,N_6665,N_6987);
and U7327 (N_7327,N_6997,N_6846);
nand U7328 (N_7328,N_6733,N_6860);
nor U7329 (N_7329,N_6656,N_6786);
nand U7330 (N_7330,N_6835,N_6765);
nor U7331 (N_7331,N_6567,N_6760);
nand U7332 (N_7332,N_6658,N_6926);
nor U7333 (N_7333,N_6615,N_6785);
and U7334 (N_7334,N_6796,N_6614);
nand U7335 (N_7335,N_6721,N_6826);
or U7336 (N_7336,N_6910,N_6620);
and U7337 (N_7337,N_6708,N_6758);
or U7338 (N_7338,N_6724,N_6642);
and U7339 (N_7339,N_6630,N_6639);
or U7340 (N_7340,N_6712,N_6812);
nand U7341 (N_7341,N_6721,N_6681);
nor U7342 (N_7342,N_6711,N_6772);
nor U7343 (N_7343,N_6608,N_6865);
xnor U7344 (N_7344,N_6585,N_6747);
and U7345 (N_7345,N_6970,N_6555);
nor U7346 (N_7346,N_6874,N_6771);
or U7347 (N_7347,N_6505,N_6589);
nand U7348 (N_7348,N_6524,N_6751);
or U7349 (N_7349,N_6671,N_6820);
or U7350 (N_7350,N_6949,N_6570);
or U7351 (N_7351,N_6956,N_6579);
nor U7352 (N_7352,N_6933,N_6942);
and U7353 (N_7353,N_6921,N_6928);
nor U7354 (N_7354,N_6600,N_6577);
nor U7355 (N_7355,N_6510,N_6893);
nor U7356 (N_7356,N_6716,N_6832);
nor U7357 (N_7357,N_6586,N_6934);
nor U7358 (N_7358,N_6810,N_6943);
or U7359 (N_7359,N_6922,N_6948);
xor U7360 (N_7360,N_6839,N_6510);
nand U7361 (N_7361,N_6535,N_6935);
and U7362 (N_7362,N_6972,N_6833);
nor U7363 (N_7363,N_6949,N_6953);
and U7364 (N_7364,N_6516,N_6951);
nor U7365 (N_7365,N_6976,N_6990);
xnor U7366 (N_7366,N_6691,N_6861);
or U7367 (N_7367,N_6981,N_6946);
or U7368 (N_7368,N_6912,N_6616);
and U7369 (N_7369,N_6514,N_6505);
nand U7370 (N_7370,N_6663,N_6576);
nor U7371 (N_7371,N_6511,N_6641);
xnor U7372 (N_7372,N_6882,N_6692);
and U7373 (N_7373,N_6871,N_6744);
and U7374 (N_7374,N_6709,N_6997);
nor U7375 (N_7375,N_6895,N_6593);
nor U7376 (N_7376,N_6924,N_6553);
and U7377 (N_7377,N_6638,N_6535);
or U7378 (N_7378,N_6741,N_6643);
or U7379 (N_7379,N_6631,N_6878);
and U7380 (N_7380,N_6540,N_6554);
xor U7381 (N_7381,N_6725,N_6783);
and U7382 (N_7382,N_6819,N_6563);
or U7383 (N_7383,N_6630,N_6681);
xnor U7384 (N_7384,N_6711,N_6530);
nor U7385 (N_7385,N_6579,N_6743);
xor U7386 (N_7386,N_6883,N_6890);
or U7387 (N_7387,N_6860,N_6853);
nand U7388 (N_7388,N_6694,N_6910);
and U7389 (N_7389,N_6716,N_6690);
and U7390 (N_7390,N_6702,N_6819);
or U7391 (N_7391,N_6504,N_6766);
nand U7392 (N_7392,N_6687,N_6925);
xnor U7393 (N_7393,N_6777,N_6719);
and U7394 (N_7394,N_6688,N_6904);
nand U7395 (N_7395,N_6670,N_6824);
and U7396 (N_7396,N_6946,N_6972);
and U7397 (N_7397,N_6687,N_6767);
or U7398 (N_7398,N_6901,N_6971);
nand U7399 (N_7399,N_6523,N_6778);
nand U7400 (N_7400,N_6956,N_6605);
nor U7401 (N_7401,N_6536,N_6864);
nor U7402 (N_7402,N_6917,N_6790);
nand U7403 (N_7403,N_6992,N_6903);
and U7404 (N_7404,N_6827,N_6800);
xnor U7405 (N_7405,N_6984,N_6518);
nand U7406 (N_7406,N_6527,N_6816);
nor U7407 (N_7407,N_6756,N_6835);
or U7408 (N_7408,N_6950,N_6671);
nor U7409 (N_7409,N_6748,N_6862);
nand U7410 (N_7410,N_6794,N_6531);
or U7411 (N_7411,N_6590,N_6686);
nand U7412 (N_7412,N_6946,N_6601);
nand U7413 (N_7413,N_6913,N_6812);
or U7414 (N_7414,N_6625,N_6871);
nand U7415 (N_7415,N_6961,N_6756);
nand U7416 (N_7416,N_6872,N_6546);
xor U7417 (N_7417,N_6692,N_6928);
or U7418 (N_7418,N_6536,N_6885);
nand U7419 (N_7419,N_6795,N_6746);
nand U7420 (N_7420,N_6758,N_6836);
and U7421 (N_7421,N_6901,N_6874);
nor U7422 (N_7422,N_6572,N_6509);
nand U7423 (N_7423,N_6814,N_6754);
and U7424 (N_7424,N_6939,N_6550);
nor U7425 (N_7425,N_6667,N_6591);
and U7426 (N_7426,N_6622,N_6768);
nor U7427 (N_7427,N_6586,N_6693);
nor U7428 (N_7428,N_6662,N_6833);
or U7429 (N_7429,N_6545,N_6944);
and U7430 (N_7430,N_6942,N_6605);
xnor U7431 (N_7431,N_6931,N_6648);
or U7432 (N_7432,N_6817,N_6801);
and U7433 (N_7433,N_6700,N_6995);
nand U7434 (N_7434,N_6644,N_6654);
or U7435 (N_7435,N_6619,N_6513);
xnor U7436 (N_7436,N_6974,N_6729);
or U7437 (N_7437,N_6818,N_6539);
nand U7438 (N_7438,N_6708,N_6968);
nor U7439 (N_7439,N_6841,N_6825);
nand U7440 (N_7440,N_6642,N_6703);
nor U7441 (N_7441,N_6511,N_6796);
and U7442 (N_7442,N_6823,N_6972);
or U7443 (N_7443,N_6528,N_6657);
nor U7444 (N_7444,N_6684,N_6600);
and U7445 (N_7445,N_6766,N_6722);
and U7446 (N_7446,N_6632,N_6825);
nand U7447 (N_7447,N_6640,N_6654);
nor U7448 (N_7448,N_6730,N_6902);
nor U7449 (N_7449,N_6804,N_6892);
nand U7450 (N_7450,N_6843,N_6523);
or U7451 (N_7451,N_6900,N_6647);
or U7452 (N_7452,N_6900,N_6651);
xnor U7453 (N_7453,N_6690,N_6633);
and U7454 (N_7454,N_6901,N_6818);
nand U7455 (N_7455,N_6783,N_6515);
and U7456 (N_7456,N_6739,N_6809);
nor U7457 (N_7457,N_6781,N_6771);
nor U7458 (N_7458,N_6857,N_6927);
xor U7459 (N_7459,N_6926,N_6949);
and U7460 (N_7460,N_6949,N_6637);
and U7461 (N_7461,N_6995,N_6529);
nor U7462 (N_7462,N_6764,N_6501);
xnor U7463 (N_7463,N_6772,N_6983);
nor U7464 (N_7464,N_6746,N_6825);
nand U7465 (N_7465,N_6599,N_6960);
nor U7466 (N_7466,N_6997,N_6751);
or U7467 (N_7467,N_6711,N_6790);
nand U7468 (N_7468,N_6710,N_6722);
nor U7469 (N_7469,N_6633,N_6915);
or U7470 (N_7470,N_6594,N_6761);
nand U7471 (N_7471,N_6645,N_6713);
nand U7472 (N_7472,N_6967,N_6934);
xnor U7473 (N_7473,N_6554,N_6950);
or U7474 (N_7474,N_6571,N_6582);
and U7475 (N_7475,N_6952,N_6691);
and U7476 (N_7476,N_6650,N_6787);
nor U7477 (N_7477,N_6769,N_6826);
nor U7478 (N_7478,N_6855,N_6988);
and U7479 (N_7479,N_6966,N_6578);
and U7480 (N_7480,N_6566,N_6732);
nor U7481 (N_7481,N_6709,N_6918);
or U7482 (N_7482,N_6753,N_6575);
or U7483 (N_7483,N_6991,N_6949);
and U7484 (N_7484,N_6770,N_6708);
nand U7485 (N_7485,N_6864,N_6503);
nor U7486 (N_7486,N_6945,N_6583);
and U7487 (N_7487,N_6979,N_6744);
nor U7488 (N_7488,N_6930,N_6531);
and U7489 (N_7489,N_6955,N_6594);
nand U7490 (N_7490,N_6772,N_6980);
nor U7491 (N_7491,N_6527,N_6605);
nor U7492 (N_7492,N_6978,N_6622);
nand U7493 (N_7493,N_6681,N_6916);
nor U7494 (N_7494,N_6829,N_6790);
or U7495 (N_7495,N_6828,N_6511);
or U7496 (N_7496,N_6985,N_6547);
or U7497 (N_7497,N_6548,N_6542);
and U7498 (N_7498,N_6895,N_6921);
nor U7499 (N_7499,N_6818,N_6957);
nand U7500 (N_7500,N_7423,N_7165);
and U7501 (N_7501,N_7109,N_7075);
and U7502 (N_7502,N_7212,N_7311);
nor U7503 (N_7503,N_7187,N_7202);
or U7504 (N_7504,N_7105,N_7484);
nand U7505 (N_7505,N_7067,N_7370);
and U7506 (N_7506,N_7084,N_7376);
nand U7507 (N_7507,N_7314,N_7008);
nor U7508 (N_7508,N_7498,N_7272);
nand U7509 (N_7509,N_7375,N_7141);
and U7510 (N_7510,N_7255,N_7177);
or U7511 (N_7511,N_7443,N_7065);
nand U7512 (N_7512,N_7028,N_7249);
nor U7513 (N_7513,N_7230,N_7362);
or U7514 (N_7514,N_7137,N_7303);
and U7515 (N_7515,N_7466,N_7035);
nand U7516 (N_7516,N_7167,N_7422);
nand U7517 (N_7517,N_7124,N_7479);
nor U7518 (N_7518,N_7203,N_7300);
and U7519 (N_7519,N_7435,N_7321);
or U7520 (N_7520,N_7259,N_7106);
xnor U7521 (N_7521,N_7011,N_7493);
and U7522 (N_7522,N_7049,N_7308);
or U7523 (N_7523,N_7029,N_7357);
nand U7524 (N_7524,N_7407,N_7116);
nand U7525 (N_7525,N_7061,N_7318);
nand U7526 (N_7526,N_7434,N_7379);
nor U7527 (N_7527,N_7487,N_7398);
nand U7528 (N_7528,N_7283,N_7056);
and U7529 (N_7529,N_7309,N_7485);
or U7530 (N_7530,N_7140,N_7437);
or U7531 (N_7531,N_7339,N_7333);
nor U7532 (N_7532,N_7136,N_7334);
and U7533 (N_7533,N_7150,N_7051);
and U7534 (N_7534,N_7367,N_7256);
and U7535 (N_7535,N_7468,N_7054);
nor U7536 (N_7536,N_7316,N_7144);
and U7537 (N_7537,N_7342,N_7095);
or U7538 (N_7538,N_7151,N_7260);
and U7539 (N_7539,N_7343,N_7129);
and U7540 (N_7540,N_7415,N_7097);
nand U7541 (N_7541,N_7414,N_7023);
and U7542 (N_7542,N_7385,N_7472);
or U7543 (N_7543,N_7459,N_7228);
or U7544 (N_7544,N_7045,N_7350);
nand U7545 (N_7545,N_7178,N_7440);
nand U7546 (N_7546,N_7491,N_7015);
or U7547 (N_7547,N_7231,N_7469);
xnor U7548 (N_7548,N_7489,N_7436);
and U7549 (N_7549,N_7041,N_7274);
and U7550 (N_7550,N_7326,N_7232);
or U7551 (N_7551,N_7060,N_7224);
nand U7552 (N_7552,N_7133,N_7306);
or U7553 (N_7553,N_7025,N_7410);
and U7554 (N_7554,N_7413,N_7372);
xnor U7555 (N_7555,N_7176,N_7315);
nor U7556 (N_7556,N_7009,N_7438);
nor U7557 (N_7557,N_7252,N_7233);
nor U7558 (N_7558,N_7348,N_7180);
and U7559 (N_7559,N_7155,N_7445);
or U7560 (N_7560,N_7001,N_7000);
nor U7561 (N_7561,N_7142,N_7301);
nand U7562 (N_7562,N_7477,N_7210);
nand U7563 (N_7563,N_7014,N_7125);
and U7564 (N_7564,N_7346,N_7033);
and U7565 (N_7565,N_7206,N_7366);
and U7566 (N_7566,N_7092,N_7122);
nor U7567 (N_7567,N_7263,N_7130);
nand U7568 (N_7568,N_7239,N_7475);
nor U7569 (N_7569,N_7026,N_7152);
nor U7570 (N_7570,N_7193,N_7369);
and U7571 (N_7571,N_7264,N_7052);
nand U7572 (N_7572,N_7280,N_7388);
and U7573 (N_7573,N_7139,N_7036);
nand U7574 (N_7574,N_7499,N_7042);
xor U7575 (N_7575,N_7135,N_7361);
nand U7576 (N_7576,N_7382,N_7409);
nand U7577 (N_7577,N_7066,N_7039);
and U7578 (N_7578,N_7021,N_7332);
nor U7579 (N_7579,N_7278,N_7148);
and U7580 (N_7580,N_7419,N_7108);
or U7581 (N_7581,N_7229,N_7310);
nor U7582 (N_7582,N_7091,N_7216);
or U7583 (N_7583,N_7380,N_7226);
nand U7584 (N_7584,N_7012,N_7497);
and U7585 (N_7585,N_7329,N_7323);
and U7586 (N_7586,N_7194,N_7374);
nor U7587 (N_7587,N_7243,N_7365);
or U7588 (N_7588,N_7392,N_7044);
or U7589 (N_7589,N_7190,N_7317);
and U7590 (N_7590,N_7421,N_7185);
nand U7591 (N_7591,N_7197,N_7441);
or U7592 (N_7592,N_7294,N_7412);
and U7593 (N_7593,N_7186,N_7387);
and U7594 (N_7594,N_7449,N_7286);
or U7595 (N_7595,N_7034,N_7113);
nand U7596 (N_7596,N_7032,N_7486);
or U7597 (N_7597,N_7099,N_7313);
nand U7598 (N_7598,N_7191,N_7364);
nand U7599 (N_7599,N_7381,N_7452);
xnor U7600 (N_7600,N_7058,N_7320);
and U7601 (N_7601,N_7235,N_7447);
and U7602 (N_7602,N_7209,N_7462);
or U7603 (N_7603,N_7335,N_7480);
nor U7604 (N_7604,N_7397,N_7022);
and U7605 (N_7605,N_7427,N_7166);
nor U7606 (N_7606,N_7199,N_7345);
nand U7607 (N_7607,N_7182,N_7161);
and U7608 (N_7608,N_7083,N_7347);
or U7609 (N_7609,N_7281,N_7006);
or U7610 (N_7610,N_7128,N_7046);
nor U7611 (N_7611,N_7063,N_7244);
and U7612 (N_7612,N_7341,N_7411);
xnor U7613 (N_7613,N_7285,N_7112);
nand U7614 (N_7614,N_7282,N_7302);
or U7615 (N_7615,N_7048,N_7170);
or U7616 (N_7616,N_7296,N_7324);
xor U7617 (N_7617,N_7117,N_7377);
nand U7618 (N_7618,N_7208,N_7246);
nand U7619 (N_7619,N_7100,N_7218);
or U7620 (N_7620,N_7353,N_7400);
and U7621 (N_7621,N_7373,N_7085);
nand U7622 (N_7622,N_7027,N_7196);
and U7623 (N_7623,N_7457,N_7164);
nand U7624 (N_7624,N_7268,N_7456);
nor U7625 (N_7625,N_7240,N_7494);
or U7626 (N_7626,N_7077,N_7204);
nor U7627 (N_7627,N_7325,N_7237);
nor U7628 (N_7628,N_7110,N_7123);
or U7629 (N_7629,N_7336,N_7024);
and U7630 (N_7630,N_7328,N_7401);
nor U7631 (N_7631,N_7262,N_7126);
nor U7632 (N_7632,N_7431,N_7453);
or U7633 (N_7633,N_7312,N_7454);
nor U7634 (N_7634,N_7471,N_7482);
nor U7635 (N_7635,N_7444,N_7173);
nor U7636 (N_7636,N_7064,N_7062);
nor U7637 (N_7637,N_7304,N_7297);
or U7638 (N_7638,N_7481,N_7254);
xnor U7639 (N_7639,N_7169,N_7354);
nor U7640 (N_7640,N_7428,N_7253);
or U7641 (N_7641,N_7340,N_7220);
nand U7642 (N_7642,N_7269,N_7082);
xnor U7643 (N_7643,N_7154,N_7219);
nand U7644 (N_7644,N_7147,N_7448);
nand U7645 (N_7645,N_7120,N_7004);
and U7646 (N_7646,N_7258,N_7030);
nor U7647 (N_7647,N_7352,N_7403);
xor U7648 (N_7648,N_7020,N_7055);
xor U7649 (N_7649,N_7071,N_7093);
nor U7650 (N_7650,N_7390,N_7273);
nand U7651 (N_7651,N_7019,N_7495);
and U7652 (N_7652,N_7201,N_7450);
xnor U7653 (N_7653,N_7211,N_7478);
or U7654 (N_7654,N_7275,N_7118);
nand U7655 (N_7655,N_7426,N_7467);
nor U7656 (N_7656,N_7356,N_7225);
nor U7657 (N_7657,N_7181,N_7163);
and U7658 (N_7658,N_7394,N_7090);
or U7659 (N_7659,N_7132,N_7358);
or U7660 (N_7660,N_7171,N_7250);
xnor U7661 (N_7661,N_7290,N_7496);
nor U7662 (N_7662,N_7406,N_7146);
and U7663 (N_7663,N_7307,N_7102);
nor U7664 (N_7664,N_7221,N_7010);
nand U7665 (N_7665,N_7289,N_7003);
nor U7666 (N_7666,N_7172,N_7198);
and U7667 (N_7667,N_7088,N_7200);
and U7668 (N_7668,N_7408,N_7295);
nand U7669 (N_7669,N_7404,N_7368);
nor U7670 (N_7670,N_7114,N_7384);
nand U7671 (N_7671,N_7465,N_7464);
nand U7672 (N_7672,N_7149,N_7002);
nor U7673 (N_7673,N_7013,N_7293);
or U7674 (N_7674,N_7127,N_7266);
nor U7675 (N_7675,N_7257,N_7395);
or U7676 (N_7676,N_7157,N_7131);
xnor U7677 (N_7677,N_7031,N_7455);
nor U7678 (N_7678,N_7214,N_7270);
xor U7679 (N_7679,N_7396,N_7371);
nand U7680 (N_7680,N_7442,N_7425);
or U7681 (N_7681,N_7305,N_7078);
and U7682 (N_7682,N_7184,N_7446);
nand U7683 (N_7683,N_7276,N_7104);
nor U7684 (N_7684,N_7195,N_7098);
or U7685 (N_7685,N_7183,N_7299);
nand U7686 (N_7686,N_7016,N_7107);
nor U7687 (N_7687,N_7330,N_7038);
or U7688 (N_7688,N_7429,N_7463);
nor U7689 (N_7689,N_7359,N_7086);
or U7690 (N_7690,N_7215,N_7072);
nor U7691 (N_7691,N_7338,N_7069);
and U7692 (N_7692,N_7430,N_7470);
and U7693 (N_7693,N_7057,N_7279);
nor U7694 (N_7694,N_7018,N_7344);
and U7695 (N_7695,N_7292,N_7159);
and U7696 (N_7696,N_7265,N_7089);
nor U7697 (N_7697,N_7433,N_7115);
nand U7698 (N_7698,N_7360,N_7079);
xor U7699 (N_7699,N_7174,N_7162);
nor U7700 (N_7700,N_7134,N_7070);
or U7701 (N_7701,N_7179,N_7068);
nand U7702 (N_7702,N_7416,N_7111);
and U7703 (N_7703,N_7432,N_7399);
or U7704 (N_7704,N_7037,N_7074);
xor U7705 (N_7705,N_7101,N_7420);
nor U7706 (N_7706,N_7322,N_7138);
and U7707 (N_7707,N_7327,N_7005);
or U7708 (N_7708,N_7059,N_7261);
and U7709 (N_7709,N_7461,N_7439);
or U7710 (N_7710,N_7158,N_7050);
or U7711 (N_7711,N_7007,N_7168);
nor U7712 (N_7712,N_7474,N_7145);
and U7713 (N_7713,N_7247,N_7103);
nor U7714 (N_7714,N_7476,N_7405);
nor U7715 (N_7715,N_7492,N_7238);
and U7716 (N_7716,N_7223,N_7188);
nand U7717 (N_7717,N_7017,N_7378);
nand U7718 (N_7718,N_7080,N_7096);
nor U7719 (N_7719,N_7043,N_7241);
and U7720 (N_7720,N_7490,N_7222);
nand U7721 (N_7721,N_7363,N_7153);
nand U7722 (N_7722,N_7242,N_7383);
nor U7723 (N_7723,N_7040,N_7349);
nand U7724 (N_7724,N_7402,N_7291);
nor U7725 (N_7725,N_7473,N_7081);
xnor U7726 (N_7726,N_7391,N_7175);
nor U7727 (N_7727,N_7458,N_7121);
nand U7728 (N_7728,N_7248,N_7298);
or U7729 (N_7729,N_7288,N_7119);
or U7730 (N_7730,N_7386,N_7424);
or U7731 (N_7731,N_7227,N_7251);
nor U7732 (N_7732,N_7418,N_7053);
or U7733 (N_7733,N_7234,N_7483);
xnor U7734 (N_7734,N_7094,N_7417);
and U7735 (N_7735,N_7160,N_7245);
and U7736 (N_7736,N_7267,N_7389);
and U7737 (N_7737,N_7488,N_7076);
xor U7738 (N_7738,N_7073,N_7284);
and U7739 (N_7739,N_7213,N_7277);
or U7740 (N_7740,N_7217,N_7287);
and U7741 (N_7741,N_7156,N_7143);
nor U7742 (N_7742,N_7351,N_7319);
and U7743 (N_7743,N_7087,N_7460);
nor U7744 (N_7744,N_7393,N_7192);
nor U7745 (N_7745,N_7331,N_7355);
xor U7746 (N_7746,N_7047,N_7271);
nor U7747 (N_7747,N_7205,N_7207);
nand U7748 (N_7748,N_7236,N_7337);
nand U7749 (N_7749,N_7189,N_7451);
nand U7750 (N_7750,N_7353,N_7062);
and U7751 (N_7751,N_7448,N_7404);
or U7752 (N_7752,N_7300,N_7216);
or U7753 (N_7753,N_7171,N_7021);
nor U7754 (N_7754,N_7214,N_7324);
nand U7755 (N_7755,N_7401,N_7416);
nor U7756 (N_7756,N_7149,N_7292);
and U7757 (N_7757,N_7035,N_7482);
or U7758 (N_7758,N_7223,N_7368);
nand U7759 (N_7759,N_7180,N_7222);
nand U7760 (N_7760,N_7250,N_7490);
nor U7761 (N_7761,N_7482,N_7276);
or U7762 (N_7762,N_7106,N_7124);
or U7763 (N_7763,N_7221,N_7137);
and U7764 (N_7764,N_7230,N_7451);
or U7765 (N_7765,N_7403,N_7140);
nor U7766 (N_7766,N_7309,N_7102);
or U7767 (N_7767,N_7353,N_7210);
nand U7768 (N_7768,N_7485,N_7227);
or U7769 (N_7769,N_7166,N_7123);
nand U7770 (N_7770,N_7146,N_7467);
and U7771 (N_7771,N_7103,N_7178);
and U7772 (N_7772,N_7100,N_7372);
nand U7773 (N_7773,N_7369,N_7128);
nor U7774 (N_7774,N_7323,N_7104);
nor U7775 (N_7775,N_7481,N_7437);
and U7776 (N_7776,N_7079,N_7172);
xor U7777 (N_7777,N_7160,N_7336);
xnor U7778 (N_7778,N_7103,N_7276);
or U7779 (N_7779,N_7373,N_7031);
nor U7780 (N_7780,N_7420,N_7456);
or U7781 (N_7781,N_7445,N_7416);
xor U7782 (N_7782,N_7114,N_7386);
or U7783 (N_7783,N_7347,N_7020);
nor U7784 (N_7784,N_7300,N_7409);
and U7785 (N_7785,N_7373,N_7076);
nor U7786 (N_7786,N_7187,N_7498);
and U7787 (N_7787,N_7200,N_7294);
or U7788 (N_7788,N_7017,N_7388);
nor U7789 (N_7789,N_7263,N_7239);
or U7790 (N_7790,N_7035,N_7451);
nor U7791 (N_7791,N_7140,N_7197);
or U7792 (N_7792,N_7312,N_7175);
nand U7793 (N_7793,N_7154,N_7257);
nor U7794 (N_7794,N_7106,N_7354);
and U7795 (N_7795,N_7026,N_7409);
nor U7796 (N_7796,N_7452,N_7058);
or U7797 (N_7797,N_7152,N_7443);
nand U7798 (N_7798,N_7253,N_7390);
and U7799 (N_7799,N_7464,N_7161);
and U7800 (N_7800,N_7479,N_7165);
nand U7801 (N_7801,N_7222,N_7332);
or U7802 (N_7802,N_7319,N_7349);
nor U7803 (N_7803,N_7389,N_7317);
nor U7804 (N_7804,N_7408,N_7018);
or U7805 (N_7805,N_7350,N_7012);
nand U7806 (N_7806,N_7362,N_7102);
or U7807 (N_7807,N_7301,N_7393);
nor U7808 (N_7808,N_7494,N_7187);
xor U7809 (N_7809,N_7111,N_7235);
xor U7810 (N_7810,N_7035,N_7006);
nand U7811 (N_7811,N_7232,N_7422);
nand U7812 (N_7812,N_7108,N_7444);
and U7813 (N_7813,N_7340,N_7165);
or U7814 (N_7814,N_7092,N_7148);
nor U7815 (N_7815,N_7088,N_7290);
and U7816 (N_7816,N_7403,N_7033);
nor U7817 (N_7817,N_7242,N_7210);
nor U7818 (N_7818,N_7177,N_7350);
and U7819 (N_7819,N_7119,N_7384);
xnor U7820 (N_7820,N_7121,N_7162);
xnor U7821 (N_7821,N_7016,N_7491);
xor U7822 (N_7822,N_7366,N_7151);
nor U7823 (N_7823,N_7237,N_7343);
and U7824 (N_7824,N_7422,N_7258);
or U7825 (N_7825,N_7327,N_7277);
and U7826 (N_7826,N_7087,N_7051);
nand U7827 (N_7827,N_7395,N_7062);
or U7828 (N_7828,N_7273,N_7350);
or U7829 (N_7829,N_7419,N_7268);
nand U7830 (N_7830,N_7221,N_7117);
xnor U7831 (N_7831,N_7405,N_7316);
or U7832 (N_7832,N_7006,N_7193);
nand U7833 (N_7833,N_7140,N_7418);
and U7834 (N_7834,N_7346,N_7140);
or U7835 (N_7835,N_7253,N_7231);
or U7836 (N_7836,N_7436,N_7166);
and U7837 (N_7837,N_7323,N_7359);
or U7838 (N_7838,N_7024,N_7325);
xnor U7839 (N_7839,N_7261,N_7026);
nand U7840 (N_7840,N_7203,N_7378);
nand U7841 (N_7841,N_7464,N_7309);
nor U7842 (N_7842,N_7409,N_7127);
or U7843 (N_7843,N_7484,N_7436);
nand U7844 (N_7844,N_7154,N_7113);
nor U7845 (N_7845,N_7430,N_7233);
and U7846 (N_7846,N_7005,N_7484);
or U7847 (N_7847,N_7129,N_7382);
nand U7848 (N_7848,N_7052,N_7483);
or U7849 (N_7849,N_7496,N_7213);
or U7850 (N_7850,N_7052,N_7004);
and U7851 (N_7851,N_7054,N_7258);
nor U7852 (N_7852,N_7238,N_7484);
nor U7853 (N_7853,N_7467,N_7193);
and U7854 (N_7854,N_7200,N_7260);
xnor U7855 (N_7855,N_7168,N_7228);
and U7856 (N_7856,N_7213,N_7137);
and U7857 (N_7857,N_7499,N_7129);
or U7858 (N_7858,N_7151,N_7282);
nand U7859 (N_7859,N_7475,N_7209);
and U7860 (N_7860,N_7443,N_7097);
or U7861 (N_7861,N_7267,N_7413);
nor U7862 (N_7862,N_7417,N_7100);
xnor U7863 (N_7863,N_7096,N_7110);
or U7864 (N_7864,N_7125,N_7416);
and U7865 (N_7865,N_7037,N_7013);
and U7866 (N_7866,N_7346,N_7288);
and U7867 (N_7867,N_7411,N_7041);
and U7868 (N_7868,N_7136,N_7032);
nand U7869 (N_7869,N_7434,N_7476);
xor U7870 (N_7870,N_7499,N_7319);
or U7871 (N_7871,N_7039,N_7398);
nor U7872 (N_7872,N_7394,N_7292);
nand U7873 (N_7873,N_7012,N_7052);
nor U7874 (N_7874,N_7353,N_7309);
nor U7875 (N_7875,N_7424,N_7123);
nor U7876 (N_7876,N_7396,N_7072);
nor U7877 (N_7877,N_7085,N_7070);
xor U7878 (N_7878,N_7387,N_7098);
xnor U7879 (N_7879,N_7306,N_7021);
nand U7880 (N_7880,N_7210,N_7354);
and U7881 (N_7881,N_7140,N_7287);
or U7882 (N_7882,N_7058,N_7280);
and U7883 (N_7883,N_7459,N_7210);
and U7884 (N_7884,N_7124,N_7442);
nand U7885 (N_7885,N_7197,N_7073);
or U7886 (N_7886,N_7380,N_7349);
xnor U7887 (N_7887,N_7197,N_7114);
or U7888 (N_7888,N_7411,N_7442);
and U7889 (N_7889,N_7335,N_7451);
nand U7890 (N_7890,N_7086,N_7491);
and U7891 (N_7891,N_7212,N_7402);
nand U7892 (N_7892,N_7411,N_7091);
or U7893 (N_7893,N_7179,N_7185);
nand U7894 (N_7894,N_7211,N_7317);
nor U7895 (N_7895,N_7363,N_7281);
xnor U7896 (N_7896,N_7439,N_7417);
or U7897 (N_7897,N_7186,N_7274);
or U7898 (N_7898,N_7346,N_7211);
nand U7899 (N_7899,N_7032,N_7441);
nor U7900 (N_7900,N_7035,N_7231);
xnor U7901 (N_7901,N_7483,N_7408);
xnor U7902 (N_7902,N_7030,N_7336);
or U7903 (N_7903,N_7073,N_7031);
nor U7904 (N_7904,N_7459,N_7431);
nand U7905 (N_7905,N_7260,N_7418);
or U7906 (N_7906,N_7465,N_7245);
and U7907 (N_7907,N_7497,N_7109);
and U7908 (N_7908,N_7311,N_7175);
nand U7909 (N_7909,N_7314,N_7428);
or U7910 (N_7910,N_7276,N_7275);
and U7911 (N_7911,N_7435,N_7160);
or U7912 (N_7912,N_7340,N_7078);
and U7913 (N_7913,N_7017,N_7063);
or U7914 (N_7914,N_7272,N_7115);
nor U7915 (N_7915,N_7236,N_7101);
nand U7916 (N_7916,N_7289,N_7446);
nand U7917 (N_7917,N_7198,N_7083);
or U7918 (N_7918,N_7151,N_7104);
xor U7919 (N_7919,N_7423,N_7358);
nand U7920 (N_7920,N_7088,N_7156);
xnor U7921 (N_7921,N_7303,N_7434);
and U7922 (N_7922,N_7223,N_7289);
nor U7923 (N_7923,N_7111,N_7494);
and U7924 (N_7924,N_7162,N_7133);
and U7925 (N_7925,N_7326,N_7372);
and U7926 (N_7926,N_7380,N_7187);
or U7927 (N_7927,N_7291,N_7286);
and U7928 (N_7928,N_7062,N_7309);
xor U7929 (N_7929,N_7328,N_7146);
and U7930 (N_7930,N_7278,N_7136);
or U7931 (N_7931,N_7052,N_7430);
nand U7932 (N_7932,N_7188,N_7264);
or U7933 (N_7933,N_7060,N_7086);
xnor U7934 (N_7934,N_7394,N_7088);
nor U7935 (N_7935,N_7218,N_7490);
or U7936 (N_7936,N_7429,N_7455);
nand U7937 (N_7937,N_7120,N_7228);
or U7938 (N_7938,N_7499,N_7114);
nor U7939 (N_7939,N_7366,N_7132);
xnor U7940 (N_7940,N_7168,N_7175);
nand U7941 (N_7941,N_7246,N_7483);
nor U7942 (N_7942,N_7058,N_7150);
or U7943 (N_7943,N_7012,N_7285);
and U7944 (N_7944,N_7460,N_7309);
and U7945 (N_7945,N_7008,N_7048);
nor U7946 (N_7946,N_7311,N_7222);
and U7947 (N_7947,N_7086,N_7091);
nor U7948 (N_7948,N_7422,N_7013);
and U7949 (N_7949,N_7457,N_7287);
nand U7950 (N_7950,N_7424,N_7180);
nand U7951 (N_7951,N_7107,N_7001);
nand U7952 (N_7952,N_7330,N_7260);
and U7953 (N_7953,N_7267,N_7309);
xor U7954 (N_7954,N_7022,N_7204);
xor U7955 (N_7955,N_7470,N_7047);
and U7956 (N_7956,N_7411,N_7281);
nor U7957 (N_7957,N_7294,N_7120);
or U7958 (N_7958,N_7012,N_7027);
nand U7959 (N_7959,N_7323,N_7368);
and U7960 (N_7960,N_7256,N_7316);
and U7961 (N_7961,N_7349,N_7361);
and U7962 (N_7962,N_7277,N_7043);
nand U7963 (N_7963,N_7069,N_7168);
nand U7964 (N_7964,N_7136,N_7071);
nor U7965 (N_7965,N_7479,N_7154);
and U7966 (N_7966,N_7109,N_7423);
nand U7967 (N_7967,N_7169,N_7448);
nor U7968 (N_7968,N_7318,N_7100);
nand U7969 (N_7969,N_7382,N_7384);
and U7970 (N_7970,N_7262,N_7414);
nor U7971 (N_7971,N_7499,N_7287);
xor U7972 (N_7972,N_7454,N_7361);
and U7973 (N_7973,N_7283,N_7058);
and U7974 (N_7974,N_7217,N_7206);
nand U7975 (N_7975,N_7221,N_7068);
nor U7976 (N_7976,N_7040,N_7380);
xor U7977 (N_7977,N_7320,N_7182);
and U7978 (N_7978,N_7470,N_7097);
and U7979 (N_7979,N_7361,N_7172);
xor U7980 (N_7980,N_7384,N_7377);
xor U7981 (N_7981,N_7085,N_7254);
and U7982 (N_7982,N_7394,N_7386);
and U7983 (N_7983,N_7421,N_7109);
nand U7984 (N_7984,N_7283,N_7145);
and U7985 (N_7985,N_7356,N_7060);
nor U7986 (N_7986,N_7381,N_7251);
nand U7987 (N_7987,N_7142,N_7327);
or U7988 (N_7988,N_7096,N_7439);
or U7989 (N_7989,N_7134,N_7099);
and U7990 (N_7990,N_7444,N_7257);
xnor U7991 (N_7991,N_7178,N_7230);
or U7992 (N_7992,N_7460,N_7488);
nor U7993 (N_7993,N_7271,N_7066);
nor U7994 (N_7994,N_7168,N_7070);
or U7995 (N_7995,N_7231,N_7432);
nand U7996 (N_7996,N_7269,N_7404);
nor U7997 (N_7997,N_7138,N_7161);
or U7998 (N_7998,N_7131,N_7392);
nand U7999 (N_7999,N_7275,N_7295);
and U8000 (N_8000,N_7826,N_7561);
nor U8001 (N_8001,N_7611,N_7981);
nor U8002 (N_8002,N_7557,N_7502);
and U8003 (N_8003,N_7857,N_7830);
or U8004 (N_8004,N_7515,N_7840);
nand U8005 (N_8005,N_7945,N_7705);
nor U8006 (N_8006,N_7684,N_7745);
nand U8007 (N_8007,N_7694,N_7687);
nand U8008 (N_8008,N_7585,N_7696);
nand U8009 (N_8009,N_7772,N_7971);
or U8010 (N_8010,N_7781,N_7630);
and U8011 (N_8011,N_7609,N_7800);
or U8012 (N_8012,N_7583,N_7839);
nor U8013 (N_8013,N_7523,N_7841);
or U8014 (N_8014,N_7579,N_7511);
or U8015 (N_8015,N_7681,N_7550);
nor U8016 (N_8016,N_7596,N_7657);
or U8017 (N_8017,N_7899,N_7816);
xor U8018 (N_8018,N_7728,N_7984);
and U8019 (N_8019,N_7709,N_7675);
nand U8020 (N_8020,N_7559,N_7973);
or U8021 (N_8021,N_7567,N_7608);
and U8022 (N_8022,N_7940,N_7530);
and U8023 (N_8023,N_7995,N_7967);
or U8024 (N_8024,N_7729,N_7814);
xor U8025 (N_8025,N_7996,N_7999);
xnor U8026 (N_8026,N_7663,N_7507);
and U8027 (N_8027,N_7722,N_7914);
and U8028 (N_8028,N_7635,N_7524);
and U8029 (N_8029,N_7812,N_7662);
xor U8030 (N_8030,N_7606,N_7831);
or U8031 (N_8031,N_7793,N_7885);
xnor U8032 (N_8032,N_7939,N_7604);
nand U8033 (N_8033,N_7680,N_7510);
nor U8034 (N_8034,N_7732,N_7886);
nor U8035 (N_8035,N_7955,N_7884);
and U8036 (N_8036,N_7533,N_7925);
nand U8037 (N_8037,N_7874,N_7811);
or U8038 (N_8038,N_7624,N_7572);
and U8039 (N_8039,N_7862,N_7948);
or U8040 (N_8040,N_7855,N_7716);
and U8041 (N_8041,N_7828,N_7619);
nand U8042 (N_8042,N_7626,N_7843);
or U8043 (N_8043,N_7938,N_7654);
and U8044 (N_8044,N_7879,N_7763);
nor U8045 (N_8045,N_7752,N_7861);
or U8046 (N_8046,N_7864,N_7564);
or U8047 (N_8047,N_7695,N_7650);
and U8048 (N_8048,N_7771,N_7897);
nand U8049 (N_8049,N_7570,N_7892);
nor U8050 (N_8050,N_7637,N_7944);
and U8051 (N_8051,N_7943,N_7714);
nor U8052 (N_8052,N_7634,N_7631);
and U8053 (N_8053,N_7903,N_7615);
and U8054 (N_8054,N_7983,N_7571);
nor U8055 (N_8055,N_7736,N_7738);
nor U8056 (N_8056,N_7954,N_7715);
nor U8057 (N_8057,N_7718,N_7780);
nand U8058 (N_8058,N_7527,N_7549);
nand U8059 (N_8059,N_7930,N_7742);
xnor U8060 (N_8060,N_7829,N_7825);
and U8061 (N_8061,N_7649,N_7907);
and U8062 (N_8062,N_7777,N_7882);
nand U8063 (N_8063,N_7591,N_7856);
xor U8064 (N_8064,N_7685,N_7957);
nand U8065 (N_8065,N_7574,N_7669);
and U8066 (N_8066,N_7540,N_7946);
xor U8067 (N_8067,N_7976,N_7818);
and U8068 (N_8068,N_7547,N_7850);
or U8069 (N_8069,N_7833,N_7985);
or U8070 (N_8070,N_7783,N_7689);
nand U8071 (N_8071,N_7911,N_7798);
or U8072 (N_8072,N_7620,N_7791);
nand U8073 (N_8073,N_7751,N_7865);
nor U8074 (N_8074,N_7670,N_7852);
and U8075 (N_8075,N_7704,N_7809);
or U8076 (N_8076,N_7951,N_7597);
or U8077 (N_8077,N_7817,N_7851);
and U8078 (N_8078,N_7933,N_7614);
or U8079 (N_8079,N_7541,N_7847);
nand U8080 (N_8080,N_7928,N_7878);
nor U8081 (N_8081,N_7845,N_7994);
or U8082 (N_8082,N_7896,N_7827);
or U8083 (N_8083,N_7532,N_7893);
or U8084 (N_8084,N_7774,N_7628);
nor U8085 (N_8085,N_7953,N_7554);
xor U8086 (N_8086,N_7539,N_7796);
xor U8087 (N_8087,N_7848,N_7921);
nand U8088 (N_8088,N_7970,N_7587);
and U8089 (N_8089,N_7590,N_7602);
and U8090 (N_8090,N_7759,N_7807);
nor U8091 (N_8091,N_7918,N_7639);
nor U8092 (N_8092,N_7778,N_7671);
nand U8093 (N_8093,N_7720,N_7676);
or U8094 (N_8094,N_7659,N_7989);
or U8095 (N_8095,N_7645,N_7834);
nand U8096 (N_8096,N_7575,N_7813);
nand U8097 (N_8097,N_7883,N_7797);
nor U8098 (N_8098,N_7627,N_7652);
nor U8099 (N_8099,N_7688,N_7859);
nand U8100 (N_8100,N_7867,N_7528);
nand U8101 (N_8101,N_7516,N_7525);
nand U8102 (N_8102,N_7513,N_7677);
and U8103 (N_8103,N_7599,N_7594);
nor U8104 (N_8104,N_7543,N_7629);
nand U8105 (N_8105,N_7582,N_7692);
xnor U8106 (N_8106,N_7673,N_7821);
nand U8107 (N_8107,N_7832,N_7711);
or U8108 (N_8108,N_7501,N_7666);
or U8109 (N_8109,N_7668,N_7558);
xor U8110 (N_8110,N_7690,N_7785);
nand U8111 (N_8111,N_7642,N_7991);
xnor U8112 (N_8112,N_7929,N_7963);
or U8113 (N_8113,N_7717,N_7647);
and U8114 (N_8114,N_7782,N_7779);
or U8115 (N_8115,N_7701,N_7721);
or U8116 (N_8116,N_7888,N_7735);
nand U8117 (N_8117,N_7758,N_7544);
nor U8118 (N_8118,N_7693,N_7998);
xor U8119 (N_8119,N_7926,N_7952);
and U8120 (N_8120,N_7706,N_7902);
nand U8121 (N_8121,N_7880,N_7801);
and U8122 (N_8122,N_7870,N_7868);
nor U8123 (N_8123,N_7871,N_7968);
xor U8124 (N_8124,N_7734,N_7529);
nand U8125 (N_8125,N_7920,N_7905);
nand U8126 (N_8126,N_7860,N_7504);
nand U8127 (N_8127,N_7787,N_7912);
and U8128 (N_8128,N_7520,N_7503);
nor U8129 (N_8129,N_7962,N_7910);
nor U8130 (N_8130,N_7819,N_7678);
xnor U8131 (N_8131,N_7906,N_7723);
or U8132 (N_8132,N_7674,N_7773);
nand U8133 (N_8133,N_7784,N_7578);
or U8134 (N_8134,N_7965,N_7600);
or U8135 (N_8135,N_7537,N_7610);
nand U8136 (N_8136,N_7712,N_7508);
or U8137 (N_8137,N_7986,N_7556);
nand U8138 (N_8138,N_7514,N_7601);
and U8139 (N_8139,N_7691,N_7708);
or U8140 (N_8140,N_7802,N_7961);
nand U8141 (N_8141,N_7877,N_7838);
xnor U8142 (N_8142,N_7733,N_7740);
nand U8143 (N_8143,N_7545,N_7936);
or U8144 (N_8144,N_7552,N_7613);
nand U8145 (N_8145,N_7636,N_7869);
xor U8146 (N_8146,N_7810,N_7555);
or U8147 (N_8147,N_7788,N_7749);
and U8148 (N_8148,N_7698,N_7644);
nor U8149 (N_8149,N_7987,N_7769);
or U8150 (N_8150,N_7931,N_7947);
nand U8151 (N_8151,N_7622,N_7569);
nor U8152 (N_8152,N_7808,N_7643);
or U8153 (N_8153,N_7616,N_7731);
or U8154 (N_8154,N_7764,N_7648);
nand U8155 (N_8155,N_7739,N_7707);
nor U8156 (N_8156,N_7997,N_7993);
or U8157 (N_8157,N_7776,N_7580);
and U8158 (N_8158,N_7979,N_7744);
nor U8159 (N_8159,N_7923,N_7756);
nand U8160 (N_8160,N_7605,N_7598);
or U8161 (N_8161,N_7700,N_7950);
and U8162 (N_8162,N_7535,N_7713);
or U8163 (N_8163,N_7618,N_7534);
or U8164 (N_8164,N_7686,N_7901);
nor U8165 (N_8165,N_7762,N_7750);
xnor U8166 (N_8166,N_7978,N_7748);
and U8167 (N_8167,N_7881,N_7573);
nor U8168 (N_8168,N_7815,N_7553);
or U8169 (N_8169,N_7803,N_7625);
or U8170 (N_8170,N_7908,N_7942);
nand U8171 (N_8171,N_7934,N_7584);
or U8172 (N_8172,N_7546,N_7824);
nor U8173 (N_8173,N_7612,N_7941);
nor U8174 (N_8174,N_7702,N_7768);
nor U8175 (N_8175,N_7697,N_7623);
nor U8176 (N_8176,N_7621,N_7949);
nor U8177 (N_8177,N_7542,N_7786);
or U8178 (N_8178,N_7975,N_7724);
nand U8179 (N_8179,N_7915,N_7972);
and U8180 (N_8180,N_7683,N_7844);
xor U8181 (N_8181,N_7927,N_7651);
nor U8182 (N_8182,N_7538,N_7964);
or U8183 (N_8183,N_7770,N_7853);
nand U8184 (N_8184,N_7726,N_7522);
and U8185 (N_8185,N_7804,N_7894);
and U8186 (N_8186,N_7846,N_7757);
or U8187 (N_8187,N_7876,N_7576);
nor U8188 (N_8188,N_7937,N_7531);
nor U8189 (N_8189,N_7506,N_7753);
nor U8190 (N_8190,N_7890,N_7737);
and U8191 (N_8191,N_7895,N_7904);
or U8192 (N_8192,N_7820,N_7919);
and U8193 (N_8193,N_7887,N_7656);
or U8194 (N_8194,N_7792,N_7891);
nand U8195 (N_8195,N_7633,N_7660);
and U8196 (N_8196,N_7806,N_7754);
nand U8197 (N_8197,N_7789,N_7568);
or U8198 (N_8198,N_7900,N_7795);
or U8199 (N_8199,N_7765,N_7640);
or U8200 (N_8200,N_7641,N_7521);
nand U8201 (N_8201,N_7730,N_7517);
and U8202 (N_8202,N_7849,N_7672);
and U8203 (N_8203,N_7767,N_7500);
nor U8204 (N_8204,N_7898,N_7679);
nor U8205 (N_8205,N_7872,N_7658);
nor U8206 (N_8206,N_7766,N_7505);
or U8207 (N_8207,N_7710,N_7664);
or U8208 (N_8208,N_7836,N_7755);
nand U8209 (N_8209,N_7842,N_7746);
or U8210 (N_8210,N_7747,N_7959);
nor U8211 (N_8211,N_7592,N_7980);
nor U8212 (N_8212,N_7982,N_7835);
nand U8213 (N_8213,N_7823,N_7551);
nor U8214 (N_8214,N_7966,N_7603);
nor U8215 (N_8215,N_7595,N_7519);
nor U8216 (N_8216,N_7924,N_7593);
or U8217 (N_8217,N_7743,N_7922);
nand U8218 (N_8218,N_7653,N_7665);
or U8219 (N_8219,N_7661,N_7866);
or U8220 (N_8220,N_7858,N_7822);
nand U8221 (N_8221,N_7682,N_7794);
nor U8222 (N_8222,N_7607,N_7917);
and U8223 (N_8223,N_7932,N_7667);
and U8224 (N_8224,N_7577,N_7956);
nor U8225 (N_8225,N_7566,N_7655);
and U8226 (N_8226,N_7617,N_7719);
nand U8227 (N_8227,N_7562,N_7563);
nand U8228 (N_8228,N_7799,N_7977);
or U8229 (N_8229,N_7699,N_7588);
or U8230 (N_8230,N_7760,N_7958);
nand U8231 (N_8231,N_7969,N_7863);
and U8232 (N_8232,N_7889,N_7586);
nor U8233 (N_8233,N_7536,N_7761);
nor U8234 (N_8234,N_7992,N_7518);
xor U8235 (N_8235,N_7988,N_7854);
or U8236 (N_8236,N_7526,N_7990);
or U8237 (N_8237,N_7727,N_7632);
and U8238 (N_8238,N_7873,N_7916);
or U8239 (N_8239,N_7725,N_7589);
and U8240 (N_8240,N_7974,N_7960);
and U8241 (N_8241,N_7548,N_7509);
nand U8242 (N_8242,N_7646,N_7512);
or U8243 (N_8243,N_7790,N_7775);
nor U8244 (N_8244,N_7581,N_7805);
and U8245 (N_8245,N_7837,N_7741);
and U8246 (N_8246,N_7875,N_7909);
or U8247 (N_8247,N_7565,N_7638);
or U8248 (N_8248,N_7703,N_7560);
or U8249 (N_8249,N_7913,N_7935);
and U8250 (N_8250,N_7900,N_7885);
nand U8251 (N_8251,N_7561,N_7590);
and U8252 (N_8252,N_7714,N_7772);
and U8253 (N_8253,N_7712,N_7671);
and U8254 (N_8254,N_7516,N_7655);
or U8255 (N_8255,N_7809,N_7921);
nor U8256 (N_8256,N_7851,N_7765);
nand U8257 (N_8257,N_7794,N_7967);
nand U8258 (N_8258,N_7869,N_7722);
and U8259 (N_8259,N_7537,N_7596);
nand U8260 (N_8260,N_7973,N_7527);
nor U8261 (N_8261,N_7968,N_7544);
and U8262 (N_8262,N_7693,N_7791);
xor U8263 (N_8263,N_7713,N_7820);
nor U8264 (N_8264,N_7824,N_7523);
or U8265 (N_8265,N_7678,N_7638);
or U8266 (N_8266,N_7576,N_7732);
nor U8267 (N_8267,N_7732,N_7529);
or U8268 (N_8268,N_7774,N_7810);
or U8269 (N_8269,N_7953,N_7856);
xor U8270 (N_8270,N_7849,N_7975);
nor U8271 (N_8271,N_7789,N_7625);
or U8272 (N_8272,N_7964,N_7620);
nand U8273 (N_8273,N_7630,N_7573);
nand U8274 (N_8274,N_7576,N_7871);
nor U8275 (N_8275,N_7630,N_7737);
or U8276 (N_8276,N_7981,N_7781);
nand U8277 (N_8277,N_7709,N_7663);
and U8278 (N_8278,N_7720,N_7901);
xnor U8279 (N_8279,N_7751,N_7715);
xnor U8280 (N_8280,N_7615,N_7879);
and U8281 (N_8281,N_7896,N_7543);
or U8282 (N_8282,N_7851,N_7701);
nand U8283 (N_8283,N_7911,N_7825);
nand U8284 (N_8284,N_7584,N_7901);
and U8285 (N_8285,N_7616,N_7994);
or U8286 (N_8286,N_7912,N_7529);
xor U8287 (N_8287,N_7968,N_7521);
nor U8288 (N_8288,N_7729,N_7658);
or U8289 (N_8289,N_7505,N_7657);
nor U8290 (N_8290,N_7618,N_7733);
nor U8291 (N_8291,N_7879,N_7811);
and U8292 (N_8292,N_7837,N_7873);
nor U8293 (N_8293,N_7969,N_7834);
xor U8294 (N_8294,N_7889,N_7843);
and U8295 (N_8295,N_7510,N_7627);
or U8296 (N_8296,N_7580,N_7721);
nand U8297 (N_8297,N_7657,N_7985);
xnor U8298 (N_8298,N_7849,N_7816);
and U8299 (N_8299,N_7665,N_7912);
or U8300 (N_8300,N_7650,N_7772);
or U8301 (N_8301,N_7864,N_7742);
and U8302 (N_8302,N_7629,N_7732);
and U8303 (N_8303,N_7646,N_7722);
nor U8304 (N_8304,N_7808,N_7565);
or U8305 (N_8305,N_7542,N_7919);
and U8306 (N_8306,N_7990,N_7507);
nor U8307 (N_8307,N_7889,N_7759);
and U8308 (N_8308,N_7735,N_7897);
or U8309 (N_8309,N_7662,N_7975);
nor U8310 (N_8310,N_7755,N_7817);
nor U8311 (N_8311,N_7730,N_7851);
or U8312 (N_8312,N_7694,N_7939);
or U8313 (N_8313,N_7695,N_7611);
nor U8314 (N_8314,N_7856,N_7749);
or U8315 (N_8315,N_7612,N_7664);
or U8316 (N_8316,N_7774,N_7899);
and U8317 (N_8317,N_7800,N_7671);
nand U8318 (N_8318,N_7814,N_7828);
nand U8319 (N_8319,N_7688,N_7852);
xor U8320 (N_8320,N_7898,N_7549);
nor U8321 (N_8321,N_7687,N_7610);
or U8322 (N_8322,N_7922,N_7939);
or U8323 (N_8323,N_7720,N_7695);
nand U8324 (N_8324,N_7954,N_7915);
nor U8325 (N_8325,N_7995,N_7856);
nand U8326 (N_8326,N_7743,N_7805);
or U8327 (N_8327,N_7895,N_7626);
nand U8328 (N_8328,N_7702,N_7852);
nor U8329 (N_8329,N_7837,N_7745);
nor U8330 (N_8330,N_7637,N_7570);
and U8331 (N_8331,N_7514,N_7538);
and U8332 (N_8332,N_7602,N_7620);
xor U8333 (N_8333,N_7792,N_7794);
or U8334 (N_8334,N_7926,N_7755);
or U8335 (N_8335,N_7913,N_7856);
nor U8336 (N_8336,N_7522,N_7523);
nand U8337 (N_8337,N_7607,N_7700);
and U8338 (N_8338,N_7564,N_7625);
xor U8339 (N_8339,N_7965,N_7971);
nor U8340 (N_8340,N_7558,N_7799);
and U8341 (N_8341,N_7965,N_7826);
or U8342 (N_8342,N_7868,N_7820);
or U8343 (N_8343,N_7538,N_7552);
and U8344 (N_8344,N_7900,N_7666);
nor U8345 (N_8345,N_7942,N_7780);
or U8346 (N_8346,N_7680,N_7847);
and U8347 (N_8347,N_7834,N_7749);
nor U8348 (N_8348,N_7852,N_7919);
or U8349 (N_8349,N_7725,N_7570);
nor U8350 (N_8350,N_7651,N_7757);
nor U8351 (N_8351,N_7506,N_7634);
nor U8352 (N_8352,N_7536,N_7640);
or U8353 (N_8353,N_7732,N_7566);
nor U8354 (N_8354,N_7762,N_7655);
nor U8355 (N_8355,N_7679,N_7745);
nand U8356 (N_8356,N_7732,N_7579);
nand U8357 (N_8357,N_7933,N_7663);
nand U8358 (N_8358,N_7591,N_7903);
nand U8359 (N_8359,N_7874,N_7697);
nand U8360 (N_8360,N_7519,N_7838);
or U8361 (N_8361,N_7824,N_7792);
xor U8362 (N_8362,N_7513,N_7880);
nor U8363 (N_8363,N_7839,N_7571);
or U8364 (N_8364,N_7854,N_7866);
or U8365 (N_8365,N_7781,N_7943);
nor U8366 (N_8366,N_7512,N_7980);
nand U8367 (N_8367,N_7817,N_7836);
nand U8368 (N_8368,N_7727,N_7830);
and U8369 (N_8369,N_7921,N_7542);
and U8370 (N_8370,N_7875,N_7958);
nor U8371 (N_8371,N_7718,N_7663);
and U8372 (N_8372,N_7589,N_7890);
nor U8373 (N_8373,N_7504,N_7972);
nand U8374 (N_8374,N_7524,N_7766);
nand U8375 (N_8375,N_7630,N_7652);
nand U8376 (N_8376,N_7715,N_7683);
nand U8377 (N_8377,N_7859,N_7758);
nand U8378 (N_8378,N_7909,N_7678);
or U8379 (N_8379,N_7584,N_7892);
or U8380 (N_8380,N_7767,N_7873);
nand U8381 (N_8381,N_7785,N_7867);
nor U8382 (N_8382,N_7574,N_7934);
or U8383 (N_8383,N_7765,N_7520);
and U8384 (N_8384,N_7588,N_7834);
and U8385 (N_8385,N_7535,N_7508);
and U8386 (N_8386,N_7799,N_7791);
nor U8387 (N_8387,N_7809,N_7900);
or U8388 (N_8388,N_7582,N_7956);
nor U8389 (N_8389,N_7862,N_7990);
or U8390 (N_8390,N_7535,N_7935);
or U8391 (N_8391,N_7573,N_7997);
or U8392 (N_8392,N_7738,N_7794);
or U8393 (N_8393,N_7656,N_7832);
or U8394 (N_8394,N_7648,N_7726);
xnor U8395 (N_8395,N_7838,N_7855);
xnor U8396 (N_8396,N_7724,N_7856);
nor U8397 (N_8397,N_7597,N_7702);
and U8398 (N_8398,N_7931,N_7677);
or U8399 (N_8399,N_7921,N_7974);
and U8400 (N_8400,N_7756,N_7508);
and U8401 (N_8401,N_7851,N_7626);
nor U8402 (N_8402,N_7758,N_7552);
nor U8403 (N_8403,N_7598,N_7664);
or U8404 (N_8404,N_7555,N_7794);
and U8405 (N_8405,N_7614,N_7724);
nor U8406 (N_8406,N_7879,N_7778);
nand U8407 (N_8407,N_7959,N_7553);
or U8408 (N_8408,N_7625,N_7648);
nor U8409 (N_8409,N_7866,N_7678);
xnor U8410 (N_8410,N_7617,N_7762);
nand U8411 (N_8411,N_7718,N_7684);
and U8412 (N_8412,N_7571,N_7986);
or U8413 (N_8413,N_7672,N_7806);
nand U8414 (N_8414,N_7674,N_7966);
nor U8415 (N_8415,N_7697,N_7871);
or U8416 (N_8416,N_7695,N_7840);
nor U8417 (N_8417,N_7729,N_7593);
nand U8418 (N_8418,N_7965,N_7692);
and U8419 (N_8419,N_7653,N_7749);
or U8420 (N_8420,N_7866,N_7685);
or U8421 (N_8421,N_7855,N_7701);
nor U8422 (N_8422,N_7849,N_7504);
nor U8423 (N_8423,N_7641,N_7689);
or U8424 (N_8424,N_7630,N_7506);
nor U8425 (N_8425,N_7659,N_7938);
nand U8426 (N_8426,N_7926,N_7710);
nor U8427 (N_8427,N_7851,N_7521);
or U8428 (N_8428,N_7878,N_7855);
nor U8429 (N_8429,N_7996,N_7939);
or U8430 (N_8430,N_7564,N_7735);
nor U8431 (N_8431,N_7953,N_7946);
nor U8432 (N_8432,N_7824,N_7721);
and U8433 (N_8433,N_7736,N_7631);
nand U8434 (N_8434,N_7598,N_7785);
or U8435 (N_8435,N_7692,N_7615);
nor U8436 (N_8436,N_7620,N_7857);
nand U8437 (N_8437,N_7904,N_7884);
and U8438 (N_8438,N_7815,N_7779);
or U8439 (N_8439,N_7544,N_7896);
nand U8440 (N_8440,N_7522,N_7645);
nand U8441 (N_8441,N_7746,N_7667);
xnor U8442 (N_8442,N_7906,N_7825);
nor U8443 (N_8443,N_7920,N_7990);
nor U8444 (N_8444,N_7904,N_7591);
and U8445 (N_8445,N_7950,N_7978);
or U8446 (N_8446,N_7919,N_7709);
nand U8447 (N_8447,N_7846,N_7677);
or U8448 (N_8448,N_7707,N_7856);
nand U8449 (N_8449,N_7914,N_7702);
xnor U8450 (N_8450,N_7502,N_7904);
nand U8451 (N_8451,N_7700,N_7676);
nor U8452 (N_8452,N_7632,N_7969);
and U8453 (N_8453,N_7646,N_7547);
xor U8454 (N_8454,N_7817,N_7509);
and U8455 (N_8455,N_7761,N_7941);
xor U8456 (N_8456,N_7768,N_7809);
and U8457 (N_8457,N_7837,N_7669);
nor U8458 (N_8458,N_7980,N_7798);
nand U8459 (N_8459,N_7514,N_7906);
nor U8460 (N_8460,N_7948,N_7627);
nand U8461 (N_8461,N_7621,N_7842);
or U8462 (N_8462,N_7898,N_7808);
and U8463 (N_8463,N_7775,N_7907);
and U8464 (N_8464,N_7720,N_7740);
or U8465 (N_8465,N_7759,N_7569);
or U8466 (N_8466,N_7527,N_7693);
xor U8467 (N_8467,N_7966,N_7662);
or U8468 (N_8468,N_7791,N_7696);
or U8469 (N_8469,N_7884,N_7906);
nand U8470 (N_8470,N_7699,N_7739);
or U8471 (N_8471,N_7880,N_7631);
nand U8472 (N_8472,N_7767,N_7962);
xnor U8473 (N_8473,N_7789,N_7577);
nand U8474 (N_8474,N_7758,N_7944);
nor U8475 (N_8475,N_7648,N_7843);
xnor U8476 (N_8476,N_7975,N_7887);
nand U8477 (N_8477,N_7969,N_7522);
and U8478 (N_8478,N_7587,N_7704);
nand U8479 (N_8479,N_7919,N_7646);
or U8480 (N_8480,N_7856,N_7963);
or U8481 (N_8481,N_7900,N_7627);
nand U8482 (N_8482,N_7731,N_7842);
nor U8483 (N_8483,N_7949,N_7619);
and U8484 (N_8484,N_7748,N_7592);
nor U8485 (N_8485,N_7897,N_7672);
nand U8486 (N_8486,N_7801,N_7808);
nor U8487 (N_8487,N_7502,N_7589);
and U8488 (N_8488,N_7542,N_7719);
nor U8489 (N_8489,N_7762,N_7708);
xnor U8490 (N_8490,N_7552,N_7848);
nand U8491 (N_8491,N_7611,N_7504);
and U8492 (N_8492,N_7578,N_7846);
nor U8493 (N_8493,N_7549,N_7523);
nand U8494 (N_8494,N_7634,N_7534);
and U8495 (N_8495,N_7635,N_7784);
and U8496 (N_8496,N_7616,N_7918);
and U8497 (N_8497,N_7702,N_7793);
or U8498 (N_8498,N_7544,N_7670);
and U8499 (N_8499,N_7917,N_7789);
nor U8500 (N_8500,N_8343,N_8195);
and U8501 (N_8501,N_8360,N_8319);
or U8502 (N_8502,N_8261,N_8112);
or U8503 (N_8503,N_8125,N_8329);
and U8504 (N_8504,N_8079,N_8355);
nor U8505 (N_8505,N_8048,N_8454);
xor U8506 (N_8506,N_8430,N_8259);
nor U8507 (N_8507,N_8174,N_8279);
nor U8508 (N_8508,N_8165,N_8148);
or U8509 (N_8509,N_8186,N_8235);
nor U8510 (N_8510,N_8043,N_8074);
nor U8511 (N_8511,N_8384,N_8085);
or U8512 (N_8512,N_8309,N_8059);
nand U8513 (N_8513,N_8067,N_8320);
nor U8514 (N_8514,N_8130,N_8250);
or U8515 (N_8515,N_8313,N_8167);
nor U8516 (N_8516,N_8228,N_8110);
nor U8517 (N_8517,N_8354,N_8251);
and U8518 (N_8518,N_8306,N_8489);
and U8519 (N_8519,N_8460,N_8442);
nand U8520 (N_8520,N_8202,N_8042);
nand U8521 (N_8521,N_8135,N_8453);
or U8522 (N_8522,N_8177,N_8030);
or U8523 (N_8523,N_8116,N_8459);
nand U8524 (N_8524,N_8469,N_8190);
or U8525 (N_8525,N_8111,N_8429);
xor U8526 (N_8526,N_8350,N_8367);
and U8527 (N_8527,N_8188,N_8417);
nor U8528 (N_8528,N_8396,N_8142);
and U8529 (N_8529,N_8184,N_8397);
and U8530 (N_8530,N_8164,N_8088);
and U8531 (N_8531,N_8427,N_8137);
xnor U8532 (N_8532,N_8376,N_8201);
xnor U8533 (N_8533,N_8325,N_8011);
or U8534 (N_8534,N_8096,N_8414);
nand U8535 (N_8535,N_8268,N_8041);
nand U8536 (N_8536,N_8040,N_8182);
or U8537 (N_8537,N_8327,N_8133);
xnor U8538 (N_8538,N_8117,N_8445);
xor U8539 (N_8539,N_8449,N_8022);
nand U8540 (N_8540,N_8389,N_8222);
nor U8541 (N_8541,N_8215,N_8093);
xnor U8542 (N_8542,N_8418,N_8101);
nand U8543 (N_8543,N_8070,N_8495);
or U8544 (N_8544,N_8439,N_8256);
nor U8545 (N_8545,N_8403,N_8257);
nand U8546 (N_8546,N_8365,N_8298);
nor U8547 (N_8547,N_8294,N_8039);
or U8548 (N_8548,N_8173,N_8082);
and U8549 (N_8549,N_8016,N_8193);
and U8550 (N_8550,N_8032,N_8156);
xnor U8551 (N_8551,N_8047,N_8075);
nand U8552 (N_8552,N_8468,N_8208);
and U8553 (N_8553,N_8197,N_8299);
nor U8554 (N_8554,N_8492,N_8420);
xor U8555 (N_8555,N_8436,N_8054);
or U8556 (N_8556,N_8395,N_8159);
nor U8557 (N_8557,N_8311,N_8340);
and U8558 (N_8558,N_8183,N_8273);
or U8559 (N_8559,N_8321,N_8007);
xor U8560 (N_8560,N_8451,N_8146);
or U8561 (N_8561,N_8203,N_8393);
nor U8562 (N_8562,N_8461,N_8226);
or U8563 (N_8563,N_8061,N_8058);
or U8564 (N_8564,N_8349,N_8302);
nand U8565 (N_8565,N_8045,N_8356);
and U8566 (N_8566,N_8390,N_8283);
nand U8567 (N_8567,N_8443,N_8363);
nand U8568 (N_8568,N_8267,N_8025);
and U8569 (N_8569,N_8179,N_8083);
and U8570 (N_8570,N_8081,N_8091);
and U8571 (N_8571,N_8410,N_8178);
nor U8572 (N_8572,N_8379,N_8232);
or U8573 (N_8573,N_8052,N_8108);
and U8574 (N_8574,N_8003,N_8448);
nor U8575 (N_8575,N_8286,N_8297);
xor U8576 (N_8576,N_8415,N_8467);
and U8577 (N_8577,N_8078,N_8002);
and U8578 (N_8578,N_8134,N_8225);
nor U8579 (N_8579,N_8104,N_8176);
and U8580 (N_8580,N_8324,N_8212);
and U8581 (N_8581,N_8404,N_8314);
or U8582 (N_8582,N_8457,N_8358);
or U8583 (N_8583,N_8018,N_8377);
and U8584 (N_8584,N_8281,N_8060);
nor U8585 (N_8585,N_8100,N_8333);
and U8586 (N_8586,N_8149,N_8163);
nand U8587 (N_8587,N_8316,N_8154);
xor U8588 (N_8588,N_8141,N_8441);
or U8589 (N_8589,N_8326,N_8065);
and U8590 (N_8590,N_8375,N_8383);
nand U8591 (N_8591,N_8481,N_8105);
nor U8592 (N_8592,N_8001,N_8057);
nand U8593 (N_8593,N_8493,N_8296);
nand U8594 (N_8594,N_8305,N_8006);
nor U8595 (N_8595,N_8152,N_8099);
nand U8596 (N_8596,N_8170,N_8046);
xor U8597 (N_8597,N_8408,N_8307);
and U8598 (N_8598,N_8243,N_8231);
and U8599 (N_8599,N_8247,N_8361);
or U8600 (N_8600,N_8284,N_8229);
or U8601 (N_8601,N_8400,N_8462);
nor U8602 (N_8602,N_8072,N_8474);
xor U8603 (N_8603,N_8171,N_8109);
or U8604 (N_8604,N_8373,N_8412);
nor U8605 (N_8605,N_8252,N_8388);
or U8606 (N_8606,N_8411,N_8084);
or U8607 (N_8607,N_8335,N_8103);
and U8608 (N_8608,N_8285,N_8458);
nor U8609 (N_8609,N_8200,N_8478);
or U8610 (N_8610,N_8424,N_8345);
and U8611 (N_8611,N_8308,N_8486);
or U8612 (N_8612,N_8346,N_8168);
xor U8613 (N_8613,N_8038,N_8020);
xor U8614 (N_8614,N_8207,N_8245);
nand U8615 (N_8615,N_8288,N_8000);
nand U8616 (N_8616,N_8253,N_8322);
and U8617 (N_8617,N_8416,N_8401);
and U8618 (N_8618,N_8272,N_8166);
or U8619 (N_8619,N_8063,N_8428);
or U8620 (N_8620,N_8338,N_8271);
and U8621 (N_8621,N_8336,N_8127);
nand U8622 (N_8622,N_8344,N_8248);
nor U8623 (N_8623,N_8371,N_8240);
nand U8624 (N_8624,N_8017,N_8293);
and U8625 (N_8625,N_8431,N_8419);
nand U8626 (N_8626,N_8161,N_8055);
xnor U8627 (N_8627,N_8386,N_8277);
and U8628 (N_8628,N_8269,N_8008);
and U8629 (N_8629,N_8262,N_8090);
nor U8630 (N_8630,N_8484,N_8066);
or U8631 (N_8631,N_8473,N_8398);
or U8632 (N_8632,N_8405,N_8233);
or U8633 (N_8633,N_8264,N_8351);
or U8634 (N_8634,N_8260,N_8169);
and U8635 (N_8635,N_8219,N_8132);
nor U8636 (N_8636,N_8372,N_8472);
or U8637 (N_8637,N_8255,N_8098);
nor U8638 (N_8638,N_8425,N_8214);
nand U8639 (N_8639,N_8475,N_8217);
nand U8640 (N_8640,N_8406,N_8077);
nand U8641 (N_8641,N_8227,N_8122);
nor U8642 (N_8642,N_8366,N_8402);
nand U8643 (N_8643,N_8392,N_8114);
or U8644 (N_8644,N_8120,N_8009);
nand U8645 (N_8645,N_8278,N_8050);
or U8646 (N_8646,N_8471,N_8194);
or U8647 (N_8647,N_8369,N_8004);
and U8648 (N_8648,N_8053,N_8160);
nor U8649 (N_8649,N_8455,N_8086);
and U8650 (N_8650,N_8220,N_8485);
and U8651 (N_8651,N_8238,N_8051);
and U8652 (N_8652,N_8433,N_8044);
and U8653 (N_8653,N_8056,N_8301);
nand U8654 (N_8654,N_8382,N_8282);
and U8655 (N_8655,N_8143,N_8465);
and U8656 (N_8656,N_8119,N_8466);
xnor U8657 (N_8657,N_8092,N_8036);
and U8658 (N_8658,N_8021,N_8204);
nand U8659 (N_8659,N_8437,N_8218);
nand U8660 (N_8660,N_8121,N_8378);
nor U8661 (N_8661,N_8089,N_8242);
or U8662 (N_8662,N_8026,N_8172);
xnor U8663 (N_8663,N_8380,N_8140);
nor U8664 (N_8664,N_8064,N_8499);
nor U8665 (N_8665,N_8224,N_8498);
and U8666 (N_8666,N_8071,N_8206);
or U8667 (N_8667,N_8115,N_8033);
and U8668 (N_8668,N_8423,N_8328);
xnor U8669 (N_8669,N_8292,N_8128);
or U8670 (N_8670,N_8385,N_8144);
or U8671 (N_8671,N_8432,N_8223);
nor U8672 (N_8672,N_8470,N_8024);
or U8673 (N_8673,N_8199,N_8221);
and U8674 (N_8674,N_8213,N_8106);
nor U8675 (N_8675,N_8491,N_8265);
nor U8676 (N_8676,N_8029,N_8413);
or U8677 (N_8677,N_8102,N_8145);
nor U8678 (N_8678,N_8175,N_8394);
nor U8679 (N_8679,N_8239,N_8312);
nand U8680 (N_8680,N_8069,N_8407);
and U8681 (N_8681,N_8364,N_8330);
and U8682 (N_8682,N_8434,N_8464);
or U8683 (N_8683,N_8300,N_8236);
xor U8684 (N_8684,N_8387,N_8005);
and U8685 (N_8685,N_8023,N_8216);
nand U8686 (N_8686,N_8118,N_8209);
nor U8687 (N_8687,N_8303,N_8359);
nand U8688 (N_8688,N_8129,N_8073);
nor U8689 (N_8689,N_8034,N_8241);
and U8690 (N_8690,N_8258,N_8447);
and U8691 (N_8691,N_8162,N_8124);
nand U8692 (N_8692,N_8234,N_8027);
nor U8693 (N_8693,N_8211,N_8332);
and U8694 (N_8694,N_8477,N_8347);
nand U8695 (N_8695,N_8076,N_8339);
and U8696 (N_8696,N_8341,N_8482);
nor U8697 (N_8697,N_8446,N_8494);
and U8698 (N_8698,N_8192,N_8249);
and U8699 (N_8699,N_8310,N_8035);
and U8700 (N_8700,N_8304,N_8357);
nand U8701 (N_8701,N_8014,N_8237);
nor U8702 (N_8702,N_8254,N_8374);
and U8703 (N_8703,N_8180,N_8331);
xnor U8704 (N_8704,N_8028,N_8381);
and U8705 (N_8705,N_8337,N_8113);
and U8706 (N_8706,N_8289,N_8181);
or U8707 (N_8707,N_8342,N_8210);
nor U8708 (N_8708,N_8287,N_8483);
nor U8709 (N_8709,N_8107,N_8421);
nand U8710 (N_8710,N_8391,N_8497);
and U8711 (N_8711,N_8496,N_8318);
xnor U8712 (N_8712,N_8019,N_8189);
nor U8713 (N_8713,N_8230,N_8435);
xor U8714 (N_8714,N_8094,N_8370);
or U8715 (N_8715,N_8087,N_8068);
or U8716 (N_8716,N_8476,N_8422);
or U8717 (N_8717,N_8479,N_8317);
nand U8718 (N_8718,N_8352,N_8151);
nor U8719 (N_8719,N_8037,N_8244);
nand U8720 (N_8720,N_8323,N_8097);
and U8721 (N_8721,N_8315,N_8295);
nand U8722 (N_8722,N_8487,N_8062);
and U8723 (N_8723,N_8399,N_8456);
or U8724 (N_8724,N_8353,N_8155);
nor U8725 (N_8725,N_8270,N_8280);
or U8726 (N_8726,N_8191,N_8131);
nor U8727 (N_8727,N_8015,N_8150);
or U8728 (N_8728,N_8444,N_8185);
and U8729 (N_8729,N_8013,N_8126);
nand U8730 (N_8730,N_8147,N_8274);
nor U8731 (N_8731,N_8157,N_8488);
nor U8732 (N_8732,N_8291,N_8452);
and U8733 (N_8733,N_8031,N_8139);
xor U8734 (N_8734,N_8276,N_8334);
or U8735 (N_8735,N_8368,N_8187);
nor U8736 (N_8736,N_8348,N_8136);
nor U8737 (N_8737,N_8490,N_8263);
or U8738 (N_8738,N_8080,N_8290);
nor U8739 (N_8739,N_8123,N_8362);
nand U8740 (N_8740,N_8438,N_8409);
nor U8741 (N_8741,N_8153,N_8198);
and U8742 (N_8742,N_8095,N_8480);
nor U8743 (N_8743,N_8205,N_8426);
xor U8744 (N_8744,N_8012,N_8275);
nor U8745 (N_8745,N_8196,N_8266);
nor U8746 (N_8746,N_8463,N_8138);
or U8747 (N_8747,N_8246,N_8010);
nor U8748 (N_8748,N_8450,N_8440);
and U8749 (N_8749,N_8158,N_8049);
nand U8750 (N_8750,N_8349,N_8459);
xnor U8751 (N_8751,N_8088,N_8193);
or U8752 (N_8752,N_8308,N_8482);
nor U8753 (N_8753,N_8028,N_8483);
nand U8754 (N_8754,N_8492,N_8244);
nor U8755 (N_8755,N_8162,N_8160);
and U8756 (N_8756,N_8425,N_8270);
nand U8757 (N_8757,N_8104,N_8118);
or U8758 (N_8758,N_8179,N_8388);
xnor U8759 (N_8759,N_8408,N_8105);
or U8760 (N_8760,N_8150,N_8347);
nand U8761 (N_8761,N_8121,N_8222);
and U8762 (N_8762,N_8017,N_8113);
or U8763 (N_8763,N_8241,N_8312);
or U8764 (N_8764,N_8434,N_8356);
or U8765 (N_8765,N_8459,N_8263);
xnor U8766 (N_8766,N_8066,N_8261);
or U8767 (N_8767,N_8252,N_8434);
and U8768 (N_8768,N_8004,N_8050);
xnor U8769 (N_8769,N_8230,N_8437);
nand U8770 (N_8770,N_8324,N_8168);
nor U8771 (N_8771,N_8448,N_8177);
and U8772 (N_8772,N_8130,N_8299);
nor U8773 (N_8773,N_8175,N_8055);
nand U8774 (N_8774,N_8117,N_8446);
or U8775 (N_8775,N_8471,N_8234);
nand U8776 (N_8776,N_8288,N_8260);
nand U8777 (N_8777,N_8388,N_8293);
nor U8778 (N_8778,N_8031,N_8040);
and U8779 (N_8779,N_8051,N_8232);
or U8780 (N_8780,N_8342,N_8284);
nand U8781 (N_8781,N_8443,N_8215);
nand U8782 (N_8782,N_8056,N_8467);
nand U8783 (N_8783,N_8221,N_8495);
nor U8784 (N_8784,N_8438,N_8456);
and U8785 (N_8785,N_8110,N_8470);
and U8786 (N_8786,N_8064,N_8085);
nor U8787 (N_8787,N_8447,N_8256);
and U8788 (N_8788,N_8275,N_8473);
and U8789 (N_8789,N_8000,N_8344);
nor U8790 (N_8790,N_8034,N_8320);
or U8791 (N_8791,N_8315,N_8417);
or U8792 (N_8792,N_8379,N_8305);
or U8793 (N_8793,N_8181,N_8454);
nand U8794 (N_8794,N_8054,N_8444);
or U8795 (N_8795,N_8393,N_8167);
xnor U8796 (N_8796,N_8153,N_8403);
nand U8797 (N_8797,N_8233,N_8048);
nand U8798 (N_8798,N_8126,N_8492);
nor U8799 (N_8799,N_8099,N_8220);
nor U8800 (N_8800,N_8338,N_8221);
xor U8801 (N_8801,N_8459,N_8229);
or U8802 (N_8802,N_8434,N_8193);
nor U8803 (N_8803,N_8476,N_8219);
or U8804 (N_8804,N_8376,N_8187);
or U8805 (N_8805,N_8399,N_8048);
xor U8806 (N_8806,N_8468,N_8180);
nor U8807 (N_8807,N_8049,N_8191);
nor U8808 (N_8808,N_8174,N_8452);
xnor U8809 (N_8809,N_8099,N_8108);
nand U8810 (N_8810,N_8356,N_8405);
xnor U8811 (N_8811,N_8429,N_8096);
xor U8812 (N_8812,N_8363,N_8141);
xnor U8813 (N_8813,N_8108,N_8141);
or U8814 (N_8814,N_8070,N_8187);
and U8815 (N_8815,N_8065,N_8016);
nand U8816 (N_8816,N_8419,N_8159);
xnor U8817 (N_8817,N_8250,N_8020);
or U8818 (N_8818,N_8245,N_8499);
and U8819 (N_8819,N_8004,N_8286);
xnor U8820 (N_8820,N_8015,N_8258);
nor U8821 (N_8821,N_8465,N_8046);
nand U8822 (N_8822,N_8403,N_8371);
nand U8823 (N_8823,N_8129,N_8231);
nand U8824 (N_8824,N_8386,N_8009);
or U8825 (N_8825,N_8249,N_8073);
nor U8826 (N_8826,N_8372,N_8229);
or U8827 (N_8827,N_8233,N_8455);
nor U8828 (N_8828,N_8189,N_8410);
or U8829 (N_8829,N_8249,N_8222);
nor U8830 (N_8830,N_8155,N_8415);
and U8831 (N_8831,N_8020,N_8311);
nor U8832 (N_8832,N_8468,N_8245);
nor U8833 (N_8833,N_8438,N_8411);
nand U8834 (N_8834,N_8028,N_8374);
or U8835 (N_8835,N_8016,N_8082);
nor U8836 (N_8836,N_8120,N_8159);
or U8837 (N_8837,N_8258,N_8427);
xor U8838 (N_8838,N_8313,N_8033);
or U8839 (N_8839,N_8377,N_8026);
or U8840 (N_8840,N_8347,N_8106);
or U8841 (N_8841,N_8326,N_8107);
nand U8842 (N_8842,N_8368,N_8083);
nor U8843 (N_8843,N_8325,N_8242);
and U8844 (N_8844,N_8229,N_8003);
and U8845 (N_8845,N_8369,N_8336);
xor U8846 (N_8846,N_8133,N_8263);
nor U8847 (N_8847,N_8320,N_8085);
nor U8848 (N_8848,N_8489,N_8460);
xnor U8849 (N_8849,N_8456,N_8361);
nor U8850 (N_8850,N_8418,N_8378);
and U8851 (N_8851,N_8129,N_8104);
xor U8852 (N_8852,N_8410,N_8135);
or U8853 (N_8853,N_8456,N_8290);
and U8854 (N_8854,N_8463,N_8343);
or U8855 (N_8855,N_8239,N_8195);
nor U8856 (N_8856,N_8380,N_8196);
nand U8857 (N_8857,N_8031,N_8360);
or U8858 (N_8858,N_8466,N_8246);
or U8859 (N_8859,N_8149,N_8471);
or U8860 (N_8860,N_8431,N_8185);
or U8861 (N_8861,N_8479,N_8213);
or U8862 (N_8862,N_8375,N_8418);
nor U8863 (N_8863,N_8294,N_8109);
and U8864 (N_8864,N_8141,N_8170);
nor U8865 (N_8865,N_8158,N_8351);
or U8866 (N_8866,N_8164,N_8101);
and U8867 (N_8867,N_8407,N_8364);
xor U8868 (N_8868,N_8302,N_8256);
and U8869 (N_8869,N_8478,N_8448);
nor U8870 (N_8870,N_8458,N_8374);
nor U8871 (N_8871,N_8272,N_8044);
xnor U8872 (N_8872,N_8143,N_8292);
and U8873 (N_8873,N_8337,N_8302);
nand U8874 (N_8874,N_8255,N_8229);
and U8875 (N_8875,N_8367,N_8177);
and U8876 (N_8876,N_8016,N_8376);
nand U8877 (N_8877,N_8288,N_8284);
or U8878 (N_8878,N_8490,N_8169);
nand U8879 (N_8879,N_8311,N_8307);
and U8880 (N_8880,N_8046,N_8073);
nor U8881 (N_8881,N_8030,N_8451);
nand U8882 (N_8882,N_8419,N_8187);
nor U8883 (N_8883,N_8464,N_8085);
nand U8884 (N_8884,N_8075,N_8485);
nand U8885 (N_8885,N_8243,N_8037);
nand U8886 (N_8886,N_8112,N_8467);
or U8887 (N_8887,N_8244,N_8491);
nor U8888 (N_8888,N_8195,N_8203);
or U8889 (N_8889,N_8047,N_8150);
and U8890 (N_8890,N_8172,N_8228);
nand U8891 (N_8891,N_8442,N_8296);
and U8892 (N_8892,N_8031,N_8493);
and U8893 (N_8893,N_8172,N_8049);
and U8894 (N_8894,N_8017,N_8405);
xor U8895 (N_8895,N_8054,N_8430);
xnor U8896 (N_8896,N_8486,N_8103);
nand U8897 (N_8897,N_8207,N_8407);
and U8898 (N_8898,N_8089,N_8494);
nand U8899 (N_8899,N_8109,N_8190);
or U8900 (N_8900,N_8427,N_8326);
nor U8901 (N_8901,N_8077,N_8234);
and U8902 (N_8902,N_8135,N_8002);
nand U8903 (N_8903,N_8009,N_8463);
nor U8904 (N_8904,N_8348,N_8118);
and U8905 (N_8905,N_8083,N_8314);
nand U8906 (N_8906,N_8130,N_8197);
xor U8907 (N_8907,N_8016,N_8239);
xnor U8908 (N_8908,N_8266,N_8486);
and U8909 (N_8909,N_8336,N_8393);
and U8910 (N_8910,N_8362,N_8035);
nor U8911 (N_8911,N_8391,N_8284);
xnor U8912 (N_8912,N_8116,N_8092);
nand U8913 (N_8913,N_8272,N_8471);
nor U8914 (N_8914,N_8299,N_8026);
nor U8915 (N_8915,N_8089,N_8135);
or U8916 (N_8916,N_8356,N_8208);
nand U8917 (N_8917,N_8069,N_8436);
nor U8918 (N_8918,N_8349,N_8397);
nand U8919 (N_8919,N_8409,N_8458);
and U8920 (N_8920,N_8206,N_8211);
and U8921 (N_8921,N_8383,N_8337);
nand U8922 (N_8922,N_8178,N_8331);
or U8923 (N_8923,N_8037,N_8315);
nor U8924 (N_8924,N_8232,N_8454);
nor U8925 (N_8925,N_8258,N_8087);
nor U8926 (N_8926,N_8020,N_8346);
and U8927 (N_8927,N_8480,N_8208);
and U8928 (N_8928,N_8488,N_8366);
nand U8929 (N_8929,N_8071,N_8046);
and U8930 (N_8930,N_8396,N_8083);
nor U8931 (N_8931,N_8436,N_8206);
nor U8932 (N_8932,N_8278,N_8398);
and U8933 (N_8933,N_8197,N_8160);
or U8934 (N_8934,N_8158,N_8331);
and U8935 (N_8935,N_8003,N_8043);
and U8936 (N_8936,N_8168,N_8204);
or U8937 (N_8937,N_8176,N_8451);
or U8938 (N_8938,N_8020,N_8251);
and U8939 (N_8939,N_8468,N_8496);
or U8940 (N_8940,N_8368,N_8459);
and U8941 (N_8941,N_8027,N_8291);
nor U8942 (N_8942,N_8347,N_8210);
or U8943 (N_8943,N_8344,N_8268);
or U8944 (N_8944,N_8125,N_8372);
or U8945 (N_8945,N_8121,N_8139);
and U8946 (N_8946,N_8055,N_8066);
nor U8947 (N_8947,N_8079,N_8253);
nor U8948 (N_8948,N_8036,N_8055);
or U8949 (N_8949,N_8034,N_8021);
and U8950 (N_8950,N_8430,N_8163);
and U8951 (N_8951,N_8094,N_8416);
and U8952 (N_8952,N_8038,N_8006);
and U8953 (N_8953,N_8359,N_8014);
nor U8954 (N_8954,N_8271,N_8070);
nor U8955 (N_8955,N_8227,N_8458);
nand U8956 (N_8956,N_8000,N_8014);
nand U8957 (N_8957,N_8288,N_8196);
nand U8958 (N_8958,N_8179,N_8481);
nand U8959 (N_8959,N_8321,N_8428);
xor U8960 (N_8960,N_8073,N_8357);
nand U8961 (N_8961,N_8454,N_8405);
and U8962 (N_8962,N_8422,N_8090);
and U8963 (N_8963,N_8410,N_8004);
nor U8964 (N_8964,N_8374,N_8307);
or U8965 (N_8965,N_8379,N_8495);
nor U8966 (N_8966,N_8210,N_8316);
nor U8967 (N_8967,N_8296,N_8104);
nor U8968 (N_8968,N_8363,N_8371);
nand U8969 (N_8969,N_8175,N_8207);
or U8970 (N_8970,N_8380,N_8041);
nand U8971 (N_8971,N_8396,N_8224);
and U8972 (N_8972,N_8005,N_8018);
or U8973 (N_8973,N_8120,N_8433);
nand U8974 (N_8974,N_8173,N_8160);
and U8975 (N_8975,N_8369,N_8247);
nor U8976 (N_8976,N_8004,N_8344);
nor U8977 (N_8977,N_8286,N_8439);
or U8978 (N_8978,N_8490,N_8025);
or U8979 (N_8979,N_8449,N_8439);
and U8980 (N_8980,N_8119,N_8051);
xnor U8981 (N_8981,N_8211,N_8446);
or U8982 (N_8982,N_8333,N_8378);
nor U8983 (N_8983,N_8451,N_8395);
nor U8984 (N_8984,N_8037,N_8279);
or U8985 (N_8985,N_8477,N_8428);
nand U8986 (N_8986,N_8120,N_8201);
and U8987 (N_8987,N_8322,N_8469);
nor U8988 (N_8988,N_8385,N_8020);
nor U8989 (N_8989,N_8363,N_8008);
and U8990 (N_8990,N_8077,N_8052);
nor U8991 (N_8991,N_8418,N_8435);
nand U8992 (N_8992,N_8178,N_8316);
nand U8993 (N_8993,N_8203,N_8209);
or U8994 (N_8994,N_8043,N_8168);
or U8995 (N_8995,N_8444,N_8220);
nor U8996 (N_8996,N_8200,N_8276);
nand U8997 (N_8997,N_8260,N_8270);
or U8998 (N_8998,N_8428,N_8015);
and U8999 (N_8999,N_8173,N_8473);
nor U9000 (N_9000,N_8613,N_8889);
nor U9001 (N_9001,N_8706,N_8587);
xor U9002 (N_9002,N_8981,N_8841);
xor U9003 (N_9003,N_8540,N_8669);
nor U9004 (N_9004,N_8594,N_8945);
or U9005 (N_9005,N_8748,N_8609);
and U9006 (N_9006,N_8678,N_8656);
and U9007 (N_9007,N_8936,N_8529);
nand U9008 (N_9008,N_8700,N_8780);
and U9009 (N_9009,N_8689,N_8568);
nand U9010 (N_9010,N_8640,N_8652);
nand U9011 (N_9011,N_8588,N_8851);
and U9012 (N_9012,N_8768,N_8733);
xnor U9013 (N_9013,N_8663,N_8525);
nor U9014 (N_9014,N_8759,N_8682);
and U9015 (N_9015,N_8893,N_8809);
nand U9016 (N_9016,N_8541,N_8967);
xnor U9017 (N_9017,N_8859,N_8964);
and U9018 (N_9018,N_8918,N_8935);
nor U9019 (N_9019,N_8581,N_8986);
or U9020 (N_9020,N_8886,N_8504);
or U9021 (N_9021,N_8726,N_8951);
or U9022 (N_9022,N_8840,N_8947);
nor U9023 (N_9023,N_8846,N_8916);
or U9024 (N_9024,N_8801,N_8815);
and U9025 (N_9025,N_8771,N_8928);
nor U9026 (N_9026,N_8731,N_8677);
nor U9027 (N_9027,N_8546,N_8533);
and U9028 (N_9028,N_8501,N_8969);
and U9029 (N_9029,N_8585,N_8575);
nand U9030 (N_9030,N_8686,N_8775);
or U9031 (N_9031,N_8752,N_8921);
or U9032 (N_9032,N_8881,N_8853);
nor U9033 (N_9033,N_8572,N_8611);
and U9034 (N_9034,N_8802,N_8625);
and U9035 (N_9035,N_8576,N_8646);
or U9036 (N_9036,N_8794,N_8531);
nand U9037 (N_9037,N_8719,N_8976);
nand U9038 (N_9038,N_8522,N_8797);
and U9039 (N_9039,N_8645,N_8852);
nor U9040 (N_9040,N_8811,N_8792);
and U9041 (N_9041,N_8612,N_8922);
nand U9042 (N_9042,N_8858,N_8778);
and U9043 (N_9043,N_8503,N_8785);
or U9044 (N_9044,N_8866,N_8997);
nor U9045 (N_9045,N_8972,N_8627);
and U9046 (N_9046,N_8683,N_8740);
or U9047 (N_9047,N_8717,N_8790);
nor U9048 (N_9048,N_8992,N_8774);
or U9049 (N_9049,N_8598,N_8791);
xnor U9050 (N_9050,N_8562,N_8749);
or U9051 (N_9051,N_8849,N_8615);
or U9052 (N_9052,N_8738,N_8620);
or U9053 (N_9053,N_8746,N_8532);
xnor U9054 (N_9054,N_8696,N_8855);
and U9055 (N_9055,N_8679,N_8716);
nand U9056 (N_9056,N_8727,N_8665);
nand U9057 (N_9057,N_8755,N_8825);
nand U9058 (N_9058,N_8667,N_8834);
nor U9059 (N_9059,N_8763,N_8655);
or U9060 (N_9060,N_8590,N_8711);
nor U9061 (N_9061,N_8699,N_8956);
or U9062 (N_9062,N_8984,N_8550);
nor U9063 (N_9063,N_8751,N_8897);
nor U9064 (N_9064,N_8545,N_8933);
or U9065 (N_9065,N_8870,N_8596);
nor U9066 (N_9066,N_8728,N_8556);
or U9067 (N_9067,N_8579,N_8597);
or U9068 (N_9068,N_8616,N_8779);
or U9069 (N_9069,N_8966,N_8900);
nand U9070 (N_9070,N_8657,N_8534);
xor U9071 (N_9071,N_8691,N_8906);
nand U9072 (N_9072,N_8917,N_8993);
nand U9073 (N_9073,N_8694,N_8567);
nand U9074 (N_9074,N_8549,N_8837);
nor U9075 (N_9075,N_8676,N_8784);
nor U9076 (N_9076,N_8629,N_8680);
nand U9077 (N_9077,N_8898,N_8845);
nor U9078 (N_9078,N_8807,N_8970);
or U9079 (N_9079,N_8542,N_8685);
nor U9080 (N_9080,N_8745,N_8560);
nor U9081 (N_9081,N_8661,N_8944);
or U9082 (N_9082,N_8637,N_8701);
and U9083 (N_9083,N_8658,N_8919);
and U9084 (N_9084,N_8994,N_8985);
or U9085 (N_9085,N_8589,N_8754);
or U9086 (N_9086,N_8712,N_8631);
nor U9087 (N_9087,N_8907,N_8729);
nand U9088 (N_9088,N_8724,N_8765);
and U9089 (N_9089,N_8979,N_8662);
nand U9090 (N_9090,N_8543,N_8982);
and U9091 (N_9091,N_8630,N_8887);
and U9092 (N_9092,N_8538,N_8618);
nand U9093 (N_9093,N_8721,N_8803);
nand U9094 (N_9094,N_8650,N_8806);
nor U9095 (N_9095,N_8583,N_8571);
xnor U9096 (N_9096,N_8702,N_8563);
and U9097 (N_9097,N_8939,N_8693);
nand U9098 (N_9098,N_8995,N_8737);
nor U9099 (N_9099,N_8674,N_8632);
xnor U9100 (N_9100,N_8660,N_8914);
and U9101 (N_9101,N_8783,N_8757);
nor U9102 (N_9102,N_8843,N_8805);
and U9103 (N_9103,N_8842,N_8684);
nor U9104 (N_9104,N_8690,N_8800);
and U9105 (N_9105,N_8564,N_8924);
nand U9106 (N_9106,N_8848,N_8938);
and U9107 (N_9107,N_8910,N_8518);
and U9108 (N_9108,N_8715,N_8566);
nor U9109 (N_9109,N_8673,N_8789);
and U9110 (N_9110,N_8633,N_8987);
or U9111 (N_9111,N_8623,N_8808);
xor U9112 (N_9112,N_8582,N_8890);
and U9113 (N_9113,N_8742,N_8856);
or U9114 (N_9114,N_8988,N_8941);
or U9115 (N_9115,N_8732,N_8978);
or U9116 (N_9116,N_8718,N_8530);
xor U9117 (N_9117,N_8810,N_8653);
nor U9118 (N_9118,N_8758,N_8876);
xnor U9119 (N_9119,N_8998,N_8980);
nor U9120 (N_9120,N_8601,N_8735);
or U9121 (N_9121,N_8832,N_8777);
nor U9122 (N_9122,N_8868,N_8904);
nor U9123 (N_9123,N_8912,N_8819);
nand U9124 (N_9124,N_8607,N_8734);
and U9125 (N_9125,N_8520,N_8844);
nor U9126 (N_9126,N_8670,N_8593);
nand U9127 (N_9127,N_8547,N_8750);
and U9128 (N_9128,N_8570,N_8644);
and U9129 (N_9129,N_8824,N_8603);
and U9130 (N_9130,N_8999,N_8864);
nor U9131 (N_9131,N_8595,N_8707);
or U9132 (N_9132,N_8880,N_8926);
or U9133 (N_9133,N_8574,N_8517);
nand U9134 (N_9134,N_8511,N_8884);
or U9135 (N_9135,N_8641,N_8854);
and U9136 (N_9136,N_8821,N_8879);
nand U9137 (N_9137,N_8920,N_8833);
nor U9138 (N_9138,N_8705,N_8602);
nand U9139 (N_9139,N_8599,N_8867);
nand U9140 (N_9140,N_8692,N_8513);
nor U9141 (N_9141,N_8923,N_8882);
nand U9142 (N_9142,N_8796,N_8622);
nand U9143 (N_9143,N_8666,N_8537);
and U9144 (N_9144,N_8558,N_8708);
and U9145 (N_9145,N_8799,N_8903);
or U9146 (N_9146,N_8638,N_8515);
or U9147 (N_9147,N_8937,N_8787);
or U9148 (N_9148,N_8872,N_8766);
nand U9149 (N_9149,N_8929,N_8739);
nor U9150 (N_9150,N_8839,N_8955);
and U9151 (N_9151,N_8552,N_8559);
and U9152 (N_9152,N_8639,N_8836);
or U9153 (N_9153,N_8888,N_8996);
xor U9154 (N_9154,N_8857,N_8703);
nand U9155 (N_9155,N_8909,N_8514);
and U9156 (N_9156,N_8899,N_8744);
and U9157 (N_9157,N_8949,N_8863);
nor U9158 (N_9158,N_8647,N_8636);
nand U9159 (N_9159,N_8814,N_8505);
and U9160 (N_9160,N_8643,N_8901);
nor U9161 (N_9161,N_8672,N_8827);
nand U9162 (N_9162,N_8905,N_8974);
or U9163 (N_9163,N_8885,N_8695);
or U9164 (N_9164,N_8990,N_8830);
or U9165 (N_9165,N_8942,N_8526);
nand U9166 (N_9166,N_8770,N_8975);
nor U9167 (N_9167,N_8592,N_8756);
and U9168 (N_9168,N_8730,N_8911);
and U9169 (N_9169,N_8930,N_8681);
or U9170 (N_9170,N_8826,N_8776);
nand U9171 (N_9171,N_8971,N_8753);
or U9172 (N_9172,N_8831,N_8519);
xor U9173 (N_9173,N_8961,N_8878);
or U9174 (N_9174,N_8604,N_8621);
nor U9175 (N_9175,N_8877,N_8769);
nor U9176 (N_9176,N_8506,N_8835);
and U9177 (N_9177,N_8772,N_8829);
or U9178 (N_9178,N_8940,N_8606);
nand U9179 (N_9179,N_8687,N_8816);
xor U9180 (N_9180,N_8795,N_8989);
or U9181 (N_9181,N_8817,N_8932);
nor U9182 (N_9182,N_8931,N_8654);
and U9183 (N_9183,N_8786,N_8516);
nor U9184 (N_9184,N_8600,N_8713);
and U9185 (N_9185,N_8675,N_8894);
xor U9186 (N_9186,N_8704,N_8895);
and U9187 (N_9187,N_8617,N_8523);
or U9188 (N_9188,N_8722,N_8577);
nor U9189 (N_9189,N_8862,N_8710);
nor U9190 (N_9190,N_8913,N_8813);
and U9191 (N_9191,N_8861,N_8965);
xnor U9192 (N_9192,N_8883,N_8747);
nand U9193 (N_9193,N_8902,N_8502);
nand U9194 (N_9194,N_8957,N_8544);
nor U9195 (N_9195,N_8874,N_8714);
xor U9196 (N_9196,N_8548,N_8512);
xor U9197 (N_9197,N_8962,N_8820);
xor U9198 (N_9198,N_8698,N_8952);
and U9199 (N_9199,N_8635,N_8578);
xnor U9200 (N_9200,N_8983,N_8565);
or U9201 (N_9201,N_8555,N_8950);
and U9202 (N_9202,N_8508,N_8973);
nand U9203 (N_9203,N_8850,N_8838);
or U9204 (N_9204,N_8723,N_8960);
nand U9205 (N_9205,N_8892,N_8628);
or U9206 (N_9206,N_8709,N_8948);
nor U9207 (N_9207,N_8925,N_8891);
and U9208 (N_9208,N_8573,N_8963);
nand U9209 (N_9209,N_8605,N_8865);
nor U9210 (N_9210,N_8847,N_8697);
nand U9211 (N_9211,N_8688,N_8659);
or U9212 (N_9212,N_8509,N_8619);
nor U9213 (N_9213,N_8812,N_8507);
or U9214 (N_9214,N_8569,N_8580);
nand U9215 (N_9215,N_8736,N_8557);
nand U9216 (N_9216,N_8943,N_8968);
nand U9217 (N_9217,N_8720,N_8610);
nand U9218 (N_9218,N_8927,N_8954);
or U9219 (N_9219,N_8584,N_8591);
nor U9220 (N_9220,N_8991,N_8608);
and U9221 (N_9221,N_8510,N_8934);
nand U9222 (N_9222,N_8528,N_8818);
nand U9223 (N_9223,N_8551,N_8767);
or U9224 (N_9224,N_8760,N_8782);
nor U9225 (N_9225,N_8649,N_8761);
or U9226 (N_9226,N_8959,N_8664);
and U9227 (N_9227,N_8822,N_8614);
nor U9228 (N_9228,N_8860,N_8648);
and U9229 (N_9229,N_8977,N_8741);
nor U9230 (N_9230,N_8671,N_8743);
xnor U9231 (N_9231,N_8554,N_8946);
nand U9232 (N_9232,N_8871,N_8553);
or U9233 (N_9233,N_8793,N_8668);
nor U9234 (N_9234,N_8524,N_8642);
or U9235 (N_9235,N_8958,N_8536);
nand U9236 (N_9236,N_8798,N_8873);
nor U9237 (N_9237,N_8651,N_8626);
and U9238 (N_9238,N_8896,N_8788);
xnor U9239 (N_9239,N_8869,N_8953);
or U9240 (N_9240,N_8634,N_8773);
nand U9241 (N_9241,N_8875,N_8915);
nand U9242 (N_9242,N_8764,N_8586);
nor U9243 (N_9243,N_8828,N_8521);
and U9244 (N_9244,N_8908,N_8500);
or U9245 (N_9245,N_8804,N_8823);
xnor U9246 (N_9246,N_8725,N_8781);
and U9247 (N_9247,N_8535,N_8624);
and U9248 (N_9248,N_8527,N_8561);
and U9249 (N_9249,N_8762,N_8539);
or U9250 (N_9250,N_8537,N_8629);
nand U9251 (N_9251,N_8638,N_8766);
nor U9252 (N_9252,N_8622,N_8968);
or U9253 (N_9253,N_8535,N_8618);
nand U9254 (N_9254,N_8734,N_8599);
nand U9255 (N_9255,N_8831,N_8814);
or U9256 (N_9256,N_8987,N_8853);
and U9257 (N_9257,N_8857,N_8886);
nand U9258 (N_9258,N_8837,N_8687);
nor U9259 (N_9259,N_8556,N_8697);
or U9260 (N_9260,N_8644,N_8792);
or U9261 (N_9261,N_8771,N_8909);
nor U9262 (N_9262,N_8897,N_8788);
or U9263 (N_9263,N_8524,N_8823);
nand U9264 (N_9264,N_8509,N_8755);
and U9265 (N_9265,N_8599,N_8528);
nor U9266 (N_9266,N_8605,N_8813);
nor U9267 (N_9267,N_8623,N_8842);
or U9268 (N_9268,N_8908,N_8709);
xnor U9269 (N_9269,N_8511,N_8590);
nand U9270 (N_9270,N_8612,N_8972);
nor U9271 (N_9271,N_8945,N_8729);
and U9272 (N_9272,N_8665,N_8728);
nor U9273 (N_9273,N_8807,N_8609);
or U9274 (N_9274,N_8793,N_8788);
or U9275 (N_9275,N_8675,N_8767);
nor U9276 (N_9276,N_8743,N_8919);
nor U9277 (N_9277,N_8893,N_8598);
and U9278 (N_9278,N_8963,N_8833);
nand U9279 (N_9279,N_8924,N_8585);
nor U9280 (N_9280,N_8879,N_8677);
nand U9281 (N_9281,N_8673,N_8917);
nand U9282 (N_9282,N_8758,N_8777);
or U9283 (N_9283,N_8799,N_8520);
or U9284 (N_9284,N_8640,N_8566);
nor U9285 (N_9285,N_8550,N_8565);
xnor U9286 (N_9286,N_8627,N_8509);
xor U9287 (N_9287,N_8629,N_8998);
and U9288 (N_9288,N_8675,N_8786);
nand U9289 (N_9289,N_8790,N_8585);
nand U9290 (N_9290,N_8666,N_8863);
or U9291 (N_9291,N_8552,N_8609);
nor U9292 (N_9292,N_8542,N_8971);
and U9293 (N_9293,N_8844,N_8595);
or U9294 (N_9294,N_8628,N_8669);
nor U9295 (N_9295,N_8645,N_8854);
xor U9296 (N_9296,N_8682,N_8805);
xnor U9297 (N_9297,N_8878,N_8935);
nand U9298 (N_9298,N_8525,N_8620);
and U9299 (N_9299,N_8859,N_8762);
nand U9300 (N_9300,N_8836,N_8676);
nor U9301 (N_9301,N_8996,N_8533);
nor U9302 (N_9302,N_8563,N_8643);
nand U9303 (N_9303,N_8684,N_8932);
or U9304 (N_9304,N_8737,N_8776);
and U9305 (N_9305,N_8611,N_8597);
or U9306 (N_9306,N_8801,N_8973);
nand U9307 (N_9307,N_8920,N_8883);
or U9308 (N_9308,N_8591,N_8658);
and U9309 (N_9309,N_8882,N_8693);
nand U9310 (N_9310,N_8531,N_8760);
nor U9311 (N_9311,N_8897,N_8764);
nand U9312 (N_9312,N_8699,N_8534);
nand U9313 (N_9313,N_8536,N_8557);
and U9314 (N_9314,N_8524,N_8544);
or U9315 (N_9315,N_8886,N_8601);
nor U9316 (N_9316,N_8507,N_8844);
and U9317 (N_9317,N_8555,N_8802);
nand U9318 (N_9318,N_8921,N_8861);
or U9319 (N_9319,N_8947,N_8896);
nand U9320 (N_9320,N_8729,N_8625);
or U9321 (N_9321,N_8594,N_8694);
nand U9322 (N_9322,N_8645,N_8751);
xnor U9323 (N_9323,N_8955,N_8517);
or U9324 (N_9324,N_8518,N_8857);
nand U9325 (N_9325,N_8881,N_8889);
or U9326 (N_9326,N_8544,N_8901);
nand U9327 (N_9327,N_8896,N_8911);
and U9328 (N_9328,N_8970,N_8828);
nand U9329 (N_9329,N_8734,N_8801);
or U9330 (N_9330,N_8739,N_8954);
xor U9331 (N_9331,N_8614,N_8599);
nand U9332 (N_9332,N_8774,N_8552);
and U9333 (N_9333,N_8957,N_8770);
and U9334 (N_9334,N_8992,N_8654);
and U9335 (N_9335,N_8675,N_8567);
xor U9336 (N_9336,N_8802,N_8703);
nor U9337 (N_9337,N_8870,N_8893);
nand U9338 (N_9338,N_8544,N_8984);
xnor U9339 (N_9339,N_8507,N_8632);
or U9340 (N_9340,N_8913,N_8968);
or U9341 (N_9341,N_8614,N_8721);
nor U9342 (N_9342,N_8580,N_8883);
or U9343 (N_9343,N_8971,N_8675);
or U9344 (N_9344,N_8933,N_8672);
nor U9345 (N_9345,N_8795,N_8632);
nand U9346 (N_9346,N_8583,N_8726);
nor U9347 (N_9347,N_8543,N_8814);
nor U9348 (N_9348,N_8887,N_8970);
nor U9349 (N_9349,N_8517,N_8633);
nor U9350 (N_9350,N_8976,N_8946);
or U9351 (N_9351,N_8763,N_8934);
and U9352 (N_9352,N_8543,N_8693);
nand U9353 (N_9353,N_8695,N_8775);
or U9354 (N_9354,N_8538,N_8894);
nand U9355 (N_9355,N_8975,N_8593);
nor U9356 (N_9356,N_8684,N_8931);
or U9357 (N_9357,N_8780,N_8881);
nor U9358 (N_9358,N_8956,N_8597);
and U9359 (N_9359,N_8760,N_8920);
xnor U9360 (N_9360,N_8762,N_8601);
or U9361 (N_9361,N_8578,N_8716);
or U9362 (N_9362,N_8658,N_8818);
or U9363 (N_9363,N_8966,N_8626);
nor U9364 (N_9364,N_8597,N_8863);
nand U9365 (N_9365,N_8956,N_8919);
nor U9366 (N_9366,N_8964,N_8825);
nand U9367 (N_9367,N_8538,N_8660);
and U9368 (N_9368,N_8687,N_8582);
and U9369 (N_9369,N_8644,N_8725);
nand U9370 (N_9370,N_8988,N_8916);
nor U9371 (N_9371,N_8562,N_8806);
or U9372 (N_9372,N_8510,N_8628);
xnor U9373 (N_9373,N_8828,N_8822);
nor U9374 (N_9374,N_8867,N_8733);
and U9375 (N_9375,N_8543,N_8798);
and U9376 (N_9376,N_8533,N_8581);
nor U9377 (N_9377,N_8751,N_8823);
and U9378 (N_9378,N_8622,N_8915);
and U9379 (N_9379,N_8695,N_8581);
or U9380 (N_9380,N_8665,N_8642);
nor U9381 (N_9381,N_8792,N_8861);
nor U9382 (N_9382,N_8821,N_8766);
or U9383 (N_9383,N_8541,N_8610);
and U9384 (N_9384,N_8963,N_8893);
nor U9385 (N_9385,N_8832,N_8850);
xor U9386 (N_9386,N_8991,N_8809);
and U9387 (N_9387,N_8583,N_8840);
or U9388 (N_9388,N_8782,N_8792);
or U9389 (N_9389,N_8520,N_8784);
or U9390 (N_9390,N_8847,N_8538);
nor U9391 (N_9391,N_8645,N_8792);
and U9392 (N_9392,N_8601,N_8840);
nand U9393 (N_9393,N_8830,N_8587);
nor U9394 (N_9394,N_8531,N_8514);
or U9395 (N_9395,N_8528,N_8993);
nor U9396 (N_9396,N_8957,N_8912);
or U9397 (N_9397,N_8725,N_8633);
and U9398 (N_9398,N_8684,N_8663);
and U9399 (N_9399,N_8516,N_8840);
xor U9400 (N_9400,N_8955,N_8620);
nor U9401 (N_9401,N_8746,N_8981);
nand U9402 (N_9402,N_8966,N_8601);
nand U9403 (N_9403,N_8717,N_8876);
and U9404 (N_9404,N_8942,N_8692);
nor U9405 (N_9405,N_8706,N_8790);
or U9406 (N_9406,N_8552,N_8878);
xor U9407 (N_9407,N_8577,N_8524);
nand U9408 (N_9408,N_8742,N_8841);
or U9409 (N_9409,N_8612,N_8516);
nand U9410 (N_9410,N_8729,N_8879);
nand U9411 (N_9411,N_8582,N_8549);
or U9412 (N_9412,N_8902,N_8935);
or U9413 (N_9413,N_8640,N_8879);
and U9414 (N_9414,N_8587,N_8501);
and U9415 (N_9415,N_8870,N_8915);
nor U9416 (N_9416,N_8535,N_8952);
and U9417 (N_9417,N_8844,N_8687);
nor U9418 (N_9418,N_8832,N_8587);
and U9419 (N_9419,N_8840,N_8785);
nor U9420 (N_9420,N_8555,N_8890);
or U9421 (N_9421,N_8724,N_8872);
nor U9422 (N_9422,N_8735,N_8923);
or U9423 (N_9423,N_8882,N_8998);
or U9424 (N_9424,N_8903,N_8730);
or U9425 (N_9425,N_8649,N_8608);
and U9426 (N_9426,N_8563,N_8780);
nand U9427 (N_9427,N_8601,N_8752);
and U9428 (N_9428,N_8698,N_8887);
or U9429 (N_9429,N_8689,N_8544);
nor U9430 (N_9430,N_8673,N_8644);
nand U9431 (N_9431,N_8536,N_8863);
and U9432 (N_9432,N_8507,N_8769);
nor U9433 (N_9433,N_8645,N_8679);
xnor U9434 (N_9434,N_8929,N_8975);
and U9435 (N_9435,N_8655,N_8504);
nor U9436 (N_9436,N_8888,N_8773);
and U9437 (N_9437,N_8606,N_8777);
xor U9438 (N_9438,N_8957,N_8946);
nand U9439 (N_9439,N_8984,N_8980);
nor U9440 (N_9440,N_8890,N_8857);
or U9441 (N_9441,N_8795,N_8700);
or U9442 (N_9442,N_8787,N_8751);
and U9443 (N_9443,N_8829,N_8846);
nor U9444 (N_9444,N_8625,N_8665);
xnor U9445 (N_9445,N_8745,N_8746);
xnor U9446 (N_9446,N_8900,N_8798);
and U9447 (N_9447,N_8866,N_8955);
or U9448 (N_9448,N_8649,N_8859);
nor U9449 (N_9449,N_8750,N_8590);
or U9450 (N_9450,N_8925,N_8775);
and U9451 (N_9451,N_8647,N_8993);
nor U9452 (N_9452,N_8685,N_8982);
or U9453 (N_9453,N_8618,N_8951);
and U9454 (N_9454,N_8869,N_8923);
nor U9455 (N_9455,N_8653,N_8823);
and U9456 (N_9456,N_8902,N_8940);
and U9457 (N_9457,N_8829,N_8632);
or U9458 (N_9458,N_8700,N_8672);
or U9459 (N_9459,N_8619,N_8694);
and U9460 (N_9460,N_8526,N_8889);
nor U9461 (N_9461,N_8917,N_8994);
or U9462 (N_9462,N_8844,N_8636);
nor U9463 (N_9463,N_8727,N_8723);
nand U9464 (N_9464,N_8589,N_8622);
nor U9465 (N_9465,N_8719,N_8528);
nand U9466 (N_9466,N_8797,N_8519);
or U9467 (N_9467,N_8981,N_8827);
or U9468 (N_9468,N_8664,N_8573);
nand U9469 (N_9469,N_8879,N_8652);
xor U9470 (N_9470,N_8874,N_8536);
and U9471 (N_9471,N_8888,N_8721);
xor U9472 (N_9472,N_8683,N_8717);
nor U9473 (N_9473,N_8693,N_8675);
and U9474 (N_9474,N_8656,N_8644);
nand U9475 (N_9475,N_8599,N_8653);
nand U9476 (N_9476,N_8896,N_8523);
or U9477 (N_9477,N_8973,N_8962);
and U9478 (N_9478,N_8617,N_8749);
and U9479 (N_9479,N_8638,N_8842);
and U9480 (N_9480,N_8625,N_8837);
nor U9481 (N_9481,N_8547,N_8650);
and U9482 (N_9482,N_8966,N_8854);
or U9483 (N_9483,N_8821,N_8638);
nand U9484 (N_9484,N_8528,N_8873);
or U9485 (N_9485,N_8516,N_8727);
or U9486 (N_9486,N_8933,N_8785);
and U9487 (N_9487,N_8788,N_8512);
nand U9488 (N_9488,N_8710,N_8571);
or U9489 (N_9489,N_8993,N_8522);
nor U9490 (N_9490,N_8801,N_8597);
and U9491 (N_9491,N_8698,N_8896);
nor U9492 (N_9492,N_8972,N_8772);
and U9493 (N_9493,N_8922,N_8501);
nand U9494 (N_9494,N_8509,N_8830);
and U9495 (N_9495,N_8521,N_8618);
and U9496 (N_9496,N_8891,N_8836);
nand U9497 (N_9497,N_8651,N_8505);
and U9498 (N_9498,N_8877,N_8655);
or U9499 (N_9499,N_8692,N_8969);
and U9500 (N_9500,N_9113,N_9381);
nor U9501 (N_9501,N_9120,N_9468);
or U9502 (N_9502,N_9329,N_9221);
nand U9503 (N_9503,N_9057,N_9379);
nor U9504 (N_9504,N_9439,N_9480);
or U9505 (N_9505,N_9376,N_9141);
or U9506 (N_9506,N_9344,N_9301);
nor U9507 (N_9507,N_9055,N_9046);
or U9508 (N_9508,N_9024,N_9089);
or U9509 (N_9509,N_9304,N_9289);
or U9510 (N_9510,N_9297,N_9119);
or U9511 (N_9511,N_9006,N_9201);
xnor U9512 (N_9512,N_9404,N_9343);
nor U9513 (N_9513,N_9281,N_9125);
or U9514 (N_9514,N_9476,N_9064);
and U9515 (N_9515,N_9163,N_9261);
nand U9516 (N_9516,N_9422,N_9446);
xnor U9517 (N_9517,N_9455,N_9019);
and U9518 (N_9518,N_9160,N_9454);
or U9519 (N_9519,N_9430,N_9410);
nor U9520 (N_9520,N_9115,N_9276);
nor U9521 (N_9521,N_9168,N_9274);
or U9522 (N_9522,N_9017,N_9239);
nor U9523 (N_9523,N_9365,N_9101);
or U9524 (N_9524,N_9429,N_9083);
xor U9525 (N_9525,N_9490,N_9292);
or U9526 (N_9526,N_9189,N_9387);
nand U9527 (N_9527,N_9037,N_9090);
or U9528 (N_9528,N_9245,N_9073);
nor U9529 (N_9529,N_9194,N_9009);
xor U9530 (N_9530,N_9440,N_9445);
nand U9531 (N_9531,N_9025,N_9075);
nand U9532 (N_9532,N_9299,N_9317);
or U9533 (N_9533,N_9449,N_9129);
nor U9534 (N_9534,N_9045,N_9155);
or U9535 (N_9535,N_9023,N_9103);
and U9536 (N_9536,N_9296,N_9032);
nand U9537 (N_9537,N_9213,N_9268);
nor U9538 (N_9538,N_9059,N_9166);
or U9539 (N_9539,N_9177,N_9408);
xnor U9540 (N_9540,N_9114,N_9345);
xor U9541 (N_9541,N_9054,N_9363);
or U9542 (N_9542,N_9362,N_9411);
nor U9543 (N_9543,N_9080,N_9104);
and U9544 (N_9544,N_9076,N_9447);
and U9545 (N_9545,N_9386,N_9259);
or U9546 (N_9546,N_9298,N_9224);
or U9547 (N_9547,N_9203,N_9328);
nand U9548 (N_9548,N_9414,N_9402);
nand U9549 (N_9549,N_9403,N_9242);
nand U9550 (N_9550,N_9173,N_9491);
or U9551 (N_9551,N_9319,N_9007);
xor U9552 (N_9552,N_9012,N_9358);
nor U9553 (N_9553,N_9167,N_9091);
and U9554 (N_9554,N_9196,N_9269);
nand U9555 (N_9555,N_9035,N_9394);
or U9556 (N_9556,N_9336,N_9378);
nand U9557 (N_9557,N_9033,N_9367);
nor U9558 (N_9558,N_9159,N_9240);
and U9559 (N_9559,N_9324,N_9058);
and U9560 (N_9560,N_9198,N_9353);
or U9561 (N_9561,N_9244,N_9066);
nor U9562 (N_9562,N_9249,N_9197);
xor U9563 (N_9563,N_9005,N_9275);
or U9564 (N_9564,N_9313,N_9279);
nor U9565 (N_9565,N_9265,N_9121);
or U9566 (N_9566,N_9392,N_9493);
xnor U9567 (N_9567,N_9099,N_9172);
or U9568 (N_9568,N_9337,N_9234);
nand U9569 (N_9569,N_9342,N_9288);
nand U9570 (N_9570,N_9456,N_9406);
or U9571 (N_9571,N_9095,N_9383);
or U9572 (N_9572,N_9047,N_9305);
nand U9573 (N_9573,N_9397,N_9157);
and U9574 (N_9574,N_9217,N_9021);
or U9575 (N_9575,N_9088,N_9195);
and U9576 (N_9576,N_9443,N_9393);
and U9577 (N_9577,N_9246,N_9149);
or U9578 (N_9578,N_9056,N_9048);
nand U9579 (N_9579,N_9001,N_9357);
xnor U9580 (N_9580,N_9013,N_9418);
nand U9581 (N_9581,N_9098,N_9235);
nor U9582 (N_9582,N_9368,N_9206);
xnor U9583 (N_9583,N_9228,N_9042);
or U9584 (N_9584,N_9388,N_9222);
and U9585 (N_9585,N_9251,N_9038);
or U9586 (N_9586,N_9465,N_9175);
nand U9587 (N_9587,N_9417,N_9267);
or U9588 (N_9588,N_9034,N_9231);
nand U9589 (N_9589,N_9109,N_9263);
or U9590 (N_9590,N_9286,N_9327);
nand U9591 (N_9591,N_9079,N_9134);
and U9592 (N_9592,N_9294,N_9110);
nor U9593 (N_9593,N_9105,N_9131);
nor U9594 (N_9594,N_9291,N_9499);
xnor U9595 (N_9595,N_9232,N_9252);
nor U9596 (N_9596,N_9052,N_9295);
nor U9597 (N_9597,N_9212,N_9225);
and U9598 (N_9598,N_9280,N_9302);
and U9599 (N_9599,N_9060,N_9085);
nor U9600 (N_9600,N_9000,N_9022);
nand U9601 (N_9601,N_9028,N_9176);
nor U9602 (N_9602,N_9136,N_9433);
and U9603 (N_9603,N_9184,N_9477);
nand U9604 (N_9604,N_9264,N_9472);
xnor U9605 (N_9605,N_9325,N_9162);
and U9606 (N_9606,N_9338,N_9179);
nor U9607 (N_9607,N_9215,N_9082);
nor U9608 (N_9608,N_9424,N_9236);
nor U9609 (N_9609,N_9389,N_9412);
xnor U9610 (N_9610,N_9036,N_9451);
nor U9611 (N_9611,N_9346,N_9322);
nor U9612 (N_9612,N_9314,N_9132);
and U9613 (N_9613,N_9413,N_9182);
and U9614 (N_9614,N_9373,N_9061);
and U9615 (N_9615,N_9371,N_9427);
or U9616 (N_9616,N_9180,N_9226);
xor U9617 (N_9617,N_9094,N_9356);
nand U9618 (N_9618,N_9030,N_9348);
or U9619 (N_9619,N_9209,N_9108);
and U9620 (N_9620,N_9306,N_9086);
nor U9621 (N_9621,N_9233,N_9174);
nand U9622 (N_9622,N_9241,N_9185);
nand U9623 (N_9623,N_9290,N_9485);
or U9624 (N_9624,N_9467,N_9370);
or U9625 (N_9625,N_9070,N_9254);
nand U9626 (N_9626,N_9481,N_9200);
or U9627 (N_9627,N_9323,N_9027);
or U9628 (N_9628,N_9421,N_9010);
and U9629 (N_9629,N_9355,N_9097);
and U9630 (N_9630,N_9186,N_9116);
and U9631 (N_9631,N_9014,N_9420);
or U9632 (N_9632,N_9315,N_9139);
nand U9633 (N_9633,N_9428,N_9093);
nand U9634 (N_9634,N_9257,N_9423);
and U9635 (N_9635,N_9366,N_9483);
nor U9636 (N_9636,N_9050,N_9354);
or U9637 (N_9637,N_9311,N_9407);
xor U9638 (N_9638,N_9247,N_9127);
nand U9639 (N_9639,N_9375,N_9130);
nand U9640 (N_9640,N_9069,N_9002);
xnor U9641 (N_9641,N_9148,N_9031);
or U9642 (N_9642,N_9312,N_9436);
nand U9643 (N_9643,N_9262,N_9040);
nand U9644 (N_9644,N_9395,N_9437);
xor U9645 (N_9645,N_9271,N_9208);
and U9646 (N_9646,N_9452,N_9207);
nor U9647 (N_9647,N_9448,N_9156);
nand U9648 (N_9648,N_9084,N_9391);
nor U9649 (N_9649,N_9457,N_9396);
nor U9650 (N_9650,N_9122,N_9253);
nand U9651 (N_9651,N_9255,N_9401);
and U9652 (N_9652,N_9332,N_9170);
nor U9653 (N_9653,N_9434,N_9219);
xor U9654 (N_9654,N_9248,N_9435);
and U9655 (N_9655,N_9380,N_9169);
or U9656 (N_9656,N_9441,N_9349);
nor U9657 (N_9657,N_9154,N_9308);
and U9658 (N_9658,N_9142,N_9277);
nor U9659 (N_9659,N_9321,N_9415);
or U9660 (N_9660,N_9102,N_9293);
and U9661 (N_9661,N_9146,N_9011);
xor U9662 (N_9662,N_9077,N_9347);
and U9663 (N_9663,N_9351,N_9340);
nand U9664 (N_9664,N_9137,N_9190);
nand U9665 (N_9665,N_9463,N_9081);
or U9666 (N_9666,N_9285,N_9191);
xnor U9667 (N_9667,N_9283,N_9118);
nor U9668 (N_9668,N_9220,N_9117);
or U9669 (N_9669,N_9106,N_9171);
nor U9670 (N_9670,N_9339,N_9331);
nand U9671 (N_9671,N_9111,N_9326);
and U9672 (N_9672,N_9300,N_9161);
and U9673 (N_9673,N_9330,N_9199);
and U9674 (N_9674,N_9334,N_9369);
or U9675 (N_9675,N_9147,N_9438);
and U9676 (N_9676,N_9214,N_9350);
or U9677 (N_9677,N_9488,N_9193);
and U9678 (N_9678,N_9462,N_9284);
nor U9679 (N_9679,N_9072,N_9178);
and U9680 (N_9680,N_9192,N_9495);
and U9681 (N_9681,N_9041,N_9153);
nor U9682 (N_9682,N_9364,N_9384);
or U9683 (N_9683,N_9078,N_9237);
and U9684 (N_9684,N_9444,N_9464);
nand U9685 (N_9685,N_9140,N_9377);
nor U9686 (N_9686,N_9309,N_9049);
nor U9687 (N_9687,N_9482,N_9187);
xor U9688 (N_9688,N_9202,N_9087);
nor U9689 (N_9689,N_9227,N_9020);
nand U9690 (N_9690,N_9359,N_9398);
nor U9691 (N_9691,N_9158,N_9018);
and U9692 (N_9692,N_9135,N_9218);
and U9693 (N_9693,N_9400,N_9124);
or U9694 (N_9694,N_9051,N_9029);
and U9695 (N_9695,N_9250,N_9318);
xor U9696 (N_9696,N_9063,N_9287);
nand U9697 (N_9697,N_9399,N_9223);
or U9698 (N_9698,N_9133,N_9390);
nand U9699 (N_9699,N_9307,N_9043);
nor U9700 (N_9700,N_9211,N_9039);
nor U9701 (N_9701,N_9092,N_9494);
nand U9702 (N_9702,N_9044,N_9181);
or U9703 (N_9703,N_9004,N_9230);
and U9704 (N_9704,N_9361,N_9431);
nor U9705 (N_9705,N_9183,N_9151);
nor U9706 (N_9706,N_9486,N_9100);
nand U9707 (N_9707,N_9497,N_9165);
nor U9708 (N_9708,N_9067,N_9143);
nand U9709 (N_9709,N_9484,N_9432);
nor U9710 (N_9710,N_9270,N_9107);
nor U9711 (N_9711,N_9144,N_9316);
nand U9712 (N_9712,N_9469,N_9341);
nand U9713 (N_9713,N_9475,N_9458);
nand U9714 (N_9714,N_9138,N_9204);
or U9715 (N_9715,N_9496,N_9065);
nor U9716 (N_9716,N_9074,N_9071);
and U9717 (N_9717,N_9335,N_9112);
or U9718 (N_9718,N_9382,N_9425);
or U9719 (N_9719,N_9372,N_9466);
xnor U9720 (N_9720,N_9450,N_9492);
nor U9721 (N_9721,N_9210,N_9068);
and U9722 (N_9722,N_9453,N_9152);
or U9723 (N_9723,N_9479,N_9352);
nand U9724 (N_9724,N_9126,N_9128);
or U9725 (N_9725,N_9385,N_9278);
or U9726 (N_9726,N_9461,N_9409);
nand U9727 (N_9727,N_9478,N_9123);
and U9728 (N_9728,N_9474,N_9026);
nand U9729 (N_9729,N_9360,N_9243);
nand U9730 (N_9730,N_9489,N_9188);
or U9731 (N_9731,N_9473,N_9426);
nand U9732 (N_9732,N_9164,N_9145);
or U9733 (N_9733,N_9258,N_9282);
nand U9734 (N_9734,N_9320,N_9487);
or U9735 (N_9735,N_9333,N_9374);
nor U9736 (N_9736,N_9205,N_9016);
xor U9737 (N_9737,N_9216,N_9260);
nor U9738 (N_9738,N_9273,N_9238);
nor U9739 (N_9739,N_9419,N_9229);
nor U9740 (N_9740,N_9256,N_9303);
nand U9741 (N_9741,N_9008,N_9272);
or U9742 (N_9742,N_9471,N_9096);
nand U9743 (N_9743,N_9460,N_9062);
xor U9744 (N_9744,N_9442,N_9150);
xnor U9745 (N_9745,N_9053,N_9015);
nor U9746 (N_9746,N_9470,N_9416);
and U9747 (N_9747,N_9459,N_9003);
nor U9748 (N_9748,N_9266,N_9405);
nand U9749 (N_9749,N_9498,N_9310);
nand U9750 (N_9750,N_9055,N_9275);
nand U9751 (N_9751,N_9050,N_9294);
or U9752 (N_9752,N_9019,N_9442);
xnor U9753 (N_9753,N_9282,N_9417);
and U9754 (N_9754,N_9410,N_9170);
and U9755 (N_9755,N_9203,N_9146);
and U9756 (N_9756,N_9387,N_9239);
nor U9757 (N_9757,N_9028,N_9070);
nand U9758 (N_9758,N_9081,N_9121);
nand U9759 (N_9759,N_9183,N_9227);
nor U9760 (N_9760,N_9042,N_9214);
and U9761 (N_9761,N_9204,N_9208);
and U9762 (N_9762,N_9215,N_9309);
or U9763 (N_9763,N_9061,N_9224);
xnor U9764 (N_9764,N_9305,N_9495);
nor U9765 (N_9765,N_9105,N_9496);
xor U9766 (N_9766,N_9321,N_9176);
and U9767 (N_9767,N_9466,N_9013);
and U9768 (N_9768,N_9362,N_9186);
nand U9769 (N_9769,N_9109,N_9131);
nor U9770 (N_9770,N_9094,N_9285);
nand U9771 (N_9771,N_9254,N_9093);
and U9772 (N_9772,N_9004,N_9122);
and U9773 (N_9773,N_9213,N_9309);
or U9774 (N_9774,N_9264,N_9327);
nand U9775 (N_9775,N_9418,N_9007);
and U9776 (N_9776,N_9029,N_9157);
nand U9777 (N_9777,N_9189,N_9314);
nor U9778 (N_9778,N_9182,N_9068);
nand U9779 (N_9779,N_9231,N_9280);
and U9780 (N_9780,N_9351,N_9376);
nor U9781 (N_9781,N_9366,N_9365);
nand U9782 (N_9782,N_9387,N_9489);
nor U9783 (N_9783,N_9056,N_9217);
nor U9784 (N_9784,N_9230,N_9000);
xnor U9785 (N_9785,N_9370,N_9137);
or U9786 (N_9786,N_9332,N_9107);
and U9787 (N_9787,N_9416,N_9405);
nor U9788 (N_9788,N_9319,N_9317);
nand U9789 (N_9789,N_9053,N_9142);
nand U9790 (N_9790,N_9127,N_9023);
or U9791 (N_9791,N_9427,N_9099);
nand U9792 (N_9792,N_9483,N_9475);
nor U9793 (N_9793,N_9481,N_9092);
and U9794 (N_9794,N_9420,N_9196);
or U9795 (N_9795,N_9070,N_9027);
or U9796 (N_9796,N_9290,N_9388);
nor U9797 (N_9797,N_9308,N_9008);
nand U9798 (N_9798,N_9002,N_9051);
or U9799 (N_9799,N_9116,N_9026);
xnor U9800 (N_9800,N_9464,N_9405);
or U9801 (N_9801,N_9301,N_9372);
and U9802 (N_9802,N_9224,N_9300);
nand U9803 (N_9803,N_9180,N_9414);
nand U9804 (N_9804,N_9227,N_9400);
nand U9805 (N_9805,N_9022,N_9098);
or U9806 (N_9806,N_9222,N_9232);
or U9807 (N_9807,N_9207,N_9165);
xor U9808 (N_9808,N_9282,N_9060);
xor U9809 (N_9809,N_9024,N_9141);
or U9810 (N_9810,N_9054,N_9247);
and U9811 (N_9811,N_9187,N_9417);
and U9812 (N_9812,N_9493,N_9396);
and U9813 (N_9813,N_9088,N_9105);
or U9814 (N_9814,N_9291,N_9222);
nor U9815 (N_9815,N_9130,N_9443);
and U9816 (N_9816,N_9373,N_9369);
nand U9817 (N_9817,N_9482,N_9260);
xor U9818 (N_9818,N_9456,N_9301);
and U9819 (N_9819,N_9362,N_9261);
or U9820 (N_9820,N_9320,N_9365);
or U9821 (N_9821,N_9357,N_9459);
nand U9822 (N_9822,N_9353,N_9476);
nand U9823 (N_9823,N_9010,N_9079);
nand U9824 (N_9824,N_9176,N_9019);
nor U9825 (N_9825,N_9481,N_9082);
and U9826 (N_9826,N_9172,N_9465);
or U9827 (N_9827,N_9100,N_9427);
and U9828 (N_9828,N_9147,N_9491);
nand U9829 (N_9829,N_9224,N_9370);
or U9830 (N_9830,N_9156,N_9012);
or U9831 (N_9831,N_9324,N_9084);
xor U9832 (N_9832,N_9441,N_9386);
nor U9833 (N_9833,N_9006,N_9307);
xor U9834 (N_9834,N_9484,N_9006);
nor U9835 (N_9835,N_9328,N_9444);
or U9836 (N_9836,N_9082,N_9093);
or U9837 (N_9837,N_9071,N_9100);
nor U9838 (N_9838,N_9383,N_9093);
nand U9839 (N_9839,N_9488,N_9286);
nand U9840 (N_9840,N_9173,N_9264);
nand U9841 (N_9841,N_9338,N_9250);
xor U9842 (N_9842,N_9086,N_9149);
or U9843 (N_9843,N_9118,N_9369);
nor U9844 (N_9844,N_9024,N_9247);
and U9845 (N_9845,N_9167,N_9384);
nor U9846 (N_9846,N_9419,N_9010);
nor U9847 (N_9847,N_9128,N_9221);
xor U9848 (N_9848,N_9170,N_9015);
nor U9849 (N_9849,N_9210,N_9406);
nand U9850 (N_9850,N_9391,N_9042);
nand U9851 (N_9851,N_9400,N_9496);
nand U9852 (N_9852,N_9166,N_9282);
and U9853 (N_9853,N_9312,N_9092);
nor U9854 (N_9854,N_9240,N_9058);
xor U9855 (N_9855,N_9428,N_9124);
nor U9856 (N_9856,N_9276,N_9101);
nand U9857 (N_9857,N_9123,N_9048);
and U9858 (N_9858,N_9113,N_9484);
nor U9859 (N_9859,N_9125,N_9254);
xnor U9860 (N_9860,N_9424,N_9038);
or U9861 (N_9861,N_9181,N_9334);
or U9862 (N_9862,N_9180,N_9213);
xnor U9863 (N_9863,N_9066,N_9461);
nor U9864 (N_9864,N_9346,N_9042);
nor U9865 (N_9865,N_9372,N_9216);
and U9866 (N_9866,N_9377,N_9423);
nor U9867 (N_9867,N_9027,N_9208);
and U9868 (N_9868,N_9366,N_9318);
and U9869 (N_9869,N_9017,N_9335);
nor U9870 (N_9870,N_9245,N_9348);
or U9871 (N_9871,N_9486,N_9165);
and U9872 (N_9872,N_9153,N_9486);
nand U9873 (N_9873,N_9448,N_9111);
nor U9874 (N_9874,N_9274,N_9009);
and U9875 (N_9875,N_9104,N_9484);
or U9876 (N_9876,N_9278,N_9438);
or U9877 (N_9877,N_9111,N_9259);
and U9878 (N_9878,N_9231,N_9414);
nand U9879 (N_9879,N_9374,N_9409);
nand U9880 (N_9880,N_9066,N_9203);
nand U9881 (N_9881,N_9036,N_9061);
or U9882 (N_9882,N_9298,N_9385);
xnor U9883 (N_9883,N_9054,N_9184);
xor U9884 (N_9884,N_9114,N_9125);
nand U9885 (N_9885,N_9375,N_9376);
xnor U9886 (N_9886,N_9411,N_9400);
or U9887 (N_9887,N_9183,N_9018);
or U9888 (N_9888,N_9318,N_9147);
and U9889 (N_9889,N_9258,N_9287);
xor U9890 (N_9890,N_9385,N_9492);
nor U9891 (N_9891,N_9269,N_9431);
and U9892 (N_9892,N_9280,N_9063);
xor U9893 (N_9893,N_9013,N_9182);
and U9894 (N_9894,N_9075,N_9249);
xor U9895 (N_9895,N_9095,N_9359);
nor U9896 (N_9896,N_9453,N_9194);
nor U9897 (N_9897,N_9388,N_9459);
and U9898 (N_9898,N_9291,N_9428);
nand U9899 (N_9899,N_9402,N_9468);
and U9900 (N_9900,N_9042,N_9451);
nand U9901 (N_9901,N_9035,N_9371);
and U9902 (N_9902,N_9215,N_9475);
nand U9903 (N_9903,N_9349,N_9345);
or U9904 (N_9904,N_9246,N_9289);
and U9905 (N_9905,N_9307,N_9114);
or U9906 (N_9906,N_9416,N_9191);
or U9907 (N_9907,N_9061,N_9472);
nor U9908 (N_9908,N_9164,N_9393);
and U9909 (N_9909,N_9427,N_9195);
nand U9910 (N_9910,N_9487,N_9496);
nand U9911 (N_9911,N_9443,N_9104);
xnor U9912 (N_9912,N_9136,N_9040);
nor U9913 (N_9913,N_9244,N_9031);
nand U9914 (N_9914,N_9007,N_9375);
or U9915 (N_9915,N_9169,N_9040);
or U9916 (N_9916,N_9333,N_9222);
and U9917 (N_9917,N_9124,N_9243);
or U9918 (N_9918,N_9196,N_9377);
nand U9919 (N_9919,N_9180,N_9316);
nor U9920 (N_9920,N_9046,N_9081);
nor U9921 (N_9921,N_9105,N_9421);
nor U9922 (N_9922,N_9463,N_9069);
xor U9923 (N_9923,N_9203,N_9124);
nand U9924 (N_9924,N_9124,N_9342);
and U9925 (N_9925,N_9492,N_9334);
nand U9926 (N_9926,N_9038,N_9324);
and U9927 (N_9927,N_9274,N_9079);
or U9928 (N_9928,N_9255,N_9278);
nor U9929 (N_9929,N_9380,N_9020);
and U9930 (N_9930,N_9290,N_9187);
and U9931 (N_9931,N_9396,N_9429);
and U9932 (N_9932,N_9354,N_9159);
nor U9933 (N_9933,N_9240,N_9428);
and U9934 (N_9934,N_9233,N_9320);
xnor U9935 (N_9935,N_9286,N_9385);
or U9936 (N_9936,N_9469,N_9391);
or U9937 (N_9937,N_9314,N_9080);
or U9938 (N_9938,N_9221,N_9388);
and U9939 (N_9939,N_9417,N_9146);
or U9940 (N_9940,N_9187,N_9271);
nor U9941 (N_9941,N_9174,N_9031);
nand U9942 (N_9942,N_9096,N_9093);
nor U9943 (N_9943,N_9478,N_9191);
and U9944 (N_9944,N_9056,N_9292);
or U9945 (N_9945,N_9293,N_9090);
or U9946 (N_9946,N_9212,N_9132);
nand U9947 (N_9947,N_9241,N_9212);
nand U9948 (N_9948,N_9315,N_9226);
nand U9949 (N_9949,N_9161,N_9237);
nor U9950 (N_9950,N_9001,N_9458);
nor U9951 (N_9951,N_9059,N_9237);
nor U9952 (N_9952,N_9175,N_9072);
nand U9953 (N_9953,N_9161,N_9066);
nor U9954 (N_9954,N_9106,N_9122);
or U9955 (N_9955,N_9322,N_9443);
or U9956 (N_9956,N_9283,N_9461);
nand U9957 (N_9957,N_9341,N_9380);
and U9958 (N_9958,N_9405,N_9460);
or U9959 (N_9959,N_9412,N_9446);
nor U9960 (N_9960,N_9366,N_9047);
and U9961 (N_9961,N_9314,N_9029);
xor U9962 (N_9962,N_9121,N_9281);
or U9963 (N_9963,N_9390,N_9185);
xnor U9964 (N_9964,N_9497,N_9402);
nand U9965 (N_9965,N_9077,N_9201);
nand U9966 (N_9966,N_9275,N_9032);
nand U9967 (N_9967,N_9345,N_9270);
and U9968 (N_9968,N_9299,N_9109);
xnor U9969 (N_9969,N_9104,N_9419);
nand U9970 (N_9970,N_9265,N_9447);
nor U9971 (N_9971,N_9115,N_9446);
and U9972 (N_9972,N_9332,N_9213);
nor U9973 (N_9973,N_9175,N_9029);
or U9974 (N_9974,N_9123,N_9246);
nor U9975 (N_9975,N_9260,N_9339);
or U9976 (N_9976,N_9429,N_9002);
and U9977 (N_9977,N_9446,N_9450);
or U9978 (N_9978,N_9044,N_9177);
nand U9979 (N_9979,N_9128,N_9182);
and U9980 (N_9980,N_9099,N_9231);
or U9981 (N_9981,N_9077,N_9251);
or U9982 (N_9982,N_9441,N_9296);
nor U9983 (N_9983,N_9233,N_9449);
and U9984 (N_9984,N_9025,N_9171);
nand U9985 (N_9985,N_9329,N_9365);
nand U9986 (N_9986,N_9207,N_9414);
or U9987 (N_9987,N_9398,N_9462);
and U9988 (N_9988,N_9272,N_9119);
and U9989 (N_9989,N_9285,N_9336);
nor U9990 (N_9990,N_9302,N_9090);
and U9991 (N_9991,N_9374,N_9170);
and U9992 (N_9992,N_9432,N_9120);
and U9993 (N_9993,N_9160,N_9156);
and U9994 (N_9994,N_9315,N_9463);
xor U9995 (N_9995,N_9080,N_9086);
xnor U9996 (N_9996,N_9424,N_9128);
nand U9997 (N_9997,N_9437,N_9326);
nor U9998 (N_9998,N_9100,N_9338);
or U9999 (N_9999,N_9080,N_9376);
or UO_0 (O_0,N_9502,N_9624);
and UO_1 (O_1,N_9662,N_9944);
and UO_2 (O_2,N_9891,N_9826);
nor UO_3 (O_3,N_9716,N_9909);
nand UO_4 (O_4,N_9788,N_9821);
nand UO_5 (O_5,N_9798,N_9635);
nor UO_6 (O_6,N_9593,N_9708);
and UO_7 (O_7,N_9658,N_9503);
nand UO_8 (O_8,N_9631,N_9611);
or UO_9 (O_9,N_9973,N_9992);
nand UO_10 (O_10,N_9764,N_9663);
nand UO_11 (O_11,N_9638,N_9552);
xor UO_12 (O_12,N_9728,N_9912);
xnor UO_13 (O_13,N_9633,N_9800);
nor UO_14 (O_14,N_9831,N_9991);
nand UO_15 (O_15,N_9896,N_9535);
xor UO_16 (O_16,N_9967,N_9885);
and UO_17 (O_17,N_9581,N_9639);
and UO_18 (O_18,N_9671,N_9510);
and UO_19 (O_19,N_9538,N_9590);
nor UO_20 (O_20,N_9765,N_9797);
nor UO_21 (O_21,N_9838,N_9855);
or UO_22 (O_22,N_9514,N_9999);
nand UO_23 (O_23,N_9698,N_9922);
and UO_24 (O_24,N_9720,N_9997);
nor UO_25 (O_25,N_9978,N_9890);
nor UO_26 (O_26,N_9557,N_9886);
nand UO_27 (O_27,N_9681,N_9702);
nand UO_28 (O_28,N_9583,N_9948);
and UO_29 (O_29,N_9609,N_9861);
or UO_30 (O_30,N_9814,N_9534);
xor UO_31 (O_31,N_9762,N_9938);
and UO_32 (O_32,N_9939,N_9872);
xnor UO_33 (O_33,N_9555,N_9600);
and UO_34 (O_34,N_9518,N_9526);
or UO_35 (O_35,N_9670,N_9719);
nand UO_36 (O_36,N_9956,N_9576);
or UO_37 (O_37,N_9691,N_9819);
nor UO_38 (O_38,N_9874,N_9976);
nand UO_39 (O_39,N_9884,N_9606);
nor UO_40 (O_40,N_9820,N_9647);
and UO_41 (O_41,N_9628,N_9780);
nand UO_42 (O_42,N_9676,N_9697);
or UO_43 (O_43,N_9562,N_9947);
and UO_44 (O_44,N_9942,N_9740);
xor UO_45 (O_45,N_9649,N_9607);
nand UO_46 (O_46,N_9830,N_9839);
nand UO_47 (O_47,N_9744,N_9906);
nor UO_48 (O_48,N_9806,N_9845);
nand UO_49 (O_49,N_9571,N_9955);
and UO_50 (O_50,N_9882,N_9927);
nor UO_51 (O_51,N_9563,N_9961);
and UO_52 (O_52,N_9677,N_9957);
or UO_53 (O_53,N_9959,N_9963);
and UO_54 (O_54,N_9962,N_9920);
and UO_55 (O_55,N_9507,N_9610);
nor UO_56 (O_56,N_9623,N_9717);
nor UO_57 (O_57,N_9859,N_9602);
nor UO_58 (O_58,N_9675,N_9597);
or UO_59 (O_59,N_9930,N_9827);
or UO_60 (O_60,N_9558,N_9977);
nor UO_61 (O_61,N_9810,N_9914);
or UO_62 (O_62,N_9949,N_9569);
and UO_63 (O_63,N_9684,N_9808);
nor UO_64 (O_64,N_9913,N_9735);
and UO_65 (O_65,N_9903,N_9857);
nand UO_66 (O_66,N_9616,N_9883);
nand UO_67 (O_67,N_9887,N_9974);
and UO_68 (O_68,N_9714,N_9895);
nor UO_69 (O_69,N_9692,N_9833);
nor UO_70 (O_70,N_9907,N_9792);
nand UO_71 (O_71,N_9986,N_9536);
nor UO_72 (O_72,N_9758,N_9899);
or UO_73 (O_73,N_9527,N_9984);
nand UO_74 (O_74,N_9879,N_9802);
nor UO_75 (O_75,N_9757,N_9876);
xnor UO_76 (O_76,N_9520,N_9584);
xnor UO_77 (O_77,N_9918,N_9572);
nand UO_78 (O_78,N_9897,N_9801);
or UO_79 (O_79,N_9531,N_9987);
nor UO_80 (O_80,N_9525,N_9644);
nand UO_81 (O_81,N_9811,N_9632);
or UO_82 (O_82,N_9568,N_9875);
or UO_83 (O_83,N_9878,N_9813);
and UO_84 (O_84,N_9911,N_9622);
nor UO_85 (O_85,N_9900,N_9546);
or UO_86 (O_86,N_9910,N_9881);
or UO_87 (O_87,N_9650,N_9595);
nor UO_88 (O_88,N_9799,N_9972);
nand UO_89 (O_89,N_9786,N_9693);
or UO_90 (O_90,N_9850,N_9782);
xor UO_91 (O_91,N_9713,N_9775);
or UO_92 (O_92,N_9867,N_9573);
nor UO_93 (O_93,N_9753,N_9749);
or UO_94 (O_94,N_9853,N_9580);
and UO_95 (O_95,N_9733,N_9931);
or UO_96 (O_96,N_9805,N_9582);
and UO_97 (O_97,N_9804,N_9946);
nand UO_98 (O_98,N_9812,N_9860);
or UO_99 (O_99,N_9605,N_9630);
nand UO_100 (O_100,N_9727,N_9768);
nand UO_101 (O_101,N_9791,N_9739);
nand UO_102 (O_102,N_9645,N_9705);
nor UO_103 (O_103,N_9504,N_9575);
nor UO_104 (O_104,N_9781,N_9608);
nand UO_105 (O_105,N_9653,N_9539);
or UO_106 (O_106,N_9548,N_9619);
and UO_107 (O_107,N_9851,N_9952);
nand UO_108 (O_108,N_9685,N_9660);
nand UO_109 (O_109,N_9544,N_9617);
and UO_110 (O_110,N_9869,N_9704);
or UO_111 (O_111,N_9640,N_9529);
and UO_112 (O_112,N_9642,N_9854);
or UO_113 (O_113,N_9598,N_9842);
xnor UO_114 (O_114,N_9577,N_9995);
nand UO_115 (O_115,N_9856,N_9594);
or UO_116 (O_116,N_9766,N_9919);
and UO_117 (O_117,N_9615,N_9591);
or UO_118 (O_118,N_9672,N_9769);
and UO_119 (O_119,N_9928,N_9500);
or UO_120 (O_120,N_9843,N_9866);
or UO_121 (O_121,N_9966,N_9665);
nor UO_122 (O_122,N_9840,N_9926);
or UO_123 (O_123,N_9824,N_9849);
nor UO_124 (O_124,N_9612,N_9996);
and UO_125 (O_125,N_9673,N_9679);
nand UO_126 (O_126,N_9817,N_9565);
nand UO_127 (O_127,N_9943,N_9755);
nor UO_128 (O_128,N_9793,N_9873);
nor UO_129 (O_129,N_9725,N_9542);
nor UO_130 (O_130,N_9561,N_9554);
or UO_131 (O_131,N_9550,N_9951);
and UO_132 (O_132,N_9722,N_9574);
nand UO_133 (O_133,N_9589,N_9998);
and UO_134 (O_134,N_9508,N_9969);
nor UO_135 (O_135,N_9736,N_9767);
nor UO_136 (O_136,N_9964,N_9868);
nand UO_137 (O_137,N_9668,N_9699);
nand UO_138 (O_138,N_9656,N_9711);
and UO_139 (O_139,N_9985,N_9960);
and UO_140 (O_140,N_9980,N_9924);
nand UO_141 (O_141,N_9862,N_9566);
or UO_142 (O_142,N_9950,N_9669);
nand UO_143 (O_143,N_9667,N_9965);
xnor UO_144 (O_144,N_9724,N_9784);
and UO_145 (O_145,N_9752,N_9648);
or UO_146 (O_146,N_9505,N_9709);
xor UO_147 (O_147,N_9712,N_9627);
or UO_148 (O_148,N_9601,N_9694);
nand UO_149 (O_149,N_9945,N_9773);
nand UO_150 (O_150,N_9994,N_9975);
or UO_151 (O_151,N_9528,N_9828);
and UO_152 (O_152,N_9686,N_9637);
and UO_153 (O_153,N_9829,N_9626);
nor UO_154 (O_154,N_9596,N_9683);
nand UO_155 (O_155,N_9770,N_9807);
nor UO_156 (O_156,N_9614,N_9889);
or UO_157 (O_157,N_9971,N_9754);
nand UO_158 (O_158,N_9603,N_9750);
nand UO_159 (O_159,N_9674,N_9659);
or UO_160 (O_160,N_9848,N_9916);
xnor UO_161 (O_161,N_9682,N_9501);
and UO_162 (O_162,N_9687,N_9530);
xnor UO_163 (O_163,N_9777,N_9937);
and UO_164 (O_164,N_9785,N_9513);
or UO_165 (O_165,N_9524,N_9511);
nor UO_166 (O_166,N_9816,N_9795);
nor UO_167 (O_167,N_9776,N_9979);
or UO_168 (O_168,N_9547,N_9982);
xor UO_169 (O_169,N_9690,N_9778);
or UO_170 (O_170,N_9745,N_9908);
nor UO_171 (O_171,N_9970,N_9689);
and UO_172 (O_172,N_9678,N_9981);
or UO_173 (O_173,N_9917,N_9723);
and UO_174 (O_174,N_9729,N_9864);
nor UO_175 (O_175,N_9519,N_9516);
nor UO_176 (O_176,N_9935,N_9703);
nand UO_177 (O_177,N_9634,N_9718);
and UO_178 (O_178,N_9836,N_9625);
or UO_179 (O_179,N_9664,N_9643);
nor UO_180 (O_180,N_9894,N_9763);
or UO_181 (O_181,N_9989,N_9695);
nand UO_182 (O_182,N_9771,N_9904);
nand UO_183 (O_183,N_9880,N_9738);
or UO_184 (O_184,N_9915,N_9523);
nand UO_185 (O_185,N_9892,N_9844);
or UO_186 (O_186,N_9517,N_9983);
nor UO_187 (O_187,N_9772,N_9588);
or UO_188 (O_188,N_9726,N_9958);
nand UO_189 (O_189,N_9940,N_9789);
and UO_190 (O_190,N_9654,N_9936);
or UO_191 (O_191,N_9818,N_9657);
and UO_192 (O_192,N_9515,N_9905);
nor UO_193 (O_193,N_9651,N_9925);
or UO_194 (O_194,N_9847,N_9578);
nand UO_195 (O_195,N_9929,N_9641);
xor UO_196 (O_196,N_9761,N_9743);
nand UO_197 (O_197,N_9721,N_9731);
nor UO_198 (O_198,N_9803,N_9646);
nand UO_199 (O_199,N_9710,N_9898);
or UO_200 (O_200,N_9556,N_9888);
nand UO_201 (O_201,N_9586,N_9680);
nor UO_202 (O_202,N_9621,N_9846);
or UO_203 (O_203,N_9809,N_9747);
and UO_204 (O_204,N_9707,N_9666);
nor UO_205 (O_205,N_9968,N_9730);
or UO_206 (O_206,N_9759,N_9652);
and UO_207 (O_207,N_9512,N_9532);
or UO_208 (O_208,N_9837,N_9852);
or UO_209 (O_209,N_9661,N_9823);
nor UO_210 (O_210,N_9506,N_9790);
and UO_211 (O_211,N_9988,N_9921);
or UO_212 (O_212,N_9990,N_9636);
nand UO_213 (O_213,N_9751,N_9620);
nand UO_214 (O_214,N_9834,N_9543);
xor UO_215 (O_215,N_9592,N_9587);
nand UO_216 (O_216,N_9655,N_9901);
and UO_217 (O_217,N_9559,N_9585);
xnor UO_218 (O_218,N_9787,N_9579);
and UO_219 (O_219,N_9688,N_9825);
and UO_220 (O_220,N_9794,N_9953);
nor UO_221 (O_221,N_9815,N_9941);
and UO_222 (O_222,N_9560,N_9796);
and UO_223 (O_223,N_9835,N_9549);
nand UO_224 (O_224,N_9564,N_9522);
nand UO_225 (O_225,N_9779,N_9541);
and UO_226 (O_226,N_9748,N_9570);
nand UO_227 (O_227,N_9706,N_9993);
nand UO_228 (O_228,N_9865,N_9863);
nor UO_229 (O_229,N_9760,N_9741);
or UO_230 (O_230,N_9537,N_9877);
or UO_231 (O_231,N_9893,N_9604);
and UO_232 (O_232,N_9715,N_9618);
and UO_233 (O_233,N_9783,N_9934);
nand UO_234 (O_234,N_9629,N_9521);
and UO_235 (O_235,N_9742,N_9540);
nand UO_236 (O_236,N_9696,N_9599);
xor UO_237 (O_237,N_9613,N_9553);
or UO_238 (O_238,N_9545,N_9732);
or UO_239 (O_239,N_9841,N_9923);
nand UO_240 (O_240,N_9509,N_9701);
and UO_241 (O_241,N_9858,N_9737);
and UO_242 (O_242,N_9746,N_9533);
nand UO_243 (O_243,N_9734,N_9870);
nand UO_244 (O_244,N_9954,N_9756);
xnor UO_245 (O_245,N_9822,N_9902);
and UO_246 (O_246,N_9871,N_9933);
or UO_247 (O_247,N_9774,N_9832);
nor UO_248 (O_248,N_9700,N_9567);
and UO_249 (O_249,N_9932,N_9551);
and UO_250 (O_250,N_9686,N_9635);
or UO_251 (O_251,N_9925,N_9861);
and UO_252 (O_252,N_9871,N_9981);
nand UO_253 (O_253,N_9672,N_9866);
nand UO_254 (O_254,N_9773,N_9691);
or UO_255 (O_255,N_9805,N_9668);
and UO_256 (O_256,N_9864,N_9948);
nand UO_257 (O_257,N_9758,N_9522);
nand UO_258 (O_258,N_9739,N_9653);
or UO_259 (O_259,N_9567,N_9792);
xor UO_260 (O_260,N_9692,N_9621);
nand UO_261 (O_261,N_9725,N_9792);
and UO_262 (O_262,N_9869,N_9550);
or UO_263 (O_263,N_9625,N_9805);
nand UO_264 (O_264,N_9758,N_9680);
or UO_265 (O_265,N_9883,N_9691);
and UO_266 (O_266,N_9856,N_9646);
or UO_267 (O_267,N_9729,N_9623);
nand UO_268 (O_268,N_9885,N_9733);
or UO_269 (O_269,N_9814,N_9924);
xnor UO_270 (O_270,N_9940,N_9658);
xor UO_271 (O_271,N_9923,N_9733);
xnor UO_272 (O_272,N_9595,N_9737);
nand UO_273 (O_273,N_9587,N_9994);
nand UO_274 (O_274,N_9641,N_9665);
nand UO_275 (O_275,N_9516,N_9671);
xnor UO_276 (O_276,N_9588,N_9693);
xor UO_277 (O_277,N_9884,N_9933);
nand UO_278 (O_278,N_9880,N_9587);
or UO_279 (O_279,N_9860,N_9893);
and UO_280 (O_280,N_9932,N_9739);
and UO_281 (O_281,N_9602,N_9743);
nand UO_282 (O_282,N_9837,N_9761);
nand UO_283 (O_283,N_9726,N_9789);
xnor UO_284 (O_284,N_9655,N_9539);
nand UO_285 (O_285,N_9818,N_9561);
and UO_286 (O_286,N_9943,N_9951);
or UO_287 (O_287,N_9577,N_9623);
nand UO_288 (O_288,N_9946,N_9870);
and UO_289 (O_289,N_9975,N_9966);
or UO_290 (O_290,N_9989,N_9684);
or UO_291 (O_291,N_9789,N_9675);
or UO_292 (O_292,N_9690,N_9500);
nand UO_293 (O_293,N_9985,N_9877);
and UO_294 (O_294,N_9989,N_9733);
nor UO_295 (O_295,N_9878,N_9807);
nor UO_296 (O_296,N_9689,N_9934);
and UO_297 (O_297,N_9940,N_9547);
nor UO_298 (O_298,N_9915,N_9707);
or UO_299 (O_299,N_9519,N_9693);
nand UO_300 (O_300,N_9745,N_9858);
nor UO_301 (O_301,N_9893,N_9716);
and UO_302 (O_302,N_9541,N_9619);
or UO_303 (O_303,N_9721,N_9507);
or UO_304 (O_304,N_9936,N_9550);
or UO_305 (O_305,N_9538,N_9688);
xnor UO_306 (O_306,N_9735,N_9769);
nor UO_307 (O_307,N_9828,N_9648);
nor UO_308 (O_308,N_9788,N_9665);
or UO_309 (O_309,N_9556,N_9636);
or UO_310 (O_310,N_9518,N_9900);
nor UO_311 (O_311,N_9588,N_9507);
nor UO_312 (O_312,N_9729,N_9950);
and UO_313 (O_313,N_9874,N_9631);
or UO_314 (O_314,N_9655,N_9550);
nand UO_315 (O_315,N_9919,N_9891);
nand UO_316 (O_316,N_9545,N_9974);
nor UO_317 (O_317,N_9879,N_9810);
xor UO_318 (O_318,N_9691,N_9926);
nand UO_319 (O_319,N_9543,N_9563);
nor UO_320 (O_320,N_9743,N_9544);
nand UO_321 (O_321,N_9926,N_9877);
nor UO_322 (O_322,N_9504,N_9688);
or UO_323 (O_323,N_9894,N_9618);
nand UO_324 (O_324,N_9545,N_9829);
or UO_325 (O_325,N_9681,N_9828);
and UO_326 (O_326,N_9747,N_9854);
xnor UO_327 (O_327,N_9693,N_9882);
nor UO_328 (O_328,N_9974,N_9897);
nor UO_329 (O_329,N_9781,N_9698);
nand UO_330 (O_330,N_9883,N_9935);
nand UO_331 (O_331,N_9674,N_9546);
nor UO_332 (O_332,N_9953,N_9814);
and UO_333 (O_333,N_9672,N_9915);
nand UO_334 (O_334,N_9540,N_9991);
xnor UO_335 (O_335,N_9908,N_9700);
or UO_336 (O_336,N_9761,N_9632);
or UO_337 (O_337,N_9848,N_9874);
nand UO_338 (O_338,N_9854,N_9675);
or UO_339 (O_339,N_9591,N_9745);
nand UO_340 (O_340,N_9954,N_9634);
nor UO_341 (O_341,N_9886,N_9985);
nor UO_342 (O_342,N_9611,N_9887);
nor UO_343 (O_343,N_9968,N_9675);
xor UO_344 (O_344,N_9508,N_9578);
xor UO_345 (O_345,N_9814,N_9838);
or UO_346 (O_346,N_9616,N_9930);
xor UO_347 (O_347,N_9586,N_9570);
nor UO_348 (O_348,N_9705,N_9675);
nor UO_349 (O_349,N_9619,N_9728);
nor UO_350 (O_350,N_9681,N_9785);
nand UO_351 (O_351,N_9895,N_9604);
and UO_352 (O_352,N_9787,N_9930);
and UO_353 (O_353,N_9839,N_9995);
nor UO_354 (O_354,N_9621,N_9509);
or UO_355 (O_355,N_9986,N_9508);
nor UO_356 (O_356,N_9710,N_9611);
or UO_357 (O_357,N_9701,N_9839);
and UO_358 (O_358,N_9824,N_9988);
and UO_359 (O_359,N_9731,N_9878);
nand UO_360 (O_360,N_9646,N_9721);
or UO_361 (O_361,N_9776,N_9843);
nor UO_362 (O_362,N_9755,N_9727);
and UO_363 (O_363,N_9613,N_9708);
nor UO_364 (O_364,N_9720,N_9948);
or UO_365 (O_365,N_9697,N_9808);
nand UO_366 (O_366,N_9851,N_9668);
or UO_367 (O_367,N_9860,N_9868);
and UO_368 (O_368,N_9577,N_9530);
nand UO_369 (O_369,N_9553,N_9745);
or UO_370 (O_370,N_9591,N_9515);
and UO_371 (O_371,N_9641,N_9605);
nand UO_372 (O_372,N_9675,N_9716);
or UO_373 (O_373,N_9585,N_9844);
nand UO_374 (O_374,N_9518,N_9577);
or UO_375 (O_375,N_9985,N_9742);
or UO_376 (O_376,N_9552,N_9914);
or UO_377 (O_377,N_9651,N_9727);
nand UO_378 (O_378,N_9766,N_9974);
or UO_379 (O_379,N_9648,N_9966);
or UO_380 (O_380,N_9745,N_9750);
nor UO_381 (O_381,N_9880,N_9503);
nor UO_382 (O_382,N_9972,N_9939);
nand UO_383 (O_383,N_9997,N_9635);
and UO_384 (O_384,N_9838,N_9636);
and UO_385 (O_385,N_9858,N_9930);
nor UO_386 (O_386,N_9565,N_9688);
or UO_387 (O_387,N_9918,N_9562);
nand UO_388 (O_388,N_9524,N_9830);
nor UO_389 (O_389,N_9953,N_9655);
nor UO_390 (O_390,N_9611,N_9805);
nor UO_391 (O_391,N_9562,N_9698);
or UO_392 (O_392,N_9567,N_9933);
and UO_393 (O_393,N_9649,N_9592);
or UO_394 (O_394,N_9532,N_9903);
xnor UO_395 (O_395,N_9880,N_9608);
nor UO_396 (O_396,N_9647,N_9962);
nor UO_397 (O_397,N_9592,N_9880);
xor UO_398 (O_398,N_9670,N_9794);
or UO_399 (O_399,N_9744,N_9597);
nor UO_400 (O_400,N_9544,N_9536);
nor UO_401 (O_401,N_9505,N_9627);
nand UO_402 (O_402,N_9627,N_9611);
and UO_403 (O_403,N_9693,N_9945);
or UO_404 (O_404,N_9893,N_9684);
and UO_405 (O_405,N_9863,N_9805);
nand UO_406 (O_406,N_9735,N_9809);
nor UO_407 (O_407,N_9690,N_9586);
nand UO_408 (O_408,N_9829,N_9605);
nor UO_409 (O_409,N_9975,N_9774);
nand UO_410 (O_410,N_9672,N_9848);
nand UO_411 (O_411,N_9922,N_9589);
nand UO_412 (O_412,N_9932,N_9958);
and UO_413 (O_413,N_9620,N_9958);
nand UO_414 (O_414,N_9745,N_9832);
or UO_415 (O_415,N_9626,N_9667);
or UO_416 (O_416,N_9678,N_9767);
nand UO_417 (O_417,N_9635,N_9575);
nor UO_418 (O_418,N_9664,N_9546);
nor UO_419 (O_419,N_9524,N_9761);
and UO_420 (O_420,N_9917,N_9542);
nor UO_421 (O_421,N_9636,N_9904);
and UO_422 (O_422,N_9538,N_9736);
nand UO_423 (O_423,N_9571,N_9885);
nand UO_424 (O_424,N_9660,N_9547);
nand UO_425 (O_425,N_9766,N_9889);
or UO_426 (O_426,N_9837,N_9932);
nor UO_427 (O_427,N_9704,N_9954);
or UO_428 (O_428,N_9651,N_9629);
or UO_429 (O_429,N_9688,N_9591);
nand UO_430 (O_430,N_9557,N_9898);
nand UO_431 (O_431,N_9528,N_9958);
xor UO_432 (O_432,N_9734,N_9941);
nand UO_433 (O_433,N_9637,N_9713);
nand UO_434 (O_434,N_9880,N_9948);
nand UO_435 (O_435,N_9626,N_9785);
and UO_436 (O_436,N_9829,N_9594);
nand UO_437 (O_437,N_9691,N_9720);
nand UO_438 (O_438,N_9920,N_9681);
and UO_439 (O_439,N_9764,N_9858);
or UO_440 (O_440,N_9709,N_9838);
or UO_441 (O_441,N_9629,N_9532);
or UO_442 (O_442,N_9848,N_9645);
nand UO_443 (O_443,N_9939,N_9959);
or UO_444 (O_444,N_9810,N_9859);
and UO_445 (O_445,N_9535,N_9589);
xnor UO_446 (O_446,N_9706,N_9936);
nand UO_447 (O_447,N_9822,N_9808);
and UO_448 (O_448,N_9522,N_9680);
nand UO_449 (O_449,N_9984,N_9771);
nand UO_450 (O_450,N_9558,N_9581);
and UO_451 (O_451,N_9728,N_9620);
xnor UO_452 (O_452,N_9958,N_9711);
and UO_453 (O_453,N_9763,N_9575);
or UO_454 (O_454,N_9835,N_9727);
or UO_455 (O_455,N_9943,N_9873);
or UO_456 (O_456,N_9795,N_9726);
nand UO_457 (O_457,N_9831,N_9762);
and UO_458 (O_458,N_9613,N_9957);
and UO_459 (O_459,N_9969,N_9864);
and UO_460 (O_460,N_9519,N_9723);
nor UO_461 (O_461,N_9813,N_9852);
nor UO_462 (O_462,N_9677,N_9978);
nand UO_463 (O_463,N_9649,N_9974);
nor UO_464 (O_464,N_9886,N_9805);
or UO_465 (O_465,N_9667,N_9868);
xnor UO_466 (O_466,N_9778,N_9642);
nor UO_467 (O_467,N_9702,N_9871);
nand UO_468 (O_468,N_9742,N_9869);
and UO_469 (O_469,N_9543,N_9520);
nand UO_470 (O_470,N_9715,N_9676);
nand UO_471 (O_471,N_9920,N_9640);
xnor UO_472 (O_472,N_9851,N_9835);
or UO_473 (O_473,N_9781,N_9910);
xor UO_474 (O_474,N_9536,N_9656);
or UO_475 (O_475,N_9591,N_9557);
or UO_476 (O_476,N_9571,N_9799);
nand UO_477 (O_477,N_9783,N_9887);
or UO_478 (O_478,N_9592,N_9774);
nand UO_479 (O_479,N_9860,N_9863);
and UO_480 (O_480,N_9956,N_9985);
xor UO_481 (O_481,N_9533,N_9898);
or UO_482 (O_482,N_9706,N_9921);
nor UO_483 (O_483,N_9730,N_9632);
and UO_484 (O_484,N_9508,N_9928);
or UO_485 (O_485,N_9978,N_9810);
and UO_486 (O_486,N_9983,N_9958);
nor UO_487 (O_487,N_9590,N_9964);
and UO_488 (O_488,N_9965,N_9544);
and UO_489 (O_489,N_9930,N_9504);
xor UO_490 (O_490,N_9886,N_9847);
nand UO_491 (O_491,N_9794,N_9535);
nand UO_492 (O_492,N_9873,N_9567);
and UO_493 (O_493,N_9528,N_9877);
or UO_494 (O_494,N_9605,N_9734);
nor UO_495 (O_495,N_9697,N_9896);
and UO_496 (O_496,N_9823,N_9926);
and UO_497 (O_497,N_9975,N_9690);
or UO_498 (O_498,N_9623,N_9755);
nor UO_499 (O_499,N_9725,N_9807);
nand UO_500 (O_500,N_9941,N_9750);
nor UO_501 (O_501,N_9823,N_9848);
nand UO_502 (O_502,N_9632,N_9756);
and UO_503 (O_503,N_9620,N_9664);
or UO_504 (O_504,N_9540,N_9881);
nand UO_505 (O_505,N_9866,N_9526);
nor UO_506 (O_506,N_9766,N_9797);
and UO_507 (O_507,N_9918,N_9581);
and UO_508 (O_508,N_9769,N_9773);
nand UO_509 (O_509,N_9927,N_9509);
nand UO_510 (O_510,N_9739,N_9908);
or UO_511 (O_511,N_9646,N_9808);
nand UO_512 (O_512,N_9505,N_9696);
and UO_513 (O_513,N_9704,N_9623);
or UO_514 (O_514,N_9526,N_9979);
nand UO_515 (O_515,N_9701,N_9533);
nand UO_516 (O_516,N_9695,N_9573);
or UO_517 (O_517,N_9603,N_9694);
xnor UO_518 (O_518,N_9604,N_9703);
or UO_519 (O_519,N_9593,N_9987);
or UO_520 (O_520,N_9567,N_9755);
nor UO_521 (O_521,N_9942,N_9818);
nor UO_522 (O_522,N_9908,N_9860);
nand UO_523 (O_523,N_9712,N_9715);
xnor UO_524 (O_524,N_9734,N_9805);
nand UO_525 (O_525,N_9893,N_9741);
nand UO_526 (O_526,N_9635,N_9644);
and UO_527 (O_527,N_9903,N_9646);
or UO_528 (O_528,N_9943,N_9955);
or UO_529 (O_529,N_9965,N_9811);
nor UO_530 (O_530,N_9656,N_9557);
nor UO_531 (O_531,N_9996,N_9862);
nand UO_532 (O_532,N_9655,N_9581);
xor UO_533 (O_533,N_9547,N_9625);
or UO_534 (O_534,N_9527,N_9578);
and UO_535 (O_535,N_9722,N_9530);
nor UO_536 (O_536,N_9618,N_9656);
and UO_537 (O_537,N_9785,N_9856);
and UO_538 (O_538,N_9531,N_9853);
or UO_539 (O_539,N_9976,N_9577);
xor UO_540 (O_540,N_9893,N_9561);
nor UO_541 (O_541,N_9636,N_9732);
or UO_542 (O_542,N_9633,N_9751);
nand UO_543 (O_543,N_9821,N_9985);
nor UO_544 (O_544,N_9650,N_9936);
or UO_545 (O_545,N_9624,N_9921);
xnor UO_546 (O_546,N_9858,N_9902);
and UO_547 (O_547,N_9846,N_9920);
nor UO_548 (O_548,N_9919,N_9689);
and UO_549 (O_549,N_9502,N_9627);
nand UO_550 (O_550,N_9659,N_9817);
or UO_551 (O_551,N_9689,N_9998);
or UO_552 (O_552,N_9539,N_9514);
nand UO_553 (O_553,N_9619,N_9926);
xnor UO_554 (O_554,N_9615,N_9924);
nor UO_555 (O_555,N_9741,N_9907);
or UO_556 (O_556,N_9959,N_9842);
nand UO_557 (O_557,N_9627,N_9857);
and UO_558 (O_558,N_9637,N_9928);
nor UO_559 (O_559,N_9603,N_9710);
and UO_560 (O_560,N_9604,N_9603);
nor UO_561 (O_561,N_9708,N_9860);
and UO_562 (O_562,N_9824,N_9808);
nor UO_563 (O_563,N_9599,N_9621);
and UO_564 (O_564,N_9712,N_9640);
and UO_565 (O_565,N_9713,N_9961);
and UO_566 (O_566,N_9963,N_9899);
nand UO_567 (O_567,N_9828,N_9730);
and UO_568 (O_568,N_9541,N_9684);
and UO_569 (O_569,N_9908,N_9666);
nand UO_570 (O_570,N_9596,N_9790);
or UO_571 (O_571,N_9533,N_9998);
xor UO_572 (O_572,N_9824,N_9832);
nor UO_573 (O_573,N_9594,N_9969);
or UO_574 (O_574,N_9679,N_9685);
xor UO_575 (O_575,N_9608,N_9972);
or UO_576 (O_576,N_9601,N_9917);
and UO_577 (O_577,N_9614,N_9702);
xor UO_578 (O_578,N_9875,N_9848);
or UO_579 (O_579,N_9943,N_9512);
nor UO_580 (O_580,N_9877,N_9694);
and UO_581 (O_581,N_9766,N_9888);
or UO_582 (O_582,N_9762,N_9883);
and UO_583 (O_583,N_9741,N_9840);
nor UO_584 (O_584,N_9953,N_9894);
xnor UO_585 (O_585,N_9934,N_9855);
nor UO_586 (O_586,N_9524,N_9785);
and UO_587 (O_587,N_9631,N_9605);
nand UO_588 (O_588,N_9757,N_9536);
nor UO_589 (O_589,N_9995,N_9920);
nor UO_590 (O_590,N_9769,N_9825);
nor UO_591 (O_591,N_9716,N_9750);
or UO_592 (O_592,N_9609,N_9767);
or UO_593 (O_593,N_9888,N_9564);
nand UO_594 (O_594,N_9620,N_9634);
nor UO_595 (O_595,N_9773,N_9754);
or UO_596 (O_596,N_9682,N_9762);
nor UO_597 (O_597,N_9709,N_9973);
nand UO_598 (O_598,N_9801,N_9655);
nor UO_599 (O_599,N_9629,N_9657);
or UO_600 (O_600,N_9579,N_9573);
or UO_601 (O_601,N_9853,N_9896);
nor UO_602 (O_602,N_9876,N_9686);
or UO_603 (O_603,N_9820,N_9530);
xnor UO_604 (O_604,N_9907,N_9871);
and UO_605 (O_605,N_9583,N_9978);
nor UO_606 (O_606,N_9991,N_9855);
xor UO_607 (O_607,N_9925,N_9984);
nor UO_608 (O_608,N_9508,N_9854);
and UO_609 (O_609,N_9503,N_9810);
or UO_610 (O_610,N_9954,N_9703);
nand UO_611 (O_611,N_9652,N_9852);
nor UO_612 (O_612,N_9534,N_9843);
nand UO_613 (O_613,N_9570,N_9861);
nor UO_614 (O_614,N_9968,N_9828);
nand UO_615 (O_615,N_9616,N_9687);
and UO_616 (O_616,N_9541,N_9666);
nor UO_617 (O_617,N_9885,N_9625);
or UO_618 (O_618,N_9809,N_9740);
nand UO_619 (O_619,N_9966,N_9731);
nor UO_620 (O_620,N_9507,N_9898);
and UO_621 (O_621,N_9991,N_9819);
and UO_622 (O_622,N_9673,N_9508);
nand UO_623 (O_623,N_9530,N_9711);
nand UO_624 (O_624,N_9614,N_9731);
or UO_625 (O_625,N_9785,N_9757);
and UO_626 (O_626,N_9883,N_9578);
nand UO_627 (O_627,N_9832,N_9861);
nor UO_628 (O_628,N_9609,N_9506);
nand UO_629 (O_629,N_9660,N_9862);
and UO_630 (O_630,N_9548,N_9873);
or UO_631 (O_631,N_9788,N_9540);
nor UO_632 (O_632,N_9528,N_9606);
nor UO_633 (O_633,N_9520,N_9628);
xor UO_634 (O_634,N_9703,N_9640);
or UO_635 (O_635,N_9548,N_9568);
xnor UO_636 (O_636,N_9964,N_9638);
nor UO_637 (O_637,N_9786,N_9613);
xnor UO_638 (O_638,N_9737,N_9664);
nand UO_639 (O_639,N_9851,N_9617);
nand UO_640 (O_640,N_9888,N_9987);
and UO_641 (O_641,N_9680,N_9530);
nor UO_642 (O_642,N_9760,N_9722);
and UO_643 (O_643,N_9920,N_9815);
nor UO_644 (O_644,N_9544,N_9667);
or UO_645 (O_645,N_9714,N_9713);
or UO_646 (O_646,N_9530,N_9739);
nand UO_647 (O_647,N_9730,N_9741);
nand UO_648 (O_648,N_9963,N_9648);
nand UO_649 (O_649,N_9904,N_9945);
xor UO_650 (O_650,N_9615,N_9577);
or UO_651 (O_651,N_9914,N_9519);
nor UO_652 (O_652,N_9911,N_9582);
or UO_653 (O_653,N_9551,N_9666);
nand UO_654 (O_654,N_9749,N_9544);
and UO_655 (O_655,N_9604,N_9801);
nand UO_656 (O_656,N_9653,N_9862);
xnor UO_657 (O_657,N_9545,N_9971);
and UO_658 (O_658,N_9916,N_9642);
nor UO_659 (O_659,N_9854,N_9581);
or UO_660 (O_660,N_9846,N_9830);
xor UO_661 (O_661,N_9600,N_9685);
and UO_662 (O_662,N_9887,N_9820);
nand UO_663 (O_663,N_9549,N_9696);
nand UO_664 (O_664,N_9590,N_9844);
nor UO_665 (O_665,N_9990,N_9676);
nand UO_666 (O_666,N_9805,N_9833);
or UO_667 (O_667,N_9993,N_9957);
or UO_668 (O_668,N_9844,N_9519);
and UO_669 (O_669,N_9770,N_9860);
or UO_670 (O_670,N_9698,N_9858);
and UO_671 (O_671,N_9855,N_9715);
or UO_672 (O_672,N_9664,N_9691);
xor UO_673 (O_673,N_9781,N_9949);
nor UO_674 (O_674,N_9918,N_9969);
nand UO_675 (O_675,N_9841,N_9928);
and UO_676 (O_676,N_9648,N_9822);
or UO_677 (O_677,N_9863,N_9917);
nor UO_678 (O_678,N_9627,N_9680);
or UO_679 (O_679,N_9549,N_9919);
or UO_680 (O_680,N_9747,N_9551);
nand UO_681 (O_681,N_9714,N_9822);
and UO_682 (O_682,N_9597,N_9610);
nand UO_683 (O_683,N_9594,N_9603);
or UO_684 (O_684,N_9641,N_9764);
nor UO_685 (O_685,N_9911,N_9518);
or UO_686 (O_686,N_9626,N_9723);
xnor UO_687 (O_687,N_9959,N_9750);
nor UO_688 (O_688,N_9781,N_9996);
and UO_689 (O_689,N_9977,N_9596);
and UO_690 (O_690,N_9680,N_9568);
and UO_691 (O_691,N_9781,N_9526);
xnor UO_692 (O_692,N_9806,N_9989);
and UO_693 (O_693,N_9772,N_9742);
and UO_694 (O_694,N_9694,N_9814);
nor UO_695 (O_695,N_9639,N_9573);
and UO_696 (O_696,N_9719,N_9897);
or UO_697 (O_697,N_9766,N_9805);
nor UO_698 (O_698,N_9624,N_9748);
and UO_699 (O_699,N_9537,N_9870);
and UO_700 (O_700,N_9952,N_9811);
and UO_701 (O_701,N_9596,N_9726);
and UO_702 (O_702,N_9510,N_9507);
xor UO_703 (O_703,N_9668,N_9828);
or UO_704 (O_704,N_9609,N_9557);
and UO_705 (O_705,N_9757,N_9779);
nor UO_706 (O_706,N_9645,N_9762);
nor UO_707 (O_707,N_9979,N_9695);
and UO_708 (O_708,N_9641,N_9801);
nor UO_709 (O_709,N_9615,N_9791);
nor UO_710 (O_710,N_9786,N_9937);
or UO_711 (O_711,N_9670,N_9829);
nor UO_712 (O_712,N_9869,N_9978);
nor UO_713 (O_713,N_9647,N_9535);
and UO_714 (O_714,N_9640,N_9893);
or UO_715 (O_715,N_9555,N_9725);
or UO_716 (O_716,N_9943,N_9942);
or UO_717 (O_717,N_9596,N_9788);
and UO_718 (O_718,N_9619,N_9552);
nor UO_719 (O_719,N_9749,N_9620);
or UO_720 (O_720,N_9867,N_9741);
and UO_721 (O_721,N_9821,N_9812);
and UO_722 (O_722,N_9655,N_9808);
and UO_723 (O_723,N_9781,N_9692);
xnor UO_724 (O_724,N_9612,N_9633);
xor UO_725 (O_725,N_9688,N_9696);
xor UO_726 (O_726,N_9732,N_9692);
nand UO_727 (O_727,N_9753,N_9720);
nor UO_728 (O_728,N_9996,N_9896);
or UO_729 (O_729,N_9826,N_9857);
and UO_730 (O_730,N_9579,N_9957);
and UO_731 (O_731,N_9850,N_9816);
xor UO_732 (O_732,N_9618,N_9822);
or UO_733 (O_733,N_9793,N_9969);
and UO_734 (O_734,N_9645,N_9834);
nor UO_735 (O_735,N_9539,N_9827);
nand UO_736 (O_736,N_9566,N_9541);
nand UO_737 (O_737,N_9794,N_9900);
or UO_738 (O_738,N_9569,N_9766);
or UO_739 (O_739,N_9659,N_9901);
and UO_740 (O_740,N_9637,N_9533);
nand UO_741 (O_741,N_9590,N_9867);
nand UO_742 (O_742,N_9583,N_9823);
or UO_743 (O_743,N_9950,N_9933);
nor UO_744 (O_744,N_9951,N_9790);
xor UO_745 (O_745,N_9798,N_9654);
and UO_746 (O_746,N_9567,N_9651);
nor UO_747 (O_747,N_9629,N_9501);
nor UO_748 (O_748,N_9806,N_9608);
nor UO_749 (O_749,N_9634,N_9938);
and UO_750 (O_750,N_9821,N_9588);
nor UO_751 (O_751,N_9819,N_9674);
nor UO_752 (O_752,N_9990,N_9657);
nand UO_753 (O_753,N_9832,N_9719);
and UO_754 (O_754,N_9701,N_9544);
or UO_755 (O_755,N_9761,N_9643);
and UO_756 (O_756,N_9916,N_9758);
nor UO_757 (O_757,N_9563,N_9770);
and UO_758 (O_758,N_9522,N_9862);
nand UO_759 (O_759,N_9511,N_9566);
nor UO_760 (O_760,N_9546,N_9926);
or UO_761 (O_761,N_9750,N_9553);
nor UO_762 (O_762,N_9942,N_9912);
nor UO_763 (O_763,N_9833,N_9802);
and UO_764 (O_764,N_9813,N_9677);
or UO_765 (O_765,N_9706,N_9821);
or UO_766 (O_766,N_9662,N_9723);
nand UO_767 (O_767,N_9619,N_9851);
and UO_768 (O_768,N_9572,N_9556);
or UO_769 (O_769,N_9952,N_9637);
nor UO_770 (O_770,N_9804,N_9830);
nand UO_771 (O_771,N_9564,N_9761);
or UO_772 (O_772,N_9559,N_9667);
and UO_773 (O_773,N_9564,N_9779);
nand UO_774 (O_774,N_9987,N_9610);
xnor UO_775 (O_775,N_9650,N_9947);
or UO_776 (O_776,N_9717,N_9531);
or UO_777 (O_777,N_9886,N_9642);
nand UO_778 (O_778,N_9510,N_9936);
xor UO_779 (O_779,N_9780,N_9779);
or UO_780 (O_780,N_9588,N_9665);
nand UO_781 (O_781,N_9671,N_9897);
nand UO_782 (O_782,N_9806,N_9637);
nand UO_783 (O_783,N_9628,N_9660);
or UO_784 (O_784,N_9619,N_9858);
and UO_785 (O_785,N_9581,N_9683);
or UO_786 (O_786,N_9599,N_9671);
and UO_787 (O_787,N_9939,N_9977);
or UO_788 (O_788,N_9935,N_9618);
and UO_789 (O_789,N_9608,N_9638);
xor UO_790 (O_790,N_9948,N_9955);
or UO_791 (O_791,N_9853,N_9682);
nor UO_792 (O_792,N_9811,N_9755);
and UO_793 (O_793,N_9912,N_9636);
or UO_794 (O_794,N_9915,N_9841);
nand UO_795 (O_795,N_9963,N_9638);
nand UO_796 (O_796,N_9510,N_9710);
xnor UO_797 (O_797,N_9907,N_9553);
nand UO_798 (O_798,N_9941,N_9662);
and UO_799 (O_799,N_9556,N_9836);
nand UO_800 (O_800,N_9905,N_9781);
and UO_801 (O_801,N_9613,N_9660);
and UO_802 (O_802,N_9554,N_9853);
nand UO_803 (O_803,N_9902,N_9963);
or UO_804 (O_804,N_9766,N_9612);
or UO_805 (O_805,N_9853,N_9663);
nand UO_806 (O_806,N_9534,N_9653);
nand UO_807 (O_807,N_9591,N_9571);
and UO_808 (O_808,N_9956,N_9861);
or UO_809 (O_809,N_9558,N_9765);
xnor UO_810 (O_810,N_9512,N_9538);
nor UO_811 (O_811,N_9678,N_9706);
nor UO_812 (O_812,N_9876,N_9666);
or UO_813 (O_813,N_9658,N_9599);
nand UO_814 (O_814,N_9738,N_9861);
and UO_815 (O_815,N_9864,N_9578);
nor UO_816 (O_816,N_9915,N_9761);
xor UO_817 (O_817,N_9765,N_9960);
or UO_818 (O_818,N_9916,N_9558);
nand UO_819 (O_819,N_9979,N_9614);
nor UO_820 (O_820,N_9851,N_9850);
nor UO_821 (O_821,N_9612,N_9500);
nor UO_822 (O_822,N_9927,N_9633);
xnor UO_823 (O_823,N_9911,N_9541);
xnor UO_824 (O_824,N_9765,N_9801);
or UO_825 (O_825,N_9834,N_9580);
xor UO_826 (O_826,N_9621,N_9997);
nand UO_827 (O_827,N_9923,N_9720);
nor UO_828 (O_828,N_9734,N_9929);
nand UO_829 (O_829,N_9999,N_9694);
nand UO_830 (O_830,N_9792,N_9665);
and UO_831 (O_831,N_9731,N_9759);
or UO_832 (O_832,N_9787,N_9637);
or UO_833 (O_833,N_9813,N_9673);
and UO_834 (O_834,N_9764,N_9737);
nand UO_835 (O_835,N_9785,N_9838);
nor UO_836 (O_836,N_9732,N_9884);
or UO_837 (O_837,N_9687,N_9756);
and UO_838 (O_838,N_9686,N_9924);
nand UO_839 (O_839,N_9853,N_9807);
or UO_840 (O_840,N_9906,N_9782);
or UO_841 (O_841,N_9570,N_9613);
nor UO_842 (O_842,N_9946,N_9800);
or UO_843 (O_843,N_9868,N_9782);
and UO_844 (O_844,N_9521,N_9864);
nor UO_845 (O_845,N_9760,N_9638);
or UO_846 (O_846,N_9714,N_9720);
nand UO_847 (O_847,N_9637,N_9892);
and UO_848 (O_848,N_9586,N_9580);
or UO_849 (O_849,N_9605,N_9655);
nor UO_850 (O_850,N_9859,N_9570);
nand UO_851 (O_851,N_9778,N_9910);
or UO_852 (O_852,N_9663,N_9630);
nand UO_853 (O_853,N_9769,N_9675);
nor UO_854 (O_854,N_9644,N_9824);
nor UO_855 (O_855,N_9729,N_9865);
nor UO_856 (O_856,N_9886,N_9875);
or UO_857 (O_857,N_9920,N_9598);
nand UO_858 (O_858,N_9754,N_9899);
xor UO_859 (O_859,N_9532,N_9888);
nor UO_860 (O_860,N_9575,N_9861);
and UO_861 (O_861,N_9807,N_9737);
nand UO_862 (O_862,N_9870,N_9810);
nand UO_863 (O_863,N_9944,N_9638);
nor UO_864 (O_864,N_9702,N_9503);
and UO_865 (O_865,N_9998,N_9954);
nand UO_866 (O_866,N_9905,N_9577);
nand UO_867 (O_867,N_9634,N_9680);
and UO_868 (O_868,N_9584,N_9640);
and UO_869 (O_869,N_9693,N_9678);
nor UO_870 (O_870,N_9850,N_9735);
and UO_871 (O_871,N_9600,N_9603);
nand UO_872 (O_872,N_9575,N_9529);
and UO_873 (O_873,N_9884,N_9678);
and UO_874 (O_874,N_9984,N_9504);
and UO_875 (O_875,N_9502,N_9617);
or UO_876 (O_876,N_9918,N_9863);
nand UO_877 (O_877,N_9729,N_9783);
or UO_878 (O_878,N_9776,N_9539);
nor UO_879 (O_879,N_9644,N_9806);
nor UO_880 (O_880,N_9548,N_9823);
or UO_881 (O_881,N_9697,N_9749);
or UO_882 (O_882,N_9535,N_9940);
nand UO_883 (O_883,N_9521,N_9534);
or UO_884 (O_884,N_9523,N_9709);
xnor UO_885 (O_885,N_9902,N_9885);
and UO_886 (O_886,N_9557,N_9679);
or UO_887 (O_887,N_9711,N_9580);
nand UO_888 (O_888,N_9922,N_9514);
nor UO_889 (O_889,N_9702,N_9688);
nor UO_890 (O_890,N_9527,N_9835);
and UO_891 (O_891,N_9691,N_9680);
nand UO_892 (O_892,N_9721,N_9911);
and UO_893 (O_893,N_9994,N_9682);
nor UO_894 (O_894,N_9666,N_9975);
and UO_895 (O_895,N_9812,N_9717);
nand UO_896 (O_896,N_9527,N_9894);
nand UO_897 (O_897,N_9700,N_9653);
nor UO_898 (O_898,N_9592,N_9666);
or UO_899 (O_899,N_9537,N_9676);
nand UO_900 (O_900,N_9879,N_9565);
nand UO_901 (O_901,N_9660,N_9769);
nor UO_902 (O_902,N_9728,N_9819);
nand UO_903 (O_903,N_9817,N_9728);
and UO_904 (O_904,N_9642,N_9805);
xnor UO_905 (O_905,N_9615,N_9880);
xor UO_906 (O_906,N_9603,N_9712);
nand UO_907 (O_907,N_9722,N_9597);
or UO_908 (O_908,N_9543,N_9595);
or UO_909 (O_909,N_9547,N_9695);
nand UO_910 (O_910,N_9552,N_9500);
and UO_911 (O_911,N_9608,N_9973);
and UO_912 (O_912,N_9684,N_9636);
xnor UO_913 (O_913,N_9560,N_9625);
xor UO_914 (O_914,N_9627,N_9962);
nor UO_915 (O_915,N_9619,N_9511);
nor UO_916 (O_916,N_9870,N_9729);
nand UO_917 (O_917,N_9900,N_9585);
or UO_918 (O_918,N_9961,N_9933);
xnor UO_919 (O_919,N_9721,N_9990);
xnor UO_920 (O_920,N_9648,N_9611);
and UO_921 (O_921,N_9840,N_9636);
and UO_922 (O_922,N_9770,N_9880);
xnor UO_923 (O_923,N_9649,N_9593);
or UO_924 (O_924,N_9686,N_9547);
or UO_925 (O_925,N_9959,N_9937);
or UO_926 (O_926,N_9886,N_9554);
nand UO_927 (O_927,N_9939,N_9662);
nand UO_928 (O_928,N_9658,N_9679);
or UO_929 (O_929,N_9921,N_9945);
nand UO_930 (O_930,N_9742,N_9710);
or UO_931 (O_931,N_9508,N_9552);
nand UO_932 (O_932,N_9647,N_9611);
xnor UO_933 (O_933,N_9949,N_9572);
nor UO_934 (O_934,N_9521,N_9699);
nand UO_935 (O_935,N_9571,N_9666);
xor UO_936 (O_936,N_9746,N_9666);
and UO_937 (O_937,N_9598,N_9661);
and UO_938 (O_938,N_9570,N_9665);
nor UO_939 (O_939,N_9684,N_9521);
and UO_940 (O_940,N_9865,N_9870);
or UO_941 (O_941,N_9638,N_9906);
nand UO_942 (O_942,N_9961,N_9994);
or UO_943 (O_943,N_9839,N_9854);
nand UO_944 (O_944,N_9626,N_9876);
and UO_945 (O_945,N_9513,N_9823);
or UO_946 (O_946,N_9730,N_9573);
nor UO_947 (O_947,N_9884,N_9569);
or UO_948 (O_948,N_9736,N_9780);
nand UO_949 (O_949,N_9521,N_9980);
and UO_950 (O_950,N_9678,N_9658);
xnor UO_951 (O_951,N_9825,N_9816);
nor UO_952 (O_952,N_9629,N_9739);
or UO_953 (O_953,N_9573,N_9664);
or UO_954 (O_954,N_9940,N_9977);
nor UO_955 (O_955,N_9906,N_9634);
nor UO_956 (O_956,N_9858,N_9574);
nand UO_957 (O_957,N_9679,N_9587);
or UO_958 (O_958,N_9915,N_9889);
or UO_959 (O_959,N_9818,N_9710);
nor UO_960 (O_960,N_9823,N_9516);
and UO_961 (O_961,N_9836,N_9669);
nor UO_962 (O_962,N_9732,N_9651);
nand UO_963 (O_963,N_9536,N_9803);
nor UO_964 (O_964,N_9938,N_9561);
nand UO_965 (O_965,N_9682,N_9955);
nor UO_966 (O_966,N_9823,N_9556);
and UO_967 (O_967,N_9542,N_9915);
nor UO_968 (O_968,N_9604,N_9735);
nor UO_969 (O_969,N_9792,N_9571);
nand UO_970 (O_970,N_9806,N_9793);
nand UO_971 (O_971,N_9972,N_9903);
nor UO_972 (O_972,N_9785,N_9551);
nor UO_973 (O_973,N_9586,N_9681);
nand UO_974 (O_974,N_9657,N_9980);
xnor UO_975 (O_975,N_9958,N_9995);
nor UO_976 (O_976,N_9706,N_9884);
nor UO_977 (O_977,N_9838,N_9807);
nand UO_978 (O_978,N_9774,N_9784);
xnor UO_979 (O_979,N_9928,N_9510);
nor UO_980 (O_980,N_9813,N_9850);
xnor UO_981 (O_981,N_9787,N_9961);
and UO_982 (O_982,N_9649,N_9746);
and UO_983 (O_983,N_9805,N_9741);
and UO_984 (O_984,N_9903,N_9698);
and UO_985 (O_985,N_9697,N_9919);
nor UO_986 (O_986,N_9624,N_9771);
nor UO_987 (O_987,N_9925,N_9824);
or UO_988 (O_988,N_9813,N_9877);
nand UO_989 (O_989,N_9523,N_9906);
nand UO_990 (O_990,N_9549,N_9615);
nor UO_991 (O_991,N_9526,N_9788);
nor UO_992 (O_992,N_9640,N_9624);
or UO_993 (O_993,N_9766,N_9673);
nand UO_994 (O_994,N_9685,N_9698);
or UO_995 (O_995,N_9755,N_9883);
nor UO_996 (O_996,N_9970,N_9787);
or UO_997 (O_997,N_9627,N_9549);
or UO_998 (O_998,N_9820,N_9754);
nand UO_999 (O_999,N_9782,N_9952);
xor UO_1000 (O_1000,N_9849,N_9581);
or UO_1001 (O_1001,N_9716,N_9630);
nand UO_1002 (O_1002,N_9562,N_9610);
nor UO_1003 (O_1003,N_9799,N_9675);
nand UO_1004 (O_1004,N_9861,N_9574);
nand UO_1005 (O_1005,N_9918,N_9724);
xnor UO_1006 (O_1006,N_9951,N_9901);
and UO_1007 (O_1007,N_9724,N_9711);
or UO_1008 (O_1008,N_9867,N_9780);
nand UO_1009 (O_1009,N_9633,N_9627);
or UO_1010 (O_1010,N_9523,N_9916);
nor UO_1011 (O_1011,N_9540,N_9637);
nand UO_1012 (O_1012,N_9564,N_9605);
nor UO_1013 (O_1013,N_9940,N_9686);
or UO_1014 (O_1014,N_9641,N_9689);
and UO_1015 (O_1015,N_9627,N_9934);
and UO_1016 (O_1016,N_9587,N_9517);
nor UO_1017 (O_1017,N_9518,N_9693);
nand UO_1018 (O_1018,N_9936,N_9601);
or UO_1019 (O_1019,N_9687,N_9631);
nand UO_1020 (O_1020,N_9710,N_9869);
nor UO_1021 (O_1021,N_9680,N_9989);
nand UO_1022 (O_1022,N_9898,N_9971);
nor UO_1023 (O_1023,N_9895,N_9825);
nand UO_1024 (O_1024,N_9881,N_9559);
nor UO_1025 (O_1025,N_9571,N_9721);
or UO_1026 (O_1026,N_9683,N_9707);
xnor UO_1027 (O_1027,N_9749,N_9886);
or UO_1028 (O_1028,N_9548,N_9645);
nor UO_1029 (O_1029,N_9761,N_9695);
nand UO_1030 (O_1030,N_9521,N_9717);
or UO_1031 (O_1031,N_9662,N_9714);
and UO_1032 (O_1032,N_9999,N_9805);
and UO_1033 (O_1033,N_9690,N_9638);
or UO_1034 (O_1034,N_9966,N_9877);
nor UO_1035 (O_1035,N_9637,N_9558);
or UO_1036 (O_1036,N_9592,N_9742);
or UO_1037 (O_1037,N_9889,N_9683);
nand UO_1038 (O_1038,N_9873,N_9508);
and UO_1039 (O_1039,N_9615,N_9975);
nand UO_1040 (O_1040,N_9550,N_9994);
or UO_1041 (O_1041,N_9549,N_9739);
and UO_1042 (O_1042,N_9736,N_9612);
and UO_1043 (O_1043,N_9593,N_9724);
nor UO_1044 (O_1044,N_9750,N_9568);
or UO_1045 (O_1045,N_9937,N_9705);
xnor UO_1046 (O_1046,N_9990,N_9981);
nand UO_1047 (O_1047,N_9521,N_9669);
or UO_1048 (O_1048,N_9508,N_9884);
or UO_1049 (O_1049,N_9577,N_9515);
or UO_1050 (O_1050,N_9584,N_9763);
and UO_1051 (O_1051,N_9692,N_9750);
or UO_1052 (O_1052,N_9500,N_9734);
nor UO_1053 (O_1053,N_9941,N_9899);
and UO_1054 (O_1054,N_9894,N_9847);
nand UO_1055 (O_1055,N_9759,N_9831);
or UO_1056 (O_1056,N_9856,N_9787);
or UO_1057 (O_1057,N_9725,N_9944);
nor UO_1058 (O_1058,N_9508,N_9796);
xor UO_1059 (O_1059,N_9616,N_9561);
nor UO_1060 (O_1060,N_9606,N_9983);
nand UO_1061 (O_1061,N_9720,N_9722);
and UO_1062 (O_1062,N_9922,N_9700);
or UO_1063 (O_1063,N_9964,N_9848);
or UO_1064 (O_1064,N_9875,N_9693);
nand UO_1065 (O_1065,N_9998,N_9557);
xnor UO_1066 (O_1066,N_9523,N_9734);
or UO_1067 (O_1067,N_9524,N_9877);
nor UO_1068 (O_1068,N_9715,N_9611);
and UO_1069 (O_1069,N_9897,N_9792);
nor UO_1070 (O_1070,N_9756,N_9614);
or UO_1071 (O_1071,N_9659,N_9602);
or UO_1072 (O_1072,N_9820,N_9579);
nor UO_1073 (O_1073,N_9852,N_9949);
or UO_1074 (O_1074,N_9770,N_9774);
or UO_1075 (O_1075,N_9917,N_9865);
nand UO_1076 (O_1076,N_9821,N_9824);
and UO_1077 (O_1077,N_9901,N_9530);
or UO_1078 (O_1078,N_9700,N_9855);
or UO_1079 (O_1079,N_9736,N_9755);
nand UO_1080 (O_1080,N_9990,N_9868);
or UO_1081 (O_1081,N_9662,N_9838);
and UO_1082 (O_1082,N_9564,N_9845);
nor UO_1083 (O_1083,N_9518,N_9729);
xnor UO_1084 (O_1084,N_9784,N_9951);
nand UO_1085 (O_1085,N_9501,N_9780);
nor UO_1086 (O_1086,N_9954,N_9644);
or UO_1087 (O_1087,N_9669,N_9712);
nor UO_1088 (O_1088,N_9941,N_9837);
or UO_1089 (O_1089,N_9648,N_9933);
and UO_1090 (O_1090,N_9941,N_9860);
nand UO_1091 (O_1091,N_9503,N_9980);
or UO_1092 (O_1092,N_9738,N_9930);
and UO_1093 (O_1093,N_9858,N_9986);
xnor UO_1094 (O_1094,N_9522,N_9955);
xnor UO_1095 (O_1095,N_9602,N_9919);
nor UO_1096 (O_1096,N_9702,N_9657);
nand UO_1097 (O_1097,N_9552,N_9856);
and UO_1098 (O_1098,N_9575,N_9872);
nand UO_1099 (O_1099,N_9691,N_9825);
or UO_1100 (O_1100,N_9881,N_9933);
or UO_1101 (O_1101,N_9522,N_9850);
and UO_1102 (O_1102,N_9737,N_9615);
nor UO_1103 (O_1103,N_9687,N_9859);
nand UO_1104 (O_1104,N_9935,N_9927);
nor UO_1105 (O_1105,N_9886,N_9690);
or UO_1106 (O_1106,N_9949,N_9802);
or UO_1107 (O_1107,N_9521,N_9619);
and UO_1108 (O_1108,N_9568,N_9601);
xnor UO_1109 (O_1109,N_9606,N_9659);
nand UO_1110 (O_1110,N_9554,N_9804);
and UO_1111 (O_1111,N_9609,N_9691);
and UO_1112 (O_1112,N_9517,N_9513);
nor UO_1113 (O_1113,N_9511,N_9504);
xor UO_1114 (O_1114,N_9670,N_9971);
nor UO_1115 (O_1115,N_9992,N_9551);
nor UO_1116 (O_1116,N_9621,N_9524);
and UO_1117 (O_1117,N_9526,N_9734);
or UO_1118 (O_1118,N_9863,N_9795);
or UO_1119 (O_1119,N_9577,N_9933);
or UO_1120 (O_1120,N_9550,N_9552);
nor UO_1121 (O_1121,N_9587,N_9561);
xor UO_1122 (O_1122,N_9756,N_9977);
and UO_1123 (O_1123,N_9963,N_9838);
nor UO_1124 (O_1124,N_9826,N_9901);
nand UO_1125 (O_1125,N_9989,N_9767);
or UO_1126 (O_1126,N_9657,N_9970);
nor UO_1127 (O_1127,N_9880,N_9656);
nand UO_1128 (O_1128,N_9915,N_9942);
nand UO_1129 (O_1129,N_9811,N_9921);
nor UO_1130 (O_1130,N_9656,N_9682);
and UO_1131 (O_1131,N_9531,N_9602);
nand UO_1132 (O_1132,N_9553,N_9666);
or UO_1133 (O_1133,N_9895,N_9567);
and UO_1134 (O_1134,N_9549,N_9666);
or UO_1135 (O_1135,N_9812,N_9561);
or UO_1136 (O_1136,N_9842,N_9602);
nand UO_1137 (O_1137,N_9920,N_9766);
nor UO_1138 (O_1138,N_9617,N_9832);
or UO_1139 (O_1139,N_9904,N_9910);
nand UO_1140 (O_1140,N_9713,N_9548);
nor UO_1141 (O_1141,N_9636,N_9640);
or UO_1142 (O_1142,N_9924,N_9685);
and UO_1143 (O_1143,N_9676,N_9828);
or UO_1144 (O_1144,N_9998,N_9681);
nand UO_1145 (O_1145,N_9782,N_9726);
and UO_1146 (O_1146,N_9724,N_9646);
nand UO_1147 (O_1147,N_9864,N_9852);
or UO_1148 (O_1148,N_9763,N_9789);
and UO_1149 (O_1149,N_9794,N_9875);
and UO_1150 (O_1150,N_9523,N_9708);
nand UO_1151 (O_1151,N_9518,N_9619);
xnor UO_1152 (O_1152,N_9652,N_9641);
xor UO_1153 (O_1153,N_9522,N_9559);
or UO_1154 (O_1154,N_9564,N_9648);
nand UO_1155 (O_1155,N_9927,N_9694);
nor UO_1156 (O_1156,N_9650,N_9558);
nor UO_1157 (O_1157,N_9872,N_9712);
or UO_1158 (O_1158,N_9771,N_9663);
xor UO_1159 (O_1159,N_9647,N_9960);
nand UO_1160 (O_1160,N_9762,N_9593);
xnor UO_1161 (O_1161,N_9672,N_9757);
nand UO_1162 (O_1162,N_9953,N_9881);
nand UO_1163 (O_1163,N_9821,N_9549);
nand UO_1164 (O_1164,N_9749,N_9936);
xor UO_1165 (O_1165,N_9533,N_9849);
or UO_1166 (O_1166,N_9817,N_9955);
and UO_1167 (O_1167,N_9846,N_9523);
nor UO_1168 (O_1168,N_9748,N_9657);
nor UO_1169 (O_1169,N_9899,N_9698);
and UO_1170 (O_1170,N_9890,N_9962);
nand UO_1171 (O_1171,N_9753,N_9528);
nor UO_1172 (O_1172,N_9888,N_9897);
and UO_1173 (O_1173,N_9848,N_9939);
or UO_1174 (O_1174,N_9623,N_9546);
or UO_1175 (O_1175,N_9610,N_9858);
or UO_1176 (O_1176,N_9826,N_9685);
nor UO_1177 (O_1177,N_9956,N_9837);
and UO_1178 (O_1178,N_9709,N_9719);
or UO_1179 (O_1179,N_9957,N_9614);
and UO_1180 (O_1180,N_9702,N_9669);
nand UO_1181 (O_1181,N_9754,N_9984);
nand UO_1182 (O_1182,N_9719,N_9784);
nor UO_1183 (O_1183,N_9649,N_9968);
xnor UO_1184 (O_1184,N_9651,N_9690);
and UO_1185 (O_1185,N_9980,N_9578);
nand UO_1186 (O_1186,N_9519,N_9564);
and UO_1187 (O_1187,N_9945,N_9750);
or UO_1188 (O_1188,N_9802,N_9881);
and UO_1189 (O_1189,N_9976,N_9585);
and UO_1190 (O_1190,N_9856,N_9751);
nand UO_1191 (O_1191,N_9994,N_9566);
nand UO_1192 (O_1192,N_9788,N_9795);
xnor UO_1193 (O_1193,N_9903,N_9741);
or UO_1194 (O_1194,N_9586,N_9964);
nor UO_1195 (O_1195,N_9947,N_9561);
or UO_1196 (O_1196,N_9793,N_9603);
nor UO_1197 (O_1197,N_9607,N_9951);
nor UO_1198 (O_1198,N_9512,N_9585);
xnor UO_1199 (O_1199,N_9695,N_9992);
xnor UO_1200 (O_1200,N_9912,N_9792);
nor UO_1201 (O_1201,N_9826,N_9934);
xnor UO_1202 (O_1202,N_9903,N_9813);
and UO_1203 (O_1203,N_9735,N_9789);
nor UO_1204 (O_1204,N_9942,N_9715);
xor UO_1205 (O_1205,N_9587,N_9577);
and UO_1206 (O_1206,N_9923,N_9585);
and UO_1207 (O_1207,N_9527,N_9644);
or UO_1208 (O_1208,N_9611,N_9671);
nand UO_1209 (O_1209,N_9548,N_9806);
nand UO_1210 (O_1210,N_9888,N_9604);
nor UO_1211 (O_1211,N_9994,N_9538);
and UO_1212 (O_1212,N_9679,N_9773);
nor UO_1213 (O_1213,N_9900,N_9838);
nor UO_1214 (O_1214,N_9670,N_9535);
or UO_1215 (O_1215,N_9616,N_9642);
or UO_1216 (O_1216,N_9773,N_9592);
nand UO_1217 (O_1217,N_9577,N_9794);
and UO_1218 (O_1218,N_9512,N_9673);
and UO_1219 (O_1219,N_9751,N_9831);
nor UO_1220 (O_1220,N_9543,N_9960);
and UO_1221 (O_1221,N_9680,N_9721);
and UO_1222 (O_1222,N_9741,N_9854);
nand UO_1223 (O_1223,N_9538,N_9678);
nand UO_1224 (O_1224,N_9841,N_9996);
nor UO_1225 (O_1225,N_9861,N_9774);
and UO_1226 (O_1226,N_9617,N_9752);
nand UO_1227 (O_1227,N_9747,N_9779);
or UO_1228 (O_1228,N_9570,N_9601);
xnor UO_1229 (O_1229,N_9943,N_9977);
or UO_1230 (O_1230,N_9749,N_9573);
nand UO_1231 (O_1231,N_9703,N_9947);
or UO_1232 (O_1232,N_9854,N_9562);
and UO_1233 (O_1233,N_9593,N_9913);
and UO_1234 (O_1234,N_9807,N_9577);
nand UO_1235 (O_1235,N_9550,N_9601);
or UO_1236 (O_1236,N_9654,N_9819);
xnor UO_1237 (O_1237,N_9645,N_9709);
and UO_1238 (O_1238,N_9841,N_9596);
nor UO_1239 (O_1239,N_9926,N_9881);
nand UO_1240 (O_1240,N_9927,N_9729);
nor UO_1241 (O_1241,N_9782,N_9950);
nand UO_1242 (O_1242,N_9667,N_9952);
or UO_1243 (O_1243,N_9629,N_9719);
or UO_1244 (O_1244,N_9754,N_9860);
nor UO_1245 (O_1245,N_9966,N_9976);
nand UO_1246 (O_1246,N_9680,N_9987);
xnor UO_1247 (O_1247,N_9836,N_9902);
nor UO_1248 (O_1248,N_9899,N_9877);
nor UO_1249 (O_1249,N_9775,N_9987);
or UO_1250 (O_1250,N_9626,N_9636);
nor UO_1251 (O_1251,N_9921,N_9719);
nand UO_1252 (O_1252,N_9973,N_9569);
and UO_1253 (O_1253,N_9880,N_9644);
or UO_1254 (O_1254,N_9847,N_9554);
nor UO_1255 (O_1255,N_9570,N_9649);
nor UO_1256 (O_1256,N_9707,N_9521);
nor UO_1257 (O_1257,N_9689,N_9521);
and UO_1258 (O_1258,N_9553,N_9814);
nand UO_1259 (O_1259,N_9613,N_9778);
nand UO_1260 (O_1260,N_9703,N_9762);
nor UO_1261 (O_1261,N_9737,N_9520);
nor UO_1262 (O_1262,N_9647,N_9822);
nand UO_1263 (O_1263,N_9974,N_9769);
nand UO_1264 (O_1264,N_9622,N_9864);
nand UO_1265 (O_1265,N_9672,N_9927);
or UO_1266 (O_1266,N_9627,N_9725);
nor UO_1267 (O_1267,N_9922,N_9804);
and UO_1268 (O_1268,N_9648,N_9733);
nor UO_1269 (O_1269,N_9699,N_9585);
nor UO_1270 (O_1270,N_9512,N_9947);
or UO_1271 (O_1271,N_9929,N_9791);
and UO_1272 (O_1272,N_9954,N_9641);
nand UO_1273 (O_1273,N_9925,N_9593);
or UO_1274 (O_1274,N_9749,N_9877);
and UO_1275 (O_1275,N_9977,N_9892);
nand UO_1276 (O_1276,N_9775,N_9533);
nor UO_1277 (O_1277,N_9983,N_9787);
nand UO_1278 (O_1278,N_9574,N_9560);
or UO_1279 (O_1279,N_9567,N_9506);
and UO_1280 (O_1280,N_9583,N_9734);
nor UO_1281 (O_1281,N_9518,N_9553);
and UO_1282 (O_1282,N_9689,N_9815);
nor UO_1283 (O_1283,N_9611,N_9868);
nand UO_1284 (O_1284,N_9903,N_9952);
xor UO_1285 (O_1285,N_9726,N_9796);
nand UO_1286 (O_1286,N_9884,N_9899);
nor UO_1287 (O_1287,N_9864,N_9738);
and UO_1288 (O_1288,N_9675,N_9764);
or UO_1289 (O_1289,N_9740,N_9927);
nand UO_1290 (O_1290,N_9778,N_9901);
nor UO_1291 (O_1291,N_9707,N_9595);
nor UO_1292 (O_1292,N_9540,N_9581);
and UO_1293 (O_1293,N_9729,N_9684);
and UO_1294 (O_1294,N_9675,N_9821);
and UO_1295 (O_1295,N_9988,N_9650);
or UO_1296 (O_1296,N_9504,N_9759);
xor UO_1297 (O_1297,N_9892,N_9677);
nand UO_1298 (O_1298,N_9618,N_9975);
or UO_1299 (O_1299,N_9537,N_9571);
nor UO_1300 (O_1300,N_9991,N_9792);
nor UO_1301 (O_1301,N_9660,N_9930);
nand UO_1302 (O_1302,N_9778,N_9630);
xor UO_1303 (O_1303,N_9821,N_9767);
nand UO_1304 (O_1304,N_9619,N_9774);
nand UO_1305 (O_1305,N_9831,N_9544);
nor UO_1306 (O_1306,N_9649,N_9945);
nor UO_1307 (O_1307,N_9632,N_9855);
or UO_1308 (O_1308,N_9988,N_9528);
or UO_1309 (O_1309,N_9544,N_9648);
and UO_1310 (O_1310,N_9779,N_9720);
or UO_1311 (O_1311,N_9680,N_9723);
nand UO_1312 (O_1312,N_9712,N_9794);
nand UO_1313 (O_1313,N_9818,N_9964);
nand UO_1314 (O_1314,N_9795,N_9770);
or UO_1315 (O_1315,N_9802,N_9882);
nor UO_1316 (O_1316,N_9916,N_9970);
or UO_1317 (O_1317,N_9600,N_9563);
and UO_1318 (O_1318,N_9787,N_9660);
nand UO_1319 (O_1319,N_9751,N_9880);
nor UO_1320 (O_1320,N_9662,N_9509);
and UO_1321 (O_1321,N_9861,N_9788);
nand UO_1322 (O_1322,N_9736,N_9779);
and UO_1323 (O_1323,N_9823,N_9618);
nor UO_1324 (O_1324,N_9929,N_9588);
and UO_1325 (O_1325,N_9915,N_9703);
or UO_1326 (O_1326,N_9919,N_9925);
or UO_1327 (O_1327,N_9504,N_9706);
and UO_1328 (O_1328,N_9786,N_9591);
or UO_1329 (O_1329,N_9701,N_9727);
or UO_1330 (O_1330,N_9915,N_9909);
and UO_1331 (O_1331,N_9884,N_9942);
nor UO_1332 (O_1332,N_9933,N_9586);
or UO_1333 (O_1333,N_9709,N_9599);
or UO_1334 (O_1334,N_9661,N_9794);
and UO_1335 (O_1335,N_9875,N_9504);
or UO_1336 (O_1336,N_9864,N_9951);
nand UO_1337 (O_1337,N_9811,N_9728);
or UO_1338 (O_1338,N_9695,N_9832);
nand UO_1339 (O_1339,N_9712,N_9577);
and UO_1340 (O_1340,N_9931,N_9944);
nor UO_1341 (O_1341,N_9686,N_9736);
or UO_1342 (O_1342,N_9908,N_9682);
nand UO_1343 (O_1343,N_9526,N_9935);
nand UO_1344 (O_1344,N_9578,N_9992);
nand UO_1345 (O_1345,N_9528,N_9639);
nor UO_1346 (O_1346,N_9755,N_9771);
nor UO_1347 (O_1347,N_9734,N_9589);
or UO_1348 (O_1348,N_9808,N_9754);
nor UO_1349 (O_1349,N_9908,N_9541);
and UO_1350 (O_1350,N_9612,N_9846);
nor UO_1351 (O_1351,N_9887,N_9504);
or UO_1352 (O_1352,N_9519,N_9508);
xor UO_1353 (O_1353,N_9515,N_9748);
xor UO_1354 (O_1354,N_9620,N_9904);
and UO_1355 (O_1355,N_9868,N_9900);
or UO_1356 (O_1356,N_9929,N_9795);
or UO_1357 (O_1357,N_9927,N_9939);
and UO_1358 (O_1358,N_9662,N_9850);
and UO_1359 (O_1359,N_9519,N_9577);
and UO_1360 (O_1360,N_9722,N_9629);
and UO_1361 (O_1361,N_9613,N_9963);
nor UO_1362 (O_1362,N_9791,N_9915);
nand UO_1363 (O_1363,N_9890,N_9798);
xnor UO_1364 (O_1364,N_9694,N_9530);
or UO_1365 (O_1365,N_9546,N_9685);
nand UO_1366 (O_1366,N_9655,N_9704);
or UO_1367 (O_1367,N_9668,N_9598);
or UO_1368 (O_1368,N_9913,N_9622);
and UO_1369 (O_1369,N_9717,N_9672);
or UO_1370 (O_1370,N_9557,N_9939);
and UO_1371 (O_1371,N_9785,N_9674);
nand UO_1372 (O_1372,N_9748,N_9620);
xor UO_1373 (O_1373,N_9703,N_9774);
nor UO_1374 (O_1374,N_9926,N_9729);
and UO_1375 (O_1375,N_9874,N_9598);
xor UO_1376 (O_1376,N_9541,N_9845);
nor UO_1377 (O_1377,N_9550,N_9761);
nor UO_1378 (O_1378,N_9555,N_9626);
nand UO_1379 (O_1379,N_9873,N_9984);
or UO_1380 (O_1380,N_9916,N_9549);
nand UO_1381 (O_1381,N_9923,N_9612);
nor UO_1382 (O_1382,N_9510,N_9743);
and UO_1383 (O_1383,N_9770,N_9732);
or UO_1384 (O_1384,N_9593,N_9640);
or UO_1385 (O_1385,N_9820,N_9957);
nand UO_1386 (O_1386,N_9620,N_9608);
or UO_1387 (O_1387,N_9605,N_9804);
nor UO_1388 (O_1388,N_9623,N_9874);
or UO_1389 (O_1389,N_9648,N_9519);
and UO_1390 (O_1390,N_9601,N_9987);
nor UO_1391 (O_1391,N_9683,N_9746);
and UO_1392 (O_1392,N_9535,N_9567);
nand UO_1393 (O_1393,N_9982,N_9920);
and UO_1394 (O_1394,N_9522,N_9946);
nand UO_1395 (O_1395,N_9824,N_9643);
xor UO_1396 (O_1396,N_9963,N_9663);
xor UO_1397 (O_1397,N_9806,N_9783);
and UO_1398 (O_1398,N_9711,N_9899);
or UO_1399 (O_1399,N_9567,N_9615);
nor UO_1400 (O_1400,N_9728,N_9947);
and UO_1401 (O_1401,N_9874,N_9568);
nand UO_1402 (O_1402,N_9884,N_9810);
nor UO_1403 (O_1403,N_9891,N_9706);
nor UO_1404 (O_1404,N_9687,N_9561);
nand UO_1405 (O_1405,N_9680,N_9870);
or UO_1406 (O_1406,N_9601,N_9612);
nand UO_1407 (O_1407,N_9686,N_9987);
or UO_1408 (O_1408,N_9788,N_9625);
nand UO_1409 (O_1409,N_9784,N_9555);
and UO_1410 (O_1410,N_9752,N_9534);
nor UO_1411 (O_1411,N_9512,N_9908);
nor UO_1412 (O_1412,N_9771,N_9664);
nor UO_1413 (O_1413,N_9741,N_9668);
xor UO_1414 (O_1414,N_9972,N_9616);
nor UO_1415 (O_1415,N_9775,N_9549);
nor UO_1416 (O_1416,N_9595,N_9795);
and UO_1417 (O_1417,N_9659,N_9894);
nor UO_1418 (O_1418,N_9762,N_9554);
nand UO_1419 (O_1419,N_9934,N_9571);
nor UO_1420 (O_1420,N_9746,N_9701);
nor UO_1421 (O_1421,N_9621,N_9782);
and UO_1422 (O_1422,N_9749,N_9636);
nor UO_1423 (O_1423,N_9916,N_9651);
nor UO_1424 (O_1424,N_9768,N_9967);
nand UO_1425 (O_1425,N_9937,N_9626);
nor UO_1426 (O_1426,N_9530,N_9576);
or UO_1427 (O_1427,N_9576,N_9679);
and UO_1428 (O_1428,N_9736,N_9551);
nand UO_1429 (O_1429,N_9977,N_9544);
nand UO_1430 (O_1430,N_9741,N_9729);
and UO_1431 (O_1431,N_9594,N_9710);
xor UO_1432 (O_1432,N_9541,N_9723);
or UO_1433 (O_1433,N_9516,N_9988);
xor UO_1434 (O_1434,N_9533,N_9988);
nor UO_1435 (O_1435,N_9876,N_9986);
or UO_1436 (O_1436,N_9744,N_9819);
and UO_1437 (O_1437,N_9933,N_9854);
or UO_1438 (O_1438,N_9857,N_9717);
and UO_1439 (O_1439,N_9586,N_9856);
and UO_1440 (O_1440,N_9889,N_9561);
nor UO_1441 (O_1441,N_9509,N_9783);
nand UO_1442 (O_1442,N_9579,N_9510);
or UO_1443 (O_1443,N_9757,N_9971);
and UO_1444 (O_1444,N_9915,N_9806);
xnor UO_1445 (O_1445,N_9846,N_9542);
xnor UO_1446 (O_1446,N_9513,N_9516);
nand UO_1447 (O_1447,N_9888,N_9802);
and UO_1448 (O_1448,N_9954,N_9819);
xnor UO_1449 (O_1449,N_9689,N_9670);
nand UO_1450 (O_1450,N_9838,N_9624);
nand UO_1451 (O_1451,N_9923,N_9542);
nor UO_1452 (O_1452,N_9800,N_9821);
nand UO_1453 (O_1453,N_9634,N_9750);
nor UO_1454 (O_1454,N_9512,N_9727);
nand UO_1455 (O_1455,N_9853,N_9828);
nor UO_1456 (O_1456,N_9992,N_9914);
or UO_1457 (O_1457,N_9600,N_9707);
and UO_1458 (O_1458,N_9784,N_9819);
and UO_1459 (O_1459,N_9897,N_9586);
and UO_1460 (O_1460,N_9701,N_9849);
nor UO_1461 (O_1461,N_9542,N_9844);
and UO_1462 (O_1462,N_9937,N_9845);
nand UO_1463 (O_1463,N_9997,N_9785);
or UO_1464 (O_1464,N_9813,N_9502);
and UO_1465 (O_1465,N_9577,N_9602);
and UO_1466 (O_1466,N_9617,N_9921);
nor UO_1467 (O_1467,N_9553,N_9697);
and UO_1468 (O_1468,N_9665,N_9963);
nand UO_1469 (O_1469,N_9650,N_9862);
nand UO_1470 (O_1470,N_9844,N_9550);
and UO_1471 (O_1471,N_9570,N_9992);
or UO_1472 (O_1472,N_9632,N_9923);
nand UO_1473 (O_1473,N_9812,N_9628);
and UO_1474 (O_1474,N_9712,N_9701);
xor UO_1475 (O_1475,N_9574,N_9876);
xnor UO_1476 (O_1476,N_9910,N_9872);
nor UO_1477 (O_1477,N_9915,N_9624);
and UO_1478 (O_1478,N_9932,N_9575);
xor UO_1479 (O_1479,N_9952,N_9856);
and UO_1480 (O_1480,N_9513,N_9636);
xnor UO_1481 (O_1481,N_9922,N_9602);
nor UO_1482 (O_1482,N_9861,N_9531);
nand UO_1483 (O_1483,N_9540,N_9919);
nand UO_1484 (O_1484,N_9765,N_9680);
and UO_1485 (O_1485,N_9521,N_9926);
xor UO_1486 (O_1486,N_9909,N_9703);
and UO_1487 (O_1487,N_9637,N_9500);
and UO_1488 (O_1488,N_9684,N_9865);
nor UO_1489 (O_1489,N_9603,N_9791);
and UO_1490 (O_1490,N_9634,N_9608);
or UO_1491 (O_1491,N_9650,N_9831);
nand UO_1492 (O_1492,N_9910,N_9911);
and UO_1493 (O_1493,N_9952,N_9558);
or UO_1494 (O_1494,N_9737,N_9749);
nor UO_1495 (O_1495,N_9872,N_9516);
or UO_1496 (O_1496,N_9528,N_9623);
nor UO_1497 (O_1497,N_9753,N_9726);
nor UO_1498 (O_1498,N_9864,N_9798);
nand UO_1499 (O_1499,N_9518,N_9715);
endmodule