module basic_2000_20000_2500_25_levels_10xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
xnor U0 (N_0,In_321,In_221);
and U1 (N_1,In_1960,In_1601);
xnor U2 (N_2,In_462,In_101);
xor U3 (N_3,In_6,In_446);
nor U4 (N_4,In_1616,In_661);
nor U5 (N_5,In_977,In_517);
nor U6 (N_6,In_738,In_1031);
nand U7 (N_7,In_1723,In_237);
xor U8 (N_8,In_482,In_288);
or U9 (N_9,In_1227,In_114);
or U10 (N_10,In_25,In_1921);
nand U11 (N_11,In_861,In_1225);
and U12 (N_12,In_539,In_1309);
nand U13 (N_13,In_197,In_1709);
or U14 (N_14,In_1846,In_1911);
nor U15 (N_15,In_1537,In_55);
nor U16 (N_16,In_1166,In_1107);
nor U17 (N_17,In_1974,In_1062);
and U18 (N_18,In_1705,In_1288);
nand U19 (N_19,In_502,In_790);
or U20 (N_20,In_1057,In_1777);
xor U21 (N_21,In_1794,In_1170);
xnor U22 (N_22,In_1732,In_1009);
xor U23 (N_23,In_917,In_1736);
and U24 (N_24,In_607,In_80);
xnor U25 (N_25,In_1180,In_1121);
nand U26 (N_26,In_1536,In_1204);
nor U27 (N_27,In_200,In_954);
nor U28 (N_28,In_1895,In_807);
xnor U29 (N_29,In_27,In_813);
nor U30 (N_30,In_1269,In_447);
xnor U31 (N_31,In_901,In_817);
and U32 (N_32,In_1764,In_1002);
or U33 (N_33,In_995,In_561);
nand U34 (N_34,In_1237,In_425);
xor U35 (N_35,In_26,In_501);
xnor U36 (N_36,In_318,In_1967);
and U37 (N_37,In_928,In_1560);
and U38 (N_38,In_991,In_1980);
xor U39 (N_39,In_593,In_492);
xor U40 (N_40,In_54,In_1864);
xor U41 (N_41,In_1702,In_1014);
nor U42 (N_42,In_30,In_1482);
or U43 (N_43,In_240,In_793);
nor U44 (N_44,In_435,In_192);
nor U45 (N_45,In_835,In_131);
and U46 (N_46,In_1868,In_879);
and U47 (N_47,In_1724,In_1826);
nor U48 (N_48,In_1428,In_49);
or U49 (N_49,In_1158,In_1966);
xnor U50 (N_50,In_859,In_716);
and U51 (N_51,In_1909,In_557);
nor U52 (N_52,In_1138,In_15);
xnor U53 (N_53,In_400,In_693);
nand U54 (N_54,In_1359,In_1594);
or U55 (N_55,In_1985,In_1645);
xor U56 (N_56,In_1042,In_183);
xnor U57 (N_57,In_189,In_575);
xor U58 (N_58,In_235,In_1618);
nor U59 (N_59,In_1215,In_1373);
xnor U60 (N_60,In_947,In_1169);
nand U61 (N_61,In_1573,In_1712);
xor U62 (N_62,In_1882,In_1234);
xnor U63 (N_63,In_1788,In_1001);
and U64 (N_64,In_1197,In_1916);
xor U65 (N_65,In_1684,In_249);
nor U66 (N_66,In_1174,In_338);
xor U67 (N_67,In_1605,In_1382);
xor U68 (N_68,In_1572,In_184);
xnor U69 (N_69,In_1737,In_260);
nor U70 (N_70,In_7,In_572);
xor U71 (N_71,In_128,In_1123);
nor U72 (N_72,In_1876,In_1196);
or U73 (N_73,In_463,In_215);
nor U74 (N_74,In_1703,In_1746);
or U75 (N_75,In_1642,In_1209);
nand U76 (N_76,In_914,In_246);
xor U77 (N_77,In_1155,In_1187);
and U78 (N_78,In_1790,In_1606);
and U79 (N_79,In_426,In_907);
nor U80 (N_80,In_1256,In_725);
nand U81 (N_81,In_1451,In_550);
and U82 (N_82,In_946,In_1579);
nor U83 (N_83,In_984,In_852);
nand U84 (N_84,In_353,In_284);
and U85 (N_85,In_1026,In_1816);
xnor U86 (N_86,In_1348,In_608);
nor U87 (N_87,In_1072,In_698);
and U88 (N_88,In_350,In_133);
or U89 (N_89,In_935,In_1625);
or U90 (N_90,In_826,In_1324);
nor U91 (N_91,In_831,In_1938);
or U92 (N_92,In_1964,In_589);
xor U93 (N_93,In_1937,In_733);
nor U94 (N_94,In_553,In_409);
xor U95 (N_95,In_708,In_1664);
and U96 (N_96,In_1733,In_180);
xor U97 (N_97,In_1052,In_1263);
xor U98 (N_98,In_1887,In_1784);
or U99 (N_99,In_1507,In_1306);
and U100 (N_100,In_228,In_1275);
nor U101 (N_101,In_1831,In_1884);
or U102 (N_102,In_1803,In_1167);
xnor U103 (N_103,In_1978,In_90);
nand U104 (N_104,In_1135,In_1946);
nor U105 (N_105,In_354,In_293);
or U106 (N_106,In_538,In_270);
or U107 (N_107,In_1617,In_1693);
nand U108 (N_108,In_1218,In_1115);
nor U109 (N_109,In_1294,In_1710);
and U110 (N_110,In_792,In_1929);
xnor U111 (N_111,In_1795,In_579);
nand U112 (N_112,In_691,In_66);
nor U113 (N_113,In_1731,In_808);
xor U114 (N_114,In_581,In_703);
or U115 (N_115,In_834,In_729);
or U116 (N_116,In_1436,In_412);
xor U117 (N_117,In_336,In_4);
nor U118 (N_118,In_1786,In_920);
nor U119 (N_119,In_1162,In_311);
nand U120 (N_120,In_1580,In_1700);
xor U121 (N_121,In_10,In_1674);
nor U122 (N_122,In_543,In_69);
or U123 (N_123,In_1302,In_457);
nand U124 (N_124,In_1010,In_1999);
or U125 (N_125,In_1927,In_1249);
or U126 (N_126,In_747,In_1201);
xor U127 (N_127,In_844,In_1818);
nor U128 (N_128,In_1976,In_1137);
xnor U129 (N_129,In_689,In_1182);
and U130 (N_130,In_818,In_345);
or U131 (N_131,In_194,In_1388);
nand U132 (N_132,In_1149,In_1479);
nor U133 (N_133,In_771,In_452);
nand U134 (N_134,In_1644,In_1726);
xor U135 (N_135,In_1983,In_1599);
nand U136 (N_136,In_1393,In_1379);
xnor U137 (N_137,In_1060,In_1833);
nand U138 (N_138,In_290,In_374);
or U139 (N_139,In_1638,In_81);
and U140 (N_140,In_1207,In_700);
xor U141 (N_141,In_1993,In_810);
or U142 (N_142,In_364,In_1953);
or U143 (N_143,In_1200,In_1856);
nor U144 (N_144,In_437,In_1516);
xnor U145 (N_145,In_1763,In_532);
nand U146 (N_146,In_281,In_1143);
and U147 (N_147,In_20,In_666);
xor U148 (N_148,In_76,In_198);
or U149 (N_149,In_672,In_1793);
xor U150 (N_150,In_1295,In_1087);
and U151 (N_151,In_886,In_1841);
nor U152 (N_152,In_1719,In_450);
or U153 (N_153,In_408,In_1741);
nor U154 (N_154,In_1779,In_1472);
and U155 (N_155,In_1319,In_1098);
and U156 (N_156,In_798,In_868);
or U157 (N_157,In_1040,In_1203);
xor U158 (N_158,In_85,In_784);
nor U159 (N_159,In_1963,In_781);
or U160 (N_160,In_1238,In_626);
nor U161 (N_161,In_1792,In_1270);
or U162 (N_162,In_1992,In_1695);
nor U163 (N_163,In_1478,In_829);
nand U164 (N_164,In_299,In_1609);
nor U165 (N_165,In_201,In_1535);
nor U166 (N_166,In_1036,In_1465);
xnor U167 (N_167,In_1151,In_277);
or U168 (N_168,In_420,In_331);
nand U169 (N_169,In_199,In_1340);
nand U170 (N_170,In_758,In_1758);
and U171 (N_171,In_57,In_418);
nor U172 (N_172,In_1932,In_443);
nand U173 (N_173,In_578,In_851);
xor U174 (N_174,In_778,In_948);
nor U175 (N_175,In_735,In_1076);
nor U176 (N_176,In_204,In_448);
or U177 (N_177,In_596,In_1530);
nand U178 (N_178,In_1113,In_1823);
xor U179 (N_179,In_1094,In_1520);
and U180 (N_180,In_1972,In_1007);
nor U181 (N_181,In_1564,In_349);
and U182 (N_182,In_279,In_1286);
xnor U183 (N_183,In_505,In_205);
and U184 (N_184,In_1531,In_1172);
and U185 (N_185,In_1216,In_1636);
or U186 (N_186,In_1171,In_261);
nand U187 (N_187,In_1728,In_1358);
or U188 (N_188,In_1041,In_1493);
xnor U189 (N_189,In_1752,In_60);
xor U190 (N_190,In_782,In_1517);
xor U191 (N_191,In_1232,In_148);
or U192 (N_192,In_1088,In_653);
nor U193 (N_193,In_1212,In_1033);
nand U194 (N_194,In_1375,In_348);
and U195 (N_195,In_1673,In_1631);
nand U196 (N_196,In_695,In_1523);
or U197 (N_197,In_1406,In_1059);
xnor U198 (N_198,In_777,In_820);
and U199 (N_199,In_1152,In_1103);
nand U200 (N_200,In_1308,In_1979);
and U201 (N_201,In_509,In_625);
xnor U202 (N_202,In_1017,In_187);
xnor U203 (N_203,In_1338,In_323);
or U204 (N_204,In_1192,In_1679);
nand U205 (N_205,In_1510,In_206);
and U206 (N_206,In_1205,In_1304);
nand U207 (N_207,In_1813,In_1410);
nor U208 (N_208,In_849,In_171);
nand U209 (N_209,In_874,In_507);
or U210 (N_210,In_179,In_75);
nand U211 (N_211,In_1383,In_245);
and U212 (N_212,In_1527,In_1142);
xnor U213 (N_213,In_930,In_1875);
or U214 (N_214,In_1329,In_1092);
and U215 (N_215,In_774,In_759);
and U216 (N_216,In_526,In_992);
and U217 (N_217,In_1783,In_497);
xor U218 (N_218,In_862,In_461);
and U219 (N_219,In_961,In_1716);
and U220 (N_220,In_1814,In_1854);
xor U221 (N_221,In_1504,In_150);
or U222 (N_222,In_1900,In_922);
nand U223 (N_223,In_1769,In_1988);
xnor U224 (N_224,In_117,In_306);
nand U225 (N_225,In_1903,In_1879);
nand U226 (N_226,In_938,In_393);
and U227 (N_227,In_91,In_1547);
nand U228 (N_228,In_1004,In_503);
nand U229 (N_229,In_602,In_1651);
or U230 (N_230,In_1133,In_255);
and U231 (N_231,In_1396,In_706);
nand U232 (N_232,In_756,In_540);
and U233 (N_233,In_337,In_52);
nand U234 (N_234,In_48,In_51);
xnor U235 (N_235,In_1347,In_949);
nand U236 (N_236,In_1184,In_1614);
nor U237 (N_237,In_1917,In_42);
nand U238 (N_238,In_588,In_1655);
or U239 (N_239,In_1415,In_1549);
xor U240 (N_240,In_1186,In_1633);
xnor U241 (N_241,In_1046,In_1539);
nand U242 (N_242,In_1771,In_795);
and U243 (N_243,In_865,In_259);
nor U244 (N_244,In_1146,In_1476);
or U245 (N_245,In_1409,In_944);
nand U246 (N_246,In_1420,In_79);
or U247 (N_247,In_483,In_1297);
or U248 (N_248,In_139,In_1093);
nand U249 (N_249,In_116,In_903);
or U250 (N_250,In_847,In_1247);
nand U251 (N_251,In_1449,In_713);
or U252 (N_252,In_29,In_969);
and U253 (N_253,In_833,In_1647);
or U254 (N_254,In_686,In_1397);
nor U255 (N_255,In_1807,In_1584);
and U256 (N_256,In_659,In_1267);
and U257 (N_257,In_1910,In_1110);
xnor U258 (N_258,In_772,In_508);
and U259 (N_259,In_1637,In_1598);
xor U260 (N_260,In_1429,In_1254);
nor U261 (N_261,In_1511,In_732);
nor U262 (N_262,In_1824,In_341);
xor U263 (N_263,In_1658,In_981);
nor U264 (N_264,In_1130,In_1571);
or U265 (N_265,In_803,In_86);
and U266 (N_266,In_398,In_170);
and U267 (N_267,In_1683,In_1013);
nand U268 (N_268,In_568,In_1287);
or U269 (N_269,In_639,In_1915);
nor U270 (N_270,In_1283,In_225);
and U271 (N_271,In_1284,In_1280);
and U272 (N_272,In_824,In_1939);
and U273 (N_273,In_1116,In_35);
and U274 (N_274,In_478,In_770);
or U275 (N_275,In_344,In_366);
nand U276 (N_276,In_1176,In_431);
and U277 (N_277,In_1652,In_641);
and U278 (N_278,In_1157,In_993);
nor U279 (N_279,In_1492,In_905);
nor U280 (N_280,In_1150,In_89);
nor U281 (N_281,In_728,In_178);
nand U282 (N_282,In_9,In_1320);
or U283 (N_283,In_1713,In_1643);
xnor U284 (N_284,In_1055,In_994);
xnor U285 (N_285,In_165,In_1498);
xor U286 (N_286,In_564,In_1495);
nor U287 (N_287,In_889,In_763);
xnor U288 (N_288,In_1469,In_335);
nand U289 (N_289,In_1131,In_968);
xnor U290 (N_290,In_387,In_1778);
or U291 (N_291,In_1470,In_1483);
xnor U292 (N_292,In_815,In_1889);
and U293 (N_293,In_1687,In_779);
or U294 (N_294,In_241,In_966);
nor U295 (N_295,In_796,In_1292);
nand U296 (N_296,In_1961,In_762);
and U297 (N_297,In_1563,In_1852);
xor U298 (N_298,In_1540,In_32);
nor U299 (N_299,In_1933,In_1127);
xor U300 (N_300,In_1202,In_1097);
xor U301 (N_301,In_1754,In_1872);
xor U302 (N_302,In_1159,In_1820);
nand U303 (N_303,In_748,In_326);
or U304 (N_304,In_1424,In_1117);
and U305 (N_305,In_670,In_972);
nor U306 (N_306,In_528,In_1734);
and U307 (N_307,In_811,In_1740);
or U308 (N_308,In_1252,In_1086);
nor U309 (N_309,In_1049,In_923);
nand U310 (N_310,In_1385,In_952);
xnor U311 (N_311,In_1891,In_481);
xor U312 (N_312,In_681,In_552);
xor U313 (N_313,In_1663,In_1799);
and U314 (N_314,In_357,In_1805);
and U315 (N_315,In_1995,In_702);
or U316 (N_316,In_330,In_379);
xor U317 (N_317,In_858,In_1721);
nor U318 (N_318,In_432,In_195);
or U319 (N_319,In_378,In_1370);
nand U320 (N_320,In_709,In_876);
nor U321 (N_321,In_1578,In_1084);
nand U322 (N_322,In_1914,In_814);
or U323 (N_323,In_942,In_1045);
and U324 (N_324,In_1838,In_8);
or U325 (N_325,In_1529,In_1595);
or U326 (N_326,In_1096,In_1906);
or U327 (N_327,In_268,In_1378);
nand U328 (N_328,In_1211,In_328);
xnor U329 (N_329,In_127,In_678);
nand U330 (N_330,In_904,In_263);
nor U331 (N_331,In_797,In_1800);
and U332 (N_332,In_1941,In_519);
or U333 (N_333,In_106,In_971);
nand U334 (N_334,In_253,In_1230);
or U335 (N_335,In_606,In_1522);
nor U336 (N_336,In_877,In_1812);
nor U337 (N_337,In_1859,In_989);
nor U338 (N_338,In_1969,In_612);
xor U339 (N_339,In_1890,In_1468);
or U340 (N_340,In_222,In_624);
nor U341 (N_341,In_866,In_1973);
or U342 (N_342,In_514,In_1592);
nor U343 (N_343,In_1437,In_872);
and U344 (N_344,In_1119,In_1078);
xor U345 (N_345,In_363,In_1623);
or U346 (N_346,In_1787,In_1899);
nand U347 (N_347,In_137,In_1441);
xor U348 (N_348,In_24,In_173);
or U349 (N_349,In_1989,In_1821);
nand U350 (N_350,In_0,In_878);
nand U351 (N_351,In_43,In_123);
nor U352 (N_352,In_1715,In_751);
xor U353 (N_353,In_1661,In_453);
and U354 (N_354,In_635,In_513);
and U355 (N_355,In_959,In_130);
nand U356 (N_356,In_1717,In_975);
xor U357 (N_357,In_1694,In_518);
and U358 (N_358,In_753,In_120);
nor U359 (N_359,In_682,In_1222);
xnor U360 (N_360,In_1738,In_1688);
or U361 (N_361,In_1129,In_34);
and U362 (N_362,In_1847,In_1108);
nand U363 (N_363,In_474,In_664);
nand U364 (N_364,In_812,In_1836);
nor U365 (N_365,In_1641,In_64);
nor U366 (N_366,In_498,In_303);
xor U367 (N_367,In_1317,In_1386);
nand U368 (N_368,In_1405,In_40);
nand U369 (N_369,In_719,In_111);
or U370 (N_370,In_651,In_47);
nand U371 (N_371,In_1105,In_283);
and U372 (N_372,In_58,In_1809);
nand U373 (N_373,In_1112,In_285);
nor U374 (N_374,In_848,In_599);
xnor U375 (N_375,In_1878,In_362);
nor U376 (N_376,In_207,In_1646);
or U377 (N_377,In_68,In_1902);
or U378 (N_378,In_1278,In_368);
and U379 (N_379,In_1928,In_282);
nor U380 (N_380,In_1952,In_1653);
and U381 (N_381,In_1438,In_512);
and U382 (N_382,In_990,In_1228);
or U383 (N_383,In_1426,In_309);
xor U384 (N_384,In_1491,In_609);
nand U385 (N_385,In_1568,In_1006);
nand U386 (N_386,In_98,In_1901);
nor U387 (N_387,In_718,In_1350);
and U388 (N_388,In_1926,In_669);
nand U389 (N_389,In_415,In_67);
or U390 (N_390,In_551,In_1525);
or U391 (N_391,In_1380,In_1950);
or U392 (N_392,In_622,In_1043);
nand U393 (N_393,In_1274,In_1081);
nand U394 (N_394,In_663,In_438);
nand U395 (N_395,In_1349,In_1221);
nand U396 (N_396,In_645,In_1880);
and U397 (N_397,In_1257,In_953);
nand U398 (N_398,In_1650,In_610);
nand U399 (N_399,In_1355,In_1848);
nand U400 (N_400,In_458,In_757);
or U401 (N_401,In_186,In_224);
nor U402 (N_402,In_791,In_427);
and U403 (N_403,In_843,In_1219);
or U404 (N_404,In_921,In_1016);
or U405 (N_405,In_1817,In_875);
xor U406 (N_406,In_1051,In_59);
and U407 (N_407,In_146,In_271);
nand U408 (N_408,In_915,In_1354);
and U409 (N_409,In_422,In_499);
and U410 (N_410,In_533,In_77);
nor U411 (N_411,In_1871,In_1487);
xnor U412 (N_412,In_822,In_524);
nor U413 (N_413,In_1834,In_216);
or U414 (N_414,In_188,In_740);
xor U415 (N_415,In_737,In_2);
xnor U416 (N_416,In_1789,In_830);
nor U417 (N_417,In_1070,In_1676);
xor U418 (N_418,In_1153,In_883);
and U419 (N_419,In_1815,In_1407);
nand U420 (N_420,In_573,In_1725);
nand U421 (N_421,In_1615,In_372);
xor U422 (N_422,In_1832,In_900);
xnor U423 (N_423,In_119,In_1949);
nor U424 (N_424,In_683,In_1632);
nand U425 (N_425,In_380,In_761);
nor U426 (N_426,In_857,In_684);
nand U427 (N_427,In_1067,In_21);
nor U428 (N_428,In_125,In_1444);
xnor U429 (N_429,In_244,In_1691);
xnor U430 (N_430,In_494,In_908);
xor U431 (N_431,In_1063,In_618);
xnor U432 (N_432,In_804,In_1611);
nand U433 (N_433,In_722,In_1797);
xnor U434 (N_434,In_1075,In_717);
nand U435 (N_435,In_1582,In_1554);
xnor U436 (N_436,In_1583,In_1392);
nand U437 (N_437,In_1839,In_272);
nand U438 (N_438,In_1000,In_1685);
nor U439 (N_439,In_675,In_1660);
and U440 (N_440,In_82,In_1865);
nand U441 (N_441,In_1332,In_1873);
or U442 (N_442,In_1745,In_1480);
xor U443 (N_443,In_1125,In_637);
or U444 (N_444,In_1447,In_155);
nor U445 (N_445,In_1990,In_776);
xor U446 (N_446,In_1047,In_1161);
xnor U447 (N_447,In_1048,In_1714);
nor U448 (N_448,In_162,In_1904);
nor U449 (N_449,In_118,In_247);
nor U450 (N_450,In_699,In_1253);
xnor U451 (N_451,In_296,In_1243);
xnor U452 (N_452,In_1073,In_401);
nor U453 (N_453,In_95,In_510);
xnor U454 (N_454,In_1515,In_1669);
and U455 (N_455,In_662,In_1056);
or U456 (N_456,In_1208,In_1500);
nand U457 (N_457,In_405,In_1488);
and U458 (N_458,In_1387,In_175);
xnor U459 (N_459,In_1453,In_460);
nand U460 (N_460,In_710,In_965);
and U461 (N_461,In_74,In_1240);
nand U462 (N_462,In_1178,In_151);
xnor U463 (N_463,In_1439,In_1154);
and U464 (N_464,In_1277,In_1519);
nor U465 (N_465,In_1851,In_1262);
and U466 (N_466,In_549,In_1610);
and U467 (N_467,In_18,In_369);
xor U468 (N_468,In_628,In_870);
nand U469 (N_469,In_1281,In_1279);
nand U470 (N_470,In_692,In_1066);
and U471 (N_471,In_500,In_1394);
nand U472 (N_472,In_329,In_1558);
and U473 (N_473,In_1991,In_266);
and U474 (N_474,In_99,In_1321);
nor U475 (N_475,In_1089,In_143);
nand U476 (N_476,In_102,In_1255);
xor U477 (N_477,In_160,In_1518);
nand U478 (N_478,In_613,In_1408);
and U479 (N_479,In_548,In_1160);
and U480 (N_480,In_960,In_308);
or U481 (N_481,In_230,In_227);
xor U482 (N_482,In_730,In_853);
and U483 (N_483,In_906,In_1432);
xnor U484 (N_484,In_487,In_1639);
or U485 (N_485,In_1411,In_1399);
nor U486 (N_486,In_1775,In_72);
nor U487 (N_487,In_214,In_1496);
and U488 (N_488,In_562,In_1603);
nand U489 (N_489,In_388,In_97);
and U490 (N_490,In_1862,In_1503);
xor U491 (N_491,In_600,In_712);
or U492 (N_492,In_1104,In_891);
nand U493 (N_493,In_304,In_50);
or U494 (N_494,In_5,In_1885);
nor U495 (N_495,In_373,In_773);
or U496 (N_496,In_1509,In_1682);
nor U497 (N_497,In_1260,In_1044);
nor U498 (N_498,In_367,In_1924);
xnor U499 (N_499,In_495,In_210);
nand U500 (N_500,In_1604,In_576);
nand U501 (N_501,In_1672,In_258);
or U502 (N_502,In_856,In_355);
nor U503 (N_503,In_1473,In_1220);
or U504 (N_504,In_1955,In_1090);
and U505 (N_505,In_1587,In_816);
xnor U506 (N_506,In_1414,In_141);
xor U507 (N_507,In_775,In_1445);
or U508 (N_508,In_1223,In_322);
xor U509 (N_509,In_1401,In_396);
and U510 (N_510,In_1671,In_1586);
and U511 (N_511,In_1344,In_1804);
and U512 (N_512,In_1389,In_87);
and U513 (N_513,In_752,In_1920);
nand U514 (N_514,In_1198,In_1199);
nand U515 (N_515,In_1542,In_1748);
xor U516 (N_516,In_1364,In_924);
and U517 (N_517,In_896,In_1984);
or U518 (N_518,In_1054,In_1126);
nand U519 (N_519,In_1398,In_943);
and U520 (N_520,In_1058,In_1322);
xor U521 (N_521,In_1689,In_407);
nand U522 (N_522,In_736,In_1467);
nor U523 (N_523,In_1521,In_397);
or U524 (N_524,In_636,In_1248);
xnor U525 (N_525,In_998,In_1956);
and U526 (N_526,In_174,In_1061);
nand U527 (N_527,In_1311,In_1111);
xor U528 (N_528,In_1258,In_1753);
or U529 (N_529,In_1597,In_940);
xnor U530 (N_530,In_441,In_1659);
and U531 (N_531,In_149,In_212);
or U532 (N_532,In_765,In_1231);
nand U533 (N_533,In_1,In_1464);
and U534 (N_534,In_1574,In_1942);
xor U535 (N_535,In_455,In_731);
nand U536 (N_536,In_647,In_129);
nand U537 (N_537,In_1968,In_1907);
or U538 (N_538,In_136,In_1305);
nand U539 (N_539,In_1621,In_1261);
xnor U540 (N_540,In_92,In_996);
and U541 (N_541,In_1919,In_301);
or U542 (N_542,In_332,In_384);
nand U543 (N_543,In_1886,In_100);
nand U544 (N_544,In_654,In_1139);
nor U545 (N_545,In_1893,In_1018);
or U546 (N_546,In_529,In_1629);
and U547 (N_547,In_1843,In_1801);
or U548 (N_548,In_1316,In_1341);
xor U549 (N_549,In_890,In_1772);
xor U550 (N_550,In_1471,In_142);
and U551 (N_551,In_1696,In_352);
nor U552 (N_552,In_193,In_1193);
nand U553 (N_553,In_571,In_1077);
xor U554 (N_554,In_383,In_537);
nor U555 (N_555,In_933,In_1462);
nand U556 (N_556,In_1524,In_305);
nand U557 (N_557,In_325,In_932);
xor U558 (N_558,In_931,In_1698);
nand U559 (N_559,In_46,In_287);
nand U560 (N_560,In_468,In_591);
or U561 (N_561,In_1459,In_1371);
xor U562 (N_562,In_36,In_334);
and U563 (N_563,In_1751,In_217);
and U564 (N_564,In_314,In_1352);
nand U565 (N_565,In_1704,In_1943);
nor U566 (N_566,In_749,In_410);
nand U567 (N_567,In_999,In_1484);
nor U568 (N_568,In_987,In_1226);
or U569 (N_569,In_1925,In_324);
xor U570 (N_570,In_714,In_1590);
nor U571 (N_571,In_1106,In_110);
or U572 (N_572,In_402,In_679);
and U573 (N_573,In_1315,In_1296);
nand U574 (N_574,In_1553,In_1082);
or U575 (N_575,In_899,In_1028);
nor U576 (N_576,In_1706,In_1246);
xnor U577 (N_577,In_1750,In_351);
xnor U578 (N_578,In_1217,In_1140);
nor U579 (N_579,In_1109,In_1177);
or U580 (N_580,In_1179,In_14);
and U581 (N_581,In_1034,In_1064);
nand U582 (N_582,In_1534,In_1781);
xnor U583 (N_583,In_1019,In_1577);
nand U584 (N_584,In_1293,In_1242);
nor U585 (N_585,In_799,In_436);
nand U586 (N_586,In_1742,In_11);
nand U587 (N_587,In_1767,In_1670);
or U588 (N_588,In_1124,In_640);
or U589 (N_589,In_94,In_542);
nand U590 (N_590,In_832,In_1550);
nor U591 (N_591,In_1970,In_634);
or U592 (N_592,In_1566,In_84);
xnor U593 (N_593,In_1640,In_1272);
nand U594 (N_594,In_73,In_1657);
and U595 (N_595,In_395,In_1883);
nor U596 (N_596,In_842,In_1289);
and U597 (N_597,In_745,In_361);
nand U598 (N_598,In_1635,In_769);
and U599 (N_599,In_556,In_787);
nand U600 (N_600,In_1079,In_1589);
or U601 (N_601,In_1923,In_252);
xnor U602 (N_602,In_33,In_1366);
nand U603 (N_603,In_108,In_973);
nor U604 (N_604,In_421,In_696);
and U605 (N_605,In_493,In_841);
nor U606 (N_606,In_371,In_615);
or U607 (N_607,In_504,In_208);
or U608 (N_608,In_577,In_153);
nand U609 (N_609,In_1918,In_919);
or U610 (N_610,In_232,In_658);
or U611 (N_611,In_456,In_411);
nand U612 (N_612,In_768,In_414);
xor U613 (N_613,In_694,In_544);
and U614 (N_614,In_1440,In_1877);
nor U615 (N_615,In_1330,In_1849);
or U616 (N_616,In_63,In_385);
and U617 (N_617,In_521,In_1313);
nor U618 (N_618,In_490,In_1291);
nand U619 (N_619,In_895,In_61);
or U620 (N_620,In_1457,In_825);
and U621 (N_621,In_1648,In_1023);
or U622 (N_622,In_887,In_1977);
xnor U623 (N_623,In_1335,In_1528);
xnor U624 (N_624,In_1128,In_535);
nand U625 (N_625,In_22,In_1622);
and U626 (N_626,In_1957,In_970);
nor U627 (N_627,In_1102,In_801);
xor U628 (N_628,In_780,In_677);
or U629 (N_629,In_416,In_604);
nor U630 (N_630,In_1501,In_1810);
and U631 (N_631,In_1181,In_276);
nand U632 (N_632,In_1423,In_1008);
or U633 (N_633,In_375,In_250);
xor U634 (N_634,In_925,In_264);
or U635 (N_635,In_860,In_333);
nor U636 (N_636,In_1840,In_1828);
and U637 (N_637,In_1768,In_1065);
and U638 (N_638,In_794,In_1749);
nand U639 (N_639,In_167,In_340);
xor U640 (N_640,In_65,In_121);
and U641 (N_641,In_377,In_1425);
or U642 (N_642,In_1863,In_1628);
and U643 (N_643,In_676,In_256);
or U644 (N_644,In_983,In_196);
nor U645 (N_645,In_1744,In_871);
nor U646 (N_646,In_1266,In_1376);
nand U647 (N_647,In_166,In_1756);
nor U648 (N_648,In_598,In_845);
xnor U649 (N_649,In_1761,In_1030);
and U650 (N_650,In_754,In_1191);
xor U651 (N_651,In_1585,In_1368);
or U652 (N_652,In_254,In_44);
and U653 (N_653,In_1037,In_1458);
nand U654 (N_654,In_916,In_1419);
and U655 (N_655,In_864,In_614);
xnor U656 (N_656,In_88,In_1720);
nor U657 (N_657,In_1268,In_838);
nand U658 (N_658,In_565,In_1837);
and U659 (N_659,In_1264,In_220);
and U660 (N_660,In_937,In_1548);
nor U661 (N_661,In_644,In_1497);
xor U662 (N_662,In_1858,In_1770);
and U663 (N_663,In_1325,In_1552);
and U664 (N_664,In_1224,In_957);
xor U665 (N_665,In_70,In_633);
and U666 (N_666,In_1326,In_711);
or U667 (N_667,In_1360,In_1802);
nor U668 (N_668,In_1431,In_746);
and U669 (N_669,In_819,In_1965);
xnor U670 (N_670,In_1798,In_632);
or U671 (N_671,In_1214,In_638);
nand U672 (N_672,In_1576,In_783);
or U673 (N_673,In_113,In_988);
and U674 (N_674,In_744,In_1374);
nor U675 (N_675,In_343,In_894);
xor U676 (N_676,In_1958,In_202);
nand U677 (N_677,In_1624,In_1333);
nor U678 (N_678,In_1163,In_980);
nor U679 (N_679,In_657,In_1811);
xor U680 (N_680,In_381,In_449);
nor U681 (N_681,In_1236,In_433);
and U682 (N_682,In_480,In_821);
or U683 (N_683,In_592,In_1656);
or U684 (N_684,In_419,In_1141);
or U685 (N_685,In_1541,In_1446);
nor U686 (N_686,In_1860,In_1512);
or U687 (N_687,In_1913,In_582);
nor U688 (N_688,In_1947,In_312);
nand U689 (N_689,In_1701,In_687);
and U690 (N_690,In_475,In_545);
or U691 (N_691,In_1251,In_665);
nor U692 (N_692,In_1168,In_884);
xnor U693 (N_693,In_1185,In_656);
nand U694 (N_694,In_233,In_190);
and U695 (N_695,In_484,In_1024);
and U696 (N_696,In_346,In_1194);
or U697 (N_697,In_1271,In_23);
and U698 (N_698,In_506,In_1020);
nand U699 (N_699,In_1427,In_885);
nand U700 (N_700,In_601,In_423);
or U701 (N_701,In_278,In_1912);
and U702 (N_702,In_464,In_1345);
or U703 (N_703,In_370,In_1692);
xnor U704 (N_704,In_1356,In_1759);
and U705 (N_705,In_1934,In_45);
nor U706 (N_706,In_1681,In_454);
or U707 (N_707,In_1935,In_103);
and U708 (N_708,In_1421,In_1662);
nor U709 (N_709,In_307,In_951);
xor U710 (N_710,In_1038,In_1866);
or U711 (N_711,In_38,In_1948);
or U712 (N_712,In_1250,In_580);
or U713 (N_713,In_471,In_473);
or U714 (N_714,In_570,In_1132);
and U715 (N_715,In_1080,In_929);
nand U716 (N_716,In_1627,In_603);
or U717 (N_717,In_1575,In_434);
xor U718 (N_718,In_631,In_985);
xnor U719 (N_719,In_1164,In_1892);
xnor U720 (N_720,In_203,In_1545);
and U721 (N_721,In_164,In_909);
or U722 (N_722,In_918,In_1422);
xor U723 (N_723,In_392,In_413);
xor U724 (N_724,In_1454,In_1757);
nand U725 (N_725,In_1307,In_1282);
xnor U726 (N_726,In_530,In_1450);
nor U727 (N_727,In_1300,In_152);
xor U728 (N_728,In_1791,In_486);
nand U729 (N_729,In_1418,In_1353);
and U730 (N_730,In_1114,In_1027);
nand U731 (N_731,In_289,In_1559);
and U732 (N_732,In_567,In_1190);
nand U733 (N_733,In_1461,In_739);
nand U734 (N_734,In_976,In_629);
nor U735 (N_735,In_1323,In_1678);
or U736 (N_736,In_1785,In_910);
nor U737 (N_737,In_655,In_317);
nand U738 (N_738,In_313,In_1477);
nor U739 (N_739,In_238,In_649);
xnor U740 (N_740,In_83,In_1290);
and U741 (N_741,In_1402,In_157);
nand U742 (N_742,In_1766,In_1951);
or U743 (N_743,In_1122,In_62);
nor U744 (N_744,In_721,In_1940);
xnor U745 (N_745,In_1808,In_1844);
nand U746 (N_746,In_1071,In_1613);
nor U747 (N_747,In_394,In_1012);
and U748 (N_748,In_690,In_956);
or U749 (N_749,In_1874,In_619);
nor U750 (N_750,In_667,In_958);
and U751 (N_751,In_1337,In_788);
nand U752 (N_752,In_1762,In_1612);
nor U753 (N_753,In_376,In_867);
xor U754 (N_754,In_294,In_892);
xnor U755 (N_755,In_1210,In_723);
nand U756 (N_756,In_515,In_138);
xnor U757 (N_757,In_893,In_597);
and U758 (N_758,In_1697,In_1855);
and U759 (N_759,In_1095,In_697);
or U760 (N_760,In_465,In_176);
and U761 (N_761,In_1780,In_1134);
and U762 (N_762,In_269,In_300);
nand U763 (N_763,In_124,In_1474);
and U764 (N_764,In_1416,In_316);
nor U765 (N_765,In_827,In_236);
and U766 (N_766,In_587,In_1433);
nor U767 (N_767,In_135,In_674);
nand U768 (N_768,In_1869,In_280);
or U769 (N_769,In_1032,In_292);
or U770 (N_770,In_1145,In_1630);
nor U771 (N_771,In_1025,In_1175);
nor U772 (N_772,In_1729,In_445);
or U773 (N_773,In_172,In_837);
nand U774 (N_774,In_440,In_1513);
nand U775 (N_775,In_211,In_444);
and U776 (N_776,In_1239,In_424);
xnor U777 (N_777,In_1343,In_1298);
or U778 (N_778,In_78,In_766);
nor U779 (N_779,In_584,In_56);
xnor U780 (N_780,In_93,In_181);
xor U781 (N_781,In_1413,In_1188);
or U782 (N_782,In_1314,In_559);
nand U783 (N_783,In_560,In_1565);
nand U784 (N_784,In_1739,In_1206);
nand U785 (N_785,In_1085,In_880);
and U786 (N_786,In_177,In_1508);
and U787 (N_787,In_1083,In_574);
xnor U788 (N_788,In_1665,In_941);
and U789 (N_789,In_1699,In_1245);
nand U790 (N_790,In_982,In_742);
nor U791 (N_791,In_997,In_1819);
and U792 (N_792,In_627,In_226);
nor U793 (N_793,In_1346,In_1303);
xnor U794 (N_794,In_963,In_476);
xnor U795 (N_795,In_1619,In_1945);
nand U796 (N_796,In_1722,In_1755);
or U797 (N_797,In_881,In_1543);
xnor U798 (N_798,In_1502,In_1707);
or U799 (N_799,In_132,In_430);
nor U800 (N_800,In_219,N_61);
xnor U801 (N_801,In_1908,In_1593);
or U802 (N_802,In_1544,N_553);
nand U803 (N_803,N_177,N_459);
nand U804 (N_804,N_533,N_276);
nor U805 (N_805,N_55,N_636);
and U806 (N_806,In_16,N_356);
nand U807 (N_807,N_510,N_769);
or U808 (N_808,In_140,N_236);
or U809 (N_809,In_144,In_1299);
xor U810 (N_810,N_669,N_639);
or U811 (N_811,In_642,N_255);
nand U812 (N_812,N_511,N_580);
or U813 (N_813,N_495,N_419);
xnor U814 (N_814,N_451,N_296);
nand U815 (N_815,N_171,N_300);
xor U816 (N_816,In_1774,N_583);
xnor U817 (N_817,N_575,N_563);
xnor U818 (N_818,N_329,N_7);
nor U819 (N_819,N_487,In_1998);
xnor U820 (N_820,N_269,N_114);
xor U821 (N_821,In_19,N_378);
xor U822 (N_822,In_590,N_702);
and U823 (N_823,N_469,N_656);
xor U824 (N_824,In_1898,In_1365);
xnor U825 (N_825,N_632,N_134);
and U826 (N_826,N_363,N_111);
nor U827 (N_827,N_120,In_1986);
nor U828 (N_828,In_327,In_1156);
nor U829 (N_829,In_1463,N_783);
and U830 (N_830,N_497,N_233);
nor U831 (N_831,N_388,N_226);
nor U832 (N_832,In_1853,N_274);
nand U833 (N_833,N_251,N_499);
nor U834 (N_834,N_607,N_650);
nor U835 (N_835,In_1822,N_578);
nand U836 (N_836,N_242,In_1481);
nand U837 (N_837,N_481,In_239);
and U838 (N_838,N_605,In_1514);
or U839 (N_839,N_308,N_721);
and U840 (N_840,In_451,N_453);
or U841 (N_841,N_198,N_347);
and U842 (N_842,N_180,In_1773);
or U843 (N_843,N_209,N_513);
nand U844 (N_844,In_248,N_392);
nand U845 (N_845,N_734,N_93);
xor U846 (N_846,In_897,N_596);
xor U847 (N_847,N_743,N_369);
and U848 (N_848,N_410,In_1596);
nand U849 (N_849,In_789,N_514);
nand U850 (N_850,In_1971,N_763);
nand U851 (N_851,N_711,N_586);
or U852 (N_852,In_1165,In_1395);
nor U853 (N_853,N_413,N_643);
nand U854 (N_854,N_624,N_132);
and U855 (N_855,N_475,N_28);
or U856 (N_856,N_485,In_760);
nand U857 (N_857,In_1448,In_750);
nor U858 (N_858,N_727,N_291);
nor U859 (N_859,N_434,N_465);
nand U860 (N_860,In_360,N_62);
xnor U861 (N_861,N_165,In_1557);
and U862 (N_862,N_110,In_134);
nor U863 (N_863,N_65,In_1870);
nor U864 (N_864,In_399,N_672);
nor U865 (N_865,N_256,N_447);
xnor U866 (N_866,N_57,N_278);
nor U867 (N_867,In_1718,N_33);
xnor U868 (N_868,N_701,In_523);
nand U869 (N_869,N_740,N_133);
xor U870 (N_870,N_557,N_741);
and U871 (N_871,N_364,N_208);
xor U872 (N_872,N_381,In_1195);
nand U873 (N_873,N_75,In_491);
xnor U874 (N_874,N_194,In_1649);
nor U875 (N_875,In_1148,In_1233);
or U876 (N_876,N_602,In_1827);
nor U877 (N_877,N_644,N_446);
nor U878 (N_878,In_479,N_397);
nor U879 (N_879,N_353,N_265);
and U880 (N_880,N_753,In_846);
nand U881 (N_881,In_522,In_1922);
and U882 (N_882,N_655,N_630);
and U883 (N_883,In_1668,N_642);
nand U884 (N_884,N_338,N_423);
nand U885 (N_885,N_22,In_1486);
nand U886 (N_886,In_347,N_393);
or U887 (N_887,N_791,N_773);
and U888 (N_888,In_724,In_41);
nand U889 (N_889,N_216,In_1331);
nor U890 (N_890,In_1556,In_964);
nand U891 (N_891,N_319,In_1363);
xor U892 (N_892,In_496,N_516);
and U893 (N_893,In_800,N_51);
nor U894 (N_894,In_466,N_123);
and U895 (N_895,N_606,N_472);
nand U896 (N_896,In_1259,N_354);
xnor U897 (N_897,N_215,In_913);
or U898 (N_898,N_433,In_1981);
and U899 (N_899,In_950,In_1505);
nor U900 (N_900,N_100,N_509);
or U901 (N_901,N_9,N_41);
and U902 (N_902,In_28,In_1930);
nand U903 (N_903,In_356,N_26);
or U904 (N_904,N_710,N_95);
and U905 (N_905,In_840,N_82);
nor U906 (N_906,N_762,N_418);
xor U907 (N_907,In_477,N_635);
nand U908 (N_908,In_520,In_242);
xor U909 (N_909,In_974,N_685);
and U910 (N_910,N_136,N_613);
nor U911 (N_911,N_435,N_657);
or U912 (N_912,N_12,N_705);
nor U913 (N_913,In_488,N_298);
xor U914 (N_914,N_337,N_684);
nand U915 (N_915,N_105,In_1867);
nor U916 (N_916,N_213,N_6);
and U917 (N_917,In_673,In_1485);
and U918 (N_918,N_548,N_148);
nor U919 (N_919,N_534,N_574);
or U920 (N_920,In_1842,N_653);
xor U921 (N_921,In_882,N_76);
nor U922 (N_922,N_107,N_524);
xnor U923 (N_923,In_1435,In_536);
nand U924 (N_924,In_646,N_460);
nand U925 (N_925,N_48,N_135);
nand U926 (N_926,N_567,N_144);
and U927 (N_927,N_204,N_34);
nor U928 (N_928,N_312,N_473);
nor U929 (N_929,In_459,N_390);
xor U930 (N_930,N_336,N_234);
or U931 (N_931,N_203,N_252);
nor U932 (N_932,N_221,N_678);
xor U933 (N_933,In_154,In_365);
nand U934 (N_934,N_340,In_1265);
nor U935 (N_935,In_979,N_550);
xor U936 (N_936,N_253,In_823);
and U937 (N_937,In_1888,In_1567);
or U938 (N_938,N_326,N_81);
and U939 (N_939,N_170,In_962);
or U940 (N_940,N_305,N_106);
xnor U941 (N_941,N_408,N_191);
and U942 (N_942,N_539,N_502);
or U943 (N_943,N_192,N_745);
or U944 (N_944,N_162,In_936);
or U945 (N_945,In_1626,N_748);
and U946 (N_946,N_240,N_661);
or U947 (N_947,In_1562,In_469);
nor U948 (N_948,N_610,N_155);
xor U949 (N_949,In_1743,In_1244);
or U950 (N_950,In_767,In_705);
xnor U951 (N_951,In_541,N_301);
xor U952 (N_952,N_324,N_659);
nor U953 (N_953,N_531,N_31);
xor U954 (N_954,N_152,In_1455);
or U955 (N_955,N_56,N_641);
nand U956 (N_956,N_579,N_130);
or U957 (N_957,N_621,N_102);
nor U958 (N_958,N_652,N_488);
nand U959 (N_959,In_17,In_707);
nor U960 (N_960,N_778,N_789);
nor U961 (N_961,In_1667,N_193);
nand U962 (N_962,In_1829,In_546);
xnor U963 (N_963,N_577,N_629);
nand U964 (N_964,N_19,N_492);
and U965 (N_965,N_71,In_1526);
nand U966 (N_966,N_692,In_404);
and U967 (N_967,In_1796,N_98);
nand U968 (N_968,N_645,N_235);
or U969 (N_969,N_501,N_355);
xnor U970 (N_970,In_1099,N_493);
and U971 (N_971,In_525,In_785);
nand U972 (N_972,In_1334,N_309);
and U973 (N_973,N_179,N_250);
xnor U974 (N_974,N_673,N_259);
nor U975 (N_975,In_297,N_341);
nor U976 (N_976,N_608,In_31);
nor U977 (N_977,N_68,N_582);
and U978 (N_978,N_272,In_1361);
nand U979 (N_979,N_168,N_145);
or U980 (N_980,N_658,N_63);
or U981 (N_981,N_747,N_156);
or U982 (N_982,N_342,N_345);
nand U983 (N_983,N_619,N_112);
and U984 (N_984,N_182,In_145);
and U985 (N_985,N_744,In_319);
nor U986 (N_986,N_751,In_1015);
nand U987 (N_987,N_99,N_505);
nand U988 (N_988,In_1620,In_302);
and U989 (N_989,N_87,In_1403);
nand U990 (N_990,In_122,N_104);
xnor U991 (N_991,In_1551,N_461);
or U992 (N_992,N_671,In_298);
xor U993 (N_993,In_13,N_551);
and U994 (N_994,N_750,In_1538);
or U995 (N_995,N_448,In_630);
xor U996 (N_996,N_527,N_88);
nor U997 (N_997,N_799,N_716);
or U998 (N_998,In_926,In_218);
nor U999 (N_999,In_978,N_691);
or U1000 (N_1000,In_1931,N_64);
nor U1001 (N_1001,N_626,N_58);
xnor U1002 (N_1002,N_163,In_1776);
xnor U1003 (N_1003,N_396,N_480);
nor U1004 (N_1004,N_199,In_945);
xor U1005 (N_1005,In_1381,N_764);
or U1006 (N_1006,N_176,In_107);
and U1007 (N_1007,N_260,N_289);
xnor U1008 (N_1008,N_483,N_697);
nand U1009 (N_1009,In_229,N_777);
nand U1010 (N_1010,In_755,N_84);
nor U1011 (N_1011,N_742,In_1369);
nor U1012 (N_1012,In_1003,N_520);
and U1013 (N_1013,N_212,N_733);
nand U1014 (N_1014,N_737,N_739);
nand U1015 (N_1015,N_592,In_555);
xnor U1016 (N_1016,N_189,In_1532);
nand U1017 (N_1017,N_384,N_471);
nand U1018 (N_1018,In_358,N_128);
nor U1019 (N_1019,N_703,N_795);
nor U1020 (N_1020,N_681,N_792);
nor U1021 (N_1021,N_454,N_439);
nor U1022 (N_1022,N_407,N_591);
xor U1023 (N_1023,N_699,In_1173);
nand U1024 (N_1024,In_1144,In_1183);
and U1025 (N_1025,In_467,N_333);
and U1026 (N_1026,N_108,N_297);
and U1027 (N_1027,N_774,In_485);
nor U1028 (N_1028,N_167,N_314);
or U1029 (N_1029,N_562,N_726);
nand U1030 (N_1030,N_264,N_504);
and U1031 (N_1031,N_776,In_1005);
xor U1032 (N_1032,N_515,N_50);
xor U1033 (N_1033,In_1452,N_521);
nor U1034 (N_1034,In_511,N_444);
nand U1035 (N_1035,In_37,In_902);
nor U1036 (N_1036,N_157,N_649);
nand U1037 (N_1037,In_1711,N_695);
nor U1038 (N_1038,N_129,N_536);
or U1039 (N_1039,N_13,N_282);
xor U1040 (N_1040,N_437,In_295);
nor U1041 (N_1041,N_175,N_103);
or U1042 (N_1042,N_543,N_540);
xor U1043 (N_1043,N_187,N_121);
nand U1044 (N_1044,In_547,In_159);
nor U1045 (N_1045,In_1850,In_1367);
nor U1046 (N_1046,N_637,N_782);
and U1047 (N_1047,N_67,In_583);
or U1048 (N_1048,In_1959,In_406);
and U1049 (N_1049,N_59,N_292);
nand U1050 (N_1050,N_37,N_218);
and U1051 (N_1051,N_8,N_498);
or U1052 (N_1052,In_715,In_234);
nand U1053 (N_1053,In_1835,In_472);
xnor U1054 (N_1054,In_310,In_470);
nand U1055 (N_1055,N_183,In_209);
and U1056 (N_1056,N_52,N_15);
nand U1057 (N_1057,N_542,N_394);
or U1058 (N_1058,N_478,N_738);
and U1059 (N_1059,N_595,N_125);
xnor U1060 (N_1060,N_609,In_1101);
xor U1061 (N_1061,N_224,In_1608);
xor U1062 (N_1062,In_569,N_771);
or U1063 (N_1063,N_768,In_704);
nand U1064 (N_1064,N_210,N_670);
or U1065 (N_1065,N_549,In_802);
and U1066 (N_1066,N_688,In_1881);
nand U1067 (N_1067,N_523,In_685);
or U1068 (N_1068,N_528,N_307);
xnor U1069 (N_1069,N_316,N_646);
and U1070 (N_1070,N_713,N_36);
and U1071 (N_1071,In_869,N_766);
xor U1072 (N_1072,N_66,In_911);
and U1073 (N_1073,N_164,N_529);
xor U1074 (N_1074,N_441,In_1677);
nand U1075 (N_1075,N_47,N_590);
xnor U1076 (N_1076,In_1351,N_558);
nand U1077 (N_1077,N_794,N_522);
xor U1078 (N_1078,N_53,In_1506);
xor U1079 (N_1079,N_414,In_566);
nor U1080 (N_1080,N_442,N_458);
nand U1081 (N_1081,N_266,N_587);
or U1082 (N_1082,N_761,N_466);
or U1083 (N_1083,N_137,N_91);
xor U1084 (N_1084,N_584,N_44);
nor U1085 (N_1085,In_1782,In_1825);
or U1086 (N_1086,In_231,In_257);
or U1087 (N_1087,In_1443,In_1975);
nor U1088 (N_1088,N_572,In_558);
or U1089 (N_1089,N_395,In_1357);
nand U1090 (N_1090,N_11,N_445);
nand U1091 (N_1091,N_438,N_677);
and U1092 (N_1092,N_246,In_115);
nor U1093 (N_1093,N_785,In_1021);
and U1094 (N_1094,In_1569,In_1727);
nor U1095 (N_1095,N_385,N_334);
and U1096 (N_1096,N_555,N_479);
or U1097 (N_1097,N_376,In_1339);
nor U1098 (N_1098,N_554,N_20);
or U1099 (N_1099,N_491,N_545);
or U1100 (N_1100,N_718,N_667);
and U1101 (N_1101,N_638,N_616);
or U1102 (N_1102,In_391,N_331);
xor U1103 (N_1103,N_757,In_786);
xor U1104 (N_1104,In_1591,In_267);
nand U1105 (N_1105,N_359,In_806);
and U1106 (N_1106,In_1118,In_3);
xor U1107 (N_1107,In_1533,N_796);
or U1108 (N_1108,In_585,N_32);
nand U1109 (N_1109,N_477,N_365);
nor U1110 (N_1110,N_589,N_325);
nand U1111 (N_1111,N_14,N_474);
and U1112 (N_1112,N_0,N_627);
and U1113 (N_1113,In_1735,In_898);
nand U1114 (N_1114,N_16,N_689);
nor U1115 (N_1115,N_343,N_714);
xor U1116 (N_1116,N_512,In_764);
nand U1117 (N_1117,In_934,N_780);
nand U1118 (N_1118,In_671,N_27);
nand U1119 (N_1119,N_564,N_676);
xnor U1120 (N_1120,N_77,N_350);
and U1121 (N_1121,N_273,In_1987);
xnor U1122 (N_1122,N_420,N_230);
nor U1123 (N_1123,N_223,N_346);
or U1124 (N_1124,N_1,In_389);
and U1125 (N_1125,In_169,In_1091);
and U1126 (N_1126,N_141,In_1905);
nor U1127 (N_1127,N_313,N_784);
or U1128 (N_1128,In_156,In_168);
and U1129 (N_1129,N_722,N_717);
nor U1130 (N_1130,N_581,N_793);
nand U1131 (N_1131,N_648,In_828);
or U1132 (N_1132,N_220,In_163);
nand U1133 (N_1133,In_1147,In_439);
nor U1134 (N_1134,In_1384,N_380);
and U1135 (N_1135,In_1475,N_374);
xnor U1136 (N_1136,In_1336,In_1069);
nor U1137 (N_1137,N_389,In_1561);
xor U1138 (N_1138,N_267,In_158);
and U1139 (N_1139,N_109,N_241);
and U1140 (N_1140,In_1362,In_701);
or U1141 (N_1141,N_544,N_754);
nand U1142 (N_1142,N_70,N_94);
nor U1143 (N_1143,N_304,In_1830);
nor U1144 (N_1144,N_150,In_1068);
and U1145 (N_1145,N_731,In_1372);
nand U1146 (N_1146,N_43,In_286);
or U1147 (N_1147,N_686,In_39);
xnor U1148 (N_1148,N_86,N_594);
and U1149 (N_1149,In_1634,N_622);
xor U1150 (N_1150,In_1301,In_1460);
nand U1151 (N_1151,In_595,In_986);
and U1152 (N_1152,N_406,In_1654);
xor U1153 (N_1153,In_1994,N_706);
or U1154 (N_1154,In_1690,N_690);
nor U1155 (N_1155,N_225,N_604);
and U1156 (N_1156,N_143,In_112);
nand U1157 (N_1157,N_640,N_614);
and U1158 (N_1158,N_724,In_1100);
nor U1159 (N_1159,N_732,N_665);
nor U1160 (N_1160,N_500,N_138);
xor U1161 (N_1161,In_12,N_526);
and U1162 (N_1162,N_623,N_618);
or U1163 (N_1163,N_736,In_850);
xor U1164 (N_1164,N_517,N_405);
nor U1165 (N_1165,N_118,N_593);
or U1166 (N_1166,In_489,N_401);
xor U1167 (N_1167,In_1602,In_1312);
and U1168 (N_1168,N_700,In_1894);
xor U1169 (N_1169,N_21,In_1120);
or U1170 (N_1170,N_42,In_648);
or U1171 (N_1171,N_239,N_696);
and U1172 (N_1172,In_291,In_1022);
nand U1173 (N_1173,N_597,N_456);
and U1174 (N_1174,In_1897,N_715);
and U1175 (N_1175,N_74,N_787);
nand U1176 (N_1176,N_29,N_426);
nand U1177 (N_1177,N_541,N_535);
nor U1178 (N_1178,N_537,In_660);
xor U1179 (N_1179,N_262,N_603);
and U1180 (N_1180,N_547,N_270);
nor U1181 (N_1181,N_470,N_320);
or U1182 (N_1182,N_482,N_197);
and U1183 (N_1183,In_720,N_119);
xnor U1184 (N_1184,In_1936,In_939);
or U1185 (N_1185,N_588,N_770);
nor U1186 (N_1186,In_1490,N_503);
and U1187 (N_1187,In_1342,N_755);
nand U1188 (N_1188,N_161,In_726);
and U1189 (N_1189,N_299,N_403);
nor U1190 (N_1190,N_360,N_39);
nand U1191 (N_1191,In_275,N_80);
nand U1192 (N_1192,N_200,N_45);
or U1193 (N_1193,In_320,N_790);
and U1194 (N_1194,N_723,N_600);
nand U1195 (N_1195,In_594,In_1400);
and U1196 (N_1196,N_559,N_315);
nor U1197 (N_1197,N_666,N_371);
nor U1198 (N_1198,In_182,In_1982);
nor U1199 (N_1199,N_525,N_78);
nor U1200 (N_1200,In_382,N_687);
and U1201 (N_1201,N_238,In_1954);
or U1202 (N_1202,N_344,N_449);
nor U1203 (N_1203,In_1404,N_358);
or U1204 (N_1204,N_463,N_280);
or U1205 (N_1205,In_1011,N_49);
and U1206 (N_1206,N_424,In_1489);
or U1207 (N_1207,N_569,N_281);
xor U1208 (N_1208,N_391,In_1494);
and U1209 (N_1209,N_383,N_683);
or U1210 (N_1210,N_54,N_131);
and U1211 (N_1211,In_1607,N_124);
nor U1212 (N_1212,N_96,N_576);
or U1213 (N_1213,In_1845,N_760);
nor U1214 (N_1214,In_104,In_1328);
xnor U1215 (N_1215,N_489,N_427);
nor U1216 (N_1216,N_279,In_161);
nor U1217 (N_1217,In_1273,In_863);
nor U1218 (N_1218,In_1050,In_1390);
or U1219 (N_1219,N_370,N_249);
or U1220 (N_1220,In_855,In_1434);
nor U1221 (N_1221,In_927,N_615);
nand U1222 (N_1222,N_275,In_809);
or U1223 (N_1223,N_709,N_663);
and U1224 (N_1224,In_417,In_213);
nand U1225 (N_1225,N_178,In_680);
or U1226 (N_1226,N_286,N_24);
nand U1227 (N_1227,N_283,N_462);
xnor U1228 (N_1228,In_967,In_262);
and U1229 (N_1229,N_417,In_586);
nand U1230 (N_1230,N_366,In_1896);
and U1231 (N_1231,N_92,In_1708);
and U1232 (N_1232,In_531,In_873);
and U1233 (N_1233,N_486,In_1686);
xor U1234 (N_1234,N_631,In_53);
or U1235 (N_1235,In_1430,N_18);
or U1236 (N_1236,In_1806,N_506);
nand U1237 (N_1237,N_440,In_643);
nor U1238 (N_1238,N_101,N_664);
nand U1239 (N_1239,N_348,N_323);
or U1240 (N_1240,N_402,N_127);
nand U1241 (N_1241,In_727,N_339);
nand U1242 (N_1242,In_1213,N_415);
xor U1243 (N_1243,N_328,N_349);
nor U1244 (N_1244,In_534,In_1730);
xnor U1245 (N_1245,In_1588,N_159);
nor U1246 (N_1246,N_202,N_507);
nand U1247 (N_1247,N_254,N_411);
nand U1248 (N_1248,N_248,In_516);
or U1249 (N_1249,N_83,N_496);
nor U1250 (N_1250,N_377,N_647);
nand U1251 (N_1251,N_172,N_321);
and U1252 (N_1252,N_277,N_196);
xnor U1253 (N_1253,N_431,N_295);
or U1254 (N_1254,In_1318,N_571);
nor U1255 (N_1255,In_251,N_229);
and U1256 (N_1256,N_25,N_772);
and U1257 (N_1257,N_244,N_2);
nor U1258 (N_1258,N_530,In_1600);
and U1259 (N_1259,N_169,N_399);
nor U1260 (N_1260,N_245,N_546);
or U1261 (N_1261,N_651,N_432);
xor U1262 (N_1262,N_708,N_720);
nor U1263 (N_1263,N_60,N_35);
xnor U1264 (N_1264,In_265,N_97);
xor U1265 (N_1265,In_854,N_668);
nor U1266 (N_1266,N_115,In_1581);
nor U1267 (N_1267,In_1039,N_153);
and U1268 (N_1268,In_1377,N_729);
xor U1269 (N_1269,N_38,N_758);
and U1270 (N_1270,N_147,N_552);
nor U1271 (N_1271,N_146,In_1456);
or U1272 (N_1272,N_628,N_494);
nor U1273 (N_1273,In_620,N_294);
and U1274 (N_1274,N_285,In_1310);
or U1275 (N_1275,N_306,In_888);
and U1276 (N_1276,N_181,N_452);
and U1277 (N_1277,In_839,N_756);
or U1278 (N_1278,In_741,N_330);
and U1279 (N_1279,N_425,N_69);
or U1280 (N_1280,N_404,In_1499);
xor U1281 (N_1281,N_214,N_719);
nor U1282 (N_1282,N_620,In_273);
xnor U1283 (N_1283,N_232,N_436);
xnor U1284 (N_1284,In_1417,In_1466);
nor U1285 (N_1285,N_160,N_186);
or U1286 (N_1286,N_601,N_476);
nand U1287 (N_1287,N_263,In_223);
nor U1288 (N_1288,N_565,N_211);
or U1289 (N_1289,N_154,N_362);
or U1290 (N_1290,N_767,N_288);
xnor U1291 (N_1291,In_1136,In_1035);
nand U1292 (N_1292,In_390,N_386);
xor U1293 (N_1293,N_268,In_274);
and U1294 (N_1294,In_429,In_623);
nor U1295 (N_1295,N_367,In_1997);
nand U1296 (N_1296,N_598,N_429);
nor U1297 (N_1297,N_142,N_318);
or U1298 (N_1298,N_287,In_1555);
xor U1299 (N_1299,N_634,In_315);
nand U1300 (N_1300,N_368,In_1857);
xnor U1301 (N_1301,N_728,In_126);
or U1302 (N_1302,N_217,In_955);
nand U1303 (N_1303,N_400,N_725);
nor U1304 (N_1304,In_1546,N_430);
nand U1305 (N_1305,N_361,N_679);
xor U1306 (N_1306,N_46,N_560);
or U1307 (N_1307,N_219,N_566);
nand U1308 (N_1308,In_1666,In_805);
xor U1309 (N_1309,N_40,N_662);
and U1310 (N_1310,In_912,N_335);
xnor U1311 (N_1311,In_1747,N_205);
or U1312 (N_1312,N_257,In_1053);
and U1313 (N_1313,In_836,In_1944);
nand U1314 (N_1314,N_188,N_151);
xnor U1315 (N_1315,N_693,In_386);
and U1316 (N_1316,N_654,N_247);
nor U1317 (N_1317,In_1996,In_1235);
or U1318 (N_1318,In_428,N_332);
or U1319 (N_1319,In_442,N_674);
nand U1320 (N_1320,N_311,N_781);
or U1321 (N_1321,N_310,N_798);
nor U1322 (N_1322,In_359,N_352);
nor U1323 (N_1323,N_290,In_1229);
and U1324 (N_1324,N_422,N_765);
and U1325 (N_1325,N_682,In_563);
and U1326 (N_1326,N_538,N_207);
or U1327 (N_1327,N_749,In_1074);
nor U1328 (N_1328,N_222,In_688);
nor U1329 (N_1329,In_1276,N_284);
or U1330 (N_1330,N_228,N_468);
nand U1331 (N_1331,N_625,N_735);
nor U1332 (N_1332,In_554,N_79);
nor U1333 (N_1333,N_149,N_3);
nor U1334 (N_1334,N_113,N_633);
or U1335 (N_1335,N_302,N_660);
and U1336 (N_1336,N_140,In_1412);
nor U1337 (N_1337,N_611,N_759);
nand U1338 (N_1338,In_652,In_1765);
nor U1339 (N_1339,N_443,N_357);
xnor U1340 (N_1340,N_30,N_126);
xnor U1341 (N_1341,N_195,N_190);
nand U1342 (N_1342,N_293,N_680);
nor U1343 (N_1343,N_85,N_490);
and U1344 (N_1344,N_158,N_243);
and U1345 (N_1345,N_237,In_616);
nand U1346 (N_1346,N_704,N_416);
xnor U1347 (N_1347,In_617,In_147);
and U1348 (N_1348,In_743,N_327);
nand U1349 (N_1349,N_375,N_409);
and U1350 (N_1350,N_464,In_96);
nor U1351 (N_1351,In_191,N_518);
xor U1352 (N_1352,In_1680,In_1675);
and U1353 (N_1353,N_261,In_1861);
nand U1354 (N_1354,In_1029,In_650);
and U1355 (N_1355,N_752,N_570);
or U1356 (N_1356,N_707,In_1760);
nor U1357 (N_1357,N_174,N_317);
or U1358 (N_1358,N_698,In_71);
or U1359 (N_1359,N_184,N_116);
xnor U1360 (N_1360,In_243,In_403);
nor U1361 (N_1361,N_484,In_185);
nand U1362 (N_1362,In_668,N_617);
and U1363 (N_1363,N_122,N_258);
nor U1364 (N_1364,In_605,N_746);
nor U1365 (N_1365,N_227,N_421);
nand U1366 (N_1366,N_712,N_387);
or U1367 (N_1367,N_797,N_322);
or U1368 (N_1368,In_1327,N_508);
xor U1369 (N_1369,N_457,N_519);
or U1370 (N_1370,N_382,N_450);
and U1371 (N_1371,In_1570,N_23);
nor U1372 (N_1372,N_73,N_532);
nor U1373 (N_1373,N_166,N_694);
nor U1374 (N_1374,N_788,N_373);
and U1375 (N_1375,N_10,N_231);
and U1376 (N_1376,N_599,N_303);
xor U1377 (N_1377,In_1189,In_621);
nand U1378 (N_1378,N_612,In_1962);
xor U1379 (N_1379,N_775,N_201);
nor U1380 (N_1380,In_1442,In_339);
and U1381 (N_1381,N_467,N_398);
nor U1382 (N_1382,N_173,N_455);
nor U1383 (N_1383,In_1285,In_734);
or U1384 (N_1384,In_527,N_786);
and U1385 (N_1385,In_109,N_139);
nor U1386 (N_1386,N_730,N_561);
xnor U1387 (N_1387,N_90,N_271);
xnor U1388 (N_1388,N_89,N_568);
xor U1389 (N_1389,N_675,In_611);
nor U1390 (N_1390,In_105,N_556);
or U1391 (N_1391,N_372,N_117);
or U1392 (N_1392,N_17,N_185);
or U1393 (N_1393,In_1241,N_428);
xnor U1394 (N_1394,N_779,In_342);
nor U1395 (N_1395,N_5,N_206);
nand U1396 (N_1396,N_412,N_4);
xnor U1397 (N_1397,N_351,N_573);
xnor U1398 (N_1398,N_585,In_1391);
nand U1399 (N_1399,N_72,N_379);
nand U1400 (N_1400,N_132,N_482);
nand U1401 (N_1401,In_840,N_477);
nand U1402 (N_1402,N_40,N_387);
and U1403 (N_1403,N_639,In_1351);
nand U1404 (N_1404,In_1053,N_251);
xor U1405 (N_1405,N_495,N_197);
nand U1406 (N_1406,N_75,In_1430);
or U1407 (N_1407,N_607,N_683);
nand U1408 (N_1408,N_772,N_528);
and U1409 (N_1409,In_12,N_434);
xnor U1410 (N_1410,In_404,N_291);
or U1411 (N_1411,N_604,N_657);
nand U1412 (N_1412,N_760,N_431);
xnor U1413 (N_1413,N_0,In_248);
xor U1414 (N_1414,N_589,N_330);
nor U1415 (N_1415,In_1362,N_11);
nand U1416 (N_1416,N_15,N_225);
and U1417 (N_1417,In_1463,In_1506);
nand U1418 (N_1418,N_645,N_635);
and U1419 (N_1419,N_743,N_628);
nor U1420 (N_1420,In_967,In_213);
nand U1421 (N_1421,In_267,N_578);
and U1422 (N_1422,N_376,In_566);
nor U1423 (N_1423,N_362,N_51);
nor U1424 (N_1424,N_552,In_182);
nand U1425 (N_1425,In_472,In_1556);
and U1426 (N_1426,N_679,N_513);
nor U1427 (N_1427,N_285,N_204);
and U1428 (N_1428,N_192,In_964);
or U1429 (N_1429,N_208,In_1936);
nand U1430 (N_1430,In_1494,N_629);
and U1431 (N_1431,N_558,N_287);
xor U1432 (N_1432,N_140,In_525);
or U1433 (N_1433,N_440,In_275);
nand U1434 (N_1434,In_1069,N_672);
or U1435 (N_1435,In_1675,In_273);
and U1436 (N_1436,N_174,N_764);
nor U1437 (N_1437,In_1005,In_764);
and U1438 (N_1438,In_417,N_321);
or U1439 (N_1439,In_660,N_339);
or U1440 (N_1440,N_34,N_17);
xnor U1441 (N_1441,In_1342,N_692);
nor U1442 (N_1442,N_264,In_1514);
and U1443 (N_1443,In_764,In_1551);
xnor U1444 (N_1444,In_1499,N_597);
nor U1445 (N_1445,N_594,N_40);
and U1446 (N_1446,In_1189,N_699);
xor U1447 (N_1447,In_1003,N_417);
or U1448 (N_1448,N_409,In_1372);
or U1449 (N_1449,N_681,N_509);
nand U1450 (N_1450,N_94,N_594);
nor U1451 (N_1451,N_395,N_621);
or U1452 (N_1452,N_63,N_256);
xnor U1453 (N_1453,N_90,N_423);
nor U1454 (N_1454,N_283,N_672);
and U1455 (N_1455,N_100,N_614);
and U1456 (N_1456,In_1466,In_1339);
nor U1457 (N_1457,N_234,N_471);
or U1458 (N_1458,N_669,N_1);
nand U1459 (N_1459,N_71,N_457);
xor U1460 (N_1460,In_646,N_243);
and U1461 (N_1461,In_1100,N_28);
and U1462 (N_1462,N_430,In_1365);
nand U1463 (N_1463,N_544,N_527);
or U1464 (N_1464,N_540,N_607);
nor U1465 (N_1465,N_371,In_1100);
and U1466 (N_1466,N_740,In_262);
nor U1467 (N_1467,N_535,N_496);
nand U1468 (N_1468,N_51,In_1861);
and U1469 (N_1469,N_759,N_113);
nor U1470 (N_1470,N_745,N_121);
xor U1471 (N_1471,N_270,N_308);
nor U1472 (N_1472,N_483,N_510);
and U1473 (N_1473,N_687,N_160);
nand U1474 (N_1474,N_277,N_565);
nand U1475 (N_1475,N_799,N_377);
or U1476 (N_1476,N_473,N_652);
xor U1477 (N_1477,N_273,In_1975);
nand U1478 (N_1478,N_474,N_388);
nor U1479 (N_1479,In_755,N_786);
nand U1480 (N_1480,In_1822,N_310);
or U1481 (N_1481,N_792,N_10);
nor U1482 (N_1482,N_236,N_478);
and U1483 (N_1483,N_8,N_331);
nand U1484 (N_1484,N_765,In_1773);
xor U1485 (N_1485,N_211,N_91);
nor U1486 (N_1486,N_293,In_704);
nor U1487 (N_1487,N_597,N_96);
nor U1488 (N_1488,In_522,N_789);
nor U1489 (N_1489,N_652,N_141);
nand U1490 (N_1490,In_1654,In_109);
xor U1491 (N_1491,N_328,In_16);
xnor U1492 (N_1492,N_303,In_1555);
or U1493 (N_1493,In_1339,N_229);
and U1494 (N_1494,In_643,N_158);
and U1495 (N_1495,N_710,N_737);
xnor U1496 (N_1496,N_641,In_365);
nor U1497 (N_1497,N_744,N_8);
xor U1498 (N_1498,N_183,N_706);
nand U1499 (N_1499,N_421,In_630);
xnor U1500 (N_1500,N_551,N_188);
xnor U1501 (N_1501,In_869,N_17);
xnor U1502 (N_1502,N_628,In_1600);
xnor U1503 (N_1503,N_479,In_275);
and U1504 (N_1504,In_158,N_746);
and U1505 (N_1505,N_442,N_552);
nand U1506 (N_1506,In_1546,N_632);
nor U1507 (N_1507,In_707,N_94);
xnor U1508 (N_1508,N_50,In_660);
nand U1509 (N_1509,N_728,In_327);
nor U1510 (N_1510,N_562,N_515);
and U1511 (N_1511,N_30,N_280);
and U1512 (N_1512,N_759,N_70);
and U1513 (N_1513,N_744,N_631);
xor U1514 (N_1514,N_434,In_404);
xnor U1515 (N_1515,N_707,N_223);
nand U1516 (N_1516,N_237,N_273);
nand U1517 (N_1517,N_266,N_713);
nand U1518 (N_1518,N_469,N_627);
nand U1519 (N_1519,N_75,N_181);
nor U1520 (N_1520,In_882,N_169);
and U1521 (N_1521,N_4,N_735);
nor U1522 (N_1522,N_183,N_538);
xnor U1523 (N_1523,N_538,N_369);
nor U1524 (N_1524,N_695,N_706);
xnor U1525 (N_1525,N_217,In_1233);
or U1526 (N_1526,N_87,In_1562);
nand U1527 (N_1527,N_245,In_1485);
nor U1528 (N_1528,N_297,In_806);
and U1529 (N_1529,In_391,N_798);
or U1530 (N_1530,In_467,In_869);
or U1531 (N_1531,N_605,N_363);
nand U1532 (N_1532,In_1021,N_275);
nand U1533 (N_1533,N_228,N_179);
nor U1534 (N_1534,N_170,N_215);
and U1535 (N_1535,N_402,In_19);
or U1536 (N_1536,In_648,N_756);
nand U1537 (N_1537,In_786,N_4);
xnor U1538 (N_1538,N_340,In_1039);
nand U1539 (N_1539,N_532,In_140);
xor U1540 (N_1540,In_854,In_1367);
or U1541 (N_1541,In_1718,N_336);
nand U1542 (N_1542,N_688,N_421);
nor U1543 (N_1543,N_799,In_209);
nand U1544 (N_1544,N_54,In_1842);
or U1545 (N_1545,N_542,N_783);
or U1546 (N_1546,N_431,N_360);
xor U1547 (N_1547,N_259,N_357);
nand U1548 (N_1548,N_330,N_289);
nor U1549 (N_1549,In_218,N_173);
nand U1550 (N_1550,In_1870,In_185);
nand U1551 (N_1551,N_221,N_670);
or U1552 (N_1552,N_231,N_582);
or U1553 (N_1553,N_798,In_1481);
nand U1554 (N_1554,N_547,N_309);
or U1555 (N_1555,In_122,In_1596);
nor U1556 (N_1556,N_249,N_564);
nand U1557 (N_1557,In_428,N_50);
or U1558 (N_1558,N_134,In_489);
or U1559 (N_1559,N_148,N_7);
nor U1560 (N_1560,N_579,N_67);
xnor U1561 (N_1561,N_193,In_1588);
nor U1562 (N_1562,In_1434,N_472);
nand U1563 (N_1563,In_1391,In_1195);
and U1564 (N_1564,N_686,N_424);
nand U1565 (N_1565,N_236,N_792);
nand U1566 (N_1566,N_480,N_128);
and U1567 (N_1567,In_1276,N_313);
or U1568 (N_1568,In_257,N_265);
xnor U1569 (N_1569,N_636,N_791);
or U1570 (N_1570,N_565,N_562);
and U1571 (N_1571,N_748,N_648);
xor U1572 (N_1572,N_174,In_297);
or U1573 (N_1573,In_1156,N_126);
xnor U1574 (N_1574,N_73,N_675);
nor U1575 (N_1575,In_39,N_772);
xnor U1576 (N_1576,In_1593,In_459);
or U1577 (N_1577,N_430,N_726);
or U1578 (N_1578,In_1460,N_759);
and U1579 (N_1579,N_424,N_189);
xor U1580 (N_1580,N_103,N_629);
or U1581 (N_1581,N_119,N_679);
xor U1582 (N_1582,In_1100,N_116);
xor U1583 (N_1583,N_174,N_263);
and U1584 (N_1584,In_1235,N_1);
nand U1585 (N_1585,N_753,N_356);
or U1586 (N_1586,N_614,N_270);
nor U1587 (N_1587,N_775,In_724);
nor U1588 (N_1588,N_309,N_202);
nor U1589 (N_1589,In_297,N_710);
nor U1590 (N_1590,N_26,N_198);
xnor U1591 (N_1591,N_373,N_601);
or U1592 (N_1592,In_516,N_773);
xnor U1593 (N_1593,N_601,In_646);
or U1594 (N_1594,N_175,In_1718);
xnor U1595 (N_1595,N_471,In_897);
or U1596 (N_1596,N_196,In_705);
or U1597 (N_1597,N_60,In_1944);
nor U1598 (N_1598,N_17,N_140);
nand U1599 (N_1599,In_488,In_1367);
or U1600 (N_1600,N_1089,N_1206);
and U1601 (N_1601,N_1346,N_862);
nor U1602 (N_1602,N_1496,N_1201);
or U1603 (N_1603,N_1382,N_1113);
xor U1604 (N_1604,N_891,N_1061);
or U1605 (N_1605,N_955,N_1214);
xor U1606 (N_1606,N_1151,N_1376);
or U1607 (N_1607,N_1543,N_1316);
nor U1608 (N_1608,N_1006,N_1452);
nor U1609 (N_1609,N_990,N_1259);
and U1610 (N_1610,N_1593,N_1375);
nand U1611 (N_1611,N_1031,N_1184);
nand U1612 (N_1612,N_1161,N_825);
nor U1613 (N_1613,N_962,N_1482);
and U1614 (N_1614,N_1192,N_1003);
nor U1615 (N_1615,N_1583,N_1379);
nand U1616 (N_1616,N_1404,N_1580);
or U1617 (N_1617,N_840,N_947);
xnor U1618 (N_1618,N_1314,N_1535);
nand U1619 (N_1619,N_1509,N_1473);
xnor U1620 (N_1620,N_1144,N_992);
xor U1621 (N_1621,N_1095,N_975);
xor U1622 (N_1622,N_1170,N_1524);
nand U1623 (N_1623,N_1514,N_1560);
nand U1624 (N_1624,N_1054,N_961);
nand U1625 (N_1625,N_864,N_1211);
and U1626 (N_1626,N_1532,N_1015);
xnor U1627 (N_1627,N_996,N_1133);
and U1628 (N_1628,N_1347,N_854);
and U1629 (N_1629,N_1344,N_1077);
xor U1630 (N_1630,N_1283,N_1588);
or U1631 (N_1631,N_998,N_1490);
or U1632 (N_1632,N_1020,N_1026);
nor U1633 (N_1633,N_1472,N_1393);
nor U1634 (N_1634,N_1049,N_1233);
nand U1635 (N_1635,N_1372,N_855);
nand U1636 (N_1636,N_929,N_1056);
nor U1637 (N_1637,N_969,N_1323);
and U1638 (N_1638,N_834,N_1459);
nor U1639 (N_1639,N_1226,N_1384);
nand U1640 (N_1640,N_991,N_941);
nor U1641 (N_1641,N_1348,N_832);
and U1642 (N_1642,N_1210,N_1574);
nor U1643 (N_1643,N_1145,N_1036);
xnor U1644 (N_1644,N_935,N_1505);
xnor U1645 (N_1645,N_1456,N_918);
nand U1646 (N_1646,N_1394,N_1175);
and U1647 (N_1647,N_1235,N_1292);
nand U1648 (N_1648,N_1238,N_852);
nor U1649 (N_1649,N_810,N_1446);
nand U1650 (N_1650,N_882,N_874);
nor U1651 (N_1651,N_836,N_1554);
or U1652 (N_1652,N_1017,N_1309);
xor U1653 (N_1653,N_835,N_902);
or U1654 (N_1654,N_1424,N_850);
xor U1655 (N_1655,N_1432,N_1025);
xnor U1656 (N_1656,N_1132,N_1256);
nor U1657 (N_1657,N_1082,N_921);
nand U1658 (N_1658,N_1033,N_1258);
nand U1659 (N_1659,N_1391,N_1492);
nand U1660 (N_1660,N_1172,N_1048);
and U1661 (N_1661,N_1199,N_1182);
nor U1662 (N_1662,N_1590,N_1537);
nand U1663 (N_1663,N_1115,N_1156);
and U1664 (N_1664,N_1581,N_1387);
xnor U1665 (N_1665,N_1257,N_899);
or U1666 (N_1666,N_1534,N_1203);
nor U1667 (N_1667,N_1093,N_1547);
or U1668 (N_1668,N_903,N_1110);
xor U1669 (N_1669,N_970,N_1517);
xnor U1670 (N_1670,N_1024,N_1365);
nand U1671 (N_1671,N_1569,N_1087);
xnor U1672 (N_1672,N_1291,N_988);
or U1673 (N_1673,N_1080,N_1148);
nand U1674 (N_1674,N_1248,N_1433);
nand U1675 (N_1675,N_847,N_1478);
nor U1676 (N_1676,N_1474,N_1083);
xnor U1677 (N_1677,N_1029,N_1167);
and U1678 (N_1678,N_985,N_957);
and U1679 (N_1679,N_888,N_1378);
and U1680 (N_1680,N_1198,N_1460);
xnor U1681 (N_1681,N_1403,N_1045);
xnor U1682 (N_1682,N_1555,N_1253);
or U1683 (N_1683,N_812,N_1325);
and U1684 (N_1684,N_1039,N_1032);
nor U1685 (N_1685,N_1584,N_1103);
nand U1686 (N_1686,N_1191,N_1339);
and U1687 (N_1687,N_1450,N_1240);
or U1688 (N_1688,N_827,N_1207);
or U1689 (N_1689,N_1266,N_1204);
xnor U1690 (N_1690,N_1069,N_806);
and U1691 (N_1691,N_984,N_861);
nor U1692 (N_1692,N_1053,N_946);
nand U1693 (N_1693,N_1350,N_1563);
and U1694 (N_1694,N_1298,N_1486);
or U1695 (N_1695,N_971,N_1369);
nand U1696 (N_1696,N_1466,N_1058);
nand U1697 (N_1697,N_1421,N_1343);
nor U1698 (N_1698,N_1219,N_1313);
or U1699 (N_1699,N_1042,N_1107);
or U1700 (N_1700,N_1334,N_865);
nand U1701 (N_1701,N_1352,N_1010);
or U1702 (N_1702,N_1511,N_1544);
xor U1703 (N_1703,N_1118,N_1549);
or U1704 (N_1704,N_1592,N_1075);
xnor U1705 (N_1705,N_1550,N_1150);
nand U1706 (N_1706,N_1037,N_811);
nor U1707 (N_1707,N_910,N_1169);
xnor U1708 (N_1708,N_1531,N_1162);
or U1709 (N_1709,N_940,N_948);
xor U1710 (N_1710,N_1332,N_1336);
xor U1711 (N_1711,N_1079,N_1270);
and U1712 (N_1712,N_1453,N_978);
or U1713 (N_1713,N_1500,N_1396);
nor U1714 (N_1714,N_1142,N_845);
and U1715 (N_1715,N_817,N_1143);
or U1716 (N_1716,N_1520,N_923);
nand U1717 (N_1717,N_1244,N_1242);
and U1718 (N_1718,N_1299,N_837);
nand U1719 (N_1719,N_1043,N_1488);
and U1720 (N_1720,N_1497,N_878);
and U1721 (N_1721,N_954,N_1519);
xnor U1722 (N_1722,N_1282,N_1341);
nand U1723 (N_1723,N_1567,N_959);
xor U1724 (N_1724,N_1512,N_838);
and U1725 (N_1725,N_1239,N_1457);
xnor U1726 (N_1726,N_1419,N_1023);
or U1727 (N_1727,N_1502,N_1277);
nor U1728 (N_1728,N_1001,N_1220);
nand U1729 (N_1729,N_905,N_1545);
nand U1730 (N_1730,N_1533,N_1541);
nor U1731 (N_1731,N_1262,N_1153);
xor U1732 (N_1732,N_980,N_960);
and U1733 (N_1733,N_1279,N_1418);
and U1734 (N_1734,N_1126,N_816);
xnor U1735 (N_1735,N_1129,N_890);
xnor U1736 (N_1736,N_1448,N_885);
or U1737 (N_1737,N_1152,N_1196);
or U1738 (N_1738,N_1027,N_805);
or U1739 (N_1739,N_1002,N_908);
and U1740 (N_1740,N_1134,N_883);
and U1741 (N_1741,N_1377,N_1578);
xnor U1742 (N_1742,N_814,N_1485);
and U1743 (N_1743,N_1081,N_1098);
or U1744 (N_1744,N_1504,N_1455);
nor U1745 (N_1745,N_933,N_868);
nor U1746 (N_1746,N_1057,N_1561);
or U1747 (N_1747,N_1105,N_949);
xnor U1748 (N_1748,N_880,N_872);
and U1749 (N_1749,N_1445,N_1530);
and U1750 (N_1750,N_1289,N_926);
or U1751 (N_1751,N_927,N_907);
nand U1752 (N_1752,N_1529,N_1510);
or U1753 (N_1753,N_867,N_1494);
nand U1754 (N_1754,N_1194,N_1559);
xor U1755 (N_1755,N_1227,N_1451);
nor U1756 (N_1756,N_1405,N_889);
and U1757 (N_1757,N_1104,N_1383);
or U1758 (N_1758,N_1503,N_1528);
xor U1759 (N_1759,N_1338,N_1471);
nor U1760 (N_1760,N_1094,N_829);
or U1761 (N_1761,N_1442,N_932);
or U1762 (N_1762,N_1287,N_1074);
or U1763 (N_1763,N_1189,N_1436);
or U1764 (N_1764,N_1465,N_1435);
nand U1765 (N_1765,N_1271,N_1587);
and U1766 (N_1766,N_1102,N_922);
xnor U1767 (N_1767,N_917,N_1318);
and U1768 (N_1768,N_1356,N_1484);
or U1769 (N_1769,N_1038,N_912);
or U1770 (N_1770,N_1265,N_800);
xor U1771 (N_1771,N_851,N_1360);
or U1772 (N_1772,N_1441,N_1414);
nor U1773 (N_1773,N_887,N_989);
or U1774 (N_1774,N_1430,N_1247);
nor U1775 (N_1775,N_944,N_1286);
and U1776 (N_1776,N_1558,N_1562);
nand U1777 (N_1777,N_897,N_1141);
nor U1778 (N_1778,N_1523,N_1345);
nor U1779 (N_1779,N_1586,N_1368);
and U1780 (N_1780,N_1538,N_1197);
xnor U1781 (N_1781,N_1408,N_1493);
xor U1782 (N_1782,N_987,N_876);
nor U1783 (N_1783,N_1437,N_1363);
nor U1784 (N_1784,N_924,N_1487);
and U1785 (N_1785,N_1234,N_981);
nand U1786 (N_1786,N_1333,N_1236);
or U1787 (N_1787,N_1216,N_1185);
or U1788 (N_1788,N_1221,N_1507);
and U1789 (N_1789,N_1136,N_1096);
or U1790 (N_1790,N_1426,N_1278);
xnor U1791 (N_1791,N_1138,N_1159);
or U1792 (N_1792,N_1551,N_1051);
xor U1793 (N_1793,N_1285,N_1301);
xor U1794 (N_1794,N_904,N_1546);
and U1795 (N_1795,N_1392,N_1140);
or U1796 (N_1796,N_920,N_906);
xor U1797 (N_1797,N_1386,N_1284);
nand U1798 (N_1798,N_1317,N_1335);
nand U1799 (N_1799,N_1599,N_1007);
xor U1800 (N_1800,N_826,N_1331);
nand U1801 (N_1801,N_1390,N_1373);
and U1802 (N_1802,N_1168,N_824);
nand U1803 (N_1803,N_1060,N_1388);
and U1804 (N_1804,N_1164,N_815);
nand U1805 (N_1805,N_1462,N_1326);
xor U1806 (N_1806,N_1355,N_1237);
or U1807 (N_1807,N_943,N_844);
xnor U1808 (N_1808,N_1040,N_1542);
and U1809 (N_1809,N_953,N_892);
nand U1810 (N_1810,N_1229,N_1536);
nand U1811 (N_1811,N_1028,N_958);
xor U1812 (N_1812,N_1364,N_1070);
nor U1813 (N_1813,N_1190,N_1123);
nor U1814 (N_1814,N_841,N_1109);
and U1815 (N_1815,N_1090,N_1328);
xor U1816 (N_1816,N_1508,N_1297);
or U1817 (N_1817,N_1217,N_1417);
xor U1818 (N_1818,N_1296,N_1183);
xnor U1819 (N_1819,N_863,N_1427);
or U1820 (N_1820,N_1389,N_1585);
or U1821 (N_1821,N_1085,N_977);
nor U1822 (N_1822,N_1273,N_1357);
or U1823 (N_1823,N_1186,N_1052);
nand U1824 (N_1824,N_1330,N_813);
and U1825 (N_1825,N_1411,N_1117);
or U1826 (N_1826,N_1556,N_1252);
and U1827 (N_1827,N_1425,N_1366);
and U1828 (N_1828,N_1209,N_1122);
xor U1829 (N_1829,N_1187,N_1181);
and U1830 (N_1830,N_909,N_1407);
or U1831 (N_1831,N_1106,N_1416);
xor U1832 (N_1832,N_860,N_1062);
or U1833 (N_1833,N_822,N_928);
and U1834 (N_1834,N_1385,N_1565);
xor U1835 (N_1835,N_1076,N_1063);
nor U1836 (N_1836,N_1361,N_1522);
or U1837 (N_1837,N_1557,N_1423);
nand U1838 (N_1838,N_1012,N_1513);
nor U1839 (N_1839,N_1370,N_1467);
nor U1840 (N_1840,N_1575,N_1255);
nand U1841 (N_1841,N_1254,N_1358);
nor U1842 (N_1842,N_994,N_1367);
nand U1843 (N_1843,N_893,N_1264);
nand U1844 (N_1844,N_1374,N_965);
nor U1845 (N_1845,N_1495,N_1014);
or U1846 (N_1846,N_1188,N_1163);
and U1847 (N_1847,N_913,N_1506);
nand U1848 (N_1848,N_1552,N_1195);
nor U1849 (N_1849,N_1499,N_1166);
xnor U1850 (N_1850,N_1213,N_1571);
and U1851 (N_1851,N_914,N_1073);
nand U1852 (N_1852,N_1092,N_915);
and U1853 (N_1853,N_1315,N_1398);
xor U1854 (N_1854,N_1349,N_870);
and U1855 (N_1855,N_916,N_972);
nand U1856 (N_1856,N_1594,N_1591);
nor U1857 (N_1857,N_1527,N_1570);
and U1858 (N_1858,N_1111,N_937);
xor U1859 (N_1859,N_1526,N_1000);
xnor U1860 (N_1860,N_1030,N_1274);
nor U1861 (N_1861,N_1112,N_843);
xnor U1862 (N_1862,N_1311,N_1035);
nor U1863 (N_1863,N_1130,N_1322);
nand U1864 (N_1864,N_1470,N_1034);
xor U1865 (N_1865,N_1589,N_1200);
xor U1866 (N_1866,N_1174,N_1295);
xor U1867 (N_1867,N_1097,N_1091);
xnor U1868 (N_1868,N_808,N_995);
or U1869 (N_1869,N_1165,N_1212);
and U1870 (N_1870,N_1401,N_1251);
nor U1871 (N_1871,N_895,N_1135);
or U1872 (N_1872,N_942,N_1064);
xor U1873 (N_1873,N_879,N_807);
and U1874 (N_1874,N_1149,N_1116);
and U1875 (N_1875,N_1086,N_1263);
and U1876 (N_1876,N_1171,N_1449);
nor U1877 (N_1877,N_884,N_1231);
nand U1878 (N_1878,N_1498,N_1595);
and U1879 (N_1879,N_1120,N_930);
nand U1880 (N_1880,N_1539,N_1067);
xor U1881 (N_1881,N_1268,N_925);
xor U1882 (N_1882,N_1059,N_1154);
nand U1883 (N_1883,N_1576,N_1225);
or U1884 (N_1884,N_1260,N_979);
xnor U1885 (N_1885,N_976,N_1124);
nand U1886 (N_1886,N_833,N_1463);
and U1887 (N_1887,N_1121,N_1250);
and U1888 (N_1888,N_1232,N_1308);
nand U1889 (N_1889,N_1481,N_842);
nand U1890 (N_1890,N_1516,N_1568);
nand U1891 (N_1891,N_1329,N_1267);
and U1892 (N_1892,N_1072,N_1066);
xor U1893 (N_1893,N_1397,N_1139);
or U1894 (N_1894,N_818,N_938);
nor U1895 (N_1895,N_967,N_1303);
and U1896 (N_1896,N_1005,N_1304);
nand U1897 (N_1897,N_858,N_1202);
and U1898 (N_1898,N_1249,N_1158);
nand U1899 (N_1899,N_819,N_869);
nand U1900 (N_1900,N_1055,N_974);
nor U1901 (N_1901,N_1218,N_801);
nand U1902 (N_1902,N_1479,N_911);
nand U1903 (N_1903,N_839,N_1176);
nand U1904 (N_1904,N_831,N_1359);
or U1905 (N_1905,N_871,N_931);
nor U1906 (N_1906,N_1157,N_1160);
xnor U1907 (N_1907,N_1230,N_1008);
nor U1908 (N_1908,N_1521,N_951);
nor U1909 (N_1909,N_1518,N_828);
nand U1910 (N_1910,N_1281,N_1489);
nor U1911 (N_1911,N_1119,N_1127);
nand U1912 (N_1912,N_848,N_1241);
or U1913 (N_1913,N_859,N_1553);
or U1914 (N_1914,N_986,N_1099);
xnor U1915 (N_1915,N_1572,N_1276);
xor U1916 (N_1916,N_1579,N_952);
or U1917 (N_1917,N_1422,N_1337);
nand U1918 (N_1918,N_1300,N_1320);
nand U1919 (N_1919,N_982,N_898);
xor U1920 (N_1920,N_993,N_1108);
nand U1921 (N_1921,N_1540,N_1362);
and U1922 (N_1922,N_956,N_1406);
nor U1923 (N_1923,N_1047,N_1412);
xor U1924 (N_1924,N_809,N_1454);
and U1925 (N_1925,N_1410,N_857);
and U1926 (N_1926,N_1147,N_1447);
and U1927 (N_1927,N_1215,N_919);
xor U1928 (N_1928,N_1420,N_973);
and U1929 (N_1929,N_945,N_1101);
and U1930 (N_1930,N_1193,N_1431);
nand U1931 (N_1931,N_1573,N_1475);
and U1932 (N_1932,N_1429,N_804);
nor U1933 (N_1933,N_963,N_1428);
nor U1934 (N_1934,N_1177,N_1041);
nand U1935 (N_1935,N_1018,N_1223);
or U1936 (N_1936,N_1114,N_1354);
nor U1937 (N_1937,N_1413,N_1179);
nor U1938 (N_1938,N_1071,N_873);
nor U1939 (N_1939,N_1483,N_901);
or U1940 (N_1940,N_1525,N_1065);
xnor U1941 (N_1941,N_1084,N_1324);
nand U1942 (N_1942,N_1131,N_1180);
nand U1943 (N_1943,N_1302,N_894);
and U1944 (N_1944,N_1128,N_1078);
or U1945 (N_1945,N_1477,N_1178);
xnor U1946 (N_1946,N_1501,N_1208);
or U1947 (N_1947,N_1275,N_823);
nor U1948 (N_1948,N_1443,N_1319);
and U1949 (N_1949,N_1245,N_821);
or U1950 (N_1950,N_1340,N_1269);
and U1951 (N_1951,N_964,N_1222);
xor U1952 (N_1952,N_1321,N_1310);
nor U1953 (N_1953,N_1548,N_1019);
nand U1954 (N_1954,N_968,N_966);
or U1955 (N_1955,N_999,N_1044);
nor U1956 (N_1956,N_1402,N_936);
and U1957 (N_1957,N_1125,N_1088);
or U1958 (N_1958,N_1046,N_1380);
nor U1959 (N_1959,N_1598,N_1011);
xor U1960 (N_1960,N_1137,N_849);
xor U1961 (N_1961,N_1280,N_1224);
nor U1962 (N_1962,N_1100,N_803);
xor U1963 (N_1963,N_1243,N_820);
nor U1964 (N_1964,N_1458,N_1021);
and U1965 (N_1965,N_1305,N_1342);
nand U1966 (N_1966,N_1351,N_866);
and U1967 (N_1967,N_1468,N_1272);
xor U1968 (N_1968,N_1440,N_1399);
and U1969 (N_1969,N_1327,N_1566);
nor U1970 (N_1970,N_1068,N_881);
xor U1971 (N_1971,N_856,N_1173);
or U1972 (N_1972,N_939,N_1381);
or U1973 (N_1973,N_1596,N_1438);
nor U1974 (N_1974,N_997,N_1004);
and U1975 (N_1975,N_1577,N_1461);
or U1976 (N_1976,N_877,N_1290);
nor U1977 (N_1977,N_1564,N_1371);
nor U1978 (N_1978,N_1582,N_1016);
or U1979 (N_1979,N_1261,N_1246);
nand U1980 (N_1980,N_1013,N_1307);
and U1981 (N_1981,N_1294,N_900);
or U1982 (N_1982,N_1293,N_1597);
nor U1983 (N_1983,N_853,N_1155);
and U1984 (N_1984,N_875,N_1480);
nor U1985 (N_1985,N_1515,N_1228);
nand U1986 (N_1986,N_830,N_886);
and U1987 (N_1987,N_1476,N_1415);
nand U1988 (N_1988,N_1353,N_1009);
nor U1989 (N_1989,N_950,N_983);
nand U1990 (N_1990,N_1491,N_1400);
and U1991 (N_1991,N_846,N_1444);
and U1992 (N_1992,N_1288,N_1312);
nor U1993 (N_1993,N_1409,N_1050);
nor U1994 (N_1994,N_1306,N_934);
nor U1995 (N_1995,N_1469,N_1439);
or U1996 (N_1996,N_1146,N_1205);
nor U1997 (N_1997,N_896,N_1022);
and U1998 (N_1998,N_1434,N_1464);
nand U1999 (N_1999,N_802,N_1395);
nand U2000 (N_2000,N_1546,N_1386);
or U2001 (N_2001,N_1333,N_1155);
nor U2002 (N_2002,N_1115,N_1237);
or U2003 (N_2003,N_1193,N_1159);
nor U2004 (N_2004,N_1489,N_838);
or U2005 (N_2005,N_815,N_988);
nand U2006 (N_2006,N_897,N_1466);
nand U2007 (N_2007,N_1309,N_969);
nor U2008 (N_2008,N_1180,N_1345);
xor U2009 (N_2009,N_1372,N_831);
or U2010 (N_2010,N_1308,N_1335);
or U2011 (N_2011,N_1570,N_1101);
xnor U2012 (N_2012,N_1109,N_1545);
and U2013 (N_2013,N_1010,N_1309);
or U2014 (N_2014,N_1065,N_958);
and U2015 (N_2015,N_1301,N_1087);
and U2016 (N_2016,N_1509,N_1460);
nand U2017 (N_2017,N_1057,N_823);
nor U2018 (N_2018,N_1132,N_1463);
or U2019 (N_2019,N_1289,N_1158);
or U2020 (N_2020,N_1147,N_935);
nor U2021 (N_2021,N_869,N_1386);
xor U2022 (N_2022,N_876,N_1340);
and U2023 (N_2023,N_1397,N_968);
nand U2024 (N_2024,N_1323,N_1482);
and U2025 (N_2025,N_1591,N_956);
nand U2026 (N_2026,N_1492,N_1397);
and U2027 (N_2027,N_981,N_1549);
or U2028 (N_2028,N_1385,N_1030);
and U2029 (N_2029,N_983,N_899);
xor U2030 (N_2030,N_861,N_1295);
nand U2031 (N_2031,N_1194,N_1082);
nand U2032 (N_2032,N_1425,N_1152);
nor U2033 (N_2033,N_1119,N_870);
and U2034 (N_2034,N_874,N_1511);
or U2035 (N_2035,N_965,N_819);
and U2036 (N_2036,N_872,N_1494);
xnor U2037 (N_2037,N_1013,N_1143);
nand U2038 (N_2038,N_1205,N_1098);
xor U2039 (N_2039,N_1113,N_1051);
nand U2040 (N_2040,N_1049,N_1555);
and U2041 (N_2041,N_919,N_971);
xnor U2042 (N_2042,N_1445,N_890);
and U2043 (N_2043,N_927,N_807);
nand U2044 (N_2044,N_1504,N_1053);
or U2045 (N_2045,N_1182,N_1141);
nand U2046 (N_2046,N_1370,N_1567);
nor U2047 (N_2047,N_909,N_839);
and U2048 (N_2048,N_1102,N_801);
xnor U2049 (N_2049,N_1074,N_1560);
xor U2050 (N_2050,N_1188,N_1323);
and U2051 (N_2051,N_1117,N_1165);
xor U2052 (N_2052,N_891,N_1279);
or U2053 (N_2053,N_1251,N_866);
xor U2054 (N_2054,N_1511,N_1534);
and U2055 (N_2055,N_1450,N_1383);
xnor U2056 (N_2056,N_1575,N_1519);
xnor U2057 (N_2057,N_1296,N_1266);
or U2058 (N_2058,N_1048,N_961);
and U2059 (N_2059,N_1463,N_920);
nor U2060 (N_2060,N_1564,N_1385);
or U2061 (N_2061,N_1482,N_1277);
or U2062 (N_2062,N_1164,N_1348);
nand U2063 (N_2063,N_1433,N_1278);
and U2064 (N_2064,N_1575,N_1510);
nand U2065 (N_2065,N_1480,N_937);
nor U2066 (N_2066,N_1459,N_1443);
and U2067 (N_2067,N_1541,N_865);
nand U2068 (N_2068,N_1297,N_1226);
and U2069 (N_2069,N_1497,N_1408);
xnor U2070 (N_2070,N_875,N_1281);
nand U2071 (N_2071,N_1461,N_1210);
and U2072 (N_2072,N_835,N_1403);
or U2073 (N_2073,N_1155,N_1102);
xnor U2074 (N_2074,N_1366,N_1156);
and U2075 (N_2075,N_814,N_1403);
nor U2076 (N_2076,N_922,N_1191);
xnor U2077 (N_2077,N_955,N_837);
nor U2078 (N_2078,N_1370,N_1595);
nand U2079 (N_2079,N_1248,N_1241);
or U2080 (N_2080,N_1030,N_1513);
nor U2081 (N_2081,N_1067,N_1384);
nand U2082 (N_2082,N_949,N_1309);
nor U2083 (N_2083,N_1573,N_1173);
xnor U2084 (N_2084,N_1404,N_1463);
xor U2085 (N_2085,N_1398,N_1263);
and U2086 (N_2086,N_959,N_956);
nand U2087 (N_2087,N_1293,N_1526);
xnor U2088 (N_2088,N_1521,N_1487);
xor U2089 (N_2089,N_1060,N_872);
nor U2090 (N_2090,N_993,N_1595);
xor U2091 (N_2091,N_1393,N_1300);
nand U2092 (N_2092,N_1479,N_1426);
nor U2093 (N_2093,N_1471,N_1205);
nor U2094 (N_2094,N_848,N_1030);
and U2095 (N_2095,N_1245,N_1254);
and U2096 (N_2096,N_1490,N_913);
or U2097 (N_2097,N_1245,N_1374);
nand U2098 (N_2098,N_1501,N_1131);
or U2099 (N_2099,N_1327,N_889);
xor U2100 (N_2100,N_1435,N_923);
xor U2101 (N_2101,N_1540,N_1285);
or U2102 (N_2102,N_871,N_1264);
or U2103 (N_2103,N_1324,N_1594);
nor U2104 (N_2104,N_1209,N_1380);
nor U2105 (N_2105,N_952,N_1457);
and U2106 (N_2106,N_1035,N_1247);
or U2107 (N_2107,N_1138,N_1364);
nor U2108 (N_2108,N_1148,N_1430);
nand U2109 (N_2109,N_1361,N_910);
xnor U2110 (N_2110,N_804,N_879);
nor U2111 (N_2111,N_1412,N_1536);
xor U2112 (N_2112,N_854,N_1220);
and U2113 (N_2113,N_870,N_1296);
and U2114 (N_2114,N_1163,N_1313);
xnor U2115 (N_2115,N_1362,N_1296);
xnor U2116 (N_2116,N_1155,N_1426);
nand U2117 (N_2117,N_1193,N_1367);
and U2118 (N_2118,N_1092,N_1464);
or U2119 (N_2119,N_1192,N_1046);
nor U2120 (N_2120,N_894,N_977);
nand U2121 (N_2121,N_1453,N_1190);
xnor U2122 (N_2122,N_1582,N_1481);
nand U2123 (N_2123,N_1441,N_1391);
and U2124 (N_2124,N_1257,N_1518);
nor U2125 (N_2125,N_1395,N_1155);
xnor U2126 (N_2126,N_1044,N_1111);
nand U2127 (N_2127,N_1189,N_1509);
or U2128 (N_2128,N_1024,N_1498);
nand U2129 (N_2129,N_1559,N_1518);
xnor U2130 (N_2130,N_943,N_839);
xnor U2131 (N_2131,N_962,N_1564);
nand U2132 (N_2132,N_1587,N_1368);
xor U2133 (N_2133,N_989,N_901);
nand U2134 (N_2134,N_848,N_1219);
xnor U2135 (N_2135,N_808,N_1490);
nor U2136 (N_2136,N_1154,N_959);
or U2137 (N_2137,N_1215,N_1368);
nor U2138 (N_2138,N_1543,N_1334);
and U2139 (N_2139,N_1404,N_824);
xor U2140 (N_2140,N_1324,N_1108);
nand U2141 (N_2141,N_1416,N_1356);
or U2142 (N_2142,N_1541,N_1410);
xor U2143 (N_2143,N_1289,N_1350);
and U2144 (N_2144,N_1172,N_924);
or U2145 (N_2145,N_1352,N_1473);
or U2146 (N_2146,N_818,N_1208);
nor U2147 (N_2147,N_1358,N_1195);
and U2148 (N_2148,N_1406,N_904);
or U2149 (N_2149,N_847,N_983);
nor U2150 (N_2150,N_1539,N_1319);
nand U2151 (N_2151,N_975,N_1484);
nor U2152 (N_2152,N_932,N_1542);
or U2153 (N_2153,N_934,N_1078);
nor U2154 (N_2154,N_853,N_1549);
nor U2155 (N_2155,N_1160,N_1508);
xor U2156 (N_2156,N_1295,N_1486);
or U2157 (N_2157,N_906,N_1593);
or U2158 (N_2158,N_1071,N_1390);
or U2159 (N_2159,N_1500,N_1261);
xor U2160 (N_2160,N_1403,N_1075);
nand U2161 (N_2161,N_1301,N_961);
or U2162 (N_2162,N_837,N_1312);
nand U2163 (N_2163,N_1320,N_967);
nand U2164 (N_2164,N_1072,N_903);
and U2165 (N_2165,N_1368,N_1162);
nor U2166 (N_2166,N_1347,N_1464);
nor U2167 (N_2167,N_1471,N_1303);
or U2168 (N_2168,N_947,N_1396);
xnor U2169 (N_2169,N_859,N_1267);
and U2170 (N_2170,N_1432,N_1174);
and U2171 (N_2171,N_807,N_1366);
and U2172 (N_2172,N_1326,N_1205);
nand U2173 (N_2173,N_837,N_978);
or U2174 (N_2174,N_981,N_946);
or U2175 (N_2175,N_1081,N_1263);
xor U2176 (N_2176,N_1541,N_928);
xnor U2177 (N_2177,N_1271,N_1053);
xnor U2178 (N_2178,N_1405,N_836);
nor U2179 (N_2179,N_1364,N_1473);
nand U2180 (N_2180,N_1230,N_1233);
or U2181 (N_2181,N_1269,N_1330);
xor U2182 (N_2182,N_1497,N_1003);
nor U2183 (N_2183,N_1277,N_931);
nand U2184 (N_2184,N_1541,N_1574);
and U2185 (N_2185,N_1528,N_1501);
nand U2186 (N_2186,N_1081,N_1381);
or U2187 (N_2187,N_860,N_995);
and U2188 (N_2188,N_1345,N_1037);
and U2189 (N_2189,N_1312,N_1037);
nand U2190 (N_2190,N_900,N_1332);
xnor U2191 (N_2191,N_1496,N_1358);
nand U2192 (N_2192,N_871,N_1542);
nor U2193 (N_2193,N_1025,N_1137);
nor U2194 (N_2194,N_1016,N_1378);
or U2195 (N_2195,N_1002,N_1348);
nand U2196 (N_2196,N_1173,N_807);
or U2197 (N_2197,N_1384,N_1490);
nor U2198 (N_2198,N_1509,N_1251);
nand U2199 (N_2199,N_1430,N_848);
or U2200 (N_2200,N_1007,N_1232);
nand U2201 (N_2201,N_1550,N_1406);
nor U2202 (N_2202,N_1251,N_1214);
xor U2203 (N_2203,N_1026,N_1049);
xnor U2204 (N_2204,N_1547,N_1450);
xnor U2205 (N_2205,N_841,N_1220);
nand U2206 (N_2206,N_1090,N_1122);
or U2207 (N_2207,N_1456,N_1253);
nand U2208 (N_2208,N_914,N_1438);
nand U2209 (N_2209,N_1317,N_1369);
xor U2210 (N_2210,N_1275,N_1311);
or U2211 (N_2211,N_1183,N_1200);
and U2212 (N_2212,N_809,N_1149);
and U2213 (N_2213,N_1314,N_877);
or U2214 (N_2214,N_1092,N_1127);
nand U2215 (N_2215,N_981,N_1113);
nand U2216 (N_2216,N_1135,N_1498);
or U2217 (N_2217,N_1430,N_1572);
xor U2218 (N_2218,N_1370,N_1056);
xnor U2219 (N_2219,N_918,N_1273);
or U2220 (N_2220,N_1302,N_984);
xor U2221 (N_2221,N_1204,N_867);
or U2222 (N_2222,N_1441,N_1551);
and U2223 (N_2223,N_1025,N_1254);
nand U2224 (N_2224,N_1549,N_1239);
or U2225 (N_2225,N_969,N_1136);
nor U2226 (N_2226,N_1033,N_892);
or U2227 (N_2227,N_1388,N_1058);
nand U2228 (N_2228,N_1227,N_1421);
xor U2229 (N_2229,N_1501,N_1370);
and U2230 (N_2230,N_1173,N_1267);
nand U2231 (N_2231,N_1036,N_1458);
and U2232 (N_2232,N_1391,N_1563);
nand U2233 (N_2233,N_1576,N_895);
or U2234 (N_2234,N_1132,N_1382);
nand U2235 (N_2235,N_1431,N_1340);
or U2236 (N_2236,N_1268,N_1077);
and U2237 (N_2237,N_948,N_1554);
nor U2238 (N_2238,N_923,N_948);
and U2239 (N_2239,N_1422,N_1217);
xor U2240 (N_2240,N_1532,N_986);
nor U2241 (N_2241,N_1513,N_1019);
and U2242 (N_2242,N_1571,N_974);
nor U2243 (N_2243,N_1564,N_992);
nand U2244 (N_2244,N_917,N_1320);
xnor U2245 (N_2245,N_1140,N_937);
nor U2246 (N_2246,N_1573,N_952);
nor U2247 (N_2247,N_1092,N_1525);
and U2248 (N_2248,N_1599,N_1029);
or U2249 (N_2249,N_1030,N_1473);
nand U2250 (N_2250,N_1213,N_1033);
or U2251 (N_2251,N_979,N_1127);
xnor U2252 (N_2252,N_1251,N_1479);
nor U2253 (N_2253,N_1214,N_832);
xor U2254 (N_2254,N_913,N_1535);
xor U2255 (N_2255,N_1180,N_1318);
nor U2256 (N_2256,N_833,N_1558);
nand U2257 (N_2257,N_895,N_1207);
nand U2258 (N_2258,N_1121,N_1388);
nand U2259 (N_2259,N_1512,N_916);
xor U2260 (N_2260,N_1015,N_1088);
and U2261 (N_2261,N_1082,N_831);
nand U2262 (N_2262,N_802,N_1585);
nor U2263 (N_2263,N_884,N_1576);
xor U2264 (N_2264,N_865,N_1560);
xnor U2265 (N_2265,N_1413,N_982);
and U2266 (N_2266,N_1034,N_1204);
or U2267 (N_2267,N_1574,N_1125);
nor U2268 (N_2268,N_1251,N_892);
xnor U2269 (N_2269,N_896,N_929);
xor U2270 (N_2270,N_1103,N_829);
nand U2271 (N_2271,N_1071,N_939);
or U2272 (N_2272,N_1032,N_1022);
xor U2273 (N_2273,N_1162,N_993);
and U2274 (N_2274,N_1412,N_1101);
and U2275 (N_2275,N_916,N_1073);
or U2276 (N_2276,N_1066,N_1135);
nand U2277 (N_2277,N_911,N_1578);
and U2278 (N_2278,N_860,N_1599);
or U2279 (N_2279,N_918,N_1414);
nor U2280 (N_2280,N_1093,N_1404);
nor U2281 (N_2281,N_1281,N_1577);
xor U2282 (N_2282,N_1004,N_1112);
or U2283 (N_2283,N_942,N_1195);
or U2284 (N_2284,N_1395,N_819);
and U2285 (N_2285,N_1380,N_1132);
nor U2286 (N_2286,N_1161,N_829);
and U2287 (N_2287,N_1244,N_1217);
nor U2288 (N_2288,N_825,N_1234);
and U2289 (N_2289,N_1078,N_1260);
and U2290 (N_2290,N_1417,N_1254);
and U2291 (N_2291,N_1529,N_1400);
xor U2292 (N_2292,N_1454,N_1047);
xor U2293 (N_2293,N_932,N_1402);
nor U2294 (N_2294,N_1376,N_1185);
nor U2295 (N_2295,N_1260,N_977);
and U2296 (N_2296,N_1554,N_1151);
or U2297 (N_2297,N_885,N_1023);
xor U2298 (N_2298,N_1577,N_1175);
nand U2299 (N_2299,N_1258,N_1240);
nor U2300 (N_2300,N_1072,N_1127);
nor U2301 (N_2301,N_849,N_1019);
or U2302 (N_2302,N_952,N_1464);
nand U2303 (N_2303,N_1523,N_1019);
xor U2304 (N_2304,N_1080,N_908);
and U2305 (N_2305,N_1143,N_1505);
xnor U2306 (N_2306,N_1505,N_1433);
or U2307 (N_2307,N_925,N_1532);
nand U2308 (N_2308,N_1526,N_1035);
or U2309 (N_2309,N_1289,N_1466);
and U2310 (N_2310,N_1395,N_1284);
nor U2311 (N_2311,N_1563,N_1264);
or U2312 (N_2312,N_1129,N_1217);
and U2313 (N_2313,N_1485,N_980);
or U2314 (N_2314,N_1540,N_876);
xnor U2315 (N_2315,N_1588,N_855);
or U2316 (N_2316,N_1516,N_877);
and U2317 (N_2317,N_1044,N_956);
nor U2318 (N_2318,N_1052,N_1008);
nand U2319 (N_2319,N_1016,N_1292);
nand U2320 (N_2320,N_1536,N_1035);
nand U2321 (N_2321,N_1127,N_1488);
xor U2322 (N_2322,N_1575,N_1188);
and U2323 (N_2323,N_1361,N_1202);
or U2324 (N_2324,N_1518,N_1420);
xnor U2325 (N_2325,N_1406,N_874);
nand U2326 (N_2326,N_1324,N_863);
nand U2327 (N_2327,N_820,N_914);
or U2328 (N_2328,N_1459,N_1073);
nand U2329 (N_2329,N_819,N_1357);
and U2330 (N_2330,N_1360,N_1507);
nand U2331 (N_2331,N_1438,N_1265);
nand U2332 (N_2332,N_1162,N_1282);
nand U2333 (N_2333,N_848,N_822);
or U2334 (N_2334,N_1280,N_1345);
nor U2335 (N_2335,N_906,N_1367);
nor U2336 (N_2336,N_985,N_1333);
or U2337 (N_2337,N_1454,N_1225);
xor U2338 (N_2338,N_1021,N_1118);
and U2339 (N_2339,N_1222,N_1520);
or U2340 (N_2340,N_1482,N_1295);
xor U2341 (N_2341,N_1573,N_872);
xor U2342 (N_2342,N_908,N_1444);
and U2343 (N_2343,N_1369,N_1358);
nor U2344 (N_2344,N_1230,N_885);
or U2345 (N_2345,N_1440,N_1402);
xor U2346 (N_2346,N_966,N_1012);
xor U2347 (N_2347,N_1267,N_1209);
xor U2348 (N_2348,N_1120,N_1364);
nand U2349 (N_2349,N_988,N_1425);
nor U2350 (N_2350,N_1245,N_833);
nand U2351 (N_2351,N_1432,N_1146);
or U2352 (N_2352,N_1533,N_1359);
nor U2353 (N_2353,N_1125,N_829);
nor U2354 (N_2354,N_852,N_1361);
nor U2355 (N_2355,N_1409,N_1017);
xnor U2356 (N_2356,N_1377,N_1453);
and U2357 (N_2357,N_1001,N_1076);
nand U2358 (N_2358,N_1251,N_1058);
and U2359 (N_2359,N_1336,N_1425);
xor U2360 (N_2360,N_1210,N_949);
nand U2361 (N_2361,N_964,N_1524);
or U2362 (N_2362,N_908,N_811);
xnor U2363 (N_2363,N_832,N_1552);
nor U2364 (N_2364,N_1263,N_1443);
and U2365 (N_2365,N_952,N_1538);
or U2366 (N_2366,N_1468,N_1157);
nand U2367 (N_2367,N_1484,N_1000);
or U2368 (N_2368,N_1503,N_1273);
nand U2369 (N_2369,N_1241,N_1416);
or U2370 (N_2370,N_1522,N_1050);
xnor U2371 (N_2371,N_1508,N_1137);
nor U2372 (N_2372,N_1282,N_1295);
xor U2373 (N_2373,N_943,N_1445);
or U2374 (N_2374,N_849,N_1469);
nor U2375 (N_2375,N_1540,N_822);
xnor U2376 (N_2376,N_1545,N_1572);
nor U2377 (N_2377,N_1474,N_992);
nand U2378 (N_2378,N_1363,N_1037);
xor U2379 (N_2379,N_1580,N_1570);
or U2380 (N_2380,N_1090,N_1289);
nor U2381 (N_2381,N_1411,N_1229);
nand U2382 (N_2382,N_1214,N_1365);
or U2383 (N_2383,N_1366,N_1460);
nor U2384 (N_2384,N_1283,N_1187);
or U2385 (N_2385,N_1376,N_1306);
xor U2386 (N_2386,N_1181,N_866);
or U2387 (N_2387,N_1544,N_1183);
nor U2388 (N_2388,N_993,N_1178);
nor U2389 (N_2389,N_1217,N_1596);
nand U2390 (N_2390,N_1459,N_1216);
and U2391 (N_2391,N_1279,N_1008);
nor U2392 (N_2392,N_1378,N_851);
and U2393 (N_2393,N_876,N_1044);
nand U2394 (N_2394,N_1253,N_1424);
and U2395 (N_2395,N_1235,N_1599);
xnor U2396 (N_2396,N_1037,N_1179);
and U2397 (N_2397,N_1374,N_968);
nor U2398 (N_2398,N_1308,N_823);
and U2399 (N_2399,N_891,N_1323);
nor U2400 (N_2400,N_2184,N_1832);
xor U2401 (N_2401,N_2242,N_1700);
or U2402 (N_2402,N_1677,N_1696);
xnor U2403 (N_2403,N_2110,N_2002);
or U2404 (N_2404,N_2001,N_2353);
xor U2405 (N_2405,N_2259,N_1951);
or U2406 (N_2406,N_2303,N_1955);
nand U2407 (N_2407,N_2337,N_1830);
and U2408 (N_2408,N_2027,N_1935);
nor U2409 (N_2409,N_2115,N_2061);
and U2410 (N_2410,N_1644,N_2006);
nor U2411 (N_2411,N_1980,N_2046);
xnor U2412 (N_2412,N_2397,N_1697);
and U2413 (N_2413,N_2272,N_2394);
and U2414 (N_2414,N_2200,N_2385);
and U2415 (N_2415,N_2297,N_1905);
or U2416 (N_2416,N_2372,N_2364);
and U2417 (N_2417,N_2008,N_1908);
and U2418 (N_2418,N_1606,N_2195);
nor U2419 (N_2419,N_2236,N_1671);
and U2420 (N_2420,N_2192,N_1719);
or U2421 (N_2421,N_1777,N_1919);
or U2422 (N_2422,N_2326,N_2298);
xnor U2423 (N_2423,N_2130,N_2309);
or U2424 (N_2424,N_1786,N_2112);
nor U2425 (N_2425,N_2310,N_1812);
and U2426 (N_2426,N_2087,N_1926);
or U2427 (N_2427,N_1614,N_2140);
and U2428 (N_2428,N_2370,N_1865);
and U2429 (N_2429,N_1949,N_1661);
xor U2430 (N_2430,N_2176,N_1858);
or U2431 (N_2431,N_2315,N_1669);
nor U2432 (N_2432,N_2304,N_1645);
nand U2433 (N_2433,N_2283,N_1646);
nor U2434 (N_2434,N_2237,N_2033);
nor U2435 (N_2435,N_2308,N_2345);
xor U2436 (N_2436,N_1826,N_1611);
nor U2437 (N_2437,N_2162,N_1638);
and U2438 (N_2438,N_1977,N_2264);
nand U2439 (N_2439,N_2206,N_1906);
and U2440 (N_2440,N_2211,N_1774);
and U2441 (N_2441,N_2220,N_1991);
nor U2442 (N_2442,N_1735,N_1924);
or U2443 (N_2443,N_1730,N_2302);
nand U2444 (N_2444,N_1983,N_2320);
xor U2445 (N_2445,N_1632,N_1739);
or U2446 (N_2446,N_1993,N_2399);
nand U2447 (N_2447,N_1605,N_1895);
nand U2448 (N_2448,N_2014,N_2371);
xor U2449 (N_2449,N_2123,N_1850);
nand U2450 (N_2450,N_2052,N_1925);
or U2451 (N_2451,N_1778,N_1853);
nor U2452 (N_2452,N_2156,N_2172);
nor U2453 (N_2453,N_1770,N_1887);
xnor U2454 (N_2454,N_2081,N_2148);
nand U2455 (N_2455,N_2127,N_2208);
xnor U2456 (N_2456,N_1986,N_1636);
and U2457 (N_2457,N_2383,N_1620);
nor U2458 (N_2458,N_2131,N_1999);
or U2459 (N_2459,N_1647,N_2128);
and U2460 (N_2460,N_1947,N_1664);
and U2461 (N_2461,N_1948,N_1725);
and U2462 (N_2462,N_1981,N_2384);
nand U2463 (N_2463,N_2245,N_2390);
and U2464 (N_2464,N_1615,N_1782);
and U2465 (N_2465,N_1685,N_1855);
and U2466 (N_2466,N_2392,N_1718);
xnor U2467 (N_2467,N_2020,N_1752);
and U2468 (N_2468,N_2025,N_1604);
or U2469 (N_2469,N_2181,N_2227);
nor U2470 (N_2470,N_1987,N_1975);
xnor U2471 (N_2471,N_2187,N_2028);
or U2472 (N_2472,N_2339,N_2048);
nand U2473 (N_2473,N_1819,N_2029);
and U2474 (N_2474,N_2331,N_1988);
or U2475 (N_2475,N_1747,N_1640);
nand U2476 (N_2476,N_2169,N_1787);
nor U2477 (N_2477,N_2257,N_1870);
xor U2478 (N_2478,N_2240,N_2049);
or U2479 (N_2479,N_2051,N_2362);
nor U2480 (N_2480,N_1861,N_2250);
or U2481 (N_2481,N_2102,N_2355);
or U2482 (N_2482,N_1940,N_2171);
nor U2483 (N_2483,N_2077,N_1923);
nor U2484 (N_2484,N_2328,N_2189);
nor U2485 (N_2485,N_2090,N_1963);
and U2486 (N_2486,N_1834,N_1889);
xor U2487 (N_2487,N_1868,N_2194);
or U2488 (N_2488,N_2203,N_2068);
nor U2489 (N_2489,N_2018,N_2166);
nand U2490 (N_2490,N_1880,N_2023);
and U2491 (N_2491,N_2150,N_2164);
xor U2492 (N_2492,N_1694,N_1723);
or U2493 (N_2493,N_2170,N_1613);
nor U2494 (N_2494,N_2146,N_1836);
nand U2495 (N_2495,N_2089,N_1901);
or U2496 (N_2496,N_1816,N_2108);
nand U2497 (N_2497,N_2199,N_2366);
xor U2498 (N_2498,N_2263,N_2239);
and U2499 (N_2499,N_1890,N_1629);
or U2500 (N_2500,N_1793,N_2137);
nand U2501 (N_2501,N_1864,N_1601);
nand U2502 (N_2502,N_2314,N_1839);
nor U2503 (N_2503,N_2352,N_1971);
and U2504 (N_2504,N_2009,N_2071);
nor U2505 (N_2505,N_2341,N_1892);
xor U2506 (N_2506,N_1771,N_2145);
or U2507 (N_2507,N_1713,N_1851);
and U2508 (N_2508,N_2324,N_2144);
or U2509 (N_2509,N_1728,N_1683);
xnor U2510 (N_2510,N_1922,N_1727);
and U2511 (N_2511,N_1686,N_2095);
nand U2512 (N_2512,N_2232,N_2276);
or U2513 (N_2513,N_2299,N_2300);
and U2514 (N_2514,N_2041,N_1966);
xnor U2515 (N_2515,N_2243,N_2210);
xnor U2516 (N_2516,N_1663,N_2104);
and U2517 (N_2517,N_2043,N_1693);
and U2518 (N_2518,N_1821,N_2292);
or U2519 (N_2519,N_2101,N_2114);
and U2520 (N_2520,N_1802,N_2265);
or U2521 (N_2521,N_2160,N_2225);
nor U2522 (N_2522,N_2230,N_1773);
or U2523 (N_2523,N_1765,N_2219);
or U2524 (N_2524,N_2159,N_2209);
and U2525 (N_2525,N_2057,N_1885);
nand U2526 (N_2526,N_1635,N_2360);
nor U2527 (N_2527,N_1682,N_1886);
nor U2528 (N_2528,N_2019,N_1676);
nand U2529 (N_2529,N_2030,N_2335);
nor U2530 (N_2530,N_1630,N_1933);
nor U2531 (N_2531,N_2058,N_1837);
xor U2532 (N_2532,N_1667,N_2363);
or U2533 (N_2533,N_2258,N_1825);
xor U2534 (N_2534,N_1627,N_1884);
or U2535 (N_2535,N_1639,N_2103);
and U2536 (N_2536,N_1746,N_2218);
nor U2537 (N_2537,N_2066,N_1603);
nand U2538 (N_2538,N_1779,N_1806);
xnor U2539 (N_2539,N_2307,N_1824);
nor U2540 (N_2540,N_2388,N_1945);
xnor U2541 (N_2541,N_2247,N_1607);
nor U2542 (N_2542,N_2361,N_1659);
and U2543 (N_2543,N_1737,N_1753);
xor U2544 (N_2544,N_1952,N_2271);
nor U2545 (N_2545,N_2273,N_1929);
nor U2546 (N_2546,N_1934,N_1707);
nand U2547 (N_2547,N_1958,N_1831);
and U2548 (N_2548,N_1849,N_1762);
and U2549 (N_2549,N_2063,N_1874);
nor U2550 (N_2550,N_1982,N_2212);
and U2551 (N_2551,N_1907,N_2075);
and U2552 (N_2552,N_2099,N_2076);
and U2553 (N_2553,N_1788,N_2055);
or U2554 (N_2554,N_2064,N_2214);
xor U2555 (N_2555,N_2138,N_1767);
nor U2556 (N_2556,N_1811,N_1891);
and U2557 (N_2557,N_1876,N_2244);
or U2558 (N_2558,N_1648,N_1888);
nand U2559 (N_2559,N_1721,N_1600);
xor U2560 (N_2560,N_2161,N_1833);
or U2561 (N_2561,N_1990,N_1954);
xor U2562 (N_2562,N_2177,N_2332);
nor U2563 (N_2563,N_1931,N_1881);
xor U2564 (N_2564,N_1785,N_1909);
nor U2565 (N_2565,N_2333,N_1715);
xor U2566 (N_2566,N_1691,N_1968);
nor U2567 (N_2567,N_1916,N_2054);
nor U2568 (N_2568,N_1626,N_1871);
or U2569 (N_2569,N_2316,N_2125);
or U2570 (N_2570,N_1724,N_1791);
nor U2571 (N_2571,N_1742,N_1709);
xnor U2572 (N_2572,N_2040,N_2381);
and U2573 (N_2573,N_2317,N_1736);
nand U2574 (N_2574,N_1985,N_2261);
xor U2575 (N_2575,N_1609,N_1658);
and U2576 (N_2576,N_1859,N_1998);
nand U2577 (N_2577,N_2017,N_2238);
and U2578 (N_2578,N_1937,N_1957);
and U2579 (N_2579,N_1712,N_1757);
and U2580 (N_2580,N_2062,N_2290);
and U2581 (N_2581,N_2183,N_1867);
nand U2582 (N_2582,N_2330,N_1996);
and U2583 (N_2583,N_2178,N_1673);
or U2584 (N_2584,N_2396,N_1956);
nand U2585 (N_2585,N_1687,N_2389);
or U2586 (N_2586,N_1829,N_1672);
and U2587 (N_2587,N_2044,N_1716);
nor U2588 (N_2588,N_1936,N_1729);
or U2589 (N_2589,N_2256,N_1962);
and U2590 (N_2590,N_2031,N_1817);
or U2591 (N_2591,N_1818,N_1717);
nand U2592 (N_2592,N_1862,N_2060);
and U2593 (N_2593,N_2174,N_1848);
nand U2594 (N_2594,N_1989,N_1984);
xnor U2595 (N_2595,N_1894,N_2274);
and U2596 (N_2596,N_1660,N_2291);
nand U2597 (N_2597,N_2375,N_1841);
nor U2598 (N_2598,N_1997,N_2323);
or U2599 (N_2599,N_2312,N_2229);
and U2600 (N_2600,N_1624,N_1628);
or U2601 (N_2601,N_2142,N_1710);
or U2602 (N_2602,N_2329,N_2022);
nand U2603 (N_2603,N_2322,N_1769);
or U2604 (N_2604,N_1761,N_2338);
nor U2605 (N_2605,N_2373,N_2191);
and U2606 (N_2606,N_1801,N_2197);
nor U2607 (N_2607,N_2325,N_1708);
or U2608 (N_2608,N_1965,N_1790);
nor U2609 (N_2609,N_1610,N_2012);
or U2610 (N_2610,N_1704,N_1656);
xnor U2611 (N_2611,N_2358,N_1838);
xor U2612 (N_2612,N_2369,N_2357);
xnor U2613 (N_2613,N_1780,N_1668);
nor U2614 (N_2614,N_2205,N_1775);
and U2615 (N_2615,N_1741,N_1680);
and U2616 (N_2616,N_2069,N_1622);
nor U2617 (N_2617,N_2254,N_2217);
and U2618 (N_2618,N_1914,N_1960);
or U2619 (N_2619,N_2248,N_1665);
nor U2620 (N_2620,N_1732,N_1827);
xnor U2621 (N_2621,N_2167,N_2287);
and U2622 (N_2622,N_1808,N_2356);
nand U2623 (N_2623,N_1722,N_1804);
nand U2624 (N_2624,N_1674,N_2182);
nand U2625 (N_2625,N_1699,N_1642);
nor U2626 (N_2626,N_2306,N_2120);
nor U2627 (N_2627,N_2074,N_1842);
xor U2628 (N_2628,N_2113,N_2368);
nor U2629 (N_2629,N_2215,N_2139);
and U2630 (N_2630,N_2147,N_1797);
xor U2631 (N_2631,N_1877,N_2386);
nand U2632 (N_2632,N_2050,N_2267);
xor U2633 (N_2633,N_1634,N_1959);
nand U2634 (N_2634,N_1772,N_1678);
and U2635 (N_2635,N_1655,N_2080);
nand U2636 (N_2636,N_2284,N_1768);
nor U2637 (N_2637,N_2295,N_2059);
xor U2638 (N_2638,N_1835,N_2013);
or U2639 (N_2639,N_1856,N_2294);
xnor U2640 (N_2640,N_2269,N_2141);
xnor U2641 (N_2641,N_2000,N_2350);
nor U2642 (N_2642,N_1843,N_2085);
xnor U2643 (N_2643,N_2015,N_1612);
nand U2644 (N_2644,N_1795,N_1684);
xnor U2645 (N_2645,N_1930,N_1743);
or U2646 (N_2646,N_2107,N_1763);
nor U2647 (N_2647,N_1706,N_1800);
xnor U2648 (N_2648,N_1897,N_2151);
or U2649 (N_2649,N_1681,N_2045);
or U2650 (N_2650,N_2288,N_2078);
and U2651 (N_2651,N_2318,N_1813);
and U2652 (N_2652,N_2135,N_2279);
or U2653 (N_2653,N_2336,N_2228);
and U2654 (N_2654,N_2188,N_1695);
nand U2655 (N_2655,N_2024,N_2393);
nand U2656 (N_2656,N_1866,N_1619);
nor U2657 (N_2657,N_1738,N_2098);
nand U2658 (N_2658,N_2398,N_2165);
or U2659 (N_2659,N_2173,N_2106);
nor U2660 (N_2660,N_2129,N_1766);
xnor U2661 (N_2661,N_1776,N_1616);
nand U2662 (N_2662,N_2268,N_2136);
nor U2663 (N_2663,N_1651,N_1726);
nand U2664 (N_2664,N_2100,N_2349);
nand U2665 (N_2665,N_2305,N_1904);
and U2666 (N_2666,N_1670,N_2072);
nand U2667 (N_2667,N_2180,N_2004);
xnor U2668 (N_2668,N_2037,N_1714);
and U2669 (N_2669,N_1703,N_2124);
nor U2670 (N_2670,N_1799,N_1943);
nor U2671 (N_2671,N_2119,N_1820);
or U2672 (N_2672,N_2032,N_1992);
nand U2673 (N_2673,N_1944,N_2285);
or U2674 (N_2674,N_2374,N_2011);
nor U2675 (N_2675,N_1882,N_2380);
xor U2676 (N_2676,N_2092,N_2289);
xor U2677 (N_2677,N_1754,N_1917);
xor U2678 (N_2678,N_2234,N_2091);
nand U2679 (N_2679,N_1847,N_1852);
nor U2680 (N_2680,N_1978,N_1860);
or U2681 (N_2681,N_1720,N_1650);
or U2682 (N_2682,N_2118,N_1784);
xnor U2683 (N_2683,N_2241,N_1883);
nand U2684 (N_2684,N_1657,N_2053);
or U2685 (N_2685,N_2354,N_1617);
or U2686 (N_2686,N_2334,N_2158);
xor U2687 (N_2687,N_2094,N_1803);
and U2688 (N_2688,N_2175,N_2367);
nand U2689 (N_2689,N_1910,N_1643);
or U2690 (N_2690,N_1970,N_2378);
nor U2691 (N_2691,N_2346,N_1918);
and U2692 (N_2692,N_2036,N_2249);
and U2693 (N_2693,N_1750,N_1733);
xor U2694 (N_2694,N_1781,N_2233);
and U2695 (N_2695,N_2277,N_1995);
and U2696 (N_2696,N_2348,N_1915);
nand U2697 (N_2697,N_1872,N_2109);
and U2698 (N_2698,N_1913,N_2149);
xnor U2699 (N_2699,N_2133,N_2190);
or U2700 (N_2700,N_1637,N_2286);
xnor U2701 (N_2701,N_2185,N_1809);
xnor U2702 (N_2702,N_2035,N_1807);
nand U2703 (N_2703,N_1734,N_2005);
xnor U2704 (N_2704,N_1938,N_1961);
xor U2705 (N_2705,N_1896,N_2395);
and U2706 (N_2706,N_2253,N_1759);
nor U2707 (N_2707,N_1873,N_2067);
nor U2708 (N_2708,N_2251,N_1828);
nor U2709 (N_2709,N_2340,N_1701);
and U2710 (N_2710,N_1879,N_2260);
nor U2711 (N_2711,N_2179,N_1950);
xor U2712 (N_2712,N_1688,N_2313);
nand U2713 (N_2713,N_1869,N_2168);
xnor U2714 (N_2714,N_2387,N_1810);
xnor U2715 (N_2715,N_1755,N_1675);
and U2716 (N_2716,N_1967,N_2278);
xor U2717 (N_2717,N_1854,N_2010);
nand U2718 (N_2718,N_1745,N_1903);
xnor U2719 (N_2719,N_2255,N_1875);
nand U2720 (N_2720,N_2224,N_1798);
xnor U2721 (N_2721,N_2204,N_2132);
xnor U2722 (N_2722,N_1823,N_2042);
nand U2723 (N_2723,N_2105,N_2216);
nor U2724 (N_2724,N_2281,N_1921);
xnor U2725 (N_2725,N_1792,N_1740);
or U2726 (N_2726,N_1621,N_2246);
or U2727 (N_2727,N_1702,N_1994);
xor U2728 (N_2728,N_1625,N_1932);
xnor U2729 (N_2729,N_1760,N_2344);
and U2730 (N_2730,N_2155,N_1902);
or U2731 (N_2731,N_1633,N_2293);
and U2732 (N_2732,N_1623,N_1972);
nand U2733 (N_2733,N_1928,N_2117);
nand U2734 (N_2734,N_2266,N_2319);
or U2735 (N_2735,N_1863,N_1805);
nor U2736 (N_2736,N_2088,N_1920);
nand U2737 (N_2737,N_2351,N_1631);
nand U2738 (N_2738,N_1857,N_1964);
nor U2739 (N_2739,N_1974,N_1711);
xnor U2740 (N_2740,N_1649,N_2084);
or U2741 (N_2741,N_1749,N_2065);
and U2742 (N_2742,N_1976,N_2143);
or U2743 (N_2743,N_1946,N_2365);
nor U2744 (N_2744,N_2093,N_1941);
nor U2745 (N_2745,N_1789,N_1751);
and U2746 (N_2746,N_2122,N_2007);
or U2747 (N_2747,N_1878,N_1690);
nand U2748 (N_2748,N_1608,N_2282);
nand U2749 (N_2749,N_1705,N_2047);
nand U2750 (N_2750,N_2280,N_1698);
nor U2751 (N_2751,N_2235,N_1666);
and U2752 (N_2752,N_2376,N_2311);
and U2753 (N_2753,N_2321,N_2153);
nor U2754 (N_2754,N_1744,N_2226);
xor U2755 (N_2755,N_2342,N_1796);
or U2756 (N_2756,N_1602,N_2082);
and U2757 (N_2757,N_1653,N_2026);
and U2758 (N_2758,N_1942,N_1689);
nor U2759 (N_2759,N_1662,N_1641);
or U2760 (N_2760,N_2223,N_2073);
nor U2761 (N_2761,N_1758,N_1731);
xnor U2762 (N_2762,N_2382,N_2079);
xor U2763 (N_2763,N_1893,N_1927);
xor U2764 (N_2764,N_1898,N_2213);
nand U2765 (N_2765,N_2039,N_2231);
and U2766 (N_2766,N_2154,N_1692);
nor U2767 (N_2767,N_1764,N_2157);
or U2768 (N_2768,N_2196,N_1844);
nor U2769 (N_2769,N_2038,N_2327);
xor U2770 (N_2770,N_1969,N_2021);
nand U2771 (N_2771,N_1815,N_2070);
and U2772 (N_2772,N_1973,N_2096);
nand U2773 (N_2773,N_2347,N_1822);
or U2774 (N_2774,N_1953,N_2003);
and U2775 (N_2775,N_2377,N_2034);
nor U2776 (N_2776,N_2343,N_2202);
xor U2777 (N_2777,N_1900,N_2193);
nand U2778 (N_2778,N_2201,N_2126);
nor U2779 (N_2779,N_2359,N_2134);
nand U2780 (N_2780,N_2301,N_1783);
and U2781 (N_2781,N_1756,N_2086);
or U2782 (N_2782,N_2207,N_1899);
and U2783 (N_2783,N_1814,N_2198);
nor U2784 (N_2784,N_1912,N_1911);
or U2785 (N_2785,N_2111,N_2391);
or U2786 (N_2786,N_2252,N_1794);
and U2787 (N_2787,N_1652,N_2296);
nor U2788 (N_2788,N_2379,N_2056);
and U2789 (N_2789,N_1618,N_2016);
nor U2790 (N_2790,N_1654,N_1979);
or U2791 (N_2791,N_2221,N_2186);
nand U2792 (N_2792,N_2163,N_2083);
or U2793 (N_2793,N_1846,N_1840);
or U2794 (N_2794,N_1939,N_2262);
nor U2795 (N_2795,N_1845,N_2152);
nand U2796 (N_2796,N_1679,N_2270);
nand U2797 (N_2797,N_2121,N_2275);
or U2798 (N_2798,N_2116,N_1748);
nor U2799 (N_2799,N_2222,N_2097);
and U2800 (N_2800,N_1804,N_2119);
or U2801 (N_2801,N_2258,N_1840);
nand U2802 (N_2802,N_1977,N_2185);
nor U2803 (N_2803,N_1696,N_2281);
xor U2804 (N_2804,N_2349,N_2074);
nand U2805 (N_2805,N_1925,N_2317);
or U2806 (N_2806,N_2318,N_1986);
nand U2807 (N_2807,N_1602,N_1761);
or U2808 (N_2808,N_1802,N_1809);
and U2809 (N_2809,N_2320,N_1778);
nand U2810 (N_2810,N_2014,N_2021);
and U2811 (N_2811,N_1973,N_2229);
nand U2812 (N_2812,N_2132,N_2279);
or U2813 (N_2813,N_2018,N_1943);
nand U2814 (N_2814,N_1943,N_2172);
or U2815 (N_2815,N_2290,N_1966);
or U2816 (N_2816,N_2064,N_1703);
nand U2817 (N_2817,N_2225,N_1785);
or U2818 (N_2818,N_1921,N_1714);
and U2819 (N_2819,N_1703,N_1765);
xor U2820 (N_2820,N_2188,N_2131);
nor U2821 (N_2821,N_2339,N_1961);
xnor U2822 (N_2822,N_2285,N_2343);
nor U2823 (N_2823,N_2207,N_1763);
and U2824 (N_2824,N_1610,N_2266);
nand U2825 (N_2825,N_2357,N_1942);
or U2826 (N_2826,N_1663,N_2163);
xor U2827 (N_2827,N_1811,N_1821);
xnor U2828 (N_2828,N_2178,N_1670);
xnor U2829 (N_2829,N_2052,N_2123);
nor U2830 (N_2830,N_1796,N_1666);
or U2831 (N_2831,N_2258,N_2348);
nor U2832 (N_2832,N_2362,N_2332);
or U2833 (N_2833,N_2038,N_1807);
and U2834 (N_2834,N_1832,N_1941);
xnor U2835 (N_2835,N_2174,N_1994);
nand U2836 (N_2836,N_2227,N_1804);
nor U2837 (N_2837,N_1678,N_2115);
and U2838 (N_2838,N_2005,N_2215);
nor U2839 (N_2839,N_2369,N_2330);
nor U2840 (N_2840,N_2219,N_1881);
or U2841 (N_2841,N_1822,N_2284);
nand U2842 (N_2842,N_2295,N_2368);
nor U2843 (N_2843,N_2118,N_1851);
and U2844 (N_2844,N_1957,N_1698);
nand U2845 (N_2845,N_2032,N_1719);
or U2846 (N_2846,N_1715,N_1614);
nor U2847 (N_2847,N_2042,N_1735);
or U2848 (N_2848,N_1732,N_1770);
or U2849 (N_2849,N_2060,N_2068);
and U2850 (N_2850,N_2030,N_2258);
and U2851 (N_2851,N_1909,N_1726);
and U2852 (N_2852,N_2053,N_2356);
and U2853 (N_2853,N_2271,N_1649);
xor U2854 (N_2854,N_1964,N_2232);
nor U2855 (N_2855,N_1626,N_2163);
or U2856 (N_2856,N_2047,N_2165);
nand U2857 (N_2857,N_1932,N_1720);
and U2858 (N_2858,N_2271,N_2178);
nand U2859 (N_2859,N_1948,N_1954);
or U2860 (N_2860,N_2236,N_2228);
xor U2861 (N_2861,N_2021,N_2277);
nand U2862 (N_2862,N_2324,N_1792);
xor U2863 (N_2863,N_2305,N_1890);
nor U2864 (N_2864,N_1952,N_2004);
nand U2865 (N_2865,N_2019,N_1681);
or U2866 (N_2866,N_2288,N_1627);
nor U2867 (N_2867,N_1722,N_1811);
nor U2868 (N_2868,N_2060,N_1907);
xor U2869 (N_2869,N_1777,N_2386);
and U2870 (N_2870,N_2004,N_1613);
nor U2871 (N_2871,N_1840,N_1856);
and U2872 (N_2872,N_1692,N_2317);
and U2873 (N_2873,N_1986,N_2142);
or U2874 (N_2874,N_2279,N_2294);
nor U2875 (N_2875,N_2200,N_1931);
or U2876 (N_2876,N_2039,N_2328);
nand U2877 (N_2877,N_1802,N_1688);
xnor U2878 (N_2878,N_2121,N_1969);
nor U2879 (N_2879,N_1979,N_1789);
xor U2880 (N_2880,N_2076,N_2024);
or U2881 (N_2881,N_2098,N_2077);
or U2882 (N_2882,N_2313,N_2225);
nand U2883 (N_2883,N_2314,N_1866);
or U2884 (N_2884,N_1945,N_1698);
or U2885 (N_2885,N_2371,N_1778);
xnor U2886 (N_2886,N_1617,N_2116);
nand U2887 (N_2887,N_1950,N_1642);
nor U2888 (N_2888,N_2011,N_1966);
xnor U2889 (N_2889,N_2220,N_2062);
and U2890 (N_2890,N_1712,N_2069);
nand U2891 (N_2891,N_2240,N_2343);
xor U2892 (N_2892,N_2180,N_1603);
nand U2893 (N_2893,N_2113,N_2248);
nor U2894 (N_2894,N_1625,N_2204);
and U2895 (N_2895,N_2096,N_1649);
or U2896 (N_2896,N_2051,N_1721);
nand U2897 (N_2897,N_1797,N_1835);
xnor U2898 (N_2898,N_1707,N_1826);
or U2899 (N_2899,N_2307,N_2298);
xor U2900 (N_2900,N_1946,N_1608);
xor U2901 (N_2901,N_1964,N_2192);
nor U2902 (N_2902,N_1685,N_2354);
nand U2903 (N_2903,N_1689,N_2203);
nor U2904 (N_2904,N_2183,N_2315);
nor U2905 (N_2905,N_1726,N_2050);
nor U2906 (N_2906,N_2046,N_2050);
nand U2907 (N_2907,N_2149,N_2329);
or U2908 (N_2908,N_1644,N_2221);
and U2909 (N_2909,N_1865,N_1816);
xor U2910 (N_2910,N_1951,N_2281);
nand U2911 (N_2911,N_1671,N_1961);
nor U2912 (N_2912,N_2148,N_1673);
and U2913 (N_2913,N_2028,N_1618);
and U2914 (N_2914,N_2334,N_1661);
nand U2915 (N_2915,N_1738,N_1959);
nand U2916 (N_2916,N_1967,N_2009);
nand U2917 (N_2917,N_1999,N_2284);
and U2918 (N_2918,N_1818,N_1702);
and U2919 (N_2919,N_2142,N_1686);
or U2920 (N_2920,N_1629,N_2382);
xnor U2921 (N_2921,N_2141,N_2088);
nand U2922 (N_2922,N_2024,N_1733);
or U2923 (N_2923,N_2163,N_2099);
nand U2924 (N_2924,N_2027,N_1798);
xnor U2925 (N_2925,N_1955,N_2251);
and U2926 (N_2926,N_1910,N_2014);
nand U2927 (N_2927,N_2318,N_2074);
and U2928 (N_2928,N_1822,N_2242);
nand U2929 (N_2929,N_2287,N_2332);
and U2930 (N_2930,N_2386,N_2065);
or U2931 (N_2931,N_1682,N_2249);
or U2932 (N_2932,N_1895,N_2228);
nand U2933 (N_2933,N_1841,N_2056);
nor U2934 (N_2934,N_2126,N_2345);
nand U2935 (N_2935,N_1927,N_2000);
xor U2936 (N_2936,N_2168,N_1696);
nand U2937 (N_2937,N_1787,N_2166);
and U2938 (N_2938,N_2316,N_2149);
nand U2939 (N_2939,N_1765,N_1613);
or U2940 (N_2940,N_1695,N_1953);
nor U2941 (N_2941,N_1988,N_1709);
xnor U2942 (N_2942,N_1745,N_2058);
xor U2943 (N_2943,N_1920,N_2033);
or U2944 (N_2944,N_1958,N_2041);
xnor U2945 (N_2945,N_2342,N_1803);
nand U2946 (N_2946,N_2235,N_1761);
nor U2947 (N_2947,N_1923,N_2240);
xnor U2948 (N_2948,N_1687,N_2061);
or U2949 (N_2949,N_1990,N_1832);
or U2950 (N_2950,N_2355,N_1673);
and U2951 (N_2951,N_2349,N_2344);
and U2952 (N_2952,N_1606,N_2098);
or U2953 (N_2953,N_2176,N_1841);
and U2954 (N_2954,N_2268,N_2365);
and U2955 (N_2955,N_1611,N_1898);
nor U2956 (N_2956,N_2093,N_1844);
and U2957 (N_2957,N_1737,N_2186);
and U2958 (N_2958,N_1672,N_1770);
and U2959 (N_2959,N_1998,N_2217);
nand U2960 (N_2960,N_2178,N_1811);
and U2961 (N_2961,N_1912,N_1864);
nor U2962 (N_2962,N_2243,N_1985);
and U2963 (N_2963,N_2107,N_2226);
or U2964 (N_2964,N_2031,N_1803);
xor U2965 (N_2965,N_2323,N_1831);
and U2966 (N_2966,N_1787,N_2283);
nor U2967 (N_2967,N_1786,N_2294);
and U2968 (N_2968,N_2013,N_2294);
and U2969 (N_2969,N_1702,N_1883);
or U2970 (N_2970,N_2206,N_1719);
and U2971 (N_2971,N_1600,N_1718);
nor U2972 (N_2972,N_2095,N_1602);
xor U2973 (N_2973,N_2015,N_1767);
and U2974 (N_2974,N_2269,N_2013);
and U2975 (N_2975,N_2283,N_1890);
or U2976 (N_2976,N_1654,N_2338);
or U2977 (N_2977,N_1741,N_2281);
xnor U2978 (N_2978,N_2003,N_1704);
xnor U2979 (N_2979,N_1620,N_2223);
and U2980 (N_2980,N_1729,N_1906);
and U2981 (N_2981,N_1690,N_2106);
nor U2982 (N_2982,N_1794,N_1971);
and U2983 (N_2983,N_1872,N_2183);
xor U2984 (N_2984,N_2304,N_2106);
or U2985 (N_2985,N_1965,N_1972);
xor U2986 (N_2986,N_1740,N_1652);
nor U2987 (N_2987,N_2144,N_1643);
or U2988 (N_2988,N_2317,N_1972);
nor U2989 (N_2989,N_2353,N_2091);
nand U2990 (N_2990,N_1651,N_2366);
nand U2991 (N_2991,N_1601,N_2114);
nor U2992 (N_2992,N_2105,N_2223);
and U2993 (N_2993,N_1793,N_1763);
nor U2994 (N_2994,N_1651,N_2227);
xor U2995 (N_2995,N_1876,N_1912);
xnor U2996 (N_2996,N_1686,N_2211);
nor U2997 (N_2997,N_2057,N_2168);
and U2998 (N_2998,N_2002,N_2167);
and U2999 (N_2999,N_1930,N_1750);
and U3000 (N_3000,N_1714,N_2340);
nor U3001 (N_3001,N_2073,N_1607);
nor U3002 (N_3002,N_1691,N_1829);
xnor U3003 (N_3003,N_1686,N_2094);
and U3004 (N_3004,N_2273,N_1790);
xnor U3005 (N_3005,N_1832,N_2141);
nand U3006 (N_3006,N_2372,N_2377);
and U3007 (N_3007,N_2322,N_1659);
nor U3008 (N_3008,N_1985,N_1786);
nand U3009 (N_3009,N_1640,N_1663);
and U3010 (N_3010,N_1725,N_1912);
nand U3011 (N_3011,N_2107,N_1768);
nand U3012 (N_3012,N_2229,N_1671);
nand U3013 (N_3013,N_2334,N_1856);
nand U3014 (N_3014,N_2109,N_2245);
and U3015 (N_3015,N_2334,N_2118);
nand U3016 (N_3016,N_1718,N_2016);
nand U3017 (N_3017,N_2349,N_2018);
nor U3018 (N_3018,N_2384,N_1988);
or U3019 (N_3019,N_2134,N_2271);
or U3020 (N_3020,N_1791,N_1721);
nor U3021 (N_3021,N_2218,N_2350);
nor U3022 (N_3022,N_1605,N_1994);
nor U3023 (N_3023,N_2266,N_2165);
xor U3024 (N_3024,N_1776,N_2205);
nor U3025 (N_3025,N_2230,N_1808);
xnor U3026 (N_3026,N_1661,N_1739);
xnor U3027 (N_3027,N_2296,N_2055);
xor U3028 (N_3028,N_1908,N_2092);
or U3029 (N_3029,N_2192,N_1778);
nor U3030 (N_3030,N_2261,N_2308);
and U3031 (N_3031,N_2114,N_1691);
nor U3032 (N_3032,N_2370,N_2078);
nand U3033 (N_3033,N_1956,N_1943);
nor U3034 (N_3034,N_1879,N_2033);
nor U3035 (N_3035,N_2113,N_1813);
or U3036 (N_3036,N_2240,N_2133);
or U3037 (N_3037,N_1731,N_2304);
xnor U3038 (N_3038,N_2267,N_2045);
and U3039 (N_3039,N_2156,N_2287);
nand U3040 (N_3040,N_2356,N_2276);
xor U3041 (N_3041,N_1824,N_2216);
or U3042 (N_3042,N_2244,N_1629);
and U3043 (N_3043,N_1980,N_2350);
nor U3044 (N_3044,N_2399,N_1616);
and U3045 (N_3045,N_2164,N_1884);
and U3046 (N_3046,N_1744,N_2011);
and U3047 (N_3047,N_1865,N_2071);
nand U3048 (N_3048,N_2108,N_2269);
xor U3049 (N_3049,N_1899,N_1950);
xnor U3050 (N_3050,N_2213,N_1919);
and U3051 (N_3051,N_2264,N_2254);
nand U3052 (N_3052,N_2355,N_1828);
nand U3053 (N_3053,N_2295,N_2279);
nand U3054 (N_3054,N_2156,N_1842);
xnor U3055 (N_3055,N_2371,N_1851);
or U3056 (N_3056,N_2296,N_2212);
nand U3057 (N_3057,N_2140,N_1892);
xor U3058 (N_3058,N_2322,N_1753);
nor U3059 (N_3059,N_2116,N_1742);
nor U3060 (N_3060,N_1705,N_2249);
xnor U3061 (N_3061,N_2234,N_2192);
nor U3062 (N_3062,N_2001,N_2217);
nand U3063 (N_3063,N_2099,N_1640);
xor U3064 (N_3064,N_2258,N_1805);
xor U3065 (N_3065,N_2036,N_1729);
or U3066 (N_3066,N_1966,N_1731);
xor U3067 (N_3067,N_2228,N_2381);
nand U3068 (N_3068,N_2340,N_1773);
nor U3069 (N_3069,N_1875,N_2197);
or U3070 (N_3070,N_1607,N_1687);
or U3071 (N_3071,N_1670,N_1690);
or U3072 (N_3072,N_1989,N_1867);
nor U3073 (N_3073,N_1972,N_1712);
or U3074 (N_3074,N_1842,N_1864);
or U3075 (N_3075,N_1807,N_2338);
or U3076 (N_3076,N_1856,N_1801);
or U3077 (N_3077,N_2178,N_1950);
nor U3078 (N_3078,N_2242,N_2045);
or U3079 (N_3079,N_1696,N_2354);
nand U3080 (N_3080,N_2026,N_2174);
or U3081 (N_3081,N_1855,N_1818);
or U3082 (N_3082,N_1991,N_2073);
and U3083 (N_3083,N_1917,N_1704);
and U3084 (N_3084,N_1775,N_2181);
nor U3085 (N_3085,N_2161,N_2324);
or U3086 (N_3086,N_1794,N_1758);
or U3087 (N_3087,N_1856,N_2142);
xor U3088 (N_3088,N_2283,N_1919);
nand U3089 (N_3089,N_2234,N_2283);
or U3090 (N_3090,N_2266,N_1807);
or U3091 (N_3091,N_1645,N_1718);
xnor U3092 (N_3092,N_1779,N_1642);
and U3093 (N_3093,N_1632,N_2132);
nand U3094 (N_3094,N_2264,N_1848);
and U3095 (N_3095,N_1807,N_1774);
nand U3096 (N_3096,N_2228,N_2253);
or U3097 (N_3097,N_2373,N_2098);
or U3098 (N_3098,N_1919,N_1800);
nand U3099 (N_3099,N_1883,N_1954);
xor U3100 (N_3100,N_1665,N_2008);
or U3101 (N_3101,N_1880,N_1796);
nand U3102 (N_3102,N_2270,N_2353);
nand U3103 (N_3103,N_2355,N_1741);
or U3104 (N_3104,N_1876,N_1610);
and U3105 (N_3105,N_2342,N_2393);
or U3106 (N_3106,N_2040,N_1696);
and U3107 (N_3107,N_1751,N_1961);
and U3108 (N_3108,N_1719,N_2023);
xor U3109 (N_3109,N_2091,N_1849);
nor U3110 (N_3110,N_2244,N_2291);
nor U3111 (N_3111,N_2156,N_1671);
nand U3112 (N_3112,N_2375,N_1670);
or U3113 (N_3113,N_2256,N_2131);
nor U3114 (N_3114,N_2037,N_2372);
xnor U3115 (N_3115,N_2155,N_2188);
xor U3116 (N_3116,N_1707,N_2340);
nor U3117 (N_3117,N_1730,N_2086);
or U3118 (N_3118,N_1898,N_1989);
or U3119 (N_3119,N_1671,N_2340);
or U3120 (N_3120,N_2036,N_1912);
or U3121 (N_3121,N_1659,N_2265);
xor U3122 (N_3122,N_2128,N_1933);
xnor U3123 (N_3123,N_2197,N_1929);
xor U3124 (N_3124,N_2349,N_1714);
nor U3125 (N_3125,N_1708,N_2394);
nor U3126 (N_3126,N_2242,N_2333);
or U3127 (N_3127,N_2183,N_2247);
nor U3128 (N_3128,N_1903,N_1841);
nand U3129 (N_3129,N_1796,N_2268);
xnor U3130 (N_3130,N_2327,N_1784);
nand U3131 (N_3131,N_1805,N_1990);
and U3132 (N_3132,N_1796,N_2142);
nand U3133 (N_3133,N_2028,N_1729);
or U3134 (N_3134,N_2235,N_2296);
xnor U3135 (N_3135,N_2255,N_2357);
and U3136 (N_3136,N_1935,N_1615);
or U3137 (N_3137,N_2255,N_1986);
and U3138 (N_3138,N_2291,N_1825);
nor U3139 (N_3139,N_2153,N_2178);
or U3140 (N_3140,N_1899,N_2302);
or U3141 (N_3141,N_2298,N_2063);
xor U3142 (N_3142,N_2325,N_2097);
xor U3143 (N_3143,N_2043,N_1606);
or U3144 (N_3144,N_1799,N_1845);
nand U3145 (N_3145,N_1649,N_2298);
nand U3146 (N_3146,N_2232,N_2122);
or U3147 (N_3147,N_2392,N_2097);
or U3148 (N_3148,N_1668,N_2311);
xnor U3149 (N_3149,N_2194,N_2277);
or U3150 (N_3150,N_1695,N_2299);
or U3151 (N_3151,N_1717,N_2379);
or U3152 (N_3152,N_1857,N_1863);
or U3153 (N_3153,N_2200,N_1831);
nor U3154 (N_3154,N_2378,N_1944);
nor U3155 (N_3155,N_2309,N_2226);
xnor U3156 (N_3156,N_1943,N_2324);
nand U3157 (N_3157,N_1946,N_2101);
or U3158 (N_3158,N_1937,N_1768);
or U3159 (N_3159,N_2118,N_1887);
xnor U3160 (N_3160,N_1811,N_1707);
nand U3161 (N_3161,N_2184,N_1928);
and U3162 (N_3162,N_2269,N_1803);
nand U3163 (N_3163,N_1811,N_1799);
xor U3164 (N_3164,N_2162,N_2121);
xor U3165 (N_3165,N_1840,N_1690);
xor U3166 (N_3166,N_1745,N_2013);
nand U3167 (N_3167,N_1755,N_1696);
or U3168 (N_3168,N_1682,N_2311);
nor U3169 (N_3169,N_2203,N_2169);
xor U3170 (N_3170,N_1947,N_1795);
nand U3171 (N_3171,N_1762,N_1611);
or U3172 (N_3172,N_2249,N_1732);
nand U3173 (N_3173,N_2338,N_1760);
xnor U3174 (N_3174,N_1969,N_2298);
and U3175 (N_3175,N_2387,N_1610);
xor U3176 (N_3176,N_1992,N_1975);
nand U3177 (N_3177,N_2103,N_2278);
and U3178 (N_3178,N_1689,N_2230);
and U3179 (N_3179,N_2049,N_1628);
xnor U3180 (N_3180,N_1997,N_2143);
nand U3181 (N_3181,N_2296,N_2084);
nand U3182 (N_3182,N_2158,N_1625);
or U3183 (N_3183,N_1672,N_2373);
nor U3184 (N_3184,N_1758,N_1801);
or U3185 (N_3185,N_1656,N_2149);
xor U3186 (N_3186,N_1843,N_2339);
nand U3187 (N_3187,N_2126,N_1833);
nor U3188 (N_3188,N_2348,N_1691);
and U3189 (N_3189,N_1744,N_1774);
xnor U3190 (N_3190,N_2026,N_2305);
xnor U3191 (N_3191,N_1870,N_2045);
xor U3192 (N_3192,N_2226,N_1804);
or U3193 (N_3193,N_1832,N_1979);
and U3194 (N_3194,N_1691,N_2234);
and U3195 (N_3195,N_2131,N_2369);
or U3196 (N_3196,N_1811,N_1744);
nor U3197 (N_3197,N_2167,N_1876);
nand U3198 (N_3198,N_2173,N_1662);
xor U3199 (N_3199,N_1662,N_1906);
xor U3200 (N_3200,N_2492,N_2475);
or U3201 (N_3201,N_2546,N_3026);
nand U3202 (N_3202,N_2667,N_2531);
xor U3203 (N_3203,N_2844,N_3063);
and U3204 (N_3204,N_2505,N_2407);
nor U3205 (N_3205,N_2541,N_3138);
nand U3206 (N_3206,N_2992,N_3035);
xnor U3207 (N_3207,N_2623,N_2597);
and U3208 (N_3208,N_2534,N_2890);
or U3209 (N_3209,N_3060,N_2832);
and U3210 (N_3210,N_2604,N_2983);
nor U3211 (N_3211,N_3185,N_2767);
or U3212 (N_3212,N_2800,N_3127);
and U3213 (N_3213,N_2413,N_3122);
and U3214 (N_3214,N_2588,N_3166);
and U3215 (N_3215,N_2951,N_2509);
nand U3216 (N_3216,N_3095,N_3046);
nor U3217 (N_3217,N_3193,N_2635);
xnor U3218 (N_3218,N_3176,N_2447);
or U3219 (N_3219,N_2609,N_2560);
nand U3220 (N_3220,N_2473,N_2876);
xor U3221 (N_3221,N_2556,N_2640);
or U3222 (N_3222,N_2704,N_2986);
and U3223 (N_3223,N_2611,N_2802);
nand U3224 (N_3224,N_2994,N_2582);
xor U3225 (N_3225,N_2647,N_3098);
or U3226 (N_3226,N_3194,N_2841);
xor U3227 (N_3227,N_3120,N_2639);
or U3228 (N_3228,N_2471,N_3054);
xor U3229 (N_3229,N_2688,N_2727);
nand U3230 (N_3230,N_2420,N_2590);
or U3231 (N_3231,N_3191,N_2772);
or U3232 (N_3232,N_3057,N_2972);
nor U3233 (N_3233,N_3093,N_2621);
and U3234 (N_3234,N_2748,N_3146);
nor U3235 (N_3235,N_2962,N_3023);
xor U3236 (N_3236,N_2622,N_2960);
xnor U3237 (N_3237,N_2861,N_2789);
and U3238 (N_3238,N_3189,N_2400);
or U3239 (N_3239,N_3102,N_2818);
nand U3240 (N_3240,N_3070,N_2725);
xor U3241 (N_3241,N_2872,N_2755);
xor U3242 (N_3242,N_2865,N_2479);
nor U3243 (N_3243,N_2857,N_2858);
nand U3244 (N_3244,N_2425,N_2482);
nor U3245 (N_3245,N_2828,N_2690);
nand U3246 (N_3246,N_2599,N_2576);
and U3247 (N_3247,N_2418,N_2982);
xnor U3248 (N_3248,N_2626,N_2750);
nand U3249 (N_3249,N_2428,N_2721);
and U3250 (N_3250,N_2637,N_3171);
nand U3251 (N_3251,N_2771,N_3075);
xnor U3252 (N_3252,N_2591,N_2764);
nor U3253 (N_3253,N_2412,N_2824);
nor U3254 (N_3254,N_3184,N_2530);
nand U3255 (N_3255,N_2956,N_2804);
nor U3256 (N_3256,N_2419,N_2922);
nor U3257 (N_3257,N_3021,N_3162);
and U3258 (N_3258,N_2592,N_2964);
xnor U3259 (N_3259,N_2881,N_2803);
nor U3260 (N_3260,N_2715,N_3000);
and U3261 (N_3261,N_3016,N_2643);
and U3262 (N_3262,N_2641,N_2692);
nor U3263 (N_3263,N_2543,N_3150);
and U3264 (N_3264,N_3179,N_2866);
xor U3265 (N_3265,N_3029,N_3143);
or U3266 (N_3266,N_3056,N_3073);
xor U3267 (N_3267,N_2459,N_2625);
or U3268 (N_3268,N_2457,N_3108);
or U3269 (N_3269,N_3004,N_2779);
nor U3270 (N_3270,N_2813,N_3113);
and U3271 (N_3271,N_2993,N_2912);
or U3272 (N_3272,N_2869,N_2535);
nand U3273 (N_3273,N_3077,N_3164);
nor U3274 (N_3274,N_2568,N_2694);
xor U3275 (N_3275,N_3148,N_3043);
or U3276 (N_3276,N_2679,N_2987);
xor U3277 (N_3277,N_2415,N_2822);
nor U3278 (N_3278,N_2874,N_3022);
nor U3279 (N_3279,N_2752,N_3099);
or U3280 (N_3280,N_2706,N_3105);
nor U3281 (N_3281,N_3136,N_3066);
nor U3282 (N_3282,N_2761,N_3178);
or U3283 (N_3283,N_2527,N_2657);
nand U3284 (N_3284,N_2746,N_2633);
and U3285 (N_3285,N_2608,N_2500);
or U3286 (N_3286,N_3182,N_2435);
and U3287 (N_3287,N_2718,N_2461);
nor U3288 (N_3288,N_2408,N_3135);
nand U3289 (N_3289,N_2421,N_2554);
nand U3290 (N_3290,N_2511,N_2529);
nor U3291 (N_3291,N_2663,N_2474);
or U3292 (N_3292,N_2636,N_2891);
nand U3293 (N_3293,N_3128,N_2884);
and U3294 (N_3294,N_2953,N_2851);
nor U3295 (N_3295,N_2513,N_2770);
and U3296 (N_3296,N_2871,N_3003);
nor U3297 (N_3297,N_2615,N_3103);
nor U3298 (N_3298,N_2935,N_2579);
or U3299 (N_3299,N_2981,N_2756);
or U3300 (N_3300,N_3180,N_2423);
or U3301 (N_3301,N_2634,N_2807);
xor U3302 (N_3302,N_2754,N_2559);
nor U3303 (N_3303,N_2744,N_2817);
nand U3304 (N_3304,N_3144,N_2409);
or U3305 (N_3305,N_2602,N_2675);
and U3306 (N_3306,N_2632,N_2436);
xor U3307 (N_3307,N_3088,N_2506);
and U3308 (N_3308,N_3078,N_3013);
xor U3309 (N_3309,N_2894,N_2976);
or U3310 (N_3310,N_3030,N_3153);
nand U3311 (N_3311,N_3169,N_2619);
xnor U3312 (N_3312,N_2860,N_3062);
xnor U3313 (N_3313,N_2870,N_2508);
or U3314 (N_3314,N_2658,N_2985);
and U3315 (N_3315,N_3058,N_3042);
xnor U3316 (N_3316,N_2886,N_2426);
or U3317 (N_3317,N_2491,N_2644);
nor U3318 (N_3318,N_3160,N_2587);
or U3319 (N_3319,N_3045,N_2778);
xnor U3320 (N_3320,N_2454,N_2713);
xnor U3321 (N_3321,N_2729,N_2558);
nand U3322 (N_3322,N_2799,N_2489);
nor U3323 (N_3323,N_2946,N_2819);
and U3324 (N_3324,N_3139,N_3133);
nand U3325 (N_3325,N_3151,N_2957);
and U3326 (N_3326,N_2716,N_2443);
and U3327 (N_3327,N_2514,N_3172);
nand U3328 (N_3328,N_3027,N_2664);
nand U3329 (N_3329,N_3094,N_2990);
nor U3330 (N_3330,N_2899,N_2689);
or U3331 (N_3331,N_2855,N_2685);
nor U3332 (N_3332,N_2758,N_2584);
nor U3333 (N_3333,N_2437,N_3118);
and U3334 (N_3334,N_2979,N_3140);
nand U3335 (N_3335,N_2465,N_2785);
nand U3336 (N_3336,N_2434,N_2714);
nor U3337 (N_3337,N_2952,N_2586);
nand U3338 (N_3338,N_2787,N_2494);
and U3339 (N_3339,N_2698,N_2928);
nand U3340 (N_3340,N_2651,N_2565);
or U3341 (N_3341,N_2537,N_2653);
xor U3342 (N_3342,N_3074,N_2888);
nor U3343 (N_3343,N_2901,N_2863);
or U3344 (N_3344,N_3085,N_2549);
and U3345 (N_3345,N_2926,N_3190);
or U3346 (N_3346,N_2835,N_2984);
xor U3347 (N_3347,N_2965,N_2701);
nand U3348 (N_3348,N_2766,N_3147);
xor U3349 (N_3349,N_2788,N_2918);
or U3350 (N_3350,N_2775,N_2797);
and U3351 (N_3351,N_2665,N_2522);
and U3352 (N_3352,N_2652,N_3101);
or U3353 (N_3353,N_2973,N_2924);
nand U3354 (N_3354,N_2441,N_3051);
and U3355 (N_3355,N_2726,N_2904);
xnor U3356 (N_3356,N_3112,N_2743);
or U3357 (N_3357,N_3082,N_2596);
nand U3358 (N_3358,N_2440,N_2416);
or U3359 (N_3359,N_2963,N_3081);
or U3360 (N_3360,N_2673,N_2941);
xor U3361 (N_3361,N_2950,N_2526);
xor U3362 (N_3362,N_2921,N_2453);
xor U3363 (N_3363,N_2896,N_3050);
nand U3364 (N_3364,N_3124,N_2879);
nand U3365 (N_3365,N_2676,N_2575);
nor U3366 (N_3366,N_2859,N_2684);
nand U3367 (N_3367,N_3159,N_3008);
and U3368 (N_3368,N_2790,N_2567);
or U3369 (N_3369,N_2677,N_2936);
nand U3370 (N_3370,N_2815,N_2794);
nand U3371 (N_3371,N_2629,N_2816);
nand U3372 (N_3372,N_3096,N_2784);
xnor U3373 (N_3373,N_2613,N_3107);
xor U3374 (N_3374,N_2949,N_2631);
and U3375 (N_3375,N_2811,N_2867);
xor U3376 (N_3376,N_2929,N_3129);
or U3377 (N_3377,N_3115,N_3020);
and U3378 (N_3378,N_2814,N_2995);
nor U3379 (N_3379,N_2850,N_3131);
and U3380 (N_3380,N_3009,N_3083);
and U3381 (N_3381,N_2538,N_3068);
or U3382 (N_3382,N_3065,N_2791);
nand U3383 (N_3383,N_2833,N_2740);
nand U3384 (N_3384,N_2488,N_2660);
xnor U3385 (N_3385,N_3173,N_3034);
or U3386 (N_3386,N_2915,N_2908);
nor U3387 (N_3387,N_2823,N_2919);
and U3388 (N_3388,N_2438,N_2431);
xor U3389 (N_3389,N_2849,N_2988);
and U3390 (N_3390,N_2838,N_2691);
nand U3391 (N_3391,N_2699,N_3142);
and U3392 (N_3392,N_2997,N_3067);
xnor U3393 (N_3393,N_3123,N_2600);
and U3394 (N_3394,N_3033,N_2540);
and U3395 (N_3395,N_2745,N_3010);
xnor U3396 (N_3396,N_2452,N_3141);
or U3397 (N_3397,N_2809,N_3132);
xnor U3398 (N_3398,N_3186,N_2923);
and U3399 (N_3399,N_2446,N_2996);
or U3400 (N_3400,N_2624,N_2940);
or U3401 (N_3401,N_2810,N_2595);
and U3402 (N_3402,N_2757,N_2769);
nand U3403 (N_3403,N_3007,N_3161);
nand U3404 (N_3404,N_3187,N_2808);
or U3405 (N_3405,N_2659,N_2432);
xnor U3406 (N_3406,N_2502,N_2909);
and U3407 (N_3407,N_3061,N_2448);
nand U3408 (N_3408,N_2966,N_2630);
or U3409 (N_3409,N_2589,N_2547);
nor U3410 (N_3410,N_2478,N_2958);
nor U3411 (N_3411,N_2910,N_2734);
and U3412 (N_3412,N_2759,N_2467);
nand U3413 (N_3413,N_2539,N_2469);
and U3414 (N_3414,N_3199,N_2661);
nor U3415 (N_3415,N_2774,N_2444);
xnor U3416 (N_3416,N_3044,N_2705);
or U3417 (N_3417,N_2551,N_3149);
xnor U3418 (N_3418,N_2895,N_2462);
or U3419 (N_3419,N_2885,N_2710);
and U3420 (N_3420,N_2564,N_2864);
nand U3421 (N_3421,N_2848,N_2401);
nor U3422 (N_3422,N_3174,N_3183);
nand U3423 (N_3423,N_2998,N_2723);
nand U3424 (N_3424,N_3017,N_2424);
nand U3425 (N_3425,N_2920,N_2545);
and U3426 (N_3426,N_2411,N_3158);
xnor U3427 (N_3427,N_2836,N_2902);
nor U3428 (N_3428,N_2528,N_2476);
and U3429 (N_3429,N_2845,N_2460);
or U3430 (N_3430,N_2882,N_2593);
and U3431 (N_3431,N_2627,N_2708);
xor U3432 (N_3432,N_3049,N_2773);
xor U3433 (N_3433,N_2693,N_3137);
nand U3434 (N_3434,N_3084,N_2825);
or U3435 (N_3435,N_2776,N_2763);
or U3436 (N_3436,N_2977,N_2429);
and U3437 (N_3437,N_2617,N_2477);
nand U3438 (N_3438,N_2612,N_2486);
nor U3439 (N_3439,N_2937,N_2472);
nor U3440 (N_3440,N_2702,N_3111);
or U3441 (N_3441,N_2430,N_2762);
and U3442 (N_3442,N_3145,N_2843);
or U3443 (N_3443,N_3039,N_2422);
and U3444 (N_3444,N_2464,N_2515);
or U3445 (N_3445,N_2450,N_2846);
nor U3446 (N_3446,N_2552,N_2854);
and U3447 (N_3447,N_3195,N_2736);
nand U3448 (N_3448,N_2581,N_3126);
xor U3449 (N_3449,N_2711,N_2484);
and U3450 (N_3450,N_3091,N_3177);
xor U3451 (N_3451,N_3117,N_3019);
and U3452 (N_3452,N_3188,N_2830);
nand U3453 (N_3453,N_3104,N_3163);
and U3454 (N_3454,N_2820,N_2405);
nor U3455 (N_3455,N_2806,N_2497);
nor U3456 (N_3456,N_2686,N_3196);
xor U3457 (N_3457,N_3167,N_2842);
or U3458 (N_3458,N_2406,N_2577);
and U3459 (N_3459,N_2512,N_2483);
and U3460 (N_3460,N_2897,N_2974);
xnor U3461 (N_3461,N_2955,N_2672);
nor U3462 (N_3462,N_2470,N_2433);
nor U3463 (N_3463,N_2839,N_2829);
xnor U3464 (N_3464,N_2468,N_2533);
and U3465 (N_3465,N_3125,N_3018);
nor U3466 (N_3466,N_2670,N_2521);
or U3467 (N_3467,N_2827,N_2603);
nand U3468 (N_3468,N_2649,N_2606);
nand U3469 (N_3469,N_3048,N_2945);
nand U3470 (N_3470,N_2707,N_2703);
nand U3471 (N_3471,N_2738,N_2666);
nor U3472 (N_3472,N_2975,N_2504);
and U3473 (N_3473,N_2485,N_2944);
xor U3474 (N_3474,N_2735,N_2751);
nor U3475 (N_3475,N_2445,N_2410);
or U3476 (N_3476,N_2455,N_2959);
nand U3477 (N_3477,N_2898,N_2796);
nor U3478 (N_3478,N_2566,N_3031);
xnor U3479 (N_3479,N_2645,N_3079);
and U3480 (N_3480,N_2449,N_2680);
xnor U3481 (N_3481,N_2907,N_2496);
or U3482 (N_3482,N_3092,N_3152);
xnor U3483 (N_3483,N_2939,N_2490);
nand U3484 (N_3484,N_2557,N_2662);
or U3485 (N_3485,N_2930,N_2903);
and U3486 (N_3486,N_3100,N_2989);
and U3487 (N_3487,N_2831,N_2925);
nor U3488 (N_3488,N_2519,N_2916);
nor U3489 (N_3489,N_2906,N_2553);
and U3490 (N_3490,N_2700,N_2697);
nor U3491 (N_3491,N_2954,N_2875);
nand U3492 (N_3492,N_2463,N_2525);
and U3493 (N_3493,N_2427,N_2610);
xnor U3494 (N_3494,N_2948,N_2742);
and U3495 (N_3495,N_2487,N_2536);
and U3496 (N_3496,N_3170,N_2532);
nand U3497 (N_3497,N_2722,N_2968);
and U3498 (N_3498,N_2798,N_2913);
or U3499 (N_3499,N_2847,N_2805);
nand U3500 (N_3500,N_2733,N_2852);
or U3501 (N_3501,N_3155,N_2747);
and U3502 (N_3502,N_2786,N_3109);
xnor U3503 (N_3503,N_2520,N_2880);
xor U3504 (N_3504,N_2555,N_2970);
xnor U3505 (N_3505,N_2458,N_3192);
nor U3506 (N_3506,N_2517,N_2414);
or U3507 (N_3507,N_2868,N_2967);
or U3508 (N_3508,N_3040,N_3097);
or U3509 (N_3509,N_3130,N_3121);
xnor U3510 (N_3510,N_2498,N_2696);
xor U3511 (N_3511,N_3055,N_2516);
and U3512 (N_3512,N_2914,N_3080);
or U3513 (N_3513,N_2730,N_2862);
nor U3514 (N_3514,N_2728,N_3032);
nand U3515 (N_3515,N_2709,N_3175);
nor U3516 (N_3516,N_2731,N_2877);
xnor U3517 (N_3517,N_2493,N_2783);
and U3518 (N_3518,N_2741,N_2682);
nor U3519 (N_3519,N_3157,N_3059);
nor U3520 (N_3520,N_3002,N_2943);
and U3521 (N_3521,N_2812,N_3197);
nor U3522 (N_3522,N_2942,N_2695);
and U3523 (N_3523,N_2683,N_2451);
xor U3524 (N_3524,N_3071,N_2837);
and U3525 (N_3525,N_2887,N_2503);
nor U3526 (N_3526,N_3011,N_2971);
xnor U3527 (N_3527,N_2656,N_2598);
and U3528 (N_3528,N_2834,N_2518);
and U3529 (N_3529,N_2466,N_2607);
xor U3530 (N_3530,N_2781,N_2480);
nor U3531 (N_3531,N_3005,N_2873);
xnor U3532 (N_3532,N_3038,N_3001);
nor U3533 (N_3533,N_2544,N_2724);
and U3534 (N_3534,N_2570,N_2580);
and U3535 (N_3535,N_2905,N_2947);
nand U3536 (N_3536,N_3119,N_3052);
nor U3537 (N_3537,N_2439,N_2561);
xor U3538 (N_3538,N_2878,N_2840);
xnor U3539 (N_3539,N_3037,N_2654);
nor U3540 (N_3540,N_2574,N_3012);
or U3541 (N_3541,N_2793,N_3047);
nor U3542 (N_3542,N_3041,N_2821);
nor U3543 (N_3543,N_3014,N_3025);
nand U3544 (N_3544,N_2601,N_2594);
nor U3545 (N_3545,N_2889,N_2616);
and U3546 (N_3546,N_3116,N_2732);
xnor U3547 (N_3547,N_3198,N_3028);
nand U3548 (N_3548,N_3156,N_2999);
xnor U3549 (N_3549,N_2853,N_2883);
nand U3550 (N_3550,N_2638,N_2933);
nor U3551 (N_3551,N_2978,N_2523);
nor U3552 (N_3552,N_2980,N_2548);
or U3553 (N_3553,N_2499,N_2717);
nand U3554 (N_3554,N_2792,N_2495);
xnor U3555 (N_3555,N_3181,N_2585);
and U3556 (N_3556,N_2826,N_2991);
and U3557 (N_3557,N_2671,N_2404);
xor U3558 (N_3558,N_3076,N_2524);
nand U3559 (N_3559,N_2550,N_3064);
nor U3560 (N_3560,N_2749,N_2442);
xor U3561 (N_3561,N_2934,N_2668);
nor U3562 (N_3562,N_2563,N_2510);
nand U3563 (N_3563,N_3072,N_2739);
or U3564 (N_3564,N_2777,N_2571);
or U3565 (N_3565,N_2572,N_2765);
nor U3566 (N_3566,N_2655,N_3069);
or U3567 (N_3567,N_2648,N_2911);
nor U3568 (N_3568,N_2760,N_2507);
or U3569 (N_3569,N_3106,N_2961);
nor U3570 (N_3570,N_3090,N_2578);
xor U3571 (N_3571,N_2932,N_2562);
xnor U3572 (N_3572,N_2642,N_2481);
nand U3573 (N_3573,N_2795,N_3015);
xor U3574 (N_3574,N_2583,N_2719);
and U3575 (N_3575,N_2893,N_2678);
xor U3576 (N_3576,N_3114,N_2782);
xnor U3577 (N_3577,N_3110,N_2801);
xor U3578 (N_3578,N_2605,N_2780);
and U3579 (N_3579,N_2969,N_3154);
and U3580 (N_3580,N_2856,N_2618);
nand U3581 (N_3581,N_2614,N_3006);
or U3582 (N_3582,N_2501,N_2892);
nor U3583 (N_3583,N_3089,N_2900);
xor U3584 (N_3584,N_2620,N_3024);
nor U3585 (N_3585,N_2403,N_3165);
nor U3586 (N_3586,N_3134,N_2681);
and U3587 (N_3587,N_2456,N_2737);
nand U3588 (N_3588,N_2628,N_2712);
or U3589 (N_3589,N_2573,N_2917);
nor U3590 (N_3590,N_2417,N_3168);
or U3591 (N_3591,N_2768,N_3053);
xnor U3592 (N_3592,N_3087,N_2542);
nand U3593 (N_3593,N_2753,N_2650);
xnor U3594 (N_3594,N_2927,N_2931);
nor U3595 (N_3595,N_2669,N_2687);
nand U3596 (N_3596,N_2720,N_2402);
or U3597 (N_3597,N_2646,N_2569);
xnor U3598 (N_3598,N_3036,N_2674);
xnor U3599 (N_3599,N_2938,N_3086);
or U3600 (N_3600,N_3012,N_2606);
or U3601 (N_3601,N_2713,N_2675);
nand U3602 (N_3602,N_2499,N_2991);
nor U3603 (N_3603,N_2978,N_2625);
or U3604 (N_3604,N_2900,N_2710);
or U3605 (N_3605,N_3111,N_3171);
nand U3606 (N_3606,N_2811,N_2992);
or U3607 (N_3607,N_3081,N_3068);
nor U3608 (N_3608,N_2412,N_2956);
or U3609 (N_3609,N_3090,N_3023);
or U3610 (N_3610,N_2636,N_3041);
xnor U3611 (N_3611,N_3185,N_2656);
nand U3612 (N_3612,N_3040,N_2584);
xor U3613 (N_3613,N_2954,N_2533);
nand U3614 (N_3614,N_3044,N_3154);
or U3615 (N_3615,N_2963,N_2876);
and U3616 (N_3616,N_2910,N_3019);
and U3617 (N_3617,N_2753,N_2718);
nand U3618 (N_3618,N_2596,N_2837);
nor U3619 (N_3619,N_3076,N_2905);
nand U3620 (N_3620,N_2849,N_3125);
xor U3621 (N_3621,N_2739,N_3147);
and U3622 (N_3622,N_2745,N_2958);
and U3623 (N_3623,N_3018,N_2922);
xnor U3624 (N_3624,N_2605,N_3013);
nor U3625 (N_3625,N_3156,N_2921);
or U3626 (N_3626,N_2416,N_2530);
nand U3627 (N_3627,N_2906,N_2662);
or U3628 (N_3628,N_2977,N_3015);
or U3629 (N_3629,N_3105,N_3115);
xnor U3630 (N_3630,N_2925,N_2763);
nand U3631 (N_3631,N_3194,N_2470);
nand U3632 (N_3632,N_2893,N_2582);
nand U3633 (N_3633,N_2910,N_2792);
nor U3634 (N_3634,N_2626,N_2962);
or U3635 (N_3635,N_2755,N_2746);
nor U3636 (N_3636,N_3149,N_2753);
and U3637 (N_3637,N_2656,N_2779);
xnor U3638 (N_3638,N_2786,N_2736);
and U3639 (N_3639,N_2547,N_3166);
or U3640 (N_3640,N_2989,N_3061);
nor U3641 (N_3641,N_2509,N_2498);
nor U3642 (N_3642,N_3020,N_3189);
nor U3643 (N_3643,N_3017,N_2604);
or U3644 (N_3644,N_2932,N_2787);
or U3645 (N_3645,N_2986,N_2952);
and U3646 (N_3646,N_2597,N_2438);
nor U3647 (N_3647,N_2445,N_2599);
and U3648 (N_3648,N_2967,N_3026);
and U3649 (N_3649,N_2657,N_2636);
or U3650 (N_3650,N_2620,N_2702);
and U3651 (N_3651,N_2433,N_2748);
nor U3652 (N_3652,N_2455,N_2647);
xnor U3653 (N_3653,N_2565,N_2656);
nand U3654 (N_3654,N_2749,N_2419);
or U3655 (N_3655,N_2480,N_3047);
xnor U3656 (N_3656,N_2847,N_3130);
or U3657 (N_3657,N_2887,N_3016);
nor U3658 (N_3658,N_3062,N_3151);
or U3659 (N_3659,N_3149,N_2903);
and U3660 (N_3660,N_2615,N_2525);
or U3661 (N_3661,N_3196,N_2889);
xor U3662 (N_3662,N_2980,N_2406);
xor U3663 (N_3663,N_2799,N_2901);
or U3664 (N_3664,N_2582,N_2953);
nor U3665 (N_3665,N_2567,N_2753);
and U3666 (N_3666,N_2409,N_2521);
and U3667 (N_3667,N_3042,N_2600);
and U3668 (N_3668,N_2793,N_2931);
nand U3669 (N_3669,N_2697,N_2703);
nor U3670 (N_3670,N_3079,N_3076);
and U3671 (N_3671,N_2556,N_2774);
and U3672 (N_3672,N_2460,N_2547);
nor U3673 (N_3673,N_3056,N_2800);
and U3674 (N_3674,N_2464,N_2804);
xnor U3675 (N_3675,N_3039,N_2783);
xnor U3676 (N_3676,N_2819,N_3017);
or U3677 (N_3677,N_3093,N_2761);
nand U3678 (N_3678,N_3154,N_2887);
or U3679 (N_3679,N_2690,N_2522);
and U3680 (N_3680,N_2473,N_2754);
or U3681 (N_3681,N_2737,N_3107);
or U3682 (N_3682,N_3081,N_2708);
xor U3683 (N_3683,N_2835,N_3165);
or U3684 (N_3684,N_2890,N_2642);
or U3685 (N_3685,N_2435,N_2751);
or U3686 (N_3686,N_2818,N_2965);
xor U3687 (N_3687,N_2743,N_2929);
nand U3688 (N_3688,N_2520,N_2961);
nor U3689 (N_3689,N_2472,N_3186);
xor U3690 (N_3690,N_2630,N_2706);
and U3691 (N_3691,N_2930,N_2486);
nand U3692 (N_3692,N_3150,N_3131);
nor U3693 (N_3693,N_2508,N_2886);
nand U3694 (N_3694,N_2973,N_2534);
nand U3695 (N_3695,N_2454,N_2730);
or U3696 (N_3696,N_2722,N_2831);
and U3697 (N_3697,N_2848,N_2702);
and U3698 (N_3698,N_2675,N_2938);
or U3699 (N_3699,N_3004,N_2618);
nor U3700 (N_3700,N_2789,N_2569);
and U3701 (N_3701,N_2477,N_2676);
and U3702 (N_3702,N_2932,N_2494);
nand U3703 (N_3703,N_2561,N_2905);
xor U3704 (N_3704,N_3087,N_2534);
nand U3705 (N_3705,N_2655,N_3081);
xnor U3706 (N_3706,N_2925,N_2839);
nand U3707 (N_3707,N_2884,N_2577);
nand U3708 (N_3708,N_2631,N_2934);
or U3709 (N_3709,N_2755,N_2886);
and U3710 (N_3710,N_2596,N_2459);
nand U3711 (N_3711,N_3046,N_2806);
xor U3712 (N_3712,N_2678,N_2792);
and U3713 (N_3713,N_3036,N_2546);
or U3714 (N_3714,N_3017,N_2561);
nand U3715 (N_3715,N_2612,N_2547);
or U3716 (N_3716,N_3002,N_2716);
nor U3717 (N_3717,N_3158,N_2844);
or U3718 (N_3718,N_3153,N_2797);
or U3719 (N_3719,N_2599,N_3070);
or U3720 (N_3720,N_2544,N_2876);
and U3721 (N_3721,N_2720,N_2677);
or U3722 (N_3722,N_2568,N_3046);
xor U3723 (N_3723,N_3053,N_2970);
or U3724 (N_3724,N_2567,N_2575);
nor U3725 (N_3725,N_2927,N_2530);
xnor U3726 (N_3726,N_2614,N_2968);
nand U3727 (N_3727,N_2807,N_2989);
xnor U3728 (N_3728,N_2771,N_3144);
and U3729 (N_3729,N_2676,N_2542);
or U3730 (N_3730,N_2741,N_3105);
and U3731 (N_3731,N_2724,N_3043);
and U3732 (N_3732,N_2405,N_2467);
and U3733 (N_3733,N_2417,N_3142);
nor U3734 (N_3734,N_3187,N_2659);
or U3735 (N_3735,N_3011,N_2527);
or U3736 (N_3736,N_2531,N_2498);
or U3737 (N_3737,N_2950,N_2502);
or U3738 (N_3738,N_2989,N_2406);
nand U3739 (N_3739,N_2768,N_2951);
and U3740 (N_3740,N_2920,N_2903);
nor U3741 (N_3741,N_2891,N_2704);
nand U3742 (N_3742,N_3078,N_2789);
nand U3743 (N_3743,N_2639,N_2724);
and U3744 (N_3744,N_2667,N_2465);
and U3745 (N_3745,N_2510,N_2448);
nor U3746 (N_3746,N_3099,N_2450);
nand U3747 (N_3747,N_2753,N_2459);
and U3748 (N_3748,N_2666,N_2908);
nor U3749 (N_3749,N_2400,N_3123);
nand U3750 (N_3750,N_3090,N_2791);
and U3751 (N_3751,N_2799,N_3119);
xor U3752 (N_3752,N_3103,N_2524);
nand U3753 (N_3753,N_2967,N_2911);
nor U3754 (N_3754,N_2907,N_2760);
xnor U3755 (N_3755,N_2476,N_2495);
nand U3756 (N_3756,N_3014,N_2739);
nand U3757 (N_3757,N_2999,N_3032);
nor U3758 (N_3758,N_3066,N_2619);
nand U3759 (N_3759,N_2509,N_2521);
nor U3760 (N_3760,N_2739,N_2770);
nor U3761 (N_3761,N_3194,N_2645);
nor U3762 (N_3762,N_2581,N_2900);
xor U3763 (N_3763,N_2944,N_3120);
or U3764 (N_3764,N_2999,N_2566);
or U3765 (N_3765,N_3022,N_2501);
nand U3766 (N_3766,N_3043,N_3144);
and U3767 (N_3767,N_3125,N_2420);
or U3768 (N_3768,N_3158,N_2739);
nand U3769 (N_3769,N_2616,N_2830);
nand U3770 (N_3770,N_3158,N_2659);
and U3771 (N_3771,N_2644,N_2614);
nor U3772 (N_3772,N_2837,N_2547);
nor U3773 (N_3773,N_2578,N_3135);
xnor U3774 (N_3774,N_2870,N_3134);
and U3775 (N_3775,N_3025,N_2777);
nand U3776 (N_3776,N_2890,N_2814);
nand U3777 (N_3777,N_2723,N_2639);
nand U3778 (N_3778,N_2933,N_2986);
nand U3779 (N_3779,N_2843,N_2498);
or U3780 (N_3780,N_2631,N_3154);
nand U3781 (N_3781,N_2993,N_3106);
or U3782 (N_3782,N_2492,N_2786);
nor U3783 (N_3783,N_3068,N_2997);
nor U3784 (N_3784,N_2631,N_3135);
nor U3785 (N_3785,N_2421,N_2401);
or U3786 (N_3786,N_2843,N_3173);
and U3787 (N_3787,N_2979,N_3087);
nand U3788 (N_3788,N_3040,N_3122);
nand U3789 (N_3789,N_2726,N_3126);
and U3790 (N_3790,N_3015,N_3139);
or U3791 (N_3791,N_2681,N_2971);
and U3792 (N_3792,N_2865,N_3041);
nor U3793 (N_3793,N_2490,N_3070);
nand U3794 (N_3794,N_3069,N_2572);
nor U3795 (N_3795,N_2637,N_2666);
nand U3796 (N_3796,N_2484,N_2782);
xnor U3797 (N_3797,N_2735,N_2709);
nand U3798 (N_3798,N_3119,N_2926);
and U3799 (N_3799,N_2687,N_3031);
nor U3800 (N_3800,N_3160,N_2486);
or U3801 (N_3801,N_3000,N_2745);
and U3802 (N_3802,N_2492,N_2480);
and U3803 (N_3803,N_2451,N_2977);
nand U3804 (N_3804,N_2579,N_2758);
and U3805 (N_3805,N_2562,N_2868);
xor U3806 (N_3806,N_2851,N_2930);
or U3807 (N_3807,N_2580,N_2519);
nor U3808 (N_3808,N_2831,N_2974);
xor U3809 (N_3809,N_3010,N_2662);
or U3810 (N_3810,N_3048,N_2927);
nor U3811 (N_3811,N_2843,N_2733);
nor U3812 (N_3812,N_2975,N_2550);
nor U3813 (N_3813,N_2749,N_3128);
nand U3814 (N_3814,N_2985,N_2947);
and U3815 (N_3815,N_3065,N_2664);
xnor U3816 (N_3816,N_3027,N_2443);
nand U3817 (N_3817,N_2586,N_2836);
nor U3818 (N_3818,N_3032,N_2906);
and U3819 (N_3819,N_2764,N_3111);
nor U3820 (N_3820,N_2969,N_3183);
nand U3821 (N_3821,N_2456,N_2463);
xor U3822 (N_3822,N_2612,N_2922);
nor U3823 (N_3823,N_2714,N_3036);
nand U3824 (N_3824,N_2498,N_2996);
nor U3825 (N_3825,N_2510,N_2632);
xnor U3826 (N_3826,N_2850,N_3094);
xnor U3827 (N_3827,N_3030,N_2878);
nor U3828 (N_3828,N_2498,N_2434);
xnor U3829 (N_3829,N_2788,N_2913);
xnor U3830 (N_3830,N_2936,N_2932);
xor U3831 (N_3831,N_2598,N_3001);
xnor U3832 (N_3832,N_2777,N_2676);
nor U3833 (N_3833,N_2721,N_3039);
and U3834 (N_3834,N_2501,N_2581);
nor U3835 (N_3835,N_2767,N_3078);
nor U3836 (N_3836,N_2464,N_3059);
nand U3837 (N_3837,N_3055,N_2550);
or U3838 (N_3838,N_3155,N_3159);
nor U3839 (N_3839,N_2581,N_3125);
and U3840 (N_3840,N_3074,N_2652);
nand U3841 (N_3841,N_2633,N_2940);
or U3842 (N_3842,N_2409,N_2854);
nor U3843 (N_3843,N_3015,N_2533);
xnor U3844 (N_3844,N_2684,N_2462);
and U3845 (N_3845,N_2527,N_2957);
nor U3846 (N_3846,N_2989,N_2668);
nor U3847 (N_3847,N_2516,N_3009);
nand U3848 (N_3848,N_2628,N_2964);
xnor U3849 (N_3849,N_2430,N_2449);
nand U3850 (N_3850,N_2415,N_3011);
xnor U3851 (N_3851,N_3127,N_2447);
xnor U3852 (N_3852,N_2952,N_2529);
or U3853 (N_3853,N_2783,N_2514);
or U3854 (N_3854,N_2805,N_2894);
xnor U3855 (N_3855,N_2617,N_3059);
xor U3856 (N_3856,N_2809,N_2686);
nor U3857 (N_3857,N_2812,N_2823);
xor U3858 (N_3858,N_3186,N_3084);
and U3859 (N_3859,N_2751,N_3016);
and U3860 (N_3860,N_3049,N_2635);
and U3861 (N_3861,N_2871,N_3166);
nand U3862 (N_3862,N_3065,N_2942);
nor U3863 (N_3863,N_2795,N_2460);
xor U3864 (N_3864,N_3163,N_2883);
nor U3865 (N_3865,N_2676,N_2449);
or U3866 (N_3866,N_2478,N_2417);
and U3867 (N_3867,N_3053,N_2486);
nor U3868 (N_3868,N_2830,N_2648);
nand U3869 (N_3869,N_2559,N_3111);
nor U3870 (N_3870,N_2908,N_2626);
xor U3871 (N_3871,N_2906,N_2659);
nand U3872 (N_3872,N_2546,N_3170);
nor U3873 (N_3873,N_2735,N_2631);
nor U3874 (N_3874,N_2522,N_3052);
nand U3875 (N_3875,N_2646,N_3018);
or U3876 (N_3876,N_2624,N_2891);
and U3877 (N_3877,N_2661,N_2923);
or U3878 (N_3878,N_2721,N_2469);
xor U3879 (N_3879,N_2702,N_3069);
xor U3880 (N_3880,N_2923,N_2407);
nand U3881 (N_3881,N_2790,N_2405);
xor U3882 (N_3882,N_2607,N_2581);
xor U3883 (N_3883,N_2987,N_3002);
and U3884 (N_3884,N_2534,N_2698);
xor U3885 (N_3885,N_3169,N_2874);
or U3886 (N_3886,N_2914,N_2509);
nand U3887 (N_3887,N_3074,N_2983);
nor U3888 (N_3888,N_3063,N_2786);
xnor U3889 (N_3889,N_2799,N_2871);
nor U3890 (N_3890,N_2881,N_3082);
xnor U3891 (N_3891,N_2404,N_2853);
xor U3892 (N_3892,N_2709,N_2501);
and U3893 (N_3893,N_2680,N_2756);
or U3894 (N_3894,N_2528,N_2813);
xor U3895 (N_3895,N_2425,N_2872);
xor U3896 (N_3896,N_2991,N_2791);
and U3897 (N_3897,N_3072,N_2462);
nor U3898 (N_3898,N_2764,N_3129);
or U3899 (N_3899,N_2478,N_2859);
or U3900 (N_3900,N_2703,N_2537);
xnor U3901 (N_3901,N_2707,N_2814);
nor U3902 (N_3902,N_3037,N_2716);
nor U3903 (N_3903,N_2629,N_2849);
xor U3904 (N_3904,N_2796,N_3170);
xor U3905 (N_3905,N_2641,N_3181);
nor U3906 (N_3906,N_3067,N_3173);
and U3907 (N_3907,N_2570,N_2441);
and U3908 (N_3908,N_3047,N_2559);
or U3909 (N_3909,N_2625,N_3023);
and U3910 (N_3910,N_2800,N_2499);
nand U3911 (N_3911,N_2405,N_2950);
and U3912 (N_3912,N_2974,N_3153);
or U3913 (N_3913,N_2875,N_2773);
nor U3914 (N_3914,N_2926,N_2691);
or U3915 (N_3915,N_3198,N_3144);
nand U3916 (N_3916,N_2699,N_2624);
xnor U3917 (N_3917,N_2991,N_2616);
or U3918 (N_3918,N_2745,N_2831);
nor U3919 (N_3919,N_2446,N_2989);
nor U3920 (N_3920,N_2898,N_2763);
nor U3921 (N_3921,N_2784,N_2859);
nor U3922 (N_3922,N_3111,N_2512);
and U3923 (N_3923,N_2612,N_3024);
nand U3924 (N_3924,N_2958,N_2423);
xor U3925 (N_3925,N_2767,N_2869);
xor U3926 (N_3926,N_2672,N_3132);
xor U3927 (N_3927,N_2787,N_3032);
or U3928 (N_3928,N_2435,N_2719);
nor U3929 (N_3929,N_2929,N_2957);
or U3930 (N_3930,N_3099,N_2476);
nand U3931 (N_3931,N_2671,N_2904);
and U3932 (N_3932,N_2998,N_2925);
nor U3933 (N_3933,N_3057,N_2943);
nand U3934 (N_3934,N_2876,N_2921);
nor U3935 (N_3935,N_2802,N_2526);
or U3936 (N_3936,N_2853,N_2602);
nand U3937 (N_3937,N_2548,N_2625);
or U3938 (N_3938,N_2413,N_2752);
and U3939 (N_3939,N_2749,N_3023);
or U3940 (N_3940,N_2906,N_3039);
and U3941 (N_3941,N_3016,N_3154);
nor U3942 (N_3942,N_3123,N_3020);
or U3943 (N_3943,N_3036,N_2846);
xnor U3944 (N_3944,N_2688,N_2730);
nand U3945 (N_3945,N_2876,N_2750);
and U3946 (N_3946,N_2691,N_3170);
nand U3947 (N_3947,N_2540,N_2688);
and U3948 (N_3948,N_2789,N_3176);
nand U3949 (N_3949,N_2870,N_2988);
xor U3950 (N_3950,N_2446,N_2839);
or U3951 (N_3951,N_2979,N_2525);
nand U3952 (N_3952,N_2796,N_2975);
nor U3953 (N_3953,N_2992,N_2887);
and U3954 (N_3954,N_2864,N_3194);
nor U3955 (N_3955,N_2855,N_2794);
nand U3956 (N_3956,N_2464,N_3091);
and U3957 (N_3957,N_2451,N_2513);
xnor U3958 (N_3958,N_3039,N_2842);
and U3959 (N_3959,N_2412,N_2930);
or U3960 (N_3960,N_2993,N_2557);
xor U3961 (N_3961,N_2886,N_2947);
nor U3962 (N_3962,N_2457,N_2594);
nand U3963 (N_3963,N_3032,N_2774);
and U3964 (N_3964,N_2931,N_2764);
or U3965 (N_3965,N_2677,N_2902);
and U3966 (N_3966,N_3110,N_3102);
xnor U3967 (N_3967,N_2558,N_2925);
nor U3968 (N_3968,N_2535,N_2627);
and U3969 (N_3969,N_2771,N_2804);
nand U3970 (N_3970,N_2911,N_2852);
nand U3971 (N_3971,N_2786,N_3084);
nand U3972 (N_3972,N_2492,N_2753);
nor U3973 (N_3973,N_2532,N_2933);
nand U3974 (N_3974,N_3111,N_2455);
nor U3975 (N_3975,N_2603,N_2434);
and U3976 (N_3976,N_2742,N_3102);
and U3977 (N_3977,N_2523,N_2663);
and U3978 (N_3978,N_3068,N_2781);
xor U3979 (N_3979,N_2687,N_2447);
nand U3980 (N_3980,N_3196,N_2841);
xnor U3981 (N_3981,N_2744,N_2554);
nand U3982 (N_3982,N_2493,N_2696);
xnor U3983 (N_3983,N_2998,N_2577);
or U3984 (N_3984,N_3155,N_2475);
nor U3985 (N_3985,N_3141,N_2893);
xor U3986 (N_3986,N_2694,N_2797);
nor U3987 (N_3987,N_2414,N_2936);
nand U3988 (N_3988,N_2633,N_2779);
or U3989 (N_3989,N_2800,N_2964);
or U3990 (N_3990,N_2787,N_2623);
xnor U3991 (N_3991,N_2499,N_2978);
nor U3992 (N_3992,N_2994,N_2737);
or U3993 (N_3993,N_2928,N_2600);
and U3994 (N_3994,N_2828,N_2644);
nand U3995 (N_3995,N_2745,N_2686);
nor U3996 (N_3996,N_2969,N_3061);
nor U3997 (N_3997,N_2891,N_2845);
nor U3998 (N_3998,N_2562,N_2696);
or U3999 (N_3999,N_3169,N_2529);
nand U4000 (N_4000,N_3787,N_3582);
nand U4001 (N_4001,N_3880,N_3974);
xor U4002 (N_4002,N_3396,N_3357);
xnor U4003 (N_4003,N_3460,N_3699);
and U4004 (N_4004,N_3951,N_3482);
nand U4005 (N_4005,N_3645,N_3464);
or U4006 (N_4006,N_3430,N_3964);
nor U4007 (N_4007,N_3561,N_3719);
or U4008 (N_4008,N_3572,N_3770);
and U4009 (N_4009,N_3264,N_3305);
xnor U4010 (N_4010,N_3382,N_3437);
xnor U4011 (N_4011,N_3591,N_3671);
xor U4012 (N_4012,N_3995,N_3440);
and U4013 (N_4013,N_3481,N_3622);
xnor U4014 (N_4014,N_3748,N_3786);
or U4015 (N_4015,N_3379,N_3223);
nor U4016 (N_4016,N_3352,N_3615);
and U4017 (N_4017,N_3971,N_3638);
or U4018 (N_4018,N_3627,N_3849);
and U4019 (N_4019,N_3338,N_3530);
and U4020 (N_4020,N_3465,N_3311);
nand U4021 (N_4021,N_3563,N_3448);
nand U4022 (N_4022,N_3546,N_3273);
nand U4023 (N_4023,N_3997,N_3872);
or U4024 (N_4024,N_3905,N_3433);
nand U4025 (N_4025,N_3734,N_3867);
and U4026 (N_4026,N_3846,N_3869);
xnor U4027 (N_4027,N_3458,N_3658);
nand U4028 (N_4028,N_3996,N_3291);
or U4029 (N_4029,N_3837,N_3220);
nand U4030 (N_4030,N_3738,N_3793);
nand U4031 (N_4031,N_3657,N_3624);
nor U4032 (N_4032,N_3606,N_3652);
xor U4033 (N_4033,N_3435,N_3850);
xor U4034 (N_4034,N_3602,N_3211);
xnor U4035 (N_4035,N_3730,N_3289);
or U4036 (N_4036,N_3716,N_3826);
xor U4037 (N_4037,N_3462,N_3203);
nand U4038 (N_4038,N_3222,N_3968);
nand U4039 (N_4039,N_3982,N_3979);
and U4040 (N_4040,N_3369,N_3577);
nor U4041 (N_4041,N_3474,N_3385);
or U4042 (N_4042,N_3973,N_3442);
nor U4043 (N_4043,N_3723,N_3976);
and U4044 (N_4044,N_3950,N_3229);
nor U4045 (N_4045,N_3536,N_3443);
xor U4046 (N_4046,N_3878,N_3801);
nor U4047 (N_4047,N_3691,N_3551);
or U4048 (N_4048,N_3255,N_3509);
xor U4049 (N_4049,N_3439,N_3752);
or U4050 (N_4050,N_3947,N_3287);
and U4051 (N_4051,N_3426,N_3900);
nor U4052 (N_4052,N_3335,N_3489);
or U4053 (N_4053,N_3907,N_3854);
xor U4054 (N_4054,N_3301,N_3362);
nor U4055 (N_4055,N_3649,N_3634);
and U4056 (N_4056,N_3936,N_3844);
xor U4057 (N_4057,N_3650,N_3498);
or U4058 (N_4058,N_3596,N_3579);
or U4059 (N_4059,N_3919,N_3763);
nand U4060 (N_4060,N_3910,N_3836);
or U4061 (N_4061,N_3772,N_3932);
and U4062 (N_4062,N_3775,N_3553);
and U4063 (N_4063,N_3597,N_3575);
nand U4064 (N_4064,N_3743,N_3513);
nand U4065 (N_4065,N_3219,N_3594);
and U4066 (N_4066,N_3922,N_3717);
xnor U4067 (N_4067,N_3901,N_3685);
or U4068 (N_4068,N_3805,N_3918);
nor U4069 (N_4069,N_3384,N_3779);
nor U4070 (N_4070,N_3924,N_3340);
xor U4071 (N_4071,N_3588,N_3796);
or U4072 (N_4072,N_3893,N_3909);
nand U4073 (N_4073,N_3954,N_3480);
or U4074 (N_4074,N_3704,N_3981);
and U4075 (N_4075,N_3792,N_3527);
or U4076 (N_4076,N_3304,N_3535);
nor U4077 (N_4077,N_3232,N_3392);
and U4078 (N_4078,N_3908,N_3461);
or U4079 (N_4079,N_3816,N_3726);
xnor U4080 (N_4080,N_3928,N_3888);
xnor U4081 (N_4081,N_3560,N_3760);
or U4082 (N_4082,N_3526,N_3733);
or U4083 (N_4083,N_3576,N_3977);
nor U4084 (N_4084,N_3927,N_3274);
and U4085 (N_4085,N_3347,N_3855);
and U4086 (N_4086,N_3504,N_3445);
nand U4087 (N_4087,N_3538,N_3533);
and U4088 (N_4088,N_3324,N_3554);
xnor U4089 (N_4089,N_3923,N_3200);
xnor U4090 (N_4090,N_3410,N_3729);
nor U4091 (N_4091,N_3742,N_3544);
nor U4092 (N_4092,N_3236,N_3903);
nand U4093 (N_4093,N_3983,N_3938);
nand U4094 (N_4094,N_3988,N_3926);
nor U4095 (N_4095,N_3765,N_3686);
or U4096 (N_4096,N_3682,N_3675);
xor U4097 (N_4097,N_3952,N_3640);
nand U4098 (N_4098,N_3641,N_3722);
xor U4099 (N_4099,N_3949,N_3916);
nor U4100 (N_4100,N_3346,N_3698);
and U4101 (N_4101,N_3331,N_3688);
and U4102 (N_4102,N_3486,N_3687);
and U4103 (N_4103,N_3310,N_3522);
nand U4104 (N_4104,N_3721,N_3496);
xor U4105 (N_4105,N_3659,N_3521);
nand U4106 (N_4106,N_3380,N_3940);
xor U4107 (N_4107,N_3838,N_3703);
nor U4108 (N_4108,N_3674,N_3630);
and U4109 (N_4109,N_3366,N_3243);
nor U4110 (N_4110,N_3957,N_3555);
or U4111 (N_4111,N_3669,N_3361);
and U4112 (N_4112,N_3339,N_3316);
xnor U4113 (N_4113,N_3386,N_3904);
and U4114 (N_4114,N_3212,N_3604);
and U4115 (N_4115,N_3409,N_3913);
nor U4116 (N_4116,N_3470,N_3350);
or U4117 (N_4117,N_3363,N_3935);
nand U4118 (N_4118,N_3595,N_3663);
nand U4119 (N_4119,N_3827,N_3660);
or U4120 (N_4120,N_3795,N_3628);
and U4121 (N_4121,N_3315,N_3601);
xor U4122 (N_4122,N_3899,N_3993);
nand U4123 (N_4123,N_3268,N_3713);
or U4124 (N_4124,N_3545,N_3956);
xor U4125 (N_4125,N_3965,N_3221);
nor U4126 (N_4126,N_3874,N_3813);
or U4127 (N_4127,N_3328,N_3831);
nor U4128 (N_4128,N_3771,N_3737);
and U4129 (N_4129,N_3318,N_3325);
or U4130 (N_4130,N_3774,N_3788);
nor U4131 (N_4131,N_3485,N_3929);
and U4132 (N_4132,N_3398,N_3423);
nor U4133 (N_4133,N_3994,N_3519);
nor U4134 (N_4134,N_3414,N_3250);
nor U4135 (N_4135,N_3343,N_3808);
nand U4136 (N_4136,N_3611,N_3736);
and U4137 (N_4137,N_3677,N_3732);
and U4138 (N_4138,N_3800,N_3963);
or U4139 (N_4139,N_3987,N_3725);
nor U4140 (N_4140,N_3724,N_3507);
or U4141 (N_4141,N_3248,N_3896);
or U4142 (N_4142,N_3585,N_3978);
or U4143 (N_4143,N_3282,N_3368);
xor U4144 (N_4144,N_3502,N_3676);
and U4145 (N_4145,N_3953,N_3495);
and U4146 (N_4146,N_3281,N_3438);
nand U4147 (N_4147,N_3383,N_3541);
and U4148 (N_4148,N_3317,N_3371);
xor U4149 (N_4149,N_3537,N_3727);
nor U4150 (N_4150,N_3262,N_3895);
nand U4151 (N_4151,N_3424,N_3708);
nand U4152 (N_4152,N_3710,N_3961);
nor U4153 (N_4153,N_3868,N_3969);
and U4154 (N_4154,N_3422,N_3647);
and U4155 (N_4155,N_3493,N_3753);
nand U4156 (N_4156,N_3313,N_3984);
nand U4157 (N_4157,N_3240,N_3802);
nor U4158 (N_4158,N_3574,N_3870);
and U4159 (N_4159,N_3930,N_3889);
and U4160 (N_4160,N_3451,N_3344);
and U4161 (N_4161,N_3931,N_3680);
xnor U4162 (N_4162,N_3405,N_3299);
xnor U4163 (N_4163,N_3859,N_3623);
and U4164 (N_4164,N_3333,N_3558);
xor U4165 (N_4165,N_3683,N_3266);
nand U4166 (N_4166,N_3945,N_3702);
and U4167 (N_4167,N_3374,N_3975);
and U4168 (N_4168,N_3532,N_3202);
and U4169 (N_4169,N_3490,N_3387);
or U4170 (N_4170,N_3402,N_3825);
or U4171 (N_4171,N_3812,N_3261);
or U4172 (N_4172,N_3373,N_3308);
xnor U4173 (N_4173,N_3841,N_3799);
and U4174 (N_4174,N_3568,N_3242);
nand U4175 (N_4175,N_3972,N_3832);
or U4176 (N_4176,N_3705,N_3946);
nand U4177 (N_4177,N_3503,N_3720);
and U4178 (N_4178,N_3668,N_3436);
or U4179 (N_4179,N_3834,N_3399);
and U4180 (N_4180,N_3283,N_3619);
or U4181 (N_4181,N_3277,N_3589);
nand U4182 (N_4182,N_3731,N_3914);
xnor U4183 (N_4183,N_3866,N_3662);
nand U4184 (N_4184,N_3421,N_3512);
nand U4185 (N_4185,N_3865,N_3639);
nor U4186 (N_4186,N_3600,N_3740);
or U4187 (N_4187,N_3672,N_3523);
or U4188 (N_4188,N_3260,N_3378);
or U4189 (N_4189,N_3456,N_3487);
nand U4190 (N_4190,N_3785,N_3635);
or U4191 (N_4191,N_3225,N_3960);
and U4192 (N_4192,N_3783,N_3427);
and U4193 (N_4193,N_3891,N_3531);
and U4194 (N_4194,N_3970,N_3449);
xnor U4195 (N_4195,N_3418,N_3603);
nand U4196 (N_4196,N_3784,N_3406);
or U4197 (N_4197,N_3566,N_3718);
nand U4198 (N_4198,N_3351,N_3213);
xnor U4199 (N_4199,N_3454,N_3570);
nand U4200 (N_4200,N_3745,N_3381);
and U4201 (N_4201,N_3573,N_3839);
xor U4202 (N_4202,N_3217,N_3694);
nor U4203 (N_4203,N_3517,N_3757);
xnor U4204 (N_4204,N_3506,N_3821);
xnor U4205 (N_4205,N_3592,N_3695);
or U4206 (N_4206,N_3279,N_3894);
xnor U4207 (N_4207,N_3810,N_3394);
nand U4208 (N_4208,N_3857,N_3216);
nand U4209 (N_4209,N_3345,N_3782);
nor U4210 (N_4210,N_3468,N_3824);
and U4211 (N_4211,N_3320,N_3432);
nor U4212 (N_4212,N_3794,N_3237);
nand U4213 (N_4213,N_3471,N_3741);
or U4214 (N_4214,N_3666,N_3276);
nand U4215 (N_4215,N_3254,N_3500);
nor U4216 (N_4216,N_3707,N_3278);
xor U4217 (N_4217,N_3681,N_3986);
nand U4218 (N_4218,N_3701,N_3670);
nand U4219 (N_4219,N_3505,N_3937);
and U4220 (N_4220,N_3581,N_3776);
nand U4221 (N_4221,N_3789,N_3655);
nand U4222 (N_4222,N_3564,N_3621);
xnor U4223 (N_4223,N_3843,N_3858);
nand U4224 (N_4224,N_3637,N_3256);
nor U4225 (N_4225,N_3355,N_3319);
xnor U4226 (N_4226,N_3205,N_3542);
xnor U4227 (N_4227,N_3550,N_3851);
nand U4228 (N_4228,N_3342,N_3210);
xnor U4229 (N_4229,N_3469,N_3696);
xor U4230 (N_4230,N_3525,N_3365);
xor U4231 (N_4231,N_3845,N_3492);
nor U4232 (N_4232,N_3610,N_3390);
and U4233 (N_4233,N_3818,N_3364);
or U4234 (N_4234,N_3265,N_3511);
nand U4235 (N_4235,N_3459,N_3848);
xnor U4236 (N_4236,N_3902,N_3514);
or U4237 (N_4237,N_3943,N_3201);
and U4238 (N_4238,N_3962,N_3241);
nor U4239 (N_4239,N_3842,N_3244);
nand U4240 (N_4240,N_3215,N_3272);
or U4241 (N_4241,N_3643,N_3646);
or U4242 (N_4242,N_3270,N_3593);
and U4243 (N_4243,N_3548,N_3428);
or U4244 (N_4244,N_3915,N_3569);
or U4245 (N_4245,N_3284,N_3678);
xor U4246 (N_4246,N_3297,N_3388);
nand U4247 (N_4247,N_3617,N_3499);
nor U4248 (N_4248,N_3238,N_3955);
and U4249 (N_4249,N_3247,N_3251);
xor U4250 (N_4250,N_3989,N_3479);
or U4251 (N_4251,N_3906,N_3330);
and U4252 (N_4252,N_3648,N_3693);
or U4253 (N_4253,N_3590,N_3292);
nand U4254 (N_4254,N_3992,N_3822);
xnor U4255 (N_4255,N_3661,N_3417);
nor U4256 (N_4256,N_3933,N_3618);
nand U4257 (N_4257,N_3510,N_3208);
and U4258 (N_4258,N_3879,N_3767);
and U4259 (N_4259,N_3269,N_3966);
nor U4260 (N_4260,N_3875,N_3881);
or U4261 (N_4261,N_3609,N_3235);
nand U4262 (N_4262,N_3689,N_3897);
nand U4263 (N_4263,N_3746,N_3814);
xnor U4264 (N_4264,N_3476,N_3556);
and U4265 (N_4265,N_3777,N_3524);
xor U4266 (N_4266,N_3815,N_3651);
nand U4267 (N_4267,N_3791,N_3584);
nor U4268 (N_4268,N_3887,N_3644);
nor U4269 (N_4269,N_3258,N_3580);
xnor U4270 (N_4270,N_3377,N_3483);
nand U4271 (N_4271,N_3206,N_3882);
xnor U4272 (N_4272,N_3452,N_3985);
or U4273 (N_4273,N_3415,N_3306);
nor U4274 (N_4274,N_3959,N_3408);
nor U4275 (N_4275,N_3370,N_3376);
or U4276 (N_4276,N_3751,N_3249);
nor U4277 (N_4277,N_3226,N_3245);
nand U4278 (N_4278,N_3833,N_3497);
xor U4279 (N_4279,N_3337,N_3780);
nor U4280 (N_4280,N_3252,N_3552);
or U4281 (N_4281,N_3395,N_3472);
and U4282 (N_4282,N_3877,N_3296);
xnor U4283 (N_4283,N_3477,N_3473);
nor U4284 (N_4284,N_3665,N_3557);
or U4285 (N_4285,N_3778,N_3204);
or U4286 (N_4286,N_3214,N_3667);
nand U4287 (N_4287,N_3467,N_3697);
nand U4288 (N_4288,N_3300,N_3823);
xnor U4289 (N_4289,N_3773,N_3334);
xnor U4290 (N_4290,N_3744,N_3413);
or U4291 (N_4291,N_3709,N_3873);
nor U4292 (N_4292,N_3420,N_3755);
xnor U4293 (N_4293,N_3425,N_3890);
or U4294 (N_4294,N_3798,N_3583);
xnor U4295 (N_4295,N_3690,N_3224);
and U4296 (N_4296,N_3835,N_3664);
and U4297 (N_4297,N_3332,N_3886);
nor U4298 (N_4298,N_3326,N_3750);
nor U4299 (N_4299,N_3654,N_3920);
and U4300 (N_4300,N_3999,N_3840);
nand U4301 (N_4301,N_3620,N_3884);
nand U4302 (N_4302,N_3911,N_3389);
and U4303 (N_4303,N_3285,N_3457);
or U4304 (N_4304,N_3759,N_3271);
xnor U4305 (N_4305,N_3466,N_3820);
xor U4306 (N_4306,N_3516,N_3586);
and U4307 (N_4307,N_3700,N_3444);
or U4308 (N_4308,N_3508,N_3941);
xnor U4309 (N_4309,N_3275,N_3599);
nor U4310 (N_4310,N_3227,N_3925);
xnor U4311 (N_4311,N_3958,N_3819);
nor U4312 (N_4312,N_3806,N_3354);
nand U4313 (N_4313,N_3852,N_3441);
xnor U4314 (N_4314,N_3565,N_3863);
and U4315 (N_4315,N_3323,N_3341);
or U4316 (N_4316,N_3539,N_3478);
or U4317 (N_4317,N_3944,N_3728);
xor U4318 (N_4318,N_3797,N_3529);
and U4319 (N_4319,N_3228,N_3828);
or U4320 (N_4320,N_3607,N_3761);
or U4321 (N_4321,N_3942,N_3559);
nor U4322 (N_4322,N_3735,N_3853);
nor U4323 (N_4323,N_3488,N_3885);
xnor U4324 (N_4324,N_3401,N_3416);
xnor U4325 (N_4325,N_3967,N_3811);
or U4326 (N_4326,N_3692,N_3758);
xnor U4327 (N_4327,N_3998,N_3501);
and U4328 (N_4328,N_3290,N_3372);
xnor U4329 (N_4329,N_3817,N_3625);
or U4330 (N_4330,N_3515,N_3356);
nand U4331 (N_4331,N_3404,N_3253);
nand U4332 (N_4332,N_3327,N_3605);
and U4333 (N_4333,N_3230,N_3288);
and U4334 (N_4334,N_3948,N_3419);
or U4335 (N_4335,N_3636,N_3714);
xor U4336 (N_4336,N_3829,N_3431);
nor U4337 (N_4337,N_3939,N_3608);
and U4338 (N_4338,N_3912,N_3547);
xnor U4339 (N_4339,N_3612,N_3856);
xor U4340 (N_4340,N_3578,N_3562);
or U4341 (N_4341,N_3864,N_3980);
and U4342 (N_4342,N_3762,N_3429);
nor U4343 (N_4343,N_3233,N_3684);
or U4344 (N_4344,N_3871,N_3312);
nor U4345 (N_4345,N_3446,N_3360);
or U4346 (N_4346,N_3412,N_3598);
nor U4347 (N_4347,N_3447,N_3411);
or U4348 (N_4348,N_3484,N_3239);
nand U4349 (N_4349,N_3990,N_3883);
and U4350 (N_4350,N_3898,N_3804);
and U4351 (N_4351,N_3917,N_3207);
and U4352 (N_4352,N_3633,N_3349);
nand U4353 (N_4353,N_3455,N_3754);
nand U4354 (N_4354,N_3860,N_3375);
nand U4355 (N_4355,N_3293,N_3309);
and U4356 (N_4356,N_3491,N_3518);
nand U4357 (N_4357,N_3766,N_3453);
or U4358 (N_4358,N_3397,N_3631);
or U4359 (N_4359,N_3286,N_3781);
xnor U4360 (N_4360,N_3534,N_3711);
and U4361 (N_4361,N_3679,N_3632);
or U4362 (N_4362,N_3616,N_3209);
nor U4363 (N_4363,N_3303,N_3768);
nor U4364 (N_4364,N_3407,N_3263);
and U4365 (N_4365,N_3934,N_3626);
or U4366 (N_4366,N_3257,N_3790);
nand U4367 (N_4367,N_3991,N_3450);
and U4368 (N_4368,N_3336,N_3494);
or U4369 (N_4369,N_3712,N_3298);
xnor U4370 (N_4370,N_3393,N_3353);
nor U4371 (N_4371,N_3892,N_3715);
xnor U4372 (N_4372,N_3847,N_3259);
nand U4373 (N_4373,N_3434,N_3307);
and U4374 (N_4374,N_3642,N_3520);
nor U4375 (N_4375,N_3218,N_3769);
nor U4376 (N_4376,N_3403,N_3830);
xor U4377 (N_4377,N_3921,N_3540);
and U4378 (N_4378,N_3348,N_3549);
and U4379 (N_4379,N_3656,N_3614);
nand U4380 (N_4380,N_3673,N_3807);
nor U4381 (N_4381,N_3861,N_3756);
and U4382 (N_4382,N_3764,N_3322);
nor U4383 (N_4383,N_3747,N_3862);
and U4384 (N_4384,N_3653,N_3329);
nand U4385 (N_4385,N_3358,N_3475);
and U4386 (N_4386,N_3314,N_3400);
or U4387 (N_4387,N_3267,N_3571);
or U4388 (N_4388,N_3295,N_3629);
xor U4389 (N_4389,N_3246,N_3302);
nand U4390 (N_4390,N_3231,N_3706);
xnor U4391 (N_4391,N_3280,N_3321);
xnor U4392 (N_4392,N_3294,N_3391);
nand U4393 (N_4393,N_3803,N_3613);
xor U4394 (N_4394,N_3567,N_3359);
nor U4395 (N_4395,N_3587,N_3367);
and U4396 (N_4396,N_3749,N_3528);
nand U4397 (N_4397,N_3463,N_3809);
nand U4398 (N_4398,N_3876,N_3739);
xor U4399 (N_4399,N_3543,N_3234);
or U4400 (N_4400,N_3532,N_3605);
xnor U4401 (N_4401,N_3958,N_3956);
nor U4402 (N_4402,N_3367,N_3643);
nand U4403 (N_4403,N_3416,N_3637);
nor U4404 (N_4404,N_3299,N_3517);
nor U4405 (N_4405,N_3460,N_3477);
nand U4406 (N_4406,N_3363,N_3546);
nor U4407 (N_4407,N_3296,N_3594);
nor U4408 (N_4408,N_3374,N_3515);
and U4409 (N_4409,N_3489,N_3960);
nor U4410 (N_4410,N_3505,N_3608);
or U4411 (N_4411,N_3916,N_3989);
and U4412 (N_4412,N_3622,N_3368);
nor U4413 (N_4413,N_3745,N_3980);
or U4414 (N_4414,N_3512,N_3911);
nor U4415 (N_4415,N_3291,N_3369);
and U4416 (N_4416,N_3370,N_3932);
xor U4417 (N_4417,N_3346,N_3232);
or U4418 (N_4418,N_3739,N_3793);
xnor U4419 (N_4419,N_3695,N_3948);
nand U4420 (N_4420,N_3746,N_3407);
nand U4421 (N_4421,N_3904,N_3337);
nand U4422 (N_4422,N_3492,N_3746);
and U4423 (N_4423,N_3618,N_3742);
xnor U4424 (N_4424,N_3316,N_3454);
nor U4425 (N_4425,N_3630,N_3288);
xor U4426 (N_4426,N_3412,N_3965);
or U4427 (N_4427,N_3649,N_3285);
nand U4428 (N_4428,N_3326,N_3624);
or U4429 (N_4429,N_3940,N_3260);
nor U4430 (N_4430,N_3435,N_3746);
nand U4431 (N_4431,N_3501,N_3241);
or U4432 (N_4432,N_3470,N_3507);
xor U4433 (N_4433,N_3685,N_3849);
xnor U4434 (N_4434,N_3717,N_3359);
nor U4435 (N_4435,N_3622,N_3562);
and U4436 (N_4436,N_3336,N_3685);
nand U4437 (N_4437,N_3965,N_3666);
or U4438 (N_4438,N_3609,N_3241);
nor U4439 (N_4439,N_3928,N_3473);
xnor U4440 (N_4440,N_3363,N_3573);
and U4441 (N_4441,N_3391,N_3229);
and U4442 (N_4442,N_3819,N_3823);
nand U4443 (N_4443,N_3558,N_3725);
nor U4444 (N_4444,N_3781,N_3717);
nand U4445 (N_4445,N_3926,N_3841);
or U4446 (N_4446,N_3399,N_3717);
nand U4447 (N_4447,N_3615,N_3826);
and U4448 (N_4448,N_3953,N_3939);
xnor U4449 (N_4449,N_3407,N_3792);
nor U4450 (N_4450,N_3936,N_3796);
xor U4451 (N_4451,N_3621,N_3567);
xnor U4452 (N_4452,N_3468,N_3668);
nand U4453 (N_4453,N_3650,N_3897);
and U4454 (N_4454,N_3882,N_3503);
nand U4455 (N_4455,N_3332,N_3952);
nor U4456 (N_4456,N_3291,N_3289);
nand U4457 (N_4457,N_3861,N_3936);
nand U4458 (N_4458,N_3902,N_3475);
or U4459 (N_4459,N_3621,N_3646);
nor U4460 (N_4460,N_3748,N_3793);
nand U4461 (N_4461,N_3997,N_3977);
xor U4462 (N_4462,N_3688,N_3719);
or U4463 (N_4463,N_3284,N_3250);
nor U4464 (N_4464,N_3614,N_3583);
nor U4465 (N_4465,N_3273,N_3508);
nor U4466 (N_4466,N_3897,N_3518);
nand U4467 (N_4467,N_3630,N_3592);
and U4468 (N_4468,N_3270,N_3850);
nand U4469 (N_4469,N_3390,N_3796);
or U4470 (N_4470,N_3809,N_3674);
nand U4471 (N_4471,N_3506,N_3747);
nor U4472 (N_4472,N_3519,N_3824);
xor U4473 (N_4473,N_3680,N_3286);
nand U4474 (N_4474,N_3853,N_3983);
or U4475 (N_4475,N_3437,N_3746);
xor U4476 (N_4476,N_3946,N_3646);
xnor U4477 (N_4477,N_3534,N_3434);
xor U4478 (N_4478,N_3432,N_3700);
or U4479 (N_4479,N_3428,N_3733);
xnor U4480 (N_4480,N_3642,N_3230);
xor U4481 (N_4481,N_3865,N_3212);
nor U4482 (N_4482,N_3995,N_3506);
nor U4483 (N_4483,N_3708,N_3814);
nor U4484 (N_4484,N_3242,N_3235);
or U4485 (N_4485,N_3572,N_3300);
or U4486 (N_4486,N_3305,N_3324);
or U4487 (N_4487,N_3831,N_3948);
nand U4488 (N_4488,N_3792,N_3498);
nand U4489 (N_4489,N_3420,N_3503);
xnor U4490 (N_4490,N_3708,N_3926);
or U4491 (N_4491,N_3274,N_3445);
and U4492 (N_4492,N_3718,N_3685);
nand U4493 (N_4493,N_3964,N_3624);
or U4494 (N_4494,N_3321,N_3994);
nor U4495 (N_4495,N_3685,N_3617);
nand U4496 (N_4496,N_3358,N_3796);
nor U4497 (N_4497,N_3701,N_3852);
xor U4498 (N_4498,N_3399,N_3437);
xnor U4499 (N_4499,N_3875,N_3336);
nand U4500 (N_4500,N_3677,N_3864);
xor U4501 (N_4501,N_3743,N_3425);
xor U4502 (N_4502,N_3327,N_3905);
or U4503 (N_4503,N_3632,N_3712);
or U4504 (N_4504,N_3697,N_3302);
or U4505 (N_4505,N_3896,N_3257);
or U4506 (N_4506,N_3352,N_3860);
xnor U4507 (N_4507,N_3808,N_3527);
nor U4508 (N_4508,N_3600,N_3453);
and U4509 (N_4509,N_3399,N_3249);
or U4510 (N_4510,N_3451,N_3804);
and U4511 (N_4511,N_3682,N_3434);
or U4512 (N_4512,N_3506,N_3968);
and U4513 (N_4513,N_3688,N_3634);
xor U4514 (N_4514,N_3263,N_3300);
nand U4515 (N_4515,N_3498,N_3781);
or U4516 (N_4516,N_3696,N_3860);
nand U4517 (N_4517,N_3977,N_3446);
nor U4518 (N_4518,N_3940,N_3287);
and U4519 (N_4519,N_3797,N_3621);
or U4520 (N_4520,N_3937,N_3893);
nor U4521 (N_4521,N_3362,N_3679);
nand U4522 (N_4522,N_3293,N_3570);
and U4523 (N_4523,N_3807,N_3221);
nor U4524 (N_4524,N_3244,N_3299);
nand U4525 (N_4525,N_3235,N_3658);
xor U4526 (N_4526,N_3337,N_3607);
nand U4527 (N_4527,N_3785,N_3746);
xnor U4528 (N_4528,N_3596,N_3798);
nor U4529 (N_4529,N_3962,N_3997);
or U4530 (N_4530,N_3847,N_3707);
nand U4531 (N_4531,N_3705,N_3954);
and U4532 (N_4532,N_3582,N_3322);
or U4533 (N_4533,N_3306,N_3777);
and U4534 (N_4534,N_3615,N_3937);
nor U4535 (N_4535,N_3442,N_3794);
nor U4536 (N_4536,N_3706,N_3385);
nand U4537 (N_4537,N_3497,N_3980);
nor U4538 (N_4538,N_3911,N_3484);
or U4539 (N_4539,N_3699,N_3208);
nand U4540 (N_4540,N_3244,N_3371);
and U4541 (N_4541,N_3562,N_3929);
or U4542 (N_4542,N_3373,N_3849);
or U4543 (N_4543,N_3697,N_3738);
and U4544 (N_4544,N_3429,N_3822);
or U4545 (N_4545,N_3314,N_3358);
nand U4546 (N_4546,N_3223,N_3538);
or U4547 (N_4547,N_3448,N_3878);
xnor U4548 (N_4548,N_3334,N_3989);
nor U4549 (N_4549,N_3533,N_3318);
xor U4550 (N_4550,N_3517,N_3776);
and U4551 (N_4551,N_3306,N_3281);
and U4552 (N_4552,N_3996,N_3640);
xor U4553 (N_4553,N_3653,N_3267);
and U4554 (N_4554,N_3221,N_3999);
or U4555 (N_4555,N_3350,N_3979);
nor U4556 (N_4556,N_3727,N_3843);
xor U4557 (N_4557,N_3555,N_3681);
xnor U4558 (N_4558,N_3931,N_3879);
nor U4559 (N_4559,N_3873,N_3694);
nor U4560 (N_4560,N_3972,N_3850);
xor U4561 (N_4561,N_3689,N_3741);
nand U4562 (N_4562,N_3975,N_3564);
and U4563 (N_4563,N_3510,N_3800);
and U4564 (N_4564,N_3789,N_3626);
and U4565 (N_4565,N_3744,N_3728);
or U4566 (N_4566,N_3636,N_3520);
or U4567 (N_4567,N_3602,N_3583);
and U4568 (N_4568,N_3214,N_3479);
nand U4569 (N_4569,N_3463,N_3580);
nand U4570 (N_4570,N_3636,N_3863);
or U4571 (N_4571,N_3512,N_3561);
xor U4572 (N_4572,N_3887,N_3503);
and U4573 (N_4573,N_3557,N_3332);
and U4574 (N_4574,N_3352,N_3210);
or U4575 (N_4575,N_3774,N_3202);
xnor U4576 (N_4576,N_3350,N_3993);
and U4577 (N_4577,N_3369,N_3875);
nand U4578 (N_4578,N_3320,N_3593);
xnor U4579 (N_4579,N_3808,N_3889);
nand U4580 (N_4580,N_3671,N_3448);
or U4581 (N_4581,N_3689,N_3612);
and U4582 (N_4582,N_3587,N_3640);
xnor U4583 (N_4583,N_3951,N_3749);
or U4584 (N_4584,N_3220,N_3998);
xor U4585 (N_4585,N_3929,N_3378);
nor U4586 (N_4586,N_3377,N_3807);
and U4587 (N_4587,N_3572,N_3547);
and U4588 (N_4588,N_3383,N_3905);
nand U4589 (N_4589,N_3380,N_3707);
xnor U4590 (N_4590,N_3275,N_3333);
nor U4591 (N_4591,N_3837,N_3981);
nand U4592 (N_4592,N_3769,N_3578);
nand U4593 (N_4593,N_3904,N_3416);
xor U4594 (N_4594,N_3227,N_3494);
xnor U4595 (N_4595,N_3717,N_3508);
nor U4596 (N_4596,N_3883,N_3993);
xnor U4597 (N_4597,N_3681,N_3302);
or U4598 (N_4598,N_3580,N_3772);
nand U4599 (N_4599,N_3919,N_3530);
or U4600 (N_4600,N_3218,N_3954);
nor U4601 (N_4601,N_3477,N_3244);
xnor U4602 (N_4602,N_3691,N_3882);
xor U4603 (N_4603,N_3900,N_3802);
nor U4604 (N_4604,N_3859,N_3244);
nand U4605 (N_4605,N_3357,N_3283);
xnor U4606 (N_4606,N_3678,N_3414);
nand U4607 (N_4607,N_3390,N_3590);
and U4608 (N_4608,N_3338,N_3981);
nand U4609 (N_4609,N_3363,N_3678);
or U4610 (N_4610,N_3955,N_3571);
and U4611 (N_4611,N_3830,N_3768);
or U4612 (N_4612,N_3659,N_3272);
nand U4613 (N_4613,N_3669,N_3639);
or U4614 (N_4614,N_3690,N_3777);
or U4615 (N_4615,N_3810,N_3213);
nor U4616 (N_4616,N_3487,N_3428);
and U4617 (N_4617,N_3785,N_3620);
nand U4618 (N_4618,N_3256,N_3644);
and U4619 (N_4619,N_3446,N_3222);
or U4620 (N_4620,N_3401,N_3970);
xor U4621 (N_4621,N_3780,N_3292);
or U4622 (N_4622,N_3445,N_3272);
nand U4623 (N_4623,N_3260,N_3458);
nand U4624 (N_4624,N_3956,N_3891);
nor U4625 (N_4625,N_3882,N_3810);
xnor U4626 (N_4626,N_3407,N_3859);
or U4627 (N_4627,N_3797,N_3916);
nor U4628 (N_4628,N_3876,N_3380);
nand U4629 (N_4629,N_3983,N_3280);
nand U4630 (N_4630,N_3906,N_3482);
xor U4631 (N_4631,N_3928,N_3959);
and U4632 (N_4632,N_3938,N_3544);
nand U4633 (N_4633,N_3467,N_3942);
nor U4634 (N_4634,N_3966,N_3237);
or U4635 (N_4635,N_3229,N_3590);
xnor U4636 (N_4636,N_3961,N_3848);
and U4637 (N_4637,N_3738,N_3861);
and U4638 (N_4638,N_3766,N_3876);
or U4639 (N_4639,N_3527,N_3786);
xor U4640 (N_4640,N_3242,N_3744);
xor U4641 (N_4641,N_3348,N_3731);
nand U4642 (N_4642,N_3642,N_3576);
nor U4643 (N_4643,N_3561,N_3495);
nand U4644 (N_4644,N_3224,N_3758);
or U4645 (N_4645,N_3208,N_3847);
nor U4646 (N_4646,N_3820,N_3519);
or U4647 (N_4647,N_3384,N_3626);
nor U4648 (N_4648,N_3889,N_3986);
xor U4649 (N_4649,N_3702,N_3862);
or U4650 (N_4650,N_3667,N_3327);
or U4651 (N_4651,N_3776,N_3233);
xnor U4652 (N_4652,N_3251,N_3803);
and U4653 (N_4653,N_3379,N_3766);
and U4654 (N_4654,N_3870,N_3210);
nor U4655 (N_4655,N_3989,N_3782);
nand U4656 (N_4656,N_3360,N_3350);
xor U4657 (N_4657,N_3311,N_3213);
nand U4658 (N_4658,N_3991,N_3807);
and U4659 (N_4659,N_3764,N_3870);
nand U4660 (N_4660,N_3254,N_3416);
and U4661 (N_4661,N_3760,N_3518);
or U4662 (N_4662,N_3661,N_3952);
and U4663 (N_4663,N_3920,N_3338);
nand U4664 (N_4664,N_3432,N_3876);
nand U4665 (N_4665,N_3499,N_3574);
and U4666 (N_4666,N_3492,N_3427);
nand U4667 (N_4667,N_3919,N_3647);
and U4668 (N_4668,N_3343,N_3893);
and U4669 (N_4669,N_3581,N_3410);
nand U4670 (N_4670,N_3512,N_3737);
nor U4671 (N_4671,N_3815,N_3522);
xor U4672 (N_4672,N_3689,N_3351);
nor U4673 (N_4673,N_3791,N_3779);
and U4674 (N_4674,N_3636,N_3631);
nor U4675 (N_4675,N_3948,N_3827);
nor U4676 (N_4676,N_3803,N_3204);
nand U4677 (N_4677,N_3753,N_3807);
and U4678 (N_4678,N_3456,N_3748);
and U4679 (N_4679,N_3755,N_3869);
nor U4680 (N_4680,N_3549,N_3419);
nor U4681 (N_4681,N_3924,N_3940);
or U4682 (N_4682,N_3350,N_3534);
nor U4683 (N_4683,N_3768,N_3508);
nor U4684 (N_4684,N_3610,N_3598);
and U4685 (N_4685,N_3314,N_3495);
and U4686 (N_4686,N_3450,N_3628);
xor U4687 (N_4687,N_3834,N_3485);
nor U4688 (N_4688,N_3851,N_3291);
xor U4689 (N_4689,N_3697,N_3484);
or U4690 (N_4690,N_3804,N_3616);
nand U4691 (N_4691,N_3544,N_3592);
and U4692 (N_4692,N_3517,N_3340);
and U4693 (N_4693,N_3941,N_3831);
and U4694 (N_4694,N_3799,N_3340);
or U4695 (N_4695,N_3290,N_3722);
nor U4696 (N_4696,N_3513,N_3915);
or U4697 (N_4697,N_3787,N_3753);
nand U4698 (N_4698,N_3924,N_3235);
and U4699 (N_4699,N_3866,N_3734);
xnor U4700 (N_4700,N_3442,N_3495);
or U4701 (N_4701,N_3385,N_3222);
nand U4702 (N_4702,N_3883,N_3894);
nand U4703 (N_4703,N_3491,N_3692);
nand U4704 (N_4704,N_3811,N_3915);
and U4705 (N_4705,N_3225,N_3783);
or U4706 (N_4706,N_3253,N_3712);
or U4707 (N_4707,N_3594,N_3879);
and U4708 (N_4708,N_3915,N_3858);
nand U4709 (N_4709,N_3914,N_3695);
nor U4710 (N_4710,N_3885,N_3371);
and U4711 (N_4711,N_3230,N_3851);
and U4712 (N_4712,N_3917,N_3878);
and U4713 (N_4713,N_3447,N_3515);
xnor U4714 (N_4714,N_3274,N_3271);
nand U4715 (N_4715,N_3657,N_3945);
or U4716 (N_4716,N_3312,N_3752);
and U4717 (N_4717,N_3244,N_3675);
or U4718 (N_4718,N_3444,N_3267);
nand U4719 (N_4719,N_3225,N_3400);
nor U4720 (N_4720,N_3692,N_3559);
nand U4721 (N_4721,N_3974,N_3833);
nand U4722 (N_4722,N_3293,N_3376);
and U4723 (N_4723,N_3885,N_3416);
or U4724 (N_4724,N_3738,N_3607);
nor U4725 (N_4725,N_3268,N_3516);
or U4726 (N_4726,N_3617,N_3782);
or U4727 (N_4727,N_3846,N_3387);
and U4728 (N_4728,N_3297,N_3973);
or U4729 (N_4729,N_3827,N_3521);
or U4730 (N_4730,N_3243,N_3771);
xor U4731 (N_4731,N_3649,N_3203);
and U4732 (N_4732,N_3415,N_3468);
nand U4733 (N_4733,N_3501,N_3899);
xor U4734 (N_4734,N_3360,N_3245);
nor U4735 (N_4735,N_3528,N_3486);
nand U4736 (N_4736,N_3409,N_3450);
and U4737 (N_4737,N_3838,N_3541);
nand U4738 (N_4738,N_3724,N_3961);
nand U4739 (N_4739,N_3460,N_3618);
nor U4740 (N_4740,N_3801,N_3263);
nand U4741 (N_4741,N_3649,N_3801);
xnor U4742 (N_4742,N_3422,N_3564);
and U4743 (N_4743,N_3354,N_3909);
or U4744 (N_4744,N_3383,N_3835);
and U4745 (N_4745,N_3674,N_3537);
nor U4746 (N_4746,N_3730,N_3420);
or U4747 (N_4747,N_3643,N_3231);
nand U4748 (N_4748,N_3227,N_3768);
nor U4749 (N_4749,N_3714,N_3528);
nand U4750 (N_4750,N_3734,N_3909);
or U4751 (N_4751,N_3853,N_3697);
nand U4752 (N_4752,N_3435,N_3517);
nand U4753 (N_4753,N_3225,N_3269);
or U4754 (N_4754,N_3308,N_3888);
nand U4755 (N_4755,N_3816,N_3542);
or U4756 (N_4756,N_3498,N_3829);
and U4757 (N_4757,N_3486,N_3315);
nor U4758 (N_4758,N_3831,N_3542);
xnor U4759 (N_4759,N_3272,N_3726);
or U4760 (N_4760,N_3989,N_3865);
nand U4761 (N_4761,N_3687,N_3732);
and U4762 (N_4762,N_3387,N_3319);
nor U4763 (N_4763,N_3482,N_3235);
and U4764 (N_4764,N_3992,N_3459);
or U4765 (N_4765,N_3386,N_3451);
nor U4766 (N_4766,N_3886,N_3703);
nand U4767 (N_4767,N_3876,N_3475);
nand U4768 (N_4768,N_3539,N_3254);
nand U4769 (N_4769,N_3427,N_3961);
or U4770 (N_4770,N_3837,N_3617);
xnor U4771 (N_4771,N_3564,N_3614);
nor U4772 (N_4772,N_3230,N_3507);
nand U4773 (N_4773,N_3322,N_3440);
or U4774 (N_4774,N_3323,N_3200);
nor U4775 (N_4775,N_3720,N_3313);
and U4776 (N_4776,N_3780,N_3712);
xnor U4777 (N_4777,N_3835,N_3327);
nand U4778 (N_4778,N_3533,N_3216);
and U4779 (N_4779,N_3819,N_3501);
nand U4780 (N_4780,N_3710,N_3854);
or U4781 (N_4781,N_3295,N_3826);
and U4782 (N_4782,N_3936,N_3207);
nand U4783 (N_4783,N_3415,N_3487);
nand U4784 (N_4784,N_3466,N_3259);
or U4785 (N_4785,N_3500,N_3323);
and U4786 (N_4786,N_3567,N_3566);
or U4787 (N_4787,N_3293,N_3775);
or U4788 (N_4788,N_3634,N_3703);
nor U4789 (N_4789,N_3319,N_3753);
nand U4790 (N_4790,N_3921,N_3437);
nor U4791 (N_4791,N_3740,N_3279);
nor U4792 (N_4792,N_3498,N_3924);
xor U4793 (N_4793,N_3803,N_3944);
nand U4794 (N_4794,N_3901,N_3442);
nor U4795 (N_4795,N_3538,N_3790);
or U4796 (N_4796,N_3678,N_3437);
and U4797 (N_4797,N_3684,N_3953);
and U4798 (N_4798,N_3935,N_3461);
and U4799 (N_4799,N_3296,N_3402);
nand U4800 (N_4800,N_4696,N_4374);
nor U4801 (N_4801,N_4220,N_4723);
nor U4802 (N_4802,N_4674,N_4380);
xor U4803 (N_4803,N_4728,N_4055);
xnor U4804 (N_4804,N_4050,N_4518);
nor U4805 (N_4805,N_4252,N_4517);
xnor U4806 (N_4806,N_4030,N_4415);
nand U4807 (N_4807,N_4065,N_4604);
nand U4808 (N_4808,N_4348,N_4179);
xor U4809 (N_4809,N_4642,N_4624);
nand U4810 (N_4810,N_4231,N_4289);
nand U4811 (N_4811,N_4207,N_4101);
and U4812 (N_4812,N_4791,N_4568);
nor U4813 (N_4813,N_4532,N_4554);
xnor U4814 (N_4814,N_4106,N_4447);
nand U4815 (N_4815,N_4639,N_4197);
nand U4816 (N_4816,N_4109,N_4602);
nand U4817 (N_4817,N_4435,N_4364);
or U4818 (N_4818,N_4031,N_4796);
xor U4819 (N_4819,N_4583,N_4720);
nor U4820 (N_4820,N_4641,N_4706);
and U4821 (N_4821,N_4680,N_4499);
and U4822 (N_4822,N_4349,N_4760);
or U4823 (N_4823,N_4362,N_4779);
or U4824 (N_4824,N_4066,N_4020);
xnor U4825 (N_4825,N_4169,N_4749);
nor U4826 (N_4826,N_4300,N_4411);
xnor U4827 (N_4827,N_4438,N_4450);
nor U4828 (N_4828,N_4341,N_4318);
nand U4829 (N_4829,N_4320,N_4730);
nand U4830 (N_4830,N_4214,N_4340);
nor U4831 (N_4831,N_4594,N_4168);
or U4832 (N_4832,N_4549,N_4162);
xnor U4833 (N_4833,N_4500,N_4471);
and U4834 (N_4834,N_4607,N_4304);
xor U4835 (N_4835,N_4528,N_4539);
xnor U4836 (N_4836,N_4385,N_4427);
xnor U4837 (N_4837,N_4714,N_4482);
nand U4838 (N_4838,N_4381,N_4149);
nand U4839 (N_4839,N_4068,N_4275);
nand U4840 (N_4840,N_4461,N_4000);
xnor U4841 (N_4841,N_4196,N_4069);
or U4842 (N_4842,N_4244,N_4799);
xnor U4843 (N_4843,N_4130,N_4224);
nand U4844 (N_4844,N_4459,N_4648);
nor U4845 (N_4845,N_4748,N_4126);
or U4846 (N_4846,N_4384,N_4294);
xnor U4847 (N_4847,N_4090,N_4012);
or U4848 (N_4848,N_4710,N_4632);
or U4849 (N_4849,N_4329,N_4584);
or U4850 (N_4850,N_4394,N_4232);
and U4851 (N_4851,N_4306,N_4444);
nand U4852 (N_4852,N_4638,N_4565);
xnor U4853 (N_4853,N_4047,N_4504);
nand U4854 (N_4854,N_4228,N_4070);
nand U4855 (N_4855,N_4146,N_4413);
nand U4856 (N_4856,N_4293,N_4316);
or U4857 (N_4857,N_4110,N_4009);
or U4858 (N_4858,N_4344,N_4431);
and U4859 (N_4859,N_4650,N_4049);
nand U4860 (N_4860,N_4083,N_4789);
nand U4861 (N_4861,N_4201,N_4524);
nor U4862 (N_4862,N_4735,N_4592);
nand U4863 (N_4863,N_4614,N_4354);
nand U4864 (N_4864,N_4111,N_4682);
and U4865 (N_4865,N_4002,N_4451);
xnor U4866 (N_4866,N_4357,N_4781);
nand U4867 (N_4867,N_4376,N_4661);
nor U4868 (N_4868,N_4627,N_4597);
nor U4869 (N_4869,N_4278,N_4393);
xnor U4870 (N_4870,N_4025,N_4040);
nand U4871 (N_4871,N_4046,N_4345);
and U4872 (N_4872,N_4725,N_4460);
nand U4873 (N_4873,N_4563,N_4608);
or U4874 (N_4874,N_4474,N_4056);
and U4875 (N_4875,N_4437,N_4022);
nor U4876 (N_4876,N_4319,N_4335);
xnor U4877 (N_4877,N_4405,N_4693);
nor U4878 (N_4878,N_4519,N_4425);
nor U4879 (N_4879,N_4079,N_4062);
xor U4880 (N_4880,N_4326,N_4315);
nand U4881 (N_4881,N_4262,N_4476);
xor U4882 (N_4882,N_4314,N_4082);
or U4883 (N_4883,N_4077,N_4239);
xor U4884 (N_4884,N_4378,N_4103);
nor U4885 (N_4885,N_4338,N_4123);
xor U4886 (N_4886,N_4339,N_4057);
nor U4887 (N_4887,N_4783,N_4178);
xor U4888 (N_4888,N_4531,N_4593);
xor U4889 (N_4889,N_4147,N_4768);
and U4890 (N_4890,N_4653,N_4550);
and U4891 (N_4891,N_4193,N_4534);
nor U4892 (N_4892,N_4507,N_4671);
xnor U4893 (N_4893,N_4521,N_4657);
nand U4894 (N_4894,N_4729,N_4154);
nor U4895 (N_4895,N_4698,N_4288);
or U4896 (N_4896,N_4757,N_4449);
and U4897 (N_4897,N_4184,N_4241);
or U4898 (N_4898,N_4076,N_4173);
nand U4899 (N_4899,N_4390,N_4058);
nor U4900 (N_4900,N_4481,N_4259);
or U4901 (N_4901,N_4309,N_4677);
nor U4902 (N_4902,N_4439,N_4466);
nand U4903 (N_4903,N_4522,N_4770);
and U4904 (N_4904,N_4051,N_4436);
xor U4905 (N_4905,N_4033,N_4547);
nand U4906 (N_4906,N_4143,N_4257);
or U4907 (N_4907,N_4733,N_4701);
and U4908 (N_4908,N_4700,N_4115);
nand U4909 (N_4909,N_4406,N_4412);
or U4910 (N_4910,N_4586,N_4073);
nand U4911 (N_4911,N_4401,N_4104);
xnor U4912 (N_4912,N_4323,N_4689);
xnor U4913 (N_4913,N_4633,N_4595);
nor U4914 (N_4914,N_4129,N_4113);
or U4915 (N_4915,N_4359,N_4313);
or U4916 (N_4916,N_4067,N_4268);
xor U4917 (N_4917,N_4238,N_4330);
or U4918 (N_4918,N_4221,N_4656);
nor U4919 (N_4919,N_4777,N_4216);
nor U4920 (N_4920,N_4759,N_4208);
and U4921 (N_4921,N_4135,N_4538);
xnor U4922 (N_4922,N_4310,N_4395);
xnor U4923 (N_4923,N_4151,N_4703);
nand U4924 (N_4924,N_4236,N_4643);
nor U4925 (N_4925,N_4561,N_4285);
and U4926 (N_4926,N_4097,N_4114);
nand U4927 (N_4927,N_4276,N_4774);
nor U4928 (N_4928,N_4102,N_4631);
nand U4929 (N_4929,N_4303,N_4124);
and U4930 (N_4930,N_4765,N_4486);
and U4931 (N_4931,N_4053,N_4520);
or U4932 (N_4932,N_4496,N_4074);
nand U4933 (N_4933,N_4121,N_4613);
nor U4934 (N_4934,N_4089,N_4156);
or U4935 (N_4935,N_4694,N_4665);
and U4936 (N_4936,N_4229,N_4287);
nor U4937 (N_4937,N_4249,N_4226);
nand U4938 (N_4938,N_4211,N_4060);
xnor U4939 (N_4939,N_4098,N_4469);
nor U4940 (N_4940,N_4695,N_4599);
and U4941 (N_4941,N_4322,N_4553);
nor U4942 (N_4942,N_4297,N_4416);
or U4943 (N_4943,N_4709,N_4014);
or U4944 (N_4944,N_4574,N_4116);
nand U4945 (N_4945,N_4426,N_4576);
and U4946 (N_4946,N_4776,N_4204);
or U4947 (N_4947,N_4254,N_4533);
nand U4948 (N_4948,N_4036,N_4332);
or U4949 (N_4949,N_4095,N_4718);
and U4950 (N_4950,N_4542,N_4407);
nor U4951 (N_4951,N_4170,N_4756);
nor U4952 (N_4952,N_4564,N_4203);
nand U4953 (N_4953,N_4324,N_4778);
or U4954 (N_4954,N_4664,N_4029);
nor U4955 (N_4955,N_4468,N_4096);
nand U4956 (N_4956,N_4587,N_4446);
nand U4957 (N_4957,N_4198,N_4346);
and U4958 (N_4958,N_4152,N_4489);
or U4959 (N_4959,N_4708,N_4064);
xnor U4960 (N_4960,N_4573,N_4750);
nand U4961 (N_4961,N_4240,N_4356);
and U4962 (N_4962,N_4286,N_4045);
and U4963 (N_4963,N_4630,N_4782);
or U4964 (N_4964,N_4371,N_4589);
and U4965 (N_4965,N_4080,N_4711);
or U4966 (N_4966,N_4491,N_4141);
and U4967 (N_4967,N_4609,N_4744);
and U4968 (N_4968,N_4365,N_4127);
or U4969 (N_4969,N_4150,N_4397);
nor U4970 (N_4970,N_4277,N_4290);
and U4971 (N_4971,N_4334,N_4299);
and U4972 (N_4972,N_4495,N_4005);
nor U4973 (N_4973,N_4041,N_4336);
or U4974 (N_4974,N_4683,N_4758);
nand U4975 (N_4975,N_4190,N_4525);
nor U4976 (N_4976,N_4256,N_4235);
or U4977 (N_4977,N_4562,N_4185);
nand U4978 (N_4978,N_4699,N_4479);
or U4979 (N_4979,N_4158,N_4727);
or U4980 (N_4980,N_4516,N_4175);
or U4981 (N_4981,N_4445,N_4472);
nand U4982 (N_4982,N_4131,N_4668);
and U4983 (N_4983,N_4387,N_4086);
or U4984 (N_4984,N_4537,N_4503);
xnor U4985 (N_4985,N_4751,N_4745);
nand U4986 (N_4986,N_4477,N_4351);
xnor U4987 (N_4987,N_4579,N_4059);
or U4988 (N_4988,N_4128,N_4464);
xor U4989 (N_4989,N_4172,N_4717);
or U4990 (N_4990,N_4003,N_4629);
nand U4991 (N_4991,N_4093,N_4785);
xor U4992 (N_4992,N_4148,N_4355);
and U4993 (N_4993,N_4763,N_4429);
and U4994 (N_4994,N_4263,N_4223);
or U4995 (N_4995,N_4566,N_4155);
nor U4996 (N_4996,N_4672,N_4042);
or U4997 (N_4997,N_4456,N_4492);
nor U4998 (N_4998,N_4747,N_4467);
and U4999 (N_4999,N_4105,N_4515);
and U5000 (N_5000,N_4743,N_4205);
or U5001 (N_5001,N_4081,N_4245);
or U5002 (N_5002,N_4506,N_4398);
nand U5003 (N_5003,N_4795,N_4498);
nand U5004 (N_5004,N_4337,N_4623);
nor U5005 (N_5005,N_4494,N_4176);
or U5006 (N_5006,N_4473,N_4248);
nand U5007 (N_5007,N_4139,N_4400);
xor U5008 (N_5008,N_4659,N_4685);
or U5009 (N_5009,N_4122,N_4026);
nor U5010 (N_5010,N_4258,N_4452);
nor U5011 (N_5011,N_4389,N_4575);
nand U5012 (N_5012,N_4511,N_4626);
nor U5013 (N_5013,N_4660,N_4513);
nor U5014 (N_5014,N_4775,N_4188);
nor U5015 (N_5015,N_4048,N_4753);
or U5016 (N_5016,N_4755,N_4296);
nand U5017 (N_5017,N_4410,N_4418);
and U5018 (N_5018,N_4360,N_4582);
xnor U5019 (N_5019,N_4443,N_4577);
or U5020 (N_5020,N_4353,N_4291);
xor U5021 (N_5021,N_4737,N_4612);
xor U5022 (N_5022,N_4616,N_4430);
or U5023 (N_5023,N_4343,N_4493);
nor U5024 (N_5024,N_4132,N_4171);
nor U5025 (N_5025,N_4716,N_4075);
and U5026 (N_5026,N_4250,N_4361);
xor U5027 (N_5027,N_4502,N_4687);
and U5028 (N_5028,N_4788,N_4707);
and U5029 (N_5029,N_4219,N_4120);
xor U5030 (N_5030,N_4658,N_4217);
xnor U5031 (N_5031,N_4581,N_4637);
or U5032 (N_5032,N_4724,N_4043);
xor U5033 (N_5033,N_4536,N_4265);
and U5034 (N_5034,N_4780,N_4761);
xor U5035 (N_5035,N_4292,N_4433);
or U5036 (N_5036,N_4386,N_4237);
and U5037 (N_5037,N_4794,N_4331);
or U5038 (N_5038,N_4636,N_4600);
nand U5039 (N_5039,N_4734,N_4261);
nor U5040 (N_5040,N_4308,N_4367);
and U5041 (N_5041,N_4792,N_4571);
and U5042 (N_5042,N_4167,N_4307);
nand U5043 (N_5043,N_4557,N_4010);
xnor U5044 (N_5044,N_4015,N_4434);
nor U5045 (N_5045,N_4271,N_4166);
xor U5046 (N_5046,N_4771,N_4373);
and U5047 (N_5047,N_4181,N_4125);
or U5048 (N_5048,N_4704,N_4118);
and U5049 (N_5049,N_4117,N_4061);
nand U5050 (N_5050,N_4560,N_4305);
xnor U5051 (N_5051,N_4767,N_4325);
xor U5052 (N_5052,N_4312,N_4606);
and U5053 (N_5053,N_4580,N_4342);
nor U5054 (N_5054,N_4255,N_4282);
and U5055 (N_5055,N_4684,N_4691);
nor U5056 (N_5056,N_4501,N_4016);
xnor U5057 (N_5057,N_4423,N_4647);
xor U5058 (N_5058,N_4283,N_4454);
xnor U5059 (N_5059,N_4008,N_4243);
or U5060 (N_5060,N_4601,N_4621);
and U5061 (N_5061,N_4272,N_4402);
or U5062 (N_5062,N_4741,N_4797);
and U5063 (N_5063,N_4462,N_4508);
and U5064 (N_5064,N_4526,N_4281);
nand U5065 (N_5065,N_4414,N_4269);
or U5066 (N_5066,N_4295,N_4368);
or U5067 (N_5067,N_4620,N_4651);
or U5068 (N_5068,N_4625,N_4404);
or U5069 (N_5069,N_4654,N_4591);
nand U5070 (N_5070,N_4352,N_4037);
nor U5071 (N_5071,N_4738,N_4142);
or U5072 (N_5072,N_4182,N_4382);
nand U5073 (N_5073,N_4399,N_4543);
or U5074 (N_5074,N_4350,N_4100);
and U5075 (N_5075,N_4087,N_4273);
nor U5076 (N_5076,N_4408,N_4164);
and U5077 (N_5077,N_4686,N_4448);
nand U5078 (N_5078,N_4705,N_4676);
or U5079 (N_5079,N_4752,N_4690);
xor U5080 (N_5080,N_4212,N_4279);
and U5081 (N_5081,N_4530,N_4375);
nor U5082 (N_5082,N_4209,N_4153);
xor U5083 (N_5083,N_4596,N_4715);
and U5084 (N_5084,N_4321,N_4260);
nand U5085 (N_5085,N_4773,N_4327);
xnor U5086 (N_5086,N_4253,N_4112);
nor U5087 (N_5087,N_4731,N_4509);
nand U5088 (N_5088,N_4721,N_4719);
nor U5089 (N_5089,N_4039,N_4634);
or U5090 (N_5090,N_4044,N_4035);
and U5091 (N_5091,N_4006,N_4480);
and U5092 (N_5092,N_4535,N_4652);
nor U5093 (N_5093,N_4552,N_4617);
nand U5094 (N_5094,N_4740,N_4267);
or U5095 (N_5095,N_4163,N_4001);
and U5096 (N_5096,N_4183,N_4567);
nand U5097 (N_5097,N_4514,N_4189);
or U5098 (N_5098,N_4663,N_4284);
nand U5099 (N_5099,N_4088,N_4266);
nand U5100 (N_5100,N_4545,N_4742);
or U5101 (N_5101,N_4505,N_4546);
xor U5102 (N_5102,N_4274,N_4071);
nand U5103 (N_5103,N_4754,N_4301);
or U5104 (N_5104,N_4085,N_4165);
and U5105 (N_5105,N_4739,N_4570);
or U5106 (N_5106,N_4218,N_4442);
xnor U5107 (N_5107,N_4688,N_4569);
and U5108 (N_5108,N_4475,N_4034);
xor U5109 (N_5109,N_4157,N_4403);
nor U5110 (N_5110,N_4108,N_4007);
and U5111 (N_5111,N_4107,N_4054);
nor U5112 (N_5112,N_4619,N_4023);
nand U5113 (N_5113,N_4667,N_4424);
xnor U5114 (N_5114,N_4251,N_4497);
nand U5115 (N_5115,N_4798,N_4541);
nand U5116 (N_5116,N_4697,N_4333);
and U5117 (N_5117,N_4302,N_4644);
or U5118 (N_5118,N_4488,N_4572);
nor U5119 (N_5119,N_4366,N_4527);
nand U5120 (N_5120,N_4215,N_4038);
nor U5121 (N_5121,N_4544,N_4409);
nand U5122 (N_5122,N_4605,N_4523);
nand U5123 (N_5123,N_4463,N_4377);
or U5124 (N_5124,N_4242,N_4646);
xnor U5125 (N_5125,N_4787,N_4233);
or U5126 (N_5126,N_4793,N_4455);
and U5127 (N_5127,N_4790,N_4540);
nand U5128 (N_5128,N_4134,N_4227);
xor U5129 (N_5129,N_4712,N_4192);
nor U5130 (N_5130,N_4072,N_4666);
nand U5131 (N_5131,N_4421,N_4200);
nand U5132 (N_5132,N_4363,N_4160);
nor U5133 (N_5133,N_4032,N_4021);
xnor U5134 (N_5134,N_4432,N_4264);
xnor U5135 (N_5135,N_4191,N_4470);
nand U5136 (N_5136,N_4013,N_4487);
nand U5137 (N_5137,N_4670,N_4529);
nor U5138 (N_5138,N_4603,N_4186);
xor U5139 (N_5139,N_4512,N_4679);
or U5140 (N_5140,N_4347,N_4669);
nand U5141 (N_5141,N_4590,N_4210);
nor U5142 (N_5142,N_4772,N_4598);
nand U5143 (N_5143,N_4247,N_4556);
and U5144 (N_5144,N_4094,N_4024);
xor U5145 (N_5145,N_4372,N_4458);
and U5146 (N_5146,N_4298,N_4358);
and U5147 (N_5147,N_4769,N_4187);
and U5148 (N_5148,N_4317,N_4628);
nor U5149 (N_5149,N_4011,N_4388);
nor U5150 (N_5150,N_4091,N_4673);
xnor U5151 (N_5151,N_4180,N_4017);
xnor U5152 (N_5152,N_4052,N_4611);
or U5153 (N_5153,N_4558,N_4441);
or U5154 (N_5154,N_4280,N_4732);
and U5155 (N_5155,N_4610,N_4370);
or U5156 (N_5156,N_4174,N_4618);
and U5157 (N_5157,N_4206,N_4213);
xor U5158 (N_5158,N_4457,N_4391);
xnor U5159 (N_5159,N_4702,N_4484);
or U5160 (N_5160,N_4692,N_4551);
or U5161 (N_5161,N_4746,N_4202);
and U5162 (N_5162,N_4640,N_4225);
or U5163 (N_5163,N_4369,N_4490);
xor U5164 (N_5164,N_4027,N_4396);
or U5165 (N_5165,N_4578,N_4222);
nor U5166 (N_5166,N_4311,N_4440);
nand U5167 (N_5167,N_4028,N_4138);
and U5168 (N_5168,N_4084,N_4555);
nand U5169 (N_5169,N_4145,N_4063);
xor U5170 (N_5170,N_4655,N_4510);
nor U5171 (N_5171,N_4392,N_4133);
or U5172 (N_5172,N_4199,N_4736);
nand U5173 (N_5173,N_4328,N_4622);
xnor U5174 (N_5174,N_4270,N_4784);
nor U5175 (N_5175,N_4383,N_4675);
or U5176 (N_5176,N_4762,N_4018);
nor U5177 (N_5177,N_4478,N_4585);
nor U5178 (N_5178,N_4078,N_4194);
nand U5179 (N_5179,N_4004,N_4419);
and U5180 (N_5180,N_4649,N_4465);
or U5181 (N_5181,N_4417,N_4713);
or U5182 (N_5182,N_4483,N_4485);
or U5183 (N_5183,N_4422,N_4559);
nand U5184 (N_5184,N_4159,N_4420);
nand U5185 (N_5185,N_4678,N_4726);
nand U5186 (N_5186,N_4140,N_4766);
or U5187 (N_5187,N_4379,N_4177);
nand U5188 (N_5188,N_4230,N_4161);
or U5189 (N_5189,N_4615,N_4099);
and U5190 (N_5190,N_4092,N_4548);
or U5191 (N_5191,N_4662,N_4786);
or U5192 (N_5192,N_4136,N_4137);
xnor U5193 (N_5193,N_4195,N_4635);
nand U5194 (N_5194,N_4119,N_4428);
nand U5195 (N_5195,N_4453,N_4588);
and U5196 (N_5196,N_4722,N_4234);
and U5197 (N_5197,N_4764,N_4246);
nor U5198 (N_5198,N_4681,N_4645);
nand U5199 (N_5199,N_4019,N_4144);
nor U5200 (N_5200,N_4312,N_4333);
xor U5201 (N_5201,N_4397,N_4155);
and U5202 (N_5202,N_4567,N_4592);
or U5203 (N_5203,N_4242,N_4035);
nor U5204 (N_5204,N_4727,N_4525);
and U5205 (N_5205,N_4128,N_4100);
and U5206 (N_5206,N_4101,N_4568);
or U5207 (N_5207,N_4732,N_4657);
nand U5208 (N_5208,N_4154,N_4174);
nand U5209 (N_5209,N_4526,N_4658);
or U5210 (N_5210,N_4027,N_4435);
or U5211 (N_5211,N_4374,N_4701);
nand U5212 (N_5212,N_4295,N_4573);
xnor U5213 (N_5213,N_4324,N_4293);
or U5214 (N_5214,N_4730,N_4338);
xor U5215 (N_5215,N_4177,N_4016);
or U5216 (N_5216,N_4374,N_4664);
nand U5217 (N_5217,N_4286,N_4071);
nor U5218 (N_5218,N_4482,N_4510);
nand U5219 (N_5219,N_4638,N_4504);
xor U5220 (N_5220,N_4329,N_4121);
nor U5221 (N_5221,N_4733,N_4329);
xor U5222 (N_5222,N_4007,N_4615);
nand U5223 (N_5223,N_4342,N_4454);
nand U5224 (N_5224,N_4739,N_4453);
nand U5225 (N_5225,N_4670,N_4676);
and U5226 (N_5226,N_4090,N_4507);
nor U5227 (N_5227,N_4388,N_4035);
nand U5228 (N_5228,N_4054,N_4778);
xor U5229 (N_5229,N_4743,N_4507);
xnor U5230 (N_5230,N_4530,N_4003);
or U5231 (N_5231,N_4032,N_4400);
nand U5232 (N_5232,N_4233,N_4092);
or U5233 (N_5233,N_4573,N_4063);
or U5234 (N_5234,N_4029,N_4095);
nand U5235 (N_5235,N_4762,N_4774);
xor U5236 (N_5236,N_4729,N_4715);
nand U5237 (N_5237,N_4337,N_4363);
nor U5238 (N_5238,N_4506,N_4389);
or U5239 (N_5239,N_4034,N_4504);
xor U5240 (N_5240,N_4554,N_4147);
nand U5241 (N_5241,N_4335,N_4428);
nand U5242 (N_5242,N_4011,N_4627);
or U5243 (N_5243,N_4014,N_4451);
xor U5244 (N_5244,N_4750,N_4297);
or U5245 (N_5245,N_4754,N_4636);
or U5246 (N_5246,N_4679,N_4744);
nand U5247 (N_5247,N_4110,N_4443);
or U5248 (N_5248,N_4593,N_4123);
xor U5249 (N_5249,N_4533,N_4601);
or U5250 (N_5250,N_4316,N_4131);
or U5251 (N_5251,N_4125,N_4278);
nor U5252 (N_5252,N_4648,N_4093);
nor U5253 (N_5253,N_4324,N_4671);
nand U5254 (N_5254,N_4293,N_4069);
xnor U5255 (N_5255,N_4525,N_4462);
nand U5256 (N_5256,N_4654,N_4202);
nor U5257 (N_5257,N_4470,N_4527);
and U5258 (N_5258,N_4150,N_4712);
and U5259 (N_5259,N_4426,N_4175);
nor U5260 (N_5260,N_4387,N_4684);
nor U5261 (N_5261,N_4650,N_4129);
nor U5262 (N_5262,N_4387,N_4789);
or U5263 (N_5263,N_4774,N_4547);
nor U5264 (N_5264,N_4042,N_4242);
and U5265 (N_5265,N_4207,N_4346);
or U5266 (N_5266,N_4303,N_4126);
or U5267 (N_5267,N_4219,N_4388);
xor U5268 (N_5268,N_4364,N_4104);
xor U5269 (N_5269,N_4343,N_4446);
nand U5270 (N_5270,N_4055,N_4124);
and U5271 (N_5271,N_4317,N_4493);
or U5272 (N_5272,N_4405,N_4182);
xor U5273 (N_5273,N_4784,N_4684);
xnor U5274 (N_5274,N_4572,N_4366);
and U5275 (N_5275,N_4176,N_4547);
or U5276 (N_5276,N_4780,N_4705);
nor U5277 (N_5277,N_4085,N_4020);
xnor U5278 (N_5278,N_4384,N_4568);
and U5279 (N_5279,N_4303,N_4155);
xnor U5280 (N_5280,N_4521,N_4227);
nand U5281 (N_5281,N_4722,N_4522);
xnor U5282 (N_5282,N_4521,N_4057);
nor U5283 (N_5283,N_4035,N_4218);
or U5284 (N_5284,N_4154,N_4096);
and U5285 (N_5285,N_4056,N_4402);
nand U5286 (N_5286,N_4561,N_4292);
nor U5287 (N_5287,N_4202,N_4570);
and U5288 (N_5288,N_4188,N_4725);
and U5289 (N_5289,N_4436,N_4773);
or U5290 (N_5290,N_4107,N_4068);
and U5291 (N_5291,N_4473,N_4562);
nand U5292 (N_5292,N_4051,N_4232);
nand U5293 (N_5293,N_4033,N_4302);
nor U5294 (N_5294,N_4401,N_4177);
nor U5295 (N_5295,N_4380,N_4555);
nor U5296 (N_5296,N_4530,N_4632);
xor U5297 (N_5297,N_4659,N_4029);
nor U5298 (N_5298,N_4137,N_4695);
and U5299 (N_5299,N_4559,N_4518);
and U5300 (N_5300,N_4610,N_4751);
and U5301 (N_5301,N_4449,N_4517);
and U5302 (N_5302,N_4116,N_4277);
or U5303 (N_5303,N_4182,N_4294);
xor U5304 (N_5304,N_4094,N_4198);
xnor U5305 (N_5305,N_4109,N_4202);
nand U5306 (N_5306,N_4618,N_4513);
nor U5307 (N_5307,N_4452,N_4055);
xor U5308 (N_5308,N_4188,N_4013);
xor U5309 (N_5309,N_4234,N_4377);
xnor U5310 (N_5310,N_4463,N_4407);
xor U5311 (N_5311,N_4076,N_4534);
nor U5312 (N_5312,N_4685,N_4772);
nor U5313 (N_5313,N_4520,N_4226);
nor U5314 (N_5314,N_4629,N_4278);
and U5315 (N_5315,N_4254,N_4257);
nor U5316 (N_5316,N_4103,N_4764);
or U5317 (N_5317,N_4406,N_4321);
and U5318 (N_5318,N_4627,N_4485);
and U5319 (N_5319,N_4201,N_4000);
xor U5320 (N_5320,N_4277,N_4300);
xor U5321 (N_5321,N_4715,N_4141);
or U5322 (N_5322,N_4158,N_4539);
or U5323 (N_5323,N_4115,N_4762);
nor U5324 (N_5324,N_4400,N_4176);
and U5325 (N_5325,N_4517,N_4174);
or U5326 (N_5326,N_4194,N_4757);
xnor U5327 (N_5327,N_4289,N_4528);
or U5328 (N_5328,N_4553,N_4279);
nor U5329 (N_5329,N_4097,N_4425);
or U5330 (N_5330,N_4157,N_4488);
or U5331 (N_5331,N_4465,N_4714);
or U5332 (N_5332,N_4576,N_4577);
and U5333 (N_5333,N_4707,N_4718);
and U5334 (N_5334,N_4786,N_4080);
and U5335 (N_5335,N_4596,N_4105);
and U5336 (N_5336,N_4644,N_4260);
xor U5337 (N_5337,N_4535,N_4599);
nor U5338 (N_5338,N_4498,N_4534);
nand U5339 (N_5339,N_4659,N_4422);
nor U5340 (N_5340,N_4576,N_4104);
or U5341 (N_5341,N_4413,N_4518);
or U5342 (N_5342,N_4701,N_4698);
nand U5343 (N_5343,N_4721,N_4173);
nand U5344 (N_5344,N_4652,N_4421);
and U5345 (N_5345,N_4702,N_4796);
or U5346 (N_5346,N_4171,N_4289);
xor U5347 (N_5347,N_4733,N_4218);
nor U5348 (N_5348,N_4259,N_4307);
xor U5349 (N_5349,N_4527,N_4168);
nor U5350 (N_5350,N_4262,N_4618);
and U5351 (N_5351,N_4363,N_4146);
and U5352 (N_5352,N_4096,N_4568);
nor U5353 (N_5353,N_4062,N_4552);
nor U5354 (N_5354,N_4305,N_4681);
xnor U5355 (N_5355,N_4254,N_4754);
nand U5356 (N_5356,N_4629,N_4137);
nand U5357 (N_5357,N_4024,N_4097);
nor U5358 (N_5358,N_4335,N_4245);
or U5359 (N_5359,N_4066,N_4144);
or U5360 (N_5360,N_4404,N_4144);
or U5361 (N_5361,N_4502,N_4647);
and U5362 (N_5362,N_4188,N_4665);
nand U5363 (N_5363,N_4590,N_4068);
nor U5364 (N_5364,N_4399,N_4693);
nand U5365 (N_5365,N_4014,N_4560);
or U5366 (N_5366,N_4495,N_4375);
nand U5367 (N_5367,N_4336,N_4234);
xor U5368 (N_5368,N_4392,N_4486);
nand U5369 (N_5369,N_4662,N_4380);
nor U5370 (N_5370,N_4624,N_4579);
and U5371 (N_5371,N_4717,N_4143);
or U5372 (N_5372,N_4168,N_4178);
nand U5373 (N_5373,N_4614,N_4468);
nor U5374 (N_5374,N_4661,N_4709);
xor U5375 (N_5375,N_4553,N_4224);
nor U5376 (N_5376,N_4088,N_4663);
nor U5377 (N_5377,N_4286,N_4763);
or U5378 (N_5378,N_4288,N_4057);
or U5379 (N_5379,N_4046,N_4326);
nand U5380 (N_5380,N_4228,N_4375);
or U5381 (N_5381,N_4559,N_4162);
nor U5382 (N_5382,N_4472,N_4191);
nand U5383 (N_5383,N_4430,N_4050);
or U5384 (N_5384,N_4507,N_4136);
or U5385 (N_5385,N_4436,N_4035);
nand U5386 (N_5386,N_4642,N_4360);
and U5387 (N_5387,N_4271,N_4291);
nand U5388 (N_5388,N_4208,N_4358);
nand U5389 (N_5389,N_4479,N_4058);
and U5390 (N_5390,N_4726,N_4428);
xor U5391 (N_5391,N_4779,N_4486);
nand U5392 (N_5392,N_4669,N_4767);
and U5393 (N_5393,N_4264,N_4485);
or U5394 (N_5394,N_4076,N_4317);
or U5395 (N_5395,N_4177,N_4733);
and U5396 (N_5396,N_4179,N_4779);
or U5397 (N_5397,N_4031,N_4798);
and U5398 (N_5398,N_4097,N_4433);
and U5399 (N_5399,N_4591,N_4725);
and U5400 (N_5400,N_4135,N_4159);
or U5401 (N_5401,N_4169,N_4468);
or U5402 (N_5402,N_4258,N_4132);
nor U5403 (N_5403,N_4502,N_4514);
and U5404 (N_5404,N_4316,N_4706);
nor U5405 (N_5405,N_4286,N_4172);
nand U5406 (N_5406,N_4366,N_4580);
xor U5407 (N_5407,N_4095,N_4547);
and U5408 (N_5408,N_4237,N_4069);
or U5409 (N_5409,N_4465,N_4318);
and U5410 (N_5410,N_4105,N_4297);
xor U5411 (N_5411,N_4513,N_4009);
or U5412 (N_5412,N_4736,N_4725);
or U5413 (N_5413,N_4629,N_4222);
nand U5414 (N_5414,N_4405,N_4799);
and U5415 (N_5415,N_4530,N_4403);
or U5416 (N_5416,N_4368,N_4611);
nor U5417 (N_5417,N_4778,N_4402);
xor U5418 (N_5418,N_4459,N_4161);
or U5419 (N_5419,N_4664,N_4341);
and U5420 (N_5420,N_4585,N_4218);
xor U5421 (N_5421,N_4304,N_4107);
and U5422 (N_5422,N_4573,N_4308);
nand U5423 (N_5423,N_4514,N_4388);
nor U5424 (N_5424,N_4276,N_4119);
xnor U5425 (N_5425,N_4084,N_4706);
nor U5426 (N_5426,N_4350,N_4692);
nor U5427 (N_5427,N_4099,N_4014);
nand U5428 (N_5428,N_4718,N_4261);
and U5429 (N_5429,N_4226,N_4572);
xnor U5430 (N_5430,N_4235,N_4429);
and U5431 (N_5431,N_4493,N_4592);
and U5432 (N_5432,N_4555,N_4378);
and U5433 (N_5433,N_4382,N_4331);
nor U5434 (N_5434,N_4519,N_4769);
xnor U5435 (N_5435,N_4140,N_4797);
and U5436 (N_5436,N_4589,N_4020);
nand U5437 (N_5437,N_4052,N_4441);
or U5438 (N_5438,N_4033,N_4658);
or U5439 (N_5439,N_4361,N_4436);
xnor U5440 (N_5440,N_4761,N_4574);
and U5441 (N_5441,N_4647,N_4089);
or U5442 (N_5442,N_4104,N_4732);
nor U5443 (N_5443,N_4706,N_4666);
nor U5444 (N_5444,N_4782,N_4699);
nand U5445 (N_5445,N_4396,N_4452);
or U5446 (N_5446,N_4415,N_4199);
nand U5447 (N_5447,N_4390,N_4152);
xnor U5448 (N_5448,N_4686,N_4321);
nand U5449 (N_5449,N_4444,N_4377);
and U5450 (N_5450,N_4573,N_4644);
nor U5451 (N_5451,N_4501,N_4731);
and U5452 (N_5452,N_4328,N_4576);
and U5453 (N_5453,N_4007,N_4289);
or U5454 (N_5454,N_4523,N_4209);
nor U5455 (N_5455,N_4792,N_4464);
nor U5456 (N_5456,N_4665,N_4282);
xor U5457 (N_5457,N_4115,N_4047);
nand U5458 (N_5458,N_4570,N_4628);
nand U5459 (N_5459,N_4065,N_4282);
nor U5460 (N_5460,N_4146,N_4222);
or U5461 (N_5461,N_4499,N_4792);
xor U5462 (N_5462,N_4529,N_4244);
nor U5463 (N_5463,N_4754,N_4577);
nand U5464 (N_5464,N_4727,N_4649);
or U5465 (N_5465,N_4545,N_4033);
or U5466 (N_5466,N_4489,N_4790);
nand U5467 (N_5467,N_4515,N_4360);
and U5468 (N_5468,N_4429,N_4702);
or U5469 (N_5469,N_4556,N_4474);
or U5470 (N_5470,N_4189,N_4734);
and U5471 (N_5471,N_4183,N_4232);
nor U5472 (N_5472,N_4627,N_4234);
nand U5473 (N_5473,N_4020,N_4733);
nand U5474 (N_5474,N_4484,N_4574);
nor U5475 (N_5475,N_4383,N_4748);
xnor U5476 (N_5476,N_4576,N_4644);
xnor U5477 (N_5477,N_4097,N_4389);
or U5478 (N_5478,N_4711,N_4646);
nor U5479 (N_5479,N_4291,N_4142);
nor U5480 (N_5480,N_4256,N_4046);
and U5481 (N_5481,N_4405,N_4564);
and U5482 (N_5482,N_4046,N_4539);
and U5483 (N_5483,N_4053,N_4398);
xnor U5484 (N_5484,N_4365,N_4402);
nor U5485 (N_5485,N_4331,N_4198);
xnor U5486 (N_5486,N_4531,N_4462);
and U5487 (N_5487,N_4283,N_4677);
nor U5488 (N_5488,N_4764,N_4784);
nor U5489 (N_5489,N_4082,N_4317);
xnor U5490 (N_5490,N_4014,N_4113);
xor U5491 (N_5491,N_4464,N_4335);
xor U5492 (N_5492,N_4559,N_4479);
xor U5493 (N_5493,N_4529,N_4351);
or U5494 (N_5494,N_4202,N_4498);
and U5495 (N_5495,N_4520,N_4775);
or U5496 (N_5496,N_4269,N_4567);
nor U5497 (N_5497,N_4747,N_4440);
xor U5498 (N_5498,N_4202,N_4403);
or U5499 (N_5499,N_4241,N_4645);
and U5500 (N_5500,N_4773,N_4652);
xor U5501 (N_5501,N_4314,N_4748);
xnor U5502 (N_5502,N_4678,N_4388);
nor U5503 (N_5503,N_4249,N_4472);
xor U5504 (N_5504,N_4524,N_4297);
and U5505 (N_5505,N_4764,N_4075);
xor U5506 (N_5506,N_4005,N_4456);
nor U5507 (N_5507,N_4479,N_4048);
nor U5508 (N_5508,N_4156,N_4072);
or U5509 (N_5509,N_4379,N_4063);
xor U5510 (N_5510,N_4188,N_4322);
nand U5511 (N_5511,N_4137,N_4126);
nor U5512 (N_5512,N_4761,N_4364);
nor U5513 (N_5513,N_4441,N_4235);
nand U5514 (N_5514,N_4761,N_4330);
nand U5515 (N_5515,N_4405,N_4785);
or U5516 (N_5516,N_4315,N_4591);
nor U5517 (N_5517,N_4120,N_4261);
nor U5518 (N_5518,N_4558,N_4581);
xor U5519 (N_5519,N_4095,N_4092);
and U5520 (N_5520,N_4380,N_4794);
nor U5521 (N_5521,N_4443,N_4423);
xor U5522 (N_5522,N_4133,N_4327);
and U5523 (N_5523,N_4327,N_4206);
and U5524 (N_5524,N_4005,N_4730);
xor U5525 (N_5525,N_4693,N_4544);
nor U5526 (N_5526,N_4474,N_4696);
xnor U5527 (N_5527,N_4479,N_4694);
or U5528 (N_5528,N_4499,N_4027);
or U5529 (N_5529,N_4540,N_4582);
nand U5530 (N_5530,N_4002,N_4600);
nor U5531 (N_5531,N_4411,N_4663);
and U5532 (N_5532,N_4143,N_4256);
xnor U5533 (N_5533,N_4647,N_4037);
and U5534 (N_5534,N_4606,N_4454);
nor U5535 (N_5535,N_4524,N_4156);
nand U5536 (N_5536,N_4406,N_4346);
nand U5537 (N_5537,N_4236,N_4731);
nand U5538 (N_5538,N_4014,N_4470);
xor U5539 (N_5539,N_4753,N_4142);
xor U5540 (N_5540,N_4095,N_4226);
and U5541 (N_5541,N_4576,N_4771);
nand U5542 (N_5542,N_4763,N_4282);
nand U5543 (N_5543,N_4718,N_4274);
nand U5544 (N_5544,N_4437,N_4295);
or U5545 (N_5545,N_4014,N_4545);
nor U5546 (N_5546,N_4561,N_4145);
xnor U5547 (N_5547,N_4026,N_4093);
or U5548 (N_5548,N_4337,N_4491);
nand U5549 (N_5549,N_4003,N_4033);
or U5550 (N_5550,N_4735,N_4406);
and U5551 (N_5551,N_4388,N_4207);
or U5552 (N_5552,N_4471,N_4741);
nand U5553 (N_5553,N_4532,N_4381);
nand U5554 (N_5554,N_4410,N_4234);
xor U5555 (N_5555,N_4300,N_4572);
nand U5556 (N_5556,N_4340,N_4188);
or U5557 (N_5557,N_4722,N_4070);
or U5558 (N_5558,N_4180,N_4123);
and U5559 (N_5559,N_4252,N_4186);
nor U5560 (N_5560,N_4749,N_4755);
xor U5561 (N_5561,N_4379,N_4621);
nor U5562 (N_5562,N_4126,N_4633);
and U5563 (N_5563,N_4445,N_4189);
and U5564 (N_5564,N_4590,N_4128);
nor U5565 (N_5565,N_4313,N_4242);
nor U5566 (N_5566,N_4176,N_4020);
or U5567 (N_5567,N_4340,N_4395);
and U5568 (N_5568,N_4408,N_4542);
and U5569 (N_5569,N_4081,N_4789);
nor U5570 (N_5570,N_4676,N_4629);
and U5571 (N_5571,N_4605,N_4018);
or U5572 (N_5572,N_4104,N_4477);
nor U5573 (N_5573,N_4585,N_4756);
and U5574 (N_5574,N_4570,N_4180);
nand U5575 (N_5575,N_4197,N_4681);
xnor U5576 (N_5576,N_4646,N_4659);
nor U5577 (N_5577,N_4010,N_4524);
and U5578 (N_5578,N_4118,N_4350);
or U5579 (N_5579,N_4635,N_4708);
nor U5580 (N_5580,N_4138,N_4216);
nand U5581 (N_5581,N_4586,N_4322);
nand U5582 (N_5582,N_4630,N_4320);
nor U5583 (N_5583,N_4602,N_4084);
or U5584 (N_5584,N_4245,N_4177);
nor U5585 (N_5585,N_4767,N_4080);
nand U5586 (N_5586,N_4337,N_4138);
xor U5587 (N_5587,N_4349,N_4422);
and U5588 (N_5588,N_4377,N_4783);
xnor U5589 (N_5589,N_4604,N_4735);
xnor U5590 (N_5590,N_4196,N_4015);
or U5591 (N_5591,N_4721,N_4159);
nor U5592 (N_5592,N_4544,N_4463);
xnor U5593 (N_5593,N_4659,N_4277);
or U5594 (N_5594,N_4491,N_4666);
or U5595 (N_5595,N_4359,N_4355);
nand U5596 (N_5596,N_4723,N_4575);
nand U5597 (N_5597,N_4135,N_4470);
or U5598 (N_5598,N_4494,N_4563);
or U5599 (N_5599,N_4365,N_4772);
nor U5600 (N_5600,N_4882,N_5535);
or U5601 (N_5601,N_4930,N_5049);
or U5602 (N_5602,N_4908,N_5136);
xnor U5603 (N_5603,N_5350,N_5352);
nand U5604 (N_5604,N_4949,N_5038);
nand U5605 (N_5605,N_5158,N_5400);
nand U5606 (N_5606,N_5058,N_5391);
nor U5607 (N_5607,N_4978,N_5495);
nand U5608 (N_5608,N_5433,N_5096);
xor U5609 (N_5609,N_5159,N_5057);
nor U5610 (N_5610,N_5178,N_5563);
and U5611 (N_5611,N_4818,N_5261);
nor U5612 (N_5612,N_4961,N_4827);
or U5613 (N_5613,N_5511,N_5526);
nor U5614 (N_5614,N_5365,N_4958);
or U5615 (N_5615,N_5104,N_5434);
and U5616 (N_5616,N_5556,N_4932);
nor U5617 (N_5617,N_4803,N_5233);
and U5618 (N_5618,N_4868,N_5152);
nor U5619 (N_5619,N_5203,N_5337);
xor U5620 (N_5620,N_5361,N_5368);
xor U5621 (N_5621,N_5354,N_5311);
nand U5622 (N_5622,N_5404,N_5305);
nor U5623 (N_5623,N_5297,N_5314);
or U5624 (N_5624,N_5224,N_4913);
or U5625 (N_5625,N_5216,N_4988);
nand U5626 (N_5626,N_5172,N_5397);
or U5627 (N_5627,N_4964,N_4843);
and U5628 (N_5628,N_5595,N_5174);
and U5629 (N_5629,N_5106,N_4973);
nand U5630 (N_5630,N_5582,N_5415);
or U5631 (N_5631,N_4983,N_5037);
and U5632 (N_5632,N_4885,N_5199);
nor U5633 (N_5633,N_4902,N_5270);
xor U5634 (N_5634,N_5528,N_5088);
and U5635 (N_5635,N_5285,N_5017);
xnor U5636 (N_5636,N_5367,N_5179);
xor U5637 (N_5637,N_5259,N_4838);
xnor U5638 (N_5638,N_4982,N_4989);
nor U5639 (N_5639,N_5380,N_4872);
nand U5640 (N_5640,N_5241,N_5502);
xor U5641 (N_5641,N_5047,N_5220);
nor U5642 (N_5642,N_5485,N_5117);
nor U5643 (N_5643,N_5041,N_5575);
xnor U5644 (N_5644,N_4993,N_5018);
nand U5645 (N_5645,N_5497,N_5211);
nand U5646 (N_5646,N_4938,N_5118);
xor U5647 (N_5647,N_5020,N_5157);
or U5648 (N_5648,N_5390,N_5084);
nand U5649 (N_5649,N_4941,N_4956);
nand U5650 (N_5650,N_5009,N_5477);
and U5651 (N_5651,N_5589,N_5405);
nand U5652 (N_5652,N_4943,N_5176);
or U5653 (N_5653,N_5230,N_5122);
nor U5654 (N_5654,N_5499,N_5262);
xnor U5655 (N_5655,N_5393,N_5430);
nand U5656 (N_5656,N_5310,N_5525);
and U5657 (N_5657,N_4879,N_5232);
and U5658 (N_5658,N_5030,N_5324);
or U5659 (N_5659,N_5286,N_5353);
nand U5660 (N_5660,N_5036,N_5214);
nand U5661 (N_5661,N_5153,N_5253);
and U5662 (N_5662,N_5170,N_5467);
or U5663 (N_5663,N_5108,N_5398);
xnor U5664 (N_5664,N_4845,N_4887);
and U5665 (N_5665,N_5119,N_4821);
or U5666 (N_5666,N_5599,N_5574);
nand U5667 (N_5667,N_5161,N_4814);
or U5668 (N_5668,N_4976,N_5093);
or U5669 (N_5669,N_5309,N_4991);
nand U5670 (N_5670,N_5003,N_5204);
xor U5671 (N_5671,N_4995,N_5592);
and U5672 (N_5672,N_5385,N_4891);
nor U5673 (N_5673,N_5587,N_5533);
nor U5674 (N_5674,N_5257,N_4965);
or U5675 (N_5675,N_4892,N_5560);
and U5676 (N_5676,N_4852,N_5540);
or U5677 (N_5677,N_5323,N_5154);
nand U5678 (N_5678,N_5284,N_5322);
xnor U5679 (N_5679,N_5454,N_5193);
and U5680 (N_5680,N_5466,N_4848);
xnor U5681 (N_5681,N_5597,N_5000);
and U5682 (N_5682,N_5583,N_5210);
nor U5683 (N_5683,N_5300,N_5191);
xor U5684 (N_5684,N_4819,N_4933);
xnor U5685 (N_5685,N_5014,N_5169);
and U5686 (N_5686,N_4909,N_4824);
and U5687 (N_5687,N_5565,N_5276);
xor U5688 (N_5688,N_5277,N_5422);
xnor U5689 (N_5689,N_5140,N_5125);
nand U5690 (N_5690,N_5054,N_4897);
or U5691 (N_5691,N_4979,N_4952);
nor U5692 (N_5692,N_5334,N_5251);
nor U5693 (N_5693,N_5032,N_5135);
and U5694 (N_5694,N_4810,N_5115);
and U5695 (N_5695,N_5357,N_5111);
nand U5696 (N_5696,N_4959,N_5229);
xnor U5697 (N_5697,N_5069,N_5530);
nand U5698 (N_5698,N_4910,N_5399);
xnor U5699 (N_5699,N_5168,N_4985);
nand U5700 (N_5700,N_5320,N_5358);
xor U5701 (N_5701,N_5532,N_4966);
xnor U5702 (N_5702,N_5281,N_4969);
and U5703 (N_5703,N_5109,N_5246);
or U5704 (N_5704,N_5266,N_5022);
nor U5705 (N_5705,N_5120,N_5151);
xnor U5706 (N_5706,N_4977,N_5013);
nor U5707 (N_5707,N_5335,N_5181);
or U5708 (N_5708,N_4916,N_5483);
nand U5709 (N_5709,N_5228,N_5059);
nor U5710 (N_5710,N_4884,N_5177);
or U5711 (N_5711,N_5458,N_5571);
or U5712 (N_5712,N_5581,N_5053);
and U5713 (N_5713,N_4847,N_5275);
nor U5714 (N_5714,N_4896,N_5234);
nand U5715 (N_5715,N_5171,N_4901);
xnor U5716 (N_5716,N_4981,N_4857);
nor U5717 (N_5717,N_4984,N_5016);
or U5718 (N_5718,N_5105,N_4948);
xnor U5719 (N_5719,N_5424,N_5001);
or U5720 (N_5720,N_5040,N_5416);
nand U5721 (N_5721,N_5212,N_5260);
nor U5722 (N_5722,N_5509,N_4898);
nor U5723 (N_5723,N_4867,N_4831);
and U5724 (N_5724,N_5376,N_5061);
or U5725 (N_5725,N_5538,N_5124);
xnor U5726 (N_5726,N_5543,N_5505);
nand U5727 (N_5727,N_5313,N_5127);
nand U5728 (N_5728,N_5306,N_4955);
or U5729 (N_5729,N_5134,N_5189);
or U5730 (N_5730,N_5489,N_5156);
or U5731 (N_5731,N_4890,N_5468);
xnor U5732 (N_5732,N_5245,N_4986);
xor U5733 (N_5733,N_4883,N_4914);
nor U5734 (N_5734,N_5374,N_5312);
nand U5735 (N_5735,N_5031,N_5307);
nor U5736 (N_5736,N_4968,N_4926);
xnor U5737 (N_5737,N_5553,N_5293);
nor U5738 (N_5738,N_5409,N_5303);
nand U5739 (N_5739,N_5396,N_5420);
xor U5740 (N_5740,N_5542,N_5508);
nor U5741 (N_5741,N_5584,N_5026);
xnor U5742 (N_5742,N_4928,N_5496);
xor U5743 (N_5743,N_5244,N_4851);
nand U5744 (N_5744,N_5185,N_5449);
and U5745 (N_5745,N_5280,N_4842);
or U5746 (N_5746,N_5527,N_5484);
or U5747 (N_5747,N_5438,N_4853);
and U5748 (N_5748,N_5373,N_5146);
and U5749 (N_5749,N_5439,N_5102);
and U5750 (N_5750,N_4812,N_5055);
nand U5751 (N_5751,N_5344,N_5523);
nor U5752 (N_5752,N_4971,N_5141);
nor U5753 (N_5753,N_4809,N_5475);
nand U5754 (N_5754,N_5550,N_5272);
nor U5755 (N_5755,N_5264,N_5142);
and U5756 (N_5756,N_4828,N_5073);
nor U5757 (N_5757,N_5081,N_5225);
nand U5758 (N_5758,N_5183,N_5348);
or U5759 (N_5759,N_5488,N_5425);
nor U5760 (N_5760,N_4807,N_5343);
or U5761 (N_5761,N_5369,N_4876);
xnor U5762 (N_5762,N_5173,N_5213);
and U5763 (N_5763,N_4836,N_5063);
and U5764 (N_5764,N_5598,N_5456);
nor U5765 (N_5765,N_4905,N_5295);
nor U5766 (N_5766,N_5577,N_5524);
nor U5767 (N_5767,N_5150,N_5147);
nor U5768 (N_5768,N_5327,N_5371);
nor U5769 (N_5769,N_5062,N_5227);
nand U5770 (N_5770,N_5242,N_5331);
and U5771 (N_5771,N_5338,N_5351);
nand U5772 (N_5772,N_4974,N_4931);
or U5773 (N_5773,N_4920,N_5573);
nor U5774 (N_5774,N_5355,N_5455);
xnor U5775 (N_5775,N_4844,N_5218);
nor U5776 (N_5776,N_5594,N_5039);
nor U5777 (N_5777,N_5103,N_4833);
nand U5778 (N_5778,N_4825,N_5408);
xnor U5779 (N_5779,N_5379,N_5356);
xnor U5780 (N_5780,N_5566,N_5362);
nand U5781 (N_5781,N_5186,N_5006);
or U5782 (N_5782,N_4816,N_5474);
xnor U5783 (N_5783,N_4999,N_5507);
nand U5784 (N_5784,N_5473,N_5319);
and U5785 (N_5785,N_5591,N_5545);
and U5786 (N_5786,N_5506,N_4804);
nor U5787 (N_5787,N_5012,N_5051);
and U5788 (N_5788,N_4805,N_5070);
nand U5789 (N_5789,N_5100,N_5547);
nand U5790 (N_5790,N_5302,N_5128);
nand U5791 (N_5791,N_5282,N_5435);
nand U5792 (N_5792,N_5129,N_5513);
nand U5793 (N_5793,N_5315,N_5187);
or U5794 (N_5794,N_5023,N_5578);
nor U5795 (N_5795,N_5196,N_5098);
nor U5796 (N_5796,N_5383,N_5465);
nor U5797 (N_5797,N_5126,N_4934);
or U5798 (N_5798,N_5480,N_5349);
and U5799 (N_5799,N_5269,N_5340);
nand U5800 (N_5800,N_5562,N_4866);
nor U5801 (N_5801,N_4915,N_5490);
nor U5802 (N_5802,N_5572,N_4865);
and U5803 (N_5803,N_4947,N_5209);
and U5804 (N_5804,N_5460,N_5576);
and U5805 (N_5805,N_5028,N_5247);
nand U5806 (N_5806,N_5060,N_5043);
or U5807 (N_5807,N_5048,N_5148);
and U5808 (N_5808,N_5586,N_5278);
or U5809 (N_5809,N_5164,N_5094);
nand U5810 (N_5810,N_5316,N_5206);
or U5811 (N_5811,N_5450,N_5461);
or U5812 (N_5812,N_5101,N_5593);
nand U5813 (N_5813,N_4975,N_5263);
or U5814 (N_5814,N_4861,N_4860);
nor U5815 (N_5815,N_4954,N_5426);
or U5816 (N_5816,N_4996,N_5294);
xnor U5817 (N_5817,N_5044,N_5500);
or U5818 (N_5818,N_5341,N_4895);
and U5819 (N_5819,N_5388,N_5195);
xnor U5820 (N_5820,N_5471,N_5437);
and U5821 (N_5821,N_5075,N_5130);
and U5822 (N_5822,N_4907,N_5436);
nor U5823 (N_5823,N_5208,N_4962);
nor U5824 (N_5824,N_5010,N_5579);
or U5825 (N_5825,N_5052,N_5321);
nor U5826 (N_5826,N_4945,N_5417);
nor U5827 (N_5827,N_5021,N_5325);
nand U5828 (N_5828,N_4811,N_5386);
and U5829 (N_5829,N_5288,N_5296);
and U5830 (N_5830,N_5292,N_5166);
xor U5831 (N_5831,N_4998,N_5363);
and U5832 (N_5832,N_5382,N_5482);
and U5833 (N_5833,N_5235,N_5231);
or U5834 (N_5834,N_5451,N_5056);
and U5835 (N_5835,N_5537,N_5114);
xnor U5836 (N_5836,N_5015,N_5290);
nor U5837 (N_5837,N_5470,N_5248);
nor U5838 (N_5838,N_4939,N_5074);
or U5839 (N_5839,N_4837,N_4840);
and U5840 (N_5840,N_5182,N_5498);
nor U5841 (N_5841,N_4921,N_5567);
nor U5842 (N_5842,N_5364,N_5517);
nor U5843 (N_5843,N_5541,N_4960);
xor U5844 (N_5844,N_5078,N_4859);
nand U5845 (N_5845,N_5370,N_5123);
nand U5846 (N_5846,N_5145,N_5520);
or U5847 (N_5847,N_4899,N_5267);
and U5848 (N_5848,N_5345,N_4886);
xor U5849 (N_5849,N_5413,N_5184);
or U5850 (N_5850,N_5429,N_5360);
or U5851 (N_5851,N_4873,N_4802);
or U5852 (N_5852,N_4922,N_5561);
xor U5853 (N_5853,N_5493,N_5478);
nor U5854 (N_5854,N_5539,N_5427);
nor U5855 (N_5855,N_5463,N_5237);
nor U5856 (N_5856,N_5308,N_4829);
nand U5857 (N_5857,N_5432,N_5240);
nand U5858 (N_5858,N_4850,N_5549);
nand U5859 (N_5859,N_5559,N_5019);
nor U5860 (N_5860,N_4846,N_5428);
xor U5861 (N_5861,N_5215,N_4911);
xor U5862 (N_5862,N_5568,N_5453);
and U5863 (N_5863,N_4925,N_5112);
nand U5864 (N_5864,N_5329,N_5372);
nand U5865 (N_5865,N_5529,N_5283);
nor U5866 (N_5866,N_5445,N_5050);
nor U5867 (N_5867,N_5097,N_5298);
and U5868 (N_5868,N_5143,N_5200);
nand U5869 (N_5869,N_5419,N_5423);
or U5870 (N_5870,N_5113,N_5531);
nand U5871 (N_5871,N_5558,N_5387);
xnor U5872 (N_5872,N_5131,N_5384);
or U5873 (N_5873,N_4919,N_5442);
nand U5874 (N_5874,N_4863,N_4900);
or U5875 (N_5875,N_5236,N_5459);
nand U5876 (N_5876,N_5107,N_5160);
or U5877 (N_5877,N_4904,N_4942);
nor U5878 (N_5878,N_4830,N_5033);
and U5879 (N_5879,N_4877,N_5086);
xor U5880 (N_5880,N_5090,N_5149);
xnor U5881 (N_5881,N_5421,N_5091);
nand U5882 (N_5882,N_5065,N_5318);
and U5883 (N_5883,N_5389,N_4963);
nor U5884 (N_5884,N_5494,N_5504);
or U5885 (N_5885,N_5175,N_5027);
and U5886 (N_5886,N_4874,N_5034);
xnor U5887 (N_5887,N_5121,N_4918);
nand U5888 (N_5888,N_5431,N_4935);
and U5889 (N_5889,N_5239,N_5008);
or U5890 (N_5890,N_4880,N_5440);
and U5891 (N_5891,N_5452,N_5301);
nand U5892 (N_5892,N_5418,N_4889);
nor U5893 (N_5893,N_5446,N_5580);
nand U5894 (N_5894,N_5273,N_5274);
nand U5895 (N_5895,N_5546,N_5238);
nor U5896 (N_5896,N_5414,N_4841);
nand U5897 (N_5897,N_5378,N_4875);
or U5898 (N_5898,N_4881,N_5192);
xnor U5899 (N_5899,N_5079,N_4858);
xnor U5900 (N_5900,N_5133,N_5518);
or U5901 (N_5901,N_5443,N_5217);
nor U5902 (N_5902,N_4906,N_4815);
or U5903 (N_5903,N_5046,N_5392);
or U5904 (N_5904,N_5025,N_5085);
xor U5905 (N_5905,N_5066,N_5254);
and U5906 (N_5906,N_5342,N_5072);
nor U5907 (N_5907,N_5190,N_5472);
xnor U5908 (N_5908,N_5029,N_5110);
nand U5909 (N_5909,N_5291,N_5139);
nor U5910 (N_5910,N_5336,N_5188);
and U5911 (N_5911,N_5132,N_5333);
or U5912 (N_5912,N_5035,N_5406);
nor U5913 (N_5913,N_5083,N_5299);
nor U5914 (N_5914,N_5410,N_5194);
xor U5915 (N_5915,N_4927,N_5162);
nand U5916 (N_5916,N_5045,N_5375);
nand U5917 (N_5917,N_4854,N_5116);
nand U5918 (N_5918,N_5155,N_4871);
or U5919 (N_5919,N_5163,N_5462);
or U5920 (N_5920,N_5457,N_5481);
nor U5921 (N_5921,N_5095,N_5407);
nand U5922 (N_5922,N_5536,N_4937);
xor U5923 (N_5923,N_5180,N_5514);
nand U5924 (N_5924,N_5521,N_5570);
nand U5925 (N_5925,N_5519,N_5347);
nand U5926 (N_5926,N_5486,N_5403);
nand U5927 (N_5927,N_4869,N_5402);
xnor U5928 (N_5928,N_5252,N_4951);
nand U5929 (N_5929,N_5165,N_4888);
xnor U5930 (N_5930,N_5441,N_5339);
or U5931 (N_5931,N_5395,N_5564);
nand U5932 (N_5932,N_4970,N_5554);
xnor U5933 (N_5933,N_5287,N_5250);
nor U5934 (N_5934,N_4953,N_5555);
or U5935 (N_5935,N_4893,N_5004);
xnor U5936 (N_5936,N_5346,N_5464);
or U5937 (N_5937,N_5082,N_5219);
nand U5938 (N_5938,N_5289,N_5099);
or U5939 (N_5939,N_5201,N_4834);
and U5940 (N_5940,N_5447,N_4987);
nor U5941 (N_5941,N_5551,N_5330);
or U5942 (N_5942,N_4950,N_4957);
nor U5943 (N_5943,N_5137,N_4992);
xnor U5944 (N_5944,N_5377,N_4923);
or U5945 (N_5945,N_4944,N_5487);
nand U5946 (N_5946,N_5089,N_5544);
or U5947 (N_5947,N_4839,N_5381);
xnor U5948 (N_5948,N_5268,N_5411);
and U5949 (N_5949,N_5205,N_5510);
and U5950 (N_5950,N_4864,N_4855);
nand U5951 (N_5951,N_5076,N_5092);
or U5952 (N_5952,N_4806,N_5522);
or U5953 (N_5953,N_5255,N_5596);
or U5954 (N_5954,N_5512,N_5503);
nor U5955 (N_5955,N_5080,N_5068);
and U5956 (N_5956,N_5007,N_4862);
or U5957 (N_5957,N_5198,N_4801);
and U5958 (N_5958,N_4856,N_5590);
xor U5959 (N_5959,N_5585,N_5064);
xor U5960 (N_5960,N_5479,N_5359);
nor U5961 (N_5961,N_5271,N_5548);
or U5962 (N_5962,N_4936,N_4946);
and U5963 (N_5963,N_5448,N_4997);
and U5964 (N_5964,N_5279,N_5412);
nand U5965 (N_5965,N_5326,N_4924);
xnor U5966 (N_5966,N_5552,N_5071);
or U5967 (N_5967,N_5167,N_4917);
xnor U5968 (N_5968,N_5317,N_5249);
or U5969 (N_5969,N_5256,N_4820);
nor U5970 (N_5970,N_4835,N_5515);
xor U5971 (N_5971,N_4826,N_5516);
and U5972 (N_5972,N_5144,N_5223);
and U5973 (N_5973,N_4849,N_5588);
nand U5974 (N_5974,N_4903,N_5366);
nand U5975 (N_5975,N_4800,N_5138);
and U5976 (N_5976,N_5444,N_5024);
nor U5977 (N_5977,N_5243,N_5222);
nand U5978 (N_5978,N_5569,N_5005);
and U5979 (N_5979,N_5469,N_5491);
xor U5980 (N_5980,N_5332,N_5265);
xor U5981 (N_5981,N_5304,N_4940);
xnor U5982 (N_5982,N_4870,N_5221);
or U5983 (N_5983,N_4878,N_5077);
nor U5984 (N_5984,N_4980,N_5476);
xnor U5985 (N_5985,N_5557,N_4817);
nand U5986 (N_5986,N_5258,N_5002);
nand U5987 (N_5987,N_5011,N_5501);
xor U5988 (N_5988,N_5534,N_4967);
and U5989 (N_5989,N_4894,N_4990);
nand U5990 (N_5990,N_5207,N_5226);
xor U5991 (N_5991,N_5401,N_4813);
and U5992 (N_5992,N_4808,N_5492);
or U5993 (N_5993,N_4832,N_4823);
and U5994 (N_5994,N_4929,N_5202);
xnor U5995 (N_5995,N_5087,N_4822);
or U5996 (N_5996,N_5328,N_5067);
or U5997 (N_5997,N_4994,N_5197);
xnor U5998 (N_5998,N_5042,N_5394);
nor U5999 (N_5999,N_4912,N_4972);
or U6000 (N_6000,N_5037,N_5510);
nand U6001 (N_6001,N_5048,N_5008);
or U6002 (N_6002,N_5274,N_5126);
and U6003 (N_6003,N_4943,N_5065);
xnor U6004 (N_6004,N_5527,N_4939);
or U6005 (N_6005,N_5469,N_5479);
xor U6006 (N_6006,N_4986,N_5087);
xnor U6007 (N_6007,N_5342,N_5101);
nand U6008 (N_6008,N_5319,N_4983);
nand U6009 (N_6009,N_5532,N_5045);
nand U6010 (N_6010,N_5081,N_5593);
xnor U6011 (N_6011,N_5335,N_5154);
or U6012 (N_6012,N_5490,N_5594);
nor U6013 (N_6013,N_5356,N_4988);
nand U6014 (N_6014,N_4835,N_5215);
nor U6015 (N_6015,N_4941,N_5451);
or U6016 (N_6016,N_5262,N_5584);
xnor U6017 (N_6017,N_5377,N_5170);
and U6018 (N_6018,N_5566,N_5461);
nand U6019 (N_6019,N_5111,N_5038);
xnor U6020 (N_6020,N_5396,N_5315);
xnor U6021 (N_6021,N_4865,N_4845);
nand U6022 (N_6022,N_5317,N_5246);
nand U6023 (N_6023,N_5146,N_4964);
or U6024 (N_6024,N_4968,N_5415);
and U6025 (N_6025,N_5089,N_4957);
and U6026 (N_6026,N_5456,N_5133);
nor U6027 (N_6027,N_4944,N_5025);
xor U6028 (N_6028,N_4843,N_4840);
and U6029 (N_6029,N_4991,N_5133);
xor U6030 (N_6030,N_4842,N_5246);
nor U6031 (N_6031,N_5536,N_5301);
nor U6032 (N_6032,N_5326,N_5561);
nor U6033 (N_6033,N_5024,N_5279);
xnor U6034 (N_6034,N_5142,N_4962);
xor U6035 (N_6035,N_5599,N_4997);
and U6036 (N_6036,N_5542,N_5215);
and U6037 (N_6037,N_4888,N_5297);
or U6038 (N_6038,N_5445,N_5589);
and U6039 (N_6039,N_5494,N_5321);
nand U6040 (N_6040,N_4961,N_4876);
or U6041 (N_6041,N_5473,N_5277);
and U6042 (N_6042,N_5331,N_5050);
nand U6043 (N_6043,N_5213,N_4943);
nor U6044 (N_6044,N_4903,N_4890);
or U6045 (N_6045,N_5440,N_5572);
nand U6046 (N_6046,N_5187,N_4941);
or U6047 (N_6047,N_5086,N_5326);
nand U6048 (N_6048,N_4923,N_5380);
or U6049 (N_6049,N_4926,N_5022);
nor U6050 (N_6050,N_5286,N_5179);
and U6051 (N_6051,N_5307,N_5064);
nand U6052 (N_6052,N_5288,N_5554);
nor U6053 (N_6053,N_4901,N_5366);
nor U6054 (N_6054,N_4842,N_5175);
and U6055 (N_6055,N_5290,N_5147);
nand U6056 (N_6056,N_5470,N_5372);
and U6057 (N_6057,N_5156,N_5236);
nor U6058 (N_6058,N_5414,N_4864);
nand U6059 (N_6059,N_5401,N_4972);
xnor U6060 (N_6060,N_5228,N_4807);
nand U6061 (N_6061,N_5481,N_5149);
or U6062 (N_6062,N_5572,N_4950);
xor U6063 (N_6063,N_5118,N_5222);
nor U6064 (N_6064,N_4841,N_4969);
nor U6065 (N_6065,N_4927,N_5556);
and U6066 (N_6066,N_5513,N_5230);
nand U6067 (N_6067,N_4835,N_5597);
xnor U6068 (N_6068,N_4952,N_5226);
xor U6069 (N_6069,N_5213,N_5315);
nand U6070 (N_6070,N_5212,N_5159);
nand U6071 (N_6071,N_5123,N_4990);
or U6072 (N_6072,N_5544,N_4952);
nand U6073 (N_6073,N_4966,N_4969);
nor U6074 (N_6074,N_5555,N_5240);
xor U6075 (N_6075,N_5201,N_4874);
nand U6076 (N_6076,N_5097,N_5423);
and U6077 (N_6077,N_5033,N_5449);
nand U6078 (N_6078,N_5353,N_5381);
or U6079 (N_6079,N_5071,N_5055);
xor U6080 (N_6080,N_5429,N_4925);
nor U6081 (N_6081,N_5358,N_5325);
and U6082 (N_6082,N_5127,N_5408);
nand U6083 (N_6083,N_5422,N_4889);
and U6084 (N_6084,N_4967,N_5505);
nand U6085 (N_6085,N_5324,N_5413);
nor U6086 (N_6086,N_5568,N_5488);
nand U6087 (N_6087,N_5312,N_4838);
nand U6088 (N_6088,N_4847,N_5562);
or U6089 (N_6089,N_5492,N_5502);
xnor U6090 (N_6090,N_5382,N_5280);
nand U6091 (N_6091,N_5138,N_5032);
nand U6092 (N_6092,N_5552,N_5551);
xnor U6093 (N_6093,N_5445,N_4834);
and U6094 (N_6094,N_5459,N_5359);
xnor U6095 (N_6095,N_5144,N_5507);
nor U6096 (N_6096,N_5507,N_5352);
xnor U6097 (N_6097,N_4933,N_5593);
xor U6098 (N_6098,N_5470,N_5419);
nand U6099 (N_6099,N_5534,N_5272);
nand U6100 (N_6100,N_5404,N_5541);
nand U6101 (N_6101,N_5022,N_5301);
nor U6102 (N_6102,N_5095,N_4849);
or U6103 (N_6103,N_4896,N_5109);
xor U6104 (N_6104,N_5180,N_5150);
nor U6105 (N_6105,N_5470,N_5013);
xor U6106 (N_6106,N_5266,N_5560);
nor U6107 (N_6107,N_5121,N_4999);
and U6108 (N_6108,N_4916,N_4990);
xor U6109 (N_6109,N_4824,N_5194);
xor U6110 (N_6110,N_5406,N_5065);
nor U6111 (N_6111,N_5362,N_4806);
nand U6112 (N_6112,N_5522,N_4931);
nor U6113 (N_6113,N_5304,N_5331);
and U6114 (N_6114,N_5321,N_5366);
and U6115 (N_6115,N_4943,N_5350);
nor U6116 (N_6116,N_4854,N_5268);
nor U6117 (N_6117,N_4821,N_4890);
and U6118 (N_6118,N_4925,N_4825);
nand U6119 (N_6119,N_4883,N_5296);
xnor U6120 (N_6120,N_5356,N_5005);
nor U6121 (N_6121,N_5436,N_5279);
nand U6122 (N_6122,N_5468,N_4965);
or U6123 (N_6123,N_4851,N_5230);
or U6124 (N_6124,N_4994,N_5151);
xnor U6125 (N_6125,N_5435,N_4961);
xor U6126 (N_6126,N_4868,N_5208);
xnor U6127 (N_6127,N_5489,N_5318);
or U6128 (N_6128,N_5183,N_4879);
xnor U6129 (N_6129,N_4903,N_5086);
or U6130 (N_6130,N_5412,N_5106);
nand U6131 (N_6131,N_5460,N_5093);
and U6132 (N_6132,N_5106,N_5517);
nor U6133 (N_6133,N_5284,N_5544);
and U6134 (N_6134,N_5262,N_5009);
nand U6135 (N_6135,N_5584,N_5025);
nor U6136 (N_6136,N_5381,N_5060);
nor U6137 (N_6137,N_5520,N_5519);
nand U6138 (N_6138,N_5006,N_4917);
or U6139 (N_6139,N_5217,N_5197);
and U6140 (N_6140,N_4830,N_5401);
or U6141 (N_6141,N_5033,N_5520);
xor U6142 (N_6142,N_5597,N_5354);
and U6143 (N_6143,N_5547,N_5173);
nand U6144 (N_6144,N_4853,N_5218);
nor U6145 (N_6145,N_5074,N_5389);
xor U6146 (N_6146,N_5368,N_4901);
nand U6147 (N_6147,N_5543,N_5028);
or U6148 (N_6148,N_5277,N_5101);
and U6149 (N_6149,N_5405,N_5175);
or U6150 (N_6150,N_5088,N_5120);
and U6151 (N_6151,N_5349,N_5511);
xor U6152 (N_6152,N_5140,N_4900);
or U6153 (N_6153,N_5156,N_4966);
or U6154 (N_6154,N_5011,N_5573);
nor U6155 (N_6155,N_4969,N_5322);
or U6156 (N_6156,N_5157,N_4806);
nand U6157 (N_6157,N_4944,N_5163);
and U6158 (N_6158,N_4864,N_5058);
nor U6159 (N_6159,N_4832,N_5294);
nor U6160 (N_6160,N_5034,N_5475);
and U6161 (N_6161,N_5213,N_4906);
and U6162 (N_6162,N_4844,N_5334);
nand U6163 (N_6163,N_5526,N_5067);
and U6164 (N_6164,N_5351,N_5067);
nor U6165 (N_6165,N_4947,N_5410);
nor U6166 (N_6166,N_5542,N_5218);
xnor U6167 (N_6167,N_4823,N_5038);
nand U6168 (N_6168,N_5174,N_5302);
or U6169 (N_6169,N_5285,N_5528);
nand U6170 (N_6170,N_4929,N_4823);
nand U6171 (N_6171,N_5285,N_4872);
nor U6172 (N_6172,N_5525,N_4998);
and U6173 (N_6173,N_5422,N_4971);
nand U6174 (N_6174,N_5418,N_4979);
nor U6175 (N_6175,N_4925,N_5248);
xnor U6176 (N_6176,N_5368,N_5440);
nand U6177 (N_6177,N_4938,N_5544);
and U6178 (N_6178,N_5577,N_5299);
and U6179 (N_6179,N_5141,N_5354);
nor U6180 (N_6180,N_5567,N_5249);
nor U6181 (N_6181,N_4995,N_5353);
or U6182 (N_6182,N_5563,N_5252);
nand U6183 (N_6183,N_4830,N_5334);
nor U6184 (N_6184,N_5350,N_4817);
xnor U6185 (N_6185,N_5448,N_5567);
nand U6186 (N_6186,N_4803,N_5062);
and U6187 (N_6187,N_5096,N_5089);
nor U6188 (N_6188,N_4847,N_4886);
or U6189 (N_6189,N_5358,N_5548);
or U6190 (N_6190,N_5444,N_5088);
nand U6191 (N_6191,N_5507,N_5410);
or U6192 (N_6192,N_4940,N_4978);
xnor U6193 (N_6193,N_5599,N_5434);
nor U6194 (N_6194,N_5094,N_4897);
nor U6195 (N_6195,N_4965,N_4943);
nor U6196 (N_6196,N_5286,N_5000);
nor U6197 (N_6197,N_5450,N_4954);
and U6198 (N_6198,N_5022,N_5173);
or U6199 (N_6199,N_4904,N_5207);
nor U6200 (N_6200,N_4811,N_5474);
nor U6201 (N_6201,N_4906,N_5572);
and U6202 (N_6202,N_4904,N_4929);
and U6203 (N_6203,N_4825,N_5597);
xnor U6204 (N_6204,N_4839,N_5401);
or U6205 (N_6205,N_5498,N_5191);
and U6206 (N_6206,N_5336,N_5357);
nor U6207 (N_6207,N_5346,N_5445);
or U6208 (N_6208,N_4839,N_5226);
nand U6209 (N_6209,N_4917,N_5187);
or U6210 (N_6210,N_5502,N_5541);
and U6211 (N_6211,N_4894,N_4860);
nor U6212 (N_6212,N_5238,N_5135);
or U6213 (N_6213,N_4804,N_5144);
nor U6214 (N_6214,N_5203,N_5559);
and U6215 (N_6215,N_5427,N_5136);
xor U6216 (N_6216,N_5312,N_5492);
nor U6217 (N_6217,N_5009,N_5482);
or U6218 (N_6218,N_4930,N_5067);
and U6219 (N_6219,N_4828,N_5507);
and U6220 (N_6220,N_5211,N_4805);
xor U6221 (N_6221,N_5594,N_5353);
and U6222 (N_6222,N_5208,N_4879);
and U6223 (N_6223,N_4837,N_5114);
and U6224 (N_6224,N_5458,N_5104);
nor U6225 (N_6225,N_5376,N_4979);
nor U6226 (N_6226,N_5440,N_5151);
and U6227 (N_6227,N_4985,N_4842);
or U6228 (N_6228,N_5467,N_5405);
nand U6229 (N_6229,N_5346,N_5064);
nand U6230 (N_6230,N_5010,N_5276);
nand U6231 (N_6231,N_5502,N_5263);
and U6232 (N_6232,N_5147,N_4925);
xnor U6233 (N_6233,N_5375,N_5330);
or U6234 (N_6234,N_5484,N_5496);
and U6235 (N_6235,N_5494,N_5376);
or U6236 (N_6236,N_4818,N_5515);
nor U6237 (N_6237,N_4897,N_5164);
or U6238 (N_6238,N_5577,N_5048);
and U6239 (N_6239,N_4983,N_5502);
xor U6240 (N_6240,N_5188,N_5037);
xnor U6241 (N_6241,N_5560,N_5357);
and U6242 (N_6242,N_4861,N_5555);
and U6243 (N_6243,N_5494,N_5517);
nand U6244 (N_6244,N_5101,N_4964);
nand U6245 (N_6245,N_5389,N_5084);
nor U6246 (N_6246,N_4803,N_5385);
nand U6247 (N_6247,N_5501,N_5484);
and U6248 (N_6248,N_5297,N_5562);
nor U6249 (N_6249,N_4864,N_4898);
and U6250 (N_6250,N_5255,N_5097);
or U6251 (N_6251,N_4917,N_4844);
and U6252 (N_6252,N_5417,N_5426);
and U6253 (N_6253,N_5256,N_5003);
or U6254 (N_6254,N_4933,N_5216);
nand U6255 (N_6255,N_5012,N_5502);
nand U6256 (N_6256,N_5403,N_5374);
nand U6257 (N_6257,N_4856,N_5182);
or U6258 (N_6258,N_5594,N_4931);
nor U6259 (N_6259,N_5400,N_5196);
xnor U6260 (N_6260,N_5201,N_5133);
or U6261 (N_6261,N_5151,N_5221);
and U6262 (N_6262,N_5421,N_5088);
or U6263 (N_6263,N_5456,N_5580);
nor U6264 (N_6264,N_5183,N_4911);
or U6265 (N_6265,N_4857,N_5149);
and U6266 (N_6266,N_4804,N_4888);
or U6267 (N_6267,N_5565,N_4969);
nor U6268 (N_6268,N_5059,N_4986);
or U6269 (N_6269,N_5548,N_4816);
nand U6270 (N_6270,N_5473,N_4850);
nand U6271 (N_6271,N_5026,N_5242);
nand U6272 (N_6272,N_4919,N_4971);
nand U6273 (N_6273,N_5116,N_5519);
nand U6274 (N_6274,N_4822,N_4874);
nor U6275 (N_6275,N_5479,N_4882);
or U6276 (N_6276,N_5104,N_5079);
xor U6277 (N_6277,N_5505,N_5399);
and U6278 (N_6278,N_5006,N_5332);
or U6279 (N_6279,N_5259,N_4960);
or U6280 (N_6280,N_4834,N_5456);
nand U6281 (N_6281,N_5055,N_5264);
or U6282 (N_6282,N_5077,N_5555);
xor U6283 (N_6283,N_4918,N_5491);
and U6284 (N_6284,N_5559,N_5265);
or U6285 (N_6285,N_5004,N_5512);
and U6286 (N_6286,N_5151,N_5412);
or U6287 (N_6287,N_5398,N_5000);
nand U6288 (N_6288,N_5386,N_4995);
and U6289 (N_6289,N_5443,N_5498);
nor U6290 (N_6290,N_4801,N_5516);
nor U6291 (N_6291,N_5541,N_5456);
nor U6292 (N_6292,N_5055,N_4913);
xnor U6293 (N_6293,N_4907,N_5504);
nor U6294 (N_6294,N_4803,N_5175);
nor U6295 (N_6295,N_4989,N_5556);
nand U6296 (N_6296,N_4899,N_4804);
and U6297 (N_6297,N_5491,N_5241);
and U6298 (N_6298,N_4876,N_5518);
and U6299 (N_6299,N_5133,N_4824);
or U6300 (N_6300,N_5320,N_4907);
nor U6301 (N_6301,N_5595,N_5598);
and U6302 (N_6302,N_5121,N_5381);
nor U6303 (N_6303,N_5104,N_5001);
nand U6304 (N_6304,N_4970,N_5332);
nor U6305 (N_6305,N_5561,N_5447);
nand U6306 (N_6306,N_5434,N_5508);
or U6307 (N_6307,N_5152,N_4826);
xnor U6308 (N_6308,N_5590,N_5018);
xnor U6309 (N_6309,N_4853,N_5004);
nor U6310 (N_6310,N_5477,N_4815);
nor U6311 (N_6311,N_4806,N_5466);
and U6312 (N_6312,N_5558,N_5358);
nand U6313 (N_6313,N_5281,N_5129);
xnor U6314 (N_6314,N_5098,N_4859);
or U6315 (N_6315,N_5330,N_5246);
nor U6316 (N_6316,N_4844,N_5074);
xor U6317 (N_6317,N_5025,N_5183);
and U6318 (N_6318,N_4937,N_5019);
nand U6319 (N_6319,N_5585,N_5499);
or U6320 (N_6320,N_4837,N_5465);
and U6321 (N_6321,N_4976,N_5227);
or U6322 (N_6322,N_5217,N_5072);
nor U6323 (N_6323,N_5383,N_5371);
xnor U6324 (N_6324,N_4835,N_5194);
and U6325 (N_6325,N_5455,N_5564);
xnor U6326 (N_6326,N_5108,N_5513);
nor U6327 (N_6327,N_5035,N_5363);
nor U6328 (N_6328,N_5199,N_5153);
nor U6329 (N_6329,N_5281,N_5527);
and U6330 (N_6330,N_5583,N_5341);
nand U6331 (N_6331,N_4816,N_5398);
nand U6332 (N_6332,N_5117,N_5016);
and U6333 (N_6333,N_4902,N_5076);
nor U6334 (N_6334,N_4959,N_5014);
nand U6335 (N_6335,N_4889,N_5307);
nor U6336 (N_6336,N_5034,N_5156);
and U6337 (N_6337,N_5180,N_5434);
nor U6338 (N_6338,N_5208,N_5316);
nand U6339 (N_6339,N_5029,N_5453);
and U6340 (N_6340,N_5537,N_4808);
nor U6341 (N_6341,N_5209,N_4948);
xor U6342 (N_6342,N_5436,N_5044);
nand U6343 (N_6343,N_5110,N_4872);
nor U6344 (N_6344,N_4908,N_5363);
or U6345 (N_6345,N_5599,N_5413);
and U6346 (N_6346,N_4817,N_5429);
nor U6347 (N_6347,N_4900,N_5259);
or U6348 (N_6348,N_5017,N_5473);
nor U6349 (N_6349,N_4991,N_5111);
nand U6350 (N_6350,N_5233,N_4804);
nand U6351 (N_6351,N_5213,N_4986);
xor U6352 (N_6352,N_4955,N_5084);
nor U6353 (N_6353,N_5068,N_5016);
and U6354 (N_6354,N_5471,N_4945);
nor U6355 (N_6355,N_5099,N_5225);
nand U6356 (N_6356,N_5591,N_4893);
and U6357 (N_6357,N_5520,N_5019);
xor U6358 (N_6358,N_4966,N_4873);
or U6359 (N_6359,N_5183,N_5540);
or U6360 (N_6360,N_4902,N_4960);
nor U6361 (N_6361,N_4953,N_5503);
and U6362 (N_6362,N_4816,N_5142);
nand U6363 (N_6363,N_5355,N_4820);
xnor U6364 (N_6364,N_5377,N_5262);
nand U6365 (N_6365,N_5254,N_5063);
nand U6366 (N_6366,N_5281,N_5507);
and U6367 (N_6367,N_5109,N_4980);
and U6368 (N_6368,N_5168,N_5044);
nor U6369 (N_6369,N_5122,N_5021);
xor U6370 (N_6370,N_5252,N_5489);
xnor U6371 (N_6371,N_4895,N_5041);
or U6372 (N_6372,N_5034,N_5597);
or U6373 (N_6373,N_5045,N_5196);
xnor U6374 (N_6374,N_5437,N_5564);
nand U6375 (N_6375,N_5418,N_5300);
nor U6376 (N_6376,N_5487,N_5411);
nor U6377 (N_6377,N_5300,N_5121);
nor U6378 (N_6378,N_5317,N_4826);
xnor U6379 (N_6379,N_5310,N_5290);
nand U6380 (N_6380,N_5499,N_5107);
xnor U6381 (N_6381,N_4961,N_5398);
nor U6382 (N_6382,N_4937,N_4910);
nand U6383 (N_6383,N_5448,N_4982);
nor U6384 (N_6384,N_5587,N_5365);
nor U6385 (N_6385,N_5123,N_4872);
and U6386 (N_6386,N_5546,N_5051);
and U6387 (N_6387,N_5082,N_5387);
and U6388 (N_6388,N_4987,N_5453);
nand U6389 (N_6389,N_5255,N_5156);
nand U6390 (N_6390,N_5043,N_4815);
nand U6391 (N_6391,N_5441,N_5396);
and U6392 (N_6392,N_5436,N_5130);
nand U6393 (N_6393,N_4953,N_5268);
xnor U6394 (N_6394,N_5147,N_5423);
nor U6395 (N_6395,N_5092,N_5161);
nor U6396 (N_6396,N_5251,N_4975);
nor U6397 (N_6397,N_4866,N_5127);
xnor U6398 (N_6398,N_5343,N_5502);
or U6399 (N_6399,N_5580,N_4958);
xnor U6400 (N_6400,N_5908,N_6162);
or U6401 (N_6401,N_5726,N_6313);
xnor U6402 (N_6402,N_5684,N_6121);
or U6403 (N_6403,N_6029,N_5606);
nor U6404 (N_6404,N_6211,N_5840);
and U6405 (N_6405,N_6181,N_5627);
xor U6406 (N_6406,N_6221,N_6288);
xor U6407 (N_6407,N_6198,N_6017);
or U6408 (N_6408,N_6069,N_6280);
or U6409 (N_6409,N_6254,N_5871);
xnor U6410 (N_6410,N_5624,N_5854);
or U6411 (N_6411,N_5894,N_5966);
xor U6412 (N_6412,N_5905,N_5963);
nand U6413 (N_6413,N_6078,N_5738);
or U6414 (N_6414,N_5896,N_5798);
or U6415 (N_6415,N_6052,N_5917);
or U6416 (N_6416,N_5919,N_5828);
nor U6417 (N_6417,N_5823,N_6383);
and U6418 (N_6418,N_6243,N_5884);
or U6419 (N_6419,N_6101,N_6238);
nor U6420 (N_6420,N_5793,N_6328);
nand U6421 (N_6421,N_5682,N_5859);
nand U6422 (N_6422,N_5926,N_5845);
nand U6423 (N_6423,N_5995,N_6189);
and U6424 (N_6424,N_5763,N_5623);
xnor U6425 (N_6425,N_5640,N_6341);
or U6426 (N_6426,N_5681,N_5839);
nor U6427 (N_6427,N_6285,N_6076);
nor U6428 (N_6428,N_5625,N_6367);
or U6429 (N_6429,N_5992,N_5915);
and U6430 (N_6430,N_5900,N_6169);
nor U6431 (N_6431,N_6318,N_6389);
and U6432 (N_6432,N_5603,N_6088);
or U6433 (N_6433,N_5647,N_6342);
and U6434 (N_6434,N_6200,N_6099);
and U6435 (N_6435,N_6265,N_5614);
nand U6436 (N_6436,N_6337,N_5948);
or U6437 (N_6437,N_6115,N_6301);
nor U6438 (N_6438,N_6156,N_6290);
or U6439 (N_6439,N_6253,N_5803);
xnor U6440 (N_6440,N_5759,N_5902);
nor U6441 (N_6441,N_6353,N_5697);
nand U6442 (N_6442,N_5735,N_5967);
xnor U6443 (N_6443,N_6377,N_5925);
xor U6444 (N_6444,N_5810,N_5933);
nand U6445 (N_6445,N_5787,N_6362);
xnor U6446 (N_6446,N_5785,N_6233);
and U6447 (N_6447,N_5887,N_5686);
or U6448 (N_6448,N_6172,N_5961);
nor U6449 (N_6449,N_6270,N_6258);
or U6450 (N_6450,N_6275,N_5984);
nor U6451 (N_6451,N_6026,N_5916);
and U6452 (N_6452,N_5901,N_5633);
and U6453 (N_6453,N_5790,N_6176);
nand U6454 (N_6454,N_6369,N_5816);
nand U6455 (N_6455,N_5841,N_5931);
or U6456 (N_6456,N_6329,N_5949);
xnor U6457 (N_6457,N_5619,N_6006);
nand U6458 (N_6458,N_6074,N_5836);
or U6459 (N_6459,N_5957,N_6059);
nand U6460 (N_6460,N_6277,N_5740);
and U6461 (N_6461,N_6217,N_5978);
nor U6462 (N_6462,N_5732,N_6097);
nor U6463 (N_6463,N_6094,N_5634);
nand U6464 (N_6464,N_6366,N_6009);
or U6465 (N_6465,N_5831,N_6073);
nand U6466 (N_6466,N_6030,N_5765);
nor U6467 (N_6467,N_5731,N_5757);
xnor U6468 (N_6468,N_5891,N_6320);
nand U6469 (N_6469,N_5802,N_5741);
nand U6470 (N_6470,N_5935,N_5970);
nor U6471 (N_6471,N_5938,N_6050);
nand U6472 (N_6472,N_5833,N_6387);
and U6473 (N_6473,N_6339,N_6212);
xor U6474 (N_6474,N_6345,N_6188);
xor U6475 (N_6475,N_6118,N_5695);
nor U6476 (N_6476,N_6202,N_6027);
nor U6477 (N_6477,N_6142,N_5779);
nor U6478 (N_6478,N_5956,N_6357);
xor U6479 (N_6479,N_6042,N_6174);
and U6480 (N_6480,N_5801,N_6286);
or U6481 (N_6481,N_6252,N_6295);
xnor U6482 (N_6482,N_5600,N_6163);
and U6483 (N_6483,N_5806,N_6114);
or U6484 (N_6484,N_6239,N_6351);
and U6485 (N_6485,N_5930,N_6084);
xor U6486 (N_6486,N_5800,N_5652);
nor U6487 (N_6487,N_5872,N_5824);
xor U6488 (N_6488,N_5880,N_5855);
or U6489 (N_6489,N_6312,N_6261);
and U6490 (N_6490,N_5775,N_6186);
nor U6491 (N_6491,N_6112,N_6304);
nor U6492 (N_6492,N_6251,N_6256);
or U6493 (N_6493,N_5692,N_6116);
nand U6494 (N_6494,N_5771,N_5711);
nand U6495 (N_6495,N_6308,N_5960);
xnor U6496 (N_6496,N_5850,N_6081);
xor U6497 (N_6497,N_5700,N_5918);
xnor U6498 (N_6498,N_6259,N_5675);
nand U6499 (N_6499,N_5747,N_5821);
xor U6500 (N_6500,N_5843,N_5649);
xnor U6501 (N_6501,N_5777,N_6289);
nand U6502 (N_6502,N_6184,N_6130);
and U6503 (N_6503,N_6151,N_6071);
or U6504 (N_6504,N_6046,N_5761);
or U6505 (N_6505,N_6106,N_5687);
nor U6506 (N_6506,N_6051,N_6031);
nor U6507 (N_6507,N_6054,N_6379);
or U6508 (N_6508,N_6102,N_6144);
or U6509 (N_6509,N_6150,N_6086);
nor U6510 (N_6510,N_5705,N_6299);
and U6511 (N_6511,N_6209,N_6185);
nor U6512 (N_6512,N_5998,N_6005);
or U6513 (N_6513,N_5715,N_5764);
nand U6514 (N_6514,N_5944,N_6350);
nand U6515 (N_6515,N_6105,N_5680);
nor U6516 (N_6516,N_5994,N_6352);
xor U6517 (N_6517,N_5677,N_6010);
nor U6518 (N_6518,N_6371,N_6340);
xor U6519 (N_6519,N_6359,N_5762);
xnor U6520 (N_6520,N_5953,N_5666);
or U6521 (N_6521,N_6298,N_6262);
or U6522 (N_6522,N_5941,N_6146);
and U6523 (N_6523,N_6120,N_6336);
xnor U6524 (N_6524,N_6398,N_5753);
and U6525 (N_6525,N_6267,N_5848);
and U6526 (N_6526,N_5822,N_5674);
and U6527 (N_6527,N_6044,N_5694);
and U6528 (N_6528,N_6082,N_6249);
xor U6529 (N_6529,N_6131,N_6175);
and U6530 (N_6530,N_6002,N_6316);
and U6531 (N_6531,N_5804,N_6374);
nor U6532 (N_6532,N_5870,N_6072);
xnor U6533 (N_6533,N_6248,N_5709);
nor U6534 (N_6534,N_5751,N_5987);
nand U6535 (N_6535,N_6392,N_6376);
and U6536 (N_6536,N_6178,N_5875);
or U6537 (N_6537,N_6113,N_6048);
nor U6538 (N_6538,N_6322,N_5865);
nand U6539 (N_6539,N_6257,N_6061);
xnor U6540 (N_6540,N_5607,N_6043);
nor U6541 (N_6541,N_6075,N_5693);
or U6542 (N_6542,N_6324,N_6236);
or U6543 (N_6543,N_5886,N_6279);
and U6544 (N_6544,N_6356,N_6108);
nor U6545 (N_6545,N_5676,N_5975);
and U6546 (N_6546,N_6347,N_5645);
or U6547 (N_6547,N_6134,N_6319);
nor U6548 (N_6548,N_6370,N_6091);
or U6549 (N_6549,N_6354,N_5628);
nor U6550 (N_6550,N_5642,N_6360);
nor U6551 (N_6551,N_5609,N_5797);
xnor U6552 (N_6552,N_5621,N_6255);
and U6553 (N_6553,N_5727,N_6232);
nor U6554 (N_6554,N_5883,N_6292);
or U6555 (N_6555,N_5660,N_6396);
or U6556 (N_6556,N_5879,N_5671);
nor U6557 (N_6557,N_5838,N_5781);
nor U6558 (N_6558,N_5745,N_5728);
or U6559 (N_6559,N_6159,N_5972);
nand U6560 (N_6560,N_6068,N_5958);
nand U6561 (N_6561,N_5667,N_5849);
xor U6562 (N_6562,N_5729,N_5683);
xnor U6563 (N_6563,N_5834,N_6206);
or U6564 (N_6564,N_6220,N_5639);
and U6565 (N_6565,N_5863,N_6305);
nand U6566 (N_6566,N_6095,N_6171);
xor U6567 (N_6567,N_5983,N_5688);
or U6568 (N_6568,N_6079,N_6021);
nand U6569 (N_6569,N_5827,N_6137);
and U6570 (N_6570,N_5730,N_5610);
nor U6571 (N_6571,N_6216,N_5835);
or U6572 (N_6572,N_6037,N_5906);
and U6573 (N_6573,N_5689,N_5955);
nor U6574 (N_6574,N_5703,N_6149);
nor U6575 (N_6575,N_5862,N_5712);
or U6576 (N_6576,N_5766,N_6022);
or U6577 (N_6577,N_6293,N_5768);
nor U6578 (N_6578,N_5853,N_5723);
xor U6579 (N_6579,N_5685,N_6124);
nor U6580 (N_6580,N_6034,N_5664);
or U6581 (N_6581,N_5754,N_5721);
or U6582 (N_6582,N_5602,N_6058);
and U6583 (N_6583,N_6273,N_6090);
xnor U6584 (N_6584,N_5909,N_5878);
nor U6585 (N_6585,N_5954,N_6136);
and U6586 (N_6586,N_6140,N_6303);
nor U6587 (N_6587,N_6127,N_6160);
nand U6588 (N_6588,N_6103,N_5981);
nand U6589 (N_6589,N_5907,N_6241);
nand U6590 (N_6590,N_5959,N_5873);
nand U6591 (N_6591,N_5940,N_6065);
xnor U6592 (N_6592,N_6049,N_5661);
xor U6593 (N_6593,N_5825,N_6139);
nor U6594 (N_6594,N_5977,N_6395);
nor U6595 (N_6595,N_6035,N_5659);
nand U6596 (N_6596,N_6314,N_6197);
or U6597 (N_6597,N_6080,N_5791);
or U6598 (N_6598,N_6066,N_6348);
xor U6599 (N_6599,N_6004,N_6064);
or U6600 (N_6600,N_5943,N_6250);
nand U6601 (N_6601,N_6331,N_5805);
nor U6602 (N_6602,N_5928,N_6158);
nor U6603 (N_6603,N_5882,N_5997);
nor U6604 (N_6604,N_5876,N_5698);
nor U6605 (N_6605,N_6391,N_6297);
and U6606 (N_6606,N_6245,N_6045);
xor U6607 (N_6607,N_5734,N_5656);
or U6608 (N_6608,N_5892,N_5663);
or U6609 (N_6609,N_5820,N_5620);
nand U6610 (N_6610,N_5991,N_5910);
nor U6611 (N_6611,N_6157,N_5922);
nor U6612 (N_6612,N_6089,N_6361);
xor U6613 (N_6613,N_6179,N_5974);
or U6614 (N_6614,N_6085,N_5867);
nor U6615 (N_6615,N_6008,N_5737);
nand U6616 (N_6616,N_5914,N_5829);
and U6617 (N_6617,N_5622,N_5699);
or U6618 (N_6618,N_5783,N_5690);
or U6619 (N_6619,N_6191,N_6019);
nand U6620 (N_6620,N_5857,N_5679);
xnor U6621 (N_6621,N_5742,N_5934);
nor U6622 (N_6622,N_6218,N_6180);
nor U6623 (N_6623,N_6390,N_6016);
and U6624 (N_6624,N_6155,N_6311);
nor U6625 (N_6625,N_6083,N_6382);
or U6626 (N_6626,N_6145,N_6317);
nand U6627 (N_6627,N_6032,N_5971);
xor U6628 (N_6628,N_6111,N_6228);
and U6629 (N_6629,N_6334,N_6183);
nor U6630 (N_6630,N_6126,N_5746);
nor U6631 (N_6631,N_5912,N_6269);
nor U6632 (N_6632,N_6284,N_6307);
nor U6633 (N_6633,N_6122,N_6399);
and U6634 (N_6634,N_6325,N_6003);
and U6635 (N_6635,N_5815,N_5662);
or U6636 (N_6636,N_6274,N_6237);
and U6637 (N_6637,N_6240,N_6332);
xnor U6638 (N_6638,N_5932,N_6047);
or U6639 (N_6639,N_5691,N_6244);
or U6640 (N_6640,N_5877,N_5989);
and U6641 (N_6641,N_6190,N_5904);
and U6642 (N_6642,N_5653,N_5604);
xor U6643 (N_6643,N_6222,N_6229);
nor U6644 (N_6644,N_5672,N_5733);
and U6645 (N_6645,N_5830,N_6187);
nor U6646 (N_6646,N_5760,N_5923);
or U6647 (N_6647,N_6287,N_6384);
nor U6648 (N_6648,N_5613,N_5897);
xnor U6649 (N_6649,N_5718,N_5710);
and U6650 (N_6650,N_5655,N_6242);
nor U6651 (N_6651,N_6266,N_5950);
xnor U6652 (N_6652,N_6343,N_5920);
or U6653 (N_6653,N_5641,N_5750);
nand U6654 (N_6654,N_5993,N_6011);
nor U6655 (N_6655,N_5895,N_5658);
xnor U6656 (N_6656,N_6201,N_6378);
nand U6657 (N_6657,N_6062,N_5635);
or U6658 (N_6658,N_6087,N_5774);
and U6659 (N_6659,N_5913,N_5702);
or U6660 (N_6660,N_6271,N_6170);
nand U6661 (N_6661,N_6117,N_5748);
nand U6662 (N_6662,N_5752,N_6355);
or U6663 (N_6663,N_6349,N_5637);
and U6664 (N_6664,N_5669,N_5631);
nor U6665 (N_6665,N_5937,N_5847);
and U6666 (N_6666,N_6096,N_5965);
nor U6667 (N_6667,N_5743,N_5856);
nand U6668 (N_6668,N_5657,N_6235);
xor U6669 (N_6669,N_5713,N_6385);
xor U6670 (N_6670,N_5813,N_6055);
nand U6671 (N_6671,N_5903,N_6092);
or U6672 (N_6672,N_6335,N_6000);
xnor U6673 (N_6673,N_5969,N_5939);
and U6674 (N_6674,N_6036,N_6128);
nand U6675 (N_6675,N_5744,N_5986);
nor U6676 (N_6676,N_5722,N_6067);
nor U6677 (N_6677,N_5756,N_5874);
xor U6678 (N_6678,N_6167,N_5654);
xnor U6679 (N_6679,N_5611,N_6358);
or U6680 (N_6680,N_5638,N_5665);
nor U6681 (N_6681,N_6310,N_5786);
xor U6682 (N_6682,N_6388,N_5707);
nor U6683 (N_6683,N_5842,N_6023);
and U6684 (N_6684,N_6300,N_6213);
xnor U6685 (N_6685,N_6093,N_6132);
and U6686 (N_6686,N_6024,N_5648);
or U6687 (N_6687,N_6226,N_6135);
xor U6688 (N_6688,N_5979,N_6207);
or U6689 (N_6689,N_6306,N_6227);
nand U6690 (N_6690,N_6294,N_5826);
nor U6691 (N_6691,N_6338,N_5988);
nor U6692 (N_6692,N_5796,N_6327);
or U6693 (N_6693,N_5605,N_6038);
xnor U6694 (N_6694,N_6012,N_5899);
nand U6695 (N_6695,N_6234,N_6373);
and U6696 (N_6696,N_6153,N_6247);
and U6697 (N_6697,N_5725,N_5947);
or U6698 (N_6698,N_6015,N_6372);
and U6699 (N_6699,N_5936,N_5809);
and U6700 (N_6700,N_6100,N_5629);
nor U6701 (N_6701,N_5861,N_6214);
nand U6702 (N_6702,N_5860,N_6166);
xor U6703 (N_6703,N_6193,N_5617);
or U6704 (N_6704,N_6321,N_6177);
xnor U6705 (N_6705,N_5811,N_6315);
nor U6706 (N_6706,N_6057,N_6053);
xor U6707 (N_6707,N_5708,N_5618);
nor U6708 (N_6708,N_5792,N_5789);
xor U6709 (N_6709,N_5643,N_6386);
or U6710 (N_6710,N_5717,N_5769);
nand U6711 (N_6711,N_5837,N_6363);
or U6712 (N_6712,N_6109,N_5812);
or U6713 (N_6713,N_5819,N_6182);
nand U6714 (N_6714,N_5968,N_6224);
or U6715 (N_6715,N_6375,N_6394);
nand U6716 (N_6716,N_5990,N_6365);
nand U6717 (N_6717,N_6302,N_6060);
and U6718 (N_6718,N_6147,N_6194);
nand U6719 (N_6719,N_6039,N_5846);
xor U6720 (N_6720,N_5888,N_5818);
or U6721 (N_6721,N_6344,N_6333);
or U6722 (N_6722,N_6041,N_5852);
and U6723 (N_6723,N_5739,N_6025);
and U6724 (N_6724,N_5770,N_5630);
nand U6725 (N_6725,N_5646,N_5982);
nor U6726 (N_6726,N_5626,N_5773);
or U6727 (N_6727,N_5985,N_5898);
xnor U6728 (N_6728,N_6223,N_6393);
nor U6729 (N_6729,N_6107,N_5716);
and U6730 (N_6730,N_6323,N_6028);
nor U6731 (N_6731,N_6018,N_5881);
and U6732 (N_6732,N_5724,N_5788);
and U6733 (N_6733,N_5782,N_5636);
nor U6734 (N_6734,N_5951,N_6368);
nand U6735 (N_6735,N_5866,N_5945);
or U6736 (N_6736,N_6397,N_5851);
xnor U6737 (N_6737,N_6138,N_5670);
nor U6738 (N_6738,N_5749,N_5999);
xor U6739 (N_6739,N_6381,N_5632);
xor U6740 (N_6740,N_5885,N_5678);
xnor U6741 (N_6741,N_6119,N_5807);
nor U6742 (N_6742,N_6143,N_6281);
xnor U6743 (N_6743,N_6192,N_5844);
and U6744 (N_6744,N_6203,N_6164);
nand U6745 (N_6745,N_6141,N_6199);
and U6746 (N_6746,N_6225,N_5973);
or U6747 (N_6747,N_5736,N_6148);
nor U6748 (N_6748,N_5776,N_6070);
or U6749 (N_6749,N_5868,N_5608);
xor U6750 (N_6750,N_6364,N_5668);
nor U6751 (N_6751,N_6208,N_5927);
or U6752 (N_6752,N_5651,N_5755);
and U6753 (N_6753,N_5784,N_6276);
nand U6754 (N_6754,N_6110,N_5673);
nor U6755 (N_6755,N_6309,N_6063);
nand U6756 (N_6756,N_5615,N_5858);
and U6757 (N_6757,N_6013,N_6272);
nor U6758 (N_6758,N_6204,N_6133);
or U6759 (N_6759,N_6283,N_5893);
or U6760 (N_6760,N_5612,N_6296);
or U6761 (N_6761,N_6020,N_6291);
xnor U6762 (N_6762,N_6007,N_5929);
xor U6763 (N_6763,N_5799,N_5601);
and U6764 (N_6764,N_5864,N_6165);
and U6765 (N_6765,N_5996,N_5794);
and U6766 (N_6766,N_6040,N_6268);
nor U6767 (N_6767,N_5772,N_6173);
nand U6768 (N_6768,N_6230,N_5767);
xnor U6769 (N_6769,N_5780,N_5720);
and U6770 (N_6770,N_6098,N_5808);
or U6771 (N_6771,N_6195,N_6246);
nor U6772 (N_6772,N_6215,N_6056);
xor U6773 (N_6773,N_5650,N_5817);
xnor U6774 (N_6774,N_6219,N_6014);
nand U6775 (N_6775,N_6330,N_6380);
nor U6776 (N_6776,N_5952,N_6210);
or U6777 (N_6777,N_5890,N_5704);
xor U6778 (N_6778,N_5778,N_6263);
and U6779 (N_6779,N_5946,N_5942);
xnor U6780 (N_6780,N_5758,N_5921);
nor U6781 (N_6781,N_5616,N_5706);
and U6782 (N_6782,N_5976,N_6033);
xor U6783 (N_6783,N_6278,N_6161);
nand U6784 (N_6784,N_6346,N_5696);
or U6785 (N_6785,N_5719,N_5911);
nand U6786 (N_6786,N_6264,N_6129);
nand U6787 (N_6787,N_5889,N_6196);
or U6788 (N_6788,N_5795,N_5869);
nor U6789 (N_6789,N_5924,N_6104);
nor U6790 (N_6790,N_5714,N_5962);
and U6791 (N_6791,N_5814,N_5701);
nor U6792 (N_6792,N_6123,N_5980);
nand U6793 (N_6793,N_6260,N_5644);
or U6794 (N_6794,N_6231,N_6125);
or U6795 (N_6795,N_6077,N_6154);
xnor U6796 (N_6796,N_6205,N_6282);
nor U6797 (N_6797,N_6168,N_6152);
xnor U6798 (N_6798,N_6326,N_5832);
xnor U6799 (N_6799,N_5964,N_6001);
and U6800 (N_6800,N_6089,N_6230);
nor U6801 (N_6801,N_6331,N_5996);
or U6802 (N_6802,N_5874,N_5878);
nor U6803 (N_6803,N_6114,N_6041);
nor U6804 (N_6804,N_6243,N_6360);
and U6805 (N_6805,N_5704,N_6274);
and U6806 (N_6806,N_5896,N_5823);
nand U6807 (N_6807,N_6129,N_5826);
or U6808 (N_6808,N_6091,N_6000);
xnor U6809 (N_6809,N_6117,N_6188);
nand U6810 (N_6810,N_5991,N_5802);
and U6811 (N_6811,N_6342,N_6109);
nand U6812 (N_6812,N_5936,N_6250);
or U6813 (N_6813,N_6372,N_6389);
and U6814 (N_6814,N_6141,N_5994);
and U6815 (N_6815,N_5961,N_6128);
or U6816 (N_6816,N_5966,N_6396);
nor U6817 (N_6817,N_5893,N_6222);
or U6818 (N_6818,N_5691,N_6071);
nor U6819 (N_6819,N_6362,N_6396);
or U6820 (N_6820,N_6168,N_5780);
nor U6821 (N_6821,N_5738,N_5610);
or U6822 (N_6822,N_6079,N_6165);
nor U6823 (N_6823,N_5793,N_6350);
nand U6824 (N_6824,N_5965,N_6033);
and U6825 (N_6825,N_5991,N_6172);
and U6826 (N_6826,N_5611,N_5628);
nand U6827 (N_6827,N_5762,N_5938);
xor U6828 (N_6828,N_6265,N_6302);
nor U6829 (N_6829,N_6340,N_6381);
nor U6830 (N_6830,N_6193,N_5921);
and U6831 (N_6831,N_5697,N_5608);
and U6832 (N_6832,N_6191,N_5773);
nor U6833 (N_6833,N_5799,N_6283);
and U6834 (N_6834,N_5996,N_5881);
xor U6835 (N_6835,N_6176,N_5714);
and U6836 (N_6836,N_5978,N_5812);
or U6837 (N_6837,N_5992,N_6079);
and U6838 (N_6838,N_5741,N_5774);
and U6839 (N_6839,N_6390,N_6120);
and U6840 (N_6840,N_6024,N_6172);
nand U6841 (N_6841,N_5662,N_5817);
or U6842 (N_6842,N_6361,N_6122);
nand U6843 (N_6843,N_5699,N_5656);
nor U6844 (N_6844,N_5743,N_6158);
and U6845 (N_6845,N_5782,N_6094);
xor U6846 (N_6846,N_6088,N_6180);
nor U6847 (N_6847,N_6324,N_6001);
nand U6848 (N_6848,N_6141,N_6223);
xor U6849 (N_6849,N_6333,N_5976);
nor U6850 (N_6850,N_5798,N_5756);
and U6851 (N_6851,N_6153,N_6294);
nand U6852 (N_6852,N_6211,N_6152);
xnor U6853 (N_6853,N_6285,N_6351);
nor U6854 (N_6854,N_5660,N_6268);
xnor U6855 (N_6855,N_5780,N_5716);
xor U6856 (N_6856,N_6301,N_5696);
xor U6857 (N_6857,N_5873,N_5877);
xor U6858 (N_6858,N_5615,N_6098);
and U6859 (N_6859,N_5677,N_5849);
and U6860 (N_6860,N_5668,N_5603);
xnor U6861 (N_6861,N_6382,N_6126);
and U6862 (N_6862,N_6357,N_5686);
and U6863 (N_6863,N_6213,N_6087);
or U6864 (N_6864,N_6077,N_6201);
nor U6865 (N_6865,N_5618,N_6142);
xor U6866 (N_6866,N_6224,N_6169);
and U6867 (N_6867,N_5738,N_6342);
and U6868 (N_6868,N_6114,N_6396);
nand U6869 (N_6869,N_5644,N_6372);
xor U6870 (N_6870,N_6360,N_5904);
nand U6871 (N_6871,N_5607,N_5633);
nor U6872 (N_6872,N_6144,N_6125);
xnor U6873 (N_6873,N_5866,N_5781);
nor U6874 (N_6874,N_5835,N_6088);
nand U6875 (N_6875,N_5859,N_5896);
nand U6876 (N_6876,N_6320,N_5810);
xor U6877 (N_6877,N_6274,N_6318);
xor U6878 (N_6878,N_5823,N_6256);
nor U6879 (N_6879,N_5743,N_6379);
or U6880 (N_6880,N_5999,N_5781);
and U6881 (N_6881,N_5749,N_6254);
xnor U6882 (N_6882,N_5783,N_5982);
nand U6883 (N_6883,N_6157,N_5806);
nor U6884 (N_6884,N_6075,N_6257);
and U6885 (N_6885,N_5633,N_5707);
nand U6886 (N_6886,N_5657,N_5925);
xor U6887 (N_6887,N_6238,N_6071);
or U6888 (N_6888,N_6016,N_5818);
or U6889 (N_6889,N_5634,N_5655);
or U6890 (N_6890,N_5756,N_5994);
and U6891 (N_6891,N_5716,N_5735);
or U6892 (N_6892,N_5897,N_5951);
or U6893 (N_6893,N_5611,N_5919);
nand U6894 (N_6894,N_5753,N_5942);
or U6895 (N_6895,N_6028,N_5910);
nand U6896 (N_6896,N_5871,N_5881);
nand U6897 (N_6897,N_5898,N_6396);
xor U6898 (N_6898,N_5700,N_6334);
or U6899 (N_6899,N_6054,N_5838);
nor U6900 (N_6900,N_5749,N_6258);
nand U6901 (N_6901,N_5990,N_6136);
nand U6902 (N_6902,N_6108,N_6304);
nor U6903 (N_6903,N_6125,N_5782);
xor U6904 (N_6904,N_6165,N_5748);
xnor U6905 (N_6905,N_5996,N_6197);
and U6906 (N_6906,N_5838,N_5723);
xor U6907 (N_6907,N_5824,N_5887);
xnor U6908 (N_6908,N_6021,N_6108);
nor U6909 (N_6909,N_5739,N_6271);
xnor U6910 (N_6910,N_6149,N_5958);
nor U6911 (N_6911,N_6336,N_5923);
nand U6912 (N_6912,N_6167,N_5963);
nor U6913 (N_6913,N_5851,N_6097);
or U6914 (N_6914,N_5964,N_6135);
nand U6915 (N_6915,N_6166,N_6087);
nor U6916 (N_6916,N_6105,N_5912);
xor U6917 (N_6917,N_6118,N_5995);
and U6918 (N_6918,N_6000,N_5606);
xor U6919 (N_6919,N_6009,N_6077);
or U6920 (N_6920,N_5621,N_5899);
nor U6921 (N_6921,N_5764,N_5885);
or U6922 (N_6922,N_6234,N_6168);
nor U6923 (N_6923,N_6036,N_5923);
or U6924 (N_6924,N_6077,N_6007);
nor U6925 (N_6925,N_5612,N_5788);
nor U6926 (N_6926,N_6298,N_6127);
and U6927 (N_6927,N_5873,N_5921);
nor U6928 (N_6928,N_5968,N_6377);
nor U6929 (N_6929,N_5639,N_6139);
and U6930 (N_6930,N_6226,N_5789);
nand U6931 (N_6931,N_6274,N_6236);
or U6932 (N_6932,N_6335,N_6341);
nand U6933 (N_6933,N_6327,N_5832);
xnor U6934 (N_6934,N_6127,N_6074);
xnor U6935 (N_6935,N_5710,N_5925);
and U6936 (N_6936,N_5600,N_6378);
nor U6937 (N_6937,N_6297,N_6384);
or U6938 (N_6938,N_6108,N_5964);
xnor U6939 (N_6939,N_6132,N_5815);
and U6940 (N_6940,N_6282,N_6126);
xnor U6941 (N_6941,N_5805,N_6114);
and U6942 (N_6942,N_6025,N_5999);
nand U6943 (N_6943,N_6039,N_6158);
and U6944 (N_6944,N_5619,N_5680);
nand U6945 (N_6945,N_5698,N_6192);
nor U6946 (N_6946,N_5946,N_6055);
nor U6947 (N_6947,N_6109,N_6161);
or U6948 (N_6948,N_5642,N_5920);
and U6949 (N_6949,N_6106,N_6295);
or U6950 (N_6950,N_6386,N_5869);
or U6951 (N_6951,N_6263,N_6205);
and U6952 (N_6952,N_6314,N_6052);
or U6953 (N_6953,N_6345,N_5909);
and U6954 (N_6954,N_6282,N_6328);
and U6955 (N_6955,N_6334,N_6100);
nand U6956 (N_6956,N_5732,N_6183);
xnor U6957 (N_6957,N_5862,N_6080);
and U6958 (N_6958,N_5842,N_6049);
xnor U6959 (N_6959,N_6202,N_5671);
and U6960 (N_6960,N_5860,N_5770);
xor U6961 (N_6961,N_5779,N_5764);
and U6962 (N_6962,N_5711,N_5943);
and U6963 (N_6963,N_6357,N_6102);
and U6964 (N_6964,N_5984,N_6341);
nor U6965 (N_6965,N_6268,N_6087);
nor U6966 (N_6966,N_5858,N_5642);
nor U6967 (N_6967,N_5751,N_6268);
and U6968 (N_6968,N_5611,N_6236);
xnor U6969 (N_6969,N_6079,N_5682);
xor U6970 (N_6970,N_6304,N_5624);
and U6971 (N_6971,N_5680,N_5626);
and U6972 (N_6972,N_5998,N_6395);
nand U6973 (N_6973,N_5667,N_6182);
xnor U6974 (N_6974,N_6314,N_5933);
nor U6975 (N_6975,N_6214,N_5717);
nand U6976 (N_6976,N_5913,N_6348);
nand U6977 (N_6977,N_6116,N_5768);
and U6978 (N_6978,N_5632,N_5749);
nand U6979 (N_6979,N_6077,N_5704);
and U6980 (N_6980,N_5958,N_5648);
and U6981 (N_6981,N_6076,N_5790);
and U6982 (N_6982,N_6367,N_5778);
or U6983 (N_6983,N_5789,N_6289);
or U6984 (N_6984,N_5637,N_5762);
or U6985 (N_6985,N_5611,N_5994);
nor U6986 (N_6986,N_6229,N_6308);
or U6987 (N_6987,N_6310,N_6100);
and U6988 (N_6988,N_6172,N_6076);
nand U6989 (N_6989,N_6106,N_5881);
nor U6990 (N_6990,N_5934,N_6367);
or U6991 (N_6991,N_6081,N_5751);
xor U6992 (N_6992,N_5949,N_6159);
nor U6993 (N_6993,N_6290,N_6087);
xor U6994 (N_6994,N_6264,N_6316);
nand U6995 (N_6995,N_6255,N_5975);
nand U6996 (N_6996,N_5945,N_6371);
nor U6997 (N_6997,N_6270,N_6082);
nor U6998 (N_6998,N_5889,N_5896);
or U6999 (N_6999,N_6013,N_5688);
and U7000 (N_7000,N_6057,N_5721);
and U7001 (N_7001,N_5963,N_6215);
xnor U7002 (N_7002,N_5981,N_5855);
and U7003 (N_7003,N_6142,N_6328);
or U7004 (N_7004,N_6207,N_6262);
or U7005 (N_7005,N_6239,N_6155);
or U7006 (N_7006,N_5621,N_6204);
or U7007 (N_7007,N_5947,N_6211);
nand U7008 (N_7008,N_6217,N_5757);
or U7009 (N_7009,N_6014,N_5771);
or U7010 (N_7010,N_5795,N_6275);
xor U7011 (N_7011,N_5611,N_6028);
nand U7012 (N_7012,N_6367,N_6269);
and U7013 (N_7013,N_5981,N_5954);
xnor U7014 (N_7014,N_6261,N_5872);
nand U7015 (N_7015,N_6275,N_6258);
nor U7016 (N_7016,N_6048,N_6248);
xnor U7017 (N_7017,N_5856,N_5730);
nor U7018 (N_7018,N_5992,N_6332);
nand U7019 (N_7019,N_6154,N_6203);
nand U7020 (N_7020,N_5625,N_5950);
nor U7021 (N_7021,N_6192,N_5985);
nand U7022 (N_7022,N_6126,N_5647);
and U7023 (N_7023,N_6273,N_6245);
nand U7024 (N_7024,N_6220,N_5619);
nand U7025 (N_7025,N_6045,N_6325);
or U7026 (N_7026,N_5997,N_6176);
and U7027 (N_7027,N_5783,N_6393);
or U7028 (N_7028,N_6224,N_6073);
or U7029 (N_7029,N_6187,N_6388);
nor U7030 (N_7030,N_6205,N_5669);
nor U7031 (N_7031,N_5679,N_5759);
and U7032 (N_7032,N_5655,N_6047);
and U7033 (N_7033,N_5817,N_6027);
nor U7034 (N_7034,N_6293,N_5609);
or U7035 (N_7035,N_5741,N_5744);
xor U7036 (N_7036,N_6099,N_6067);
nor U7037 (N_7037,N_5899,N_6293);
or U7038 (N_7038,N_5931,N_5614);
and U7039 (N_7039,N_6276,N_5627);
nand U7040 (N_7040,N_5897,N_5845);
xor U7041 (N_7041,N_6041,N_5824);
nor U7042 (N_7042,N_6130,N_6330);
or U7043 (N_7043,N_6141,N_5860);
or U7044 (N_7044,N_5887,N_6154);
nor U7045 (N_7045,N_6261,N_5892);
or U7046 (N_7046,N_6301,N_6329);
or U7047 (N_7047,N_5964,N_5751);
nand U7048 (N_7048,N_5769,N_5869);
xor U7049 (N_7049,N_5887,N_6337);
and U7050 (N_7050,N_6151,N_6127);
xor U7051 (N_7051,N_5748,N_6150);
nor U7052 (N_7052,N_5798,N_6051);
nor U7053 (N_7053,N_5798,N_6018);
xor U7054 (N_7054,N_6250,N_6254);
or U7055 (N_7055,N_6251,N_6292);
or U7056 (N_7056,N_6061,N_6397);
and U7057 (N_7057,N_5799,N_6274);
xnor U7058 (N_7058,N_6228,N_5953);
nand U7059 (N_7059,N_5906,N_6088);
nand U7060 (N_7060,N_5673,N_5947);
nor U7061 (N_7061,N_5888,N_5621);
or U7062 (N_7062,N_5698,N_6375);
nor U7063 (N_7063,N_6287,N_5982);
or U7064 (N_7064,N_6101,N_5668);
or U7065 (N_7065,N_6364,N_5781);
nand U7066 (N_7066,N_6064,N_5668);
and U7067 (N_7067,N_5877,N_5692);
or U7068 (N_7068,N_6009,N_5751);
nand U7069 (N_7069,N_5769,N_5665);
xor U7070 (N_7070,N_5714,N_6141);
xnor U7071 (N_7071,N_6113,N_6075);
nand U7072 (N_7072,N_6027,N_5673);
xnor U7073 (N_7073,N_5852,N_6044);
nor U7074 (N_7074,N_6279,N_5683);
nand U7075 (N_7075,N_6345,N_5978);
or U7076 (N_7076,N_5763,N_6272);
and U7077 (N_7077,N_6257,N_6249);
xor U7078 (N_7078,N_5858,N_5838);
xnor U7079 (N_7079,N_6355,N_6157);
nor U7080 (N_7080,N_5744,N_6121);
nor U7081 (N_7081,N_5727,N_5854);
nand U7082 (N_7082,N_6331,N_5770);
nor U7083 (N_7083,N_6009,N_6311);
and U7084 (N_7084,N_5649,N_5809);
nand U7085 (N_7085,N_6039,N_5863);
nor U7086 (N_7086,N_5649,N_6148);
xnor U7087 (N_7087,N_5778,N_6271);
and U7088 (N_7088,N_6355,N_5797);
xor U7089 (N_7089,N_6253,N_5660);
nand U7090 (N_7090,N_6100,N_6369);
nor U7091 (N_7091,N_5875,N_6074);
or U7092 (N_7092,N_6016,N_6077);
nand U7093 (N_7093,N_5958,N_6339);
or U7094 (N_7094,N_6340,N_5641);
xnor U7095 (N_7095,N_5671,N_5882);
nor U7096 (N_7096,N_6338,N_5643);
nand U7097 (N_7097,N_6241,N_5767);
and U7098 (N_7098,N_6274,N_6234);
nand U7099 (N_7099,N_5789,N_6232);
xor U7100 (N_7100,N_6259,N_6087);
nor U7101 (N_7101,N_5903,N_5682);
nand U7102 (N_7102,N_6063,N_6060);
nand U7103 (N_7103,N_6396,N_6274);
nand U7104 (N_7104,N_5920,N_6387);
nand U7105 (N_7105,N_6233,N_5823);
nand U7106 (N_7106,N_5953,N_5711);
nand U7107 (N_7107,N_5946,N_5872);
and U7108 (N_7108,N_5690,N_5834);
xnor U7109 (N_7109,N_5894,N_5667);
or U7110 (N_7110,N_6059,N_6332);
nand U7111 (N_7111,N_6207,N_5699);
or U7112 (N_7112,N_5630,N_5671);
nand U7113 (N_7113,N_5772,N_6004);
nand U7114 (N_7114,N_6088,N_5778);
nor U7115 (N_7115,N_5741,N_5960);
nor U7116 (N_7116,N_5724,N_5798);
and U7117 (N_7117,N_5793,N_5938);
nand U7118 (N_7118,N_6020,N_6362);
and U7119 (N_7119,N_6080,N_5724);
and U7120 (N_7120,N_5968,N_6356);
or U7121 (N_7121,N_5612,N_6066);
xor U7122 (N_7122,N_6051,N_6223);
xor U7123 (N_7123,N_6042,N_5900);
or U7124 (N_7124,N_5683,N_6138);
nand U7125 (N_7125,N_6321,N_6145);
and U7126 (N_7126,N_5900,N_6090);
nor U7127 (N_7127,N_6034,N_5931);
or U7128 (N_7128,N_5882,N_5932);
xnor U7129 (N_7129,N_6387,N_6057);
and U7130 (N_7130,N_5899,N_5831);
or U7131 (N_7131,N_5794,N_6234);
nor U7132 (N_7132,N_6080,N_6066);
xor U7133 (N_7133,N_6398,N_6294);
and U7134 (N_7134,N_6370,N_5696);
or U7135 (N_7135,N_5841,N_5881);
or U7136 (N_7136,N_5849,N_6327);
xor U7137 (N_7137,N_5874,N_5950);
nor U7138 (N_7138,N_6072,N_6360);
and U7139 (N_7139,N_6050,N_6253);
or U7140 (N_7140,N_5829,N_6215);
xor U7141 (N_7141,N_5912,N_5829);
xor U7142 (N_7142,N_6287,N_6315);
nand U7143 (N_7143,N_5712,N_6193);
and U7144 (N_7144,N_6395,N_6329);
xnor U7145 (N_7145,N_6249,N_6203);
and U7146 (N_7146,N_6163,N_5649);
and U7147 (N_7147,N_6041,N_5912);
or U7148 (N_7148,N_6143,N_6396);
nor U7149 (N_7149,N_5789,N_6009);
nand U7150 (N_7150,N_5970,N_6377);
nand U7151 (N_7151,N_5664,N_6020);
xor U7152 (N_7152,N_5956,N_6094);
and U7153 (N_7153,N_6331,N_6359);
and U7154 (N_7154,N_6083,N_5617);
nand U7155 (N_7155,N_5947,N_5887);
nand U7156 (N_7156,N_5953,N_6239);
or U7157 (N_7157,N_6383,N_5761);
nand U7158 (N_7158,N_5837,N_5996);
nand U7159 (N_7159,N_5643,N_6259);
nor U7160 (N_7160,N_6276,N_5849);
xor U7161 (N_7161,N_5933,N_5981);
nor U7162 (N_7162,N_6085,N_5987);
nor U7163 (N_7163,N_5777,N_6188);
or U7164 (N_7164,N_6315,N_5605);
and U7165 (N_7165,N_6200,N_6345);
nor U7166 (N_7166,N_6290,N_6292);
xnor U7167 (N_7167,N_6213,N_6313);
xnor U7168 (N_7168,N_6119,N_6389);
and U7169 (N_7169,N_5852,N_6084);
and U7170 (N_7170,N_5628,N_5729);
or U7171 (N_7171,N_5657,N_6316);
nor U7172 (N_7172,N_5601,N_6381);
xor U7173 (N_7173,N_5840,N_5673);
nor U7174 (N_7174,N_5775,N_5736);
and U7175 (N_7175,N_6393,N_6076);
nor U7176 (N_7176,N_5608,N_5854);
xor U7177 (N_7177,N_6021,N_5808);
and U7178 (N_7178,N_6174,N_6260);
and U7179 (N_7179,N_6386,N_6397);
or U7180 (N_7180,N_6380,N_5845);
and U7181 (N_7181,N_6191,N_5969);
and U7182 (N_7182,N_5937,N_6192);
nor U7183 (N_7183,N_5934,N_6085);
nor U7184 (N_7184,N_5628,N_5932);
nor U7185 (N_7185,N_5802,N_5884);
xnor U7186 (N_7186,N_5771,N_5854);
or U7187 (N_7187,N_6028,N_6155);
or U7188 (N_7188,N_5685,N_6149);
and U7189 (N_7189,N_6368,N_5718);
xor U7190 (N_7190,N_5673,N_6225);
and U7191 (N_7191,N_5987,N_5835);
xor U7192 (N_7192,N_5873,N_5710);
xnor U7193 (N_7193,N_6266,N_5728);
nor U7194 (N_7194,N_6363,N_5999);
nor U7195 (N_7195,N_6111,N_6136);
nand U7196 (N_7196,N_6275,N_6310);
nor U7197 (N_7197,N_5836,N_5977);
xor U7198 (N_7198,N_5884,N_6319);
xnor U7199 (N_7199,N_6151,N_6290);
nor U7200 (N_7200,N_7098,N_6665);
and U7201 (N_7201,N_6460,N_6635);
nand U7202 (N_7202,N_6436,N_6552);
nor U7203 (N_7203,N_7180,N_6823);
and U7204 (N_7204,N_7021,N_6727);
nand U7205 (N_7205,N_6675,N_6775);
or U7206 (N_7206,N_7085,N_6414);
nand U7207 (N_7207,N_7078,N_6555);
nand U7208 (N_7208,N_6629,N_7036);
nand U7209 (N_7209,N_6982,N_7123);
xor U7210 (N_7210,N_6974,N_7013);
nor U7211 (N_7211,N_6899,N_6494);
xnor U7212 (N_7212,N_7096,N_6572);
or U7213 (N_7213,N_6706,N_6699);
or U7214 (N_7214,N_6631,N_6780);
and U7215 (N_7215,N_6554,N_6513);
or U7216 (N_7216,N_6569,N_6420);
and U7217 (N_7217,N_6924,N_6531);
xnor U7218 (N_7218,N_6789,N_6451);
nor U7219 (N_7219,N_6486,N_7110);
nand U7220 (N_7220,N_6603,N_6887);
nor U7221 (N_7221,N_6751,N_6556);
xnor U7222 (N_7222,N_6758,N_6406);
nand U7223 (N_7223,N_6830,N_7070);
or U7224 (N_7224,N_6688,N_6496);
nor U7225 (N_7225,N_6622,N_7097);
or U7226 (N_7226,N_6587,N_6841);
or U7227 (N_7227,N_6836,N_6452);
xor U7228 (N_7228,N_7064,N_6840);
nand U7229 (N_7229,N_7113,N_7145);
nand U7230 (N_7230,N_6803,N_7032);
xnor U7231 (N_7231,N_6626,N_7019);
xor U7232 (N_7232,N_6525,N_6915);
and U7233 (N_7233,N_6827,N_7191);
nor U7234 (N_7234,N_6644,N_6471);
nor U7235 (N_7235,N_6488,N_6655);
nor U7236 (N_7236,N_6870,N_6530);
or U7237 (N_7237,N_6875,N_6522);
nand U7238 (N_7238,N_6577,N_6683);
and U7239 (N_7239,N_6491,N_6457);
xor U7240 (N_7240,N_6582,N_7107);
xor U7241 (N_7241,N_7074,N_6772);
or U7242 (N_7242,N_6548,N_6692);
xnor U7243 (N_7243,N_6432,N_6740);
xor U7244 (N_7244,N_6422,N_6517);
xnor U7245 (N_7245,N_6987,N_6516);
xor U7246 (N_7246,N_6983,N_6779);
nand U7247 (N_7247,N_6431,N_6458);
and U7248 (N_7248,N_7161,N_6632);
or U7249 (N_7249,N_6979,N_6862);
nand U7250 (N_7250,N_6905,N_6616);
and U7251 (N_7251,N_6819,N_6993);
or U7252 (N_7252,N_7126,N_6508);
nor U7253 (N_7253,N_6829,N_7170);
and U7254 (N_7254,N_6636,N_6701);
or U7255 (N_7255,N_6678,N_6400);
xnor U7256 (N_7256,N_6663,N_6586);
xnor U7257 (N_7257,N_6935,N_7118);
xor U7258 (N_7258,N_6445,N_6553);
nand U7259 (N_7259,N_7017,N_6742);
nor U7260 (N_7260,N_6895,N_6746);
xnor U7261 (N_7261,N_7043,N_6575);
nand U7262 (N_7262,N_7117,N_6484);
nand U7263 (N_7263,N_6900,N_6777);
and U7264 (N_7264,N_6782,N_7060);
or U7265 (N_7265,N_6847,N_7157);
xor U7266 (N_7266,N_6704,N_6995);
xnor U7267 (N_7267,N_6628,N_6863);
and U7268 (N_7268,N_6788,N_6954);
nand U7269 (N_7269,N_6617,N_6591);
nor U7270 (N_7270,N_6401,N_6413);
and U7271 (N_7271,N_6690,N_7169);
or U7272 (N_7272,N_7094,N_6930);
xor U7273 (N_7273,N_7067,N_7027);
and U7274 (N_7274,N_6966,N_6792);
xnor U7275 (N_7275,N_6939,N_6910);
or U7276 (N_7276,N_7159,N_6957);
nand U7277 (N_7277,N_7086,N_6916);
and U7278 (N_7278,N_7024,N_7150);
nor U7279 (N_7279,N_6854,N_6456);
nand U7280 (N_7280,N_6934,N_7142);
nor U7281 (N_7281,N_7066,N_7035);
and U7282 (N_7282,N_6697,N_6927);
nor U7283 (N_7283,N_7073,N_6518);
and U7284 (N_7284,N_7090,N_7174);
or U7285 (N_7285,N_7058,N_6956);
and U7286 (N_7286,N_7114,N_6835);
nand U7287 (N_7287,N_7182,N_6909);
nand U7288 (N_7288,N_6502,N_6412);
nor U7289 (N_7289,N_6563,N_6737);
xnor U7290 (N_7290,N_7065,N_6495);
xnor U7291 (N_7291,N_6784,N_6943);
or U7292 (N_7292,N_7025,N_7130);
xor U7293 (N_7293,N_6681,N_6507);
or U7294 (N_7294,N_6756,N_6465);
and U7295 (N_7295,N_6951,N_7020);
or U7296 (N_7296,N_7111,N_6977);
or U7297 (N_7297,N_6973,N_6672);
or U7298 (N_7298,N_7038,N_7077);
or U7299 (N_7299,N_6947,N_7162);
or U7300 (N_7300,N_7015,N_7155);
nand U7301 (N_7301,N_7049,N_6748);
nand U7302 (N_7302,N_6833,N_6735);
nand U7303 (N_7303,N_6764,N_6477);
nor U7304 (N_7304,N_7028,N_6839);
and U7305 (N_7305,N_6579,N_6888);
and U7306 (N_7306,N_7132,N_6762);
nand U7307 (N_7307,N_6506,N_7047);
xnor U7308 (N_7308,N_6728,N_6892);
xor U7309 (N_7309,N_6442,N_6922);
or U7310 (N_7310,N_6882,N_6476);
or U7311 (N_7311,N_6851,N_6567);
and U7312 (N_7312,N_6886,N_6834);
or U7313 (N_7313,N_6670,N_7091);
xor U7314 (N_7314,N_7165,N_6410);
nand U7315 (N_7315,N_6593,N_7016);
xor U7316 (N_7316,N_7037,N_7102);
or U7317 (N_7317,N_6624,N_6405);
and U7318 (N_7318,N_6687,N_6529);
nand U7319 (N_7319,N_6416,N_6736);
nand U7320 (N_7320,N_6783,N_7108);
nand U7321 (N_7321,N_6913,N_6967);
or U7322 (N_7322,N_7121,N_6510);
xor U7323 (N_7323,N_6768,N_6744);
nor U7324 (N_7324,N_6489,N_6609);
nor U7325 (N_7325,N_7008,N_6565);
nand U7326 (N_7326,N_6437,N_6814);
xnor U7327 (N_7327,N_6599,N_6429);
nor U7328 (N_7328,N_6820,N_6642);
and U7329 (N_7329,N_6885,N_6997);
or U7330 (N_7330,N_6797,N_6970);
nor U7331 (N_7331,N_6485,N_6466);
and U7332 (N_7332,N_6509,N_6694);
and U7333 (N_7333,N_6448,N_6896);
nor U7334 (N_7334,N_6604,N_6868);
nand U7335 (N_7335,N_6865,N_6500);
or U7336 (N_7336,N_6972,N_7172);
nand U7337 (N_7337,N_6791,N_6621);
and U7338 (N_7338,N_6876,N_6656);
and U7339 (N_7339,N_6625,N_6950);
and U7340 (N_7340,N_6946,N_6848);
xor U7341 (N_7341,N_6686,N_7134);
nand U7342 (N_7342,N_6858,N_6707);
and U7343 (N_7343,N_7040,N_6733);
or U7344 (N_7344,N_6534,N_6535);
nor U7345 (N_7345,N_6475,N_6976);
nand U7346 (N_7346,N_6615,N_7103);
nand U7347 (N_7347,N_6594,N_7173);
nand U7348 (N_7348,N_7009,N_6754);
and U7349 (N_7349,N_6630,N_6812);
or U7350 (N_7350,N_7022,N_6454);
nor U7351 (N_7351,N_7124,N_6822);
nor U7352 (N_7352,N_6856,N_6773);
or U7353 (N_7353,N_7166,N_7087);
or U7354 (N_7354,N_7194,N_7149);
and U7355 (N_7355,N_7089,N_7072);
or U7356 (N_7356,N_6592,N_7075);
nor U7357 (N_7357,N_7154,N_6691);
nand U7358 (N_7358,N_7178,N_7081);
nor U7359 (N_7359,N_6596,N_6796);
nand U7360 (N_7360,N_7140,N_6904);
nor U7361 (N_7361,N_7125,N_6749);
and U7362 (N_7362,N_6785,N_6418);
or U7363 (N_7363,N_6880,N_6717);
nor U7364 (N_7364,N_6404,N_6597);
nor U7365 (N_7365,N_7083,N_7101);
nor U7366 (N_7366,N_7193,N_6571);
xor U7367 (N_7367,N_7186,N_6818);
and U7368 (N_7368,N_6503,N_6710);
nor U7369 (N_7369,N_6659,N_6845);
nor U7370 (N_7370,N_7129,N_6718);
and U7371 (N_7371,N_7069,N_7192);
or U7372 (N_7372,N_6719,N_6981);
xor U7373 (N_7373,N_6521,N_7007);
or U7374 (N_7374,N_6857,N_6763);
and U7375 (N_7375,N_7199,N_7099);
nand U7376 (N_7376,N_7148,N_7105);
xor U7377 (N_7377,N_6730,N_7033);
xor U7378 (N_7378,N_7136,N_6557);
or U7379 (N_7379,N_6623,N_6969);
and U7380 (N_7380,N_7018,N_6523);
and U7381 (N_7381,N_6526,N_6573);
and U7382 (N_7382,N_6520,N_6580);
nor U7383 (N_7383,N_6793,N_6980);
nand U7384 (N_7384,N_6455,N_6440);
nand U7385 (N_7385,N_7104,N_6761);
or U7386 (N_7386,N_6450,N_7002);
nand U7387 (N_7387,N_6874,N_6726);
nand U7388 (N_7388,N_7023,N_6671);
xor U7389 (N_7389,N_6963,N_7167);
nor U7390 (N_7390,N_6498,N_6729);
nand U7391 (N_7391,N_6825,N_6588);
xnor U7392 (N_7392,N_6601,N_7119);
xnor U7393 (N_7393,N_7001,N_6544);
or U7394 (N_7394,N_6795,N_6590);
nand U7395 (N_7395,N_6894,N_7039);
xor U7396 (N_7396,N_6949,N_7053);
xnor U7397 (N_7397,N_6747,N_6919);
xnor U7398 (N_7398,N_6873,N_6907);
nor U7399 (N_7399,N_7071,N_6807);
or U7400 (N_7400,N_6902,N_7106);
nor U7401 (N_7401,N_6918,N_6645);
nand U7402 (N_7402,N_7133,N_7052);
xnor U7403 (N_7403,N_6651,N_6725);
and U7404 (N_7404,N_6467,N_7059);
xor U7405 (N_7405,N_7055,N_6838);
and U7406 (N_7406,N_6473,N_6504);
nor U7407 (N_7407,N_6660,N_6443);
nand U7408 (N_7408,N_6867,N_6408);
and U7409 (N_7409,N_6734,N_7177);
and U7410 (N_7410,N_6667,N_6612);
or U7411 (N_7411,N_6770,N_6499);
and U7412 (N_7412,N_7042,N_7068);
or U7413 (N_7413,N_6669,N_6852);
and U7414 (N_7414,N_6897,N_6698);
or U7415 (N_7415,N_6619,N_6908);
nand U7416 (N_7416,N_6545,N_7062);
xor U7417 (N_7417,N_6741,N_6600);
nor U7418 (N_7418,N_6937,N_7026);
or U7419 (N_7419,N_6810,N_6549);
nand U7420 (N_7420,N_7131,N_6767);
xor U7421 (N_7421,N_6427,N_7144);
and U7422 (N_7422,N_6666,N_7115);
or U7423 (N_7423,N_6559,N_6738);
xnor U7424 (N_7424,N_6799,N_6677);
nand U7425 (N_7425,N_6444,N_6425);
xor U7426 (N_7426,N_6536,N_7011);
and U7427 (N_7427,N_6928,N_6990);
nor U7428 (N_7428,N_7120,N_6598);
and U7429 (N_7429,N_6620,N_6511);
or U7430 (N_7430,N_6716,N_7116);
nor U7431 (N_7431,N_6832,N_6505);
nor U7432 (N_7432,N_6402,N_7012);
xnor U7433 (N_7433,N_6891,N_6654);
or U7434 (N_7434,N_6844,N_6689);
nor U7435 (N_7435,N_6842,N_7138);
nor U7436 (N_7436,N_7112,N_6668);
xnor U7437 (N_7437,N_6960,N_7046);
xnor U7438 (N_7438,N_6745,N_7048);
nand U7439 (N_7439,N_7184,N_6607);
xor U7440 (N_7440,N_6715,N_6816);
and U7441 (N_7441,N_6532,N_7156);
nand U7442 (N_7442,N_7146,N_6403);
and U7443 (N_7443,N_6929,N_6986);
or U7444 (N_7444,N_6912,N_6605);
nand U7445 (N_7445,N_7152,N_7029);
nand U7446 (N_7446,N_6564,N_6472);
and U7447 (N_7447,N_6546,N_6826);
or U7448 (N_7448,N_6649,N_6942);
nand U7449 (N_7449,N_6759,N_6640);
and U7450 (N_7450,N_7163,N_6700);
or U7451 (N_7451,N_6537,N_7041);
and U7452 (N_7452,N_6648,N_7147);
or U7453 (N_7453,N_6614,N_6702);
or U7454 (N_7454,N_6547,N_6533);
xnor U7455 (N_7455,N_6992,N_6898);
nor U7456 (N_7456,N_6673,N_6643);
nand U7457 (N_7457,N_6984,N_6778);
and U7458 (N_7458,N_7004,N_6578);
or U7459 (N_7459,N_7051,N_6703);
and U7460 (N_7460,N_6562,N_6490);
and U7461 (N_7461,N_6468,N_6676);
nor U7462 (N_7462,N_7175,N_6800);
nand U7463 (N_7463,N_6664,N_6968);
or U7464 (N_7464,N_6903,N_6566);
nand U7465 (N_7465,N_6638,N_6883);
nor U7466 (N_7466,N_6480,N_6828);
nand U7467 (N_7467,N_6487,N_6541);
and U7468 (N_7468,N_6550,N_6540);
nand U7469 (N_7469,N_6627,N_6948);
or U7470 (N_7470,N_6709,N_6959);
and U7471 (N_7471,N_7076,N_6479);
or U7472 (N_7472,N_6921,N_7031);
nor U7473 (N_7473,N_6589,N_6693);
xnor U7474 (N_7474,N_7082,N_7128);
xor U7475 (N_7475,N_6864,N_6781);
or U7476 (N_7476,N_7158,N_6771);
and U7477 (N_7477,N_6953,N_6519);
or U7478 (N_7478,N_6426,N_6722);
xor U7479 (N_7479,N_6602,N_7092);
xor U7480 (N_7480,N_6815,N_6925);
or U7481 (N_7481,N_6430,N_6493);
and U7482 (N_7482,N_7151,N_6809);
and U7483 (N_7483,N_7179,N_6708);
or U7484 (N_7484,N_6750,N_6441);
nor U7485 (N_7485,N_6952,N_6637);
xnor U7486 (N_7486,N_7181,N_6855);
nor U7487 (N_7487,N_6538,N_7005);
nor U7488 (N_7488,N_6958,N_7080);
and U7489 (N_7489,N_7093,N_6911);
or U7490 (N_7490,N_6755,N_7188);
nor U7491 (N_7491,N_6438,N_6794);
nor U7492 (N_7492,N_6743,N_6711);
nor U7493 (N_7493,N_6991,N_6872);
nor U7494 (N_7494,N_7054,N_7088);
xnor U7495 (N_7495,N_6920,N_6435);
xnor U7496 (N_7496,N_7183,N_6802);
and U7497 (N_7497,N_7135,N_6945);
xnor U7498 (N_7498,N_6850,N_7164);
xor U7499 (N_7499,N_6765,N_6512);
nor U7500 (N_7500,N_6786,N_6846);
xnor U7501 (N_7501,N_6584,N_6931);
nand U7502 (N_7502,N_6662,N_7143);
xnor U7503 (N_7503,N_7079,N_6641);
nor U7504 (N_7504,N_6805,N_6890);
or U7505 (N_7505,N_6415,N_6634);
xor U7506 (N_7506,N_6806,N_6633);
nand U7507 (N_7507,N_6843,N_6714);
and U7508 (N_7508,N_6424,N_6449);
nor U7509 (N_7509,N_7141,N_6831);
nand U7510 (N_7510,N_6861,N_6433);
nor U7511 (N_7511,N_6962,N_6721);
nor U7512 (N_7512,N_6492,N_6657);
nand U7513 (N_7513,N_6923,N_6646);
or U7514 (N_7514,N_6469,N_6497);
or U7515 (N_7515,N_6712,N_7127);
nor U7516 (N_7516,N_7137,N_6470);
or U7517 (N_7517,N_6661,N_6877);
nand U7518 (N_7518,N_6583,N_6817);
xor U7519 (N_7519,N_6434,N_6824);
nor U7520 (N_7520,N_6955,N_6849);
and U7521 (N_7521,N_6515,N_6417);
nor U7522 (N_7522,N_6732,N_6879);
nor U7523 (N_7523,N_6461,N_7168);
nand U7524 (N_7524,N_6720,N_6474);
nand U7525 (N_7525,N_7063,N_6853);
nor U7526 (N_7526,N_7006,N_7000);
and U7527 (N_7527,N_6999,N_6938);
or U7528 (N_7528,N_6936,N_6653);
and U7529 (N_7529,N_6705,N_7045);
and U7530 (N_7530,N_6610,N_7189);
nor U7531 (N_7531,N_6551,N_7190);
xnor U7532 (N_7532,N_6906,N_6527);
or U7533 (N_7533,N_6696,N_6608);
xnor U7534 (N_7534,N_6570,N_7195);
and U7535 (N_7535,N_6423,N_6685);
nor U7536 (N_7536,N_6790,N_6585);
xnor U7537 (N_7537,N_7061,N_6866);
nor U7538 (N_7538,N_6568,N_6941);
or U7539 (N_7539,N_6914,N_6869);
or U7540 (N_7540,N_6965,N_6811);
xnor U7541 (N_7541,N_6419,N_6901);
xnor U7542 (N_7542,N_7003,N_6932);
nand U7543 (N_7543,N_6801,N_6446);
nor U7544 (N_7544,N_6787,N_6933);
and U7545 (N_7545,N_6884,N_7198);
nand U7546 (N_7546,N_6428,N_6926);
and U7547 (N_7547,N_7044,N_6996);
or U7548 (N_7548,N_6859,N_6611);
nand U7549 (N_7549,N_6639,N_6439);
nand U7550 (N_7550,N_6752,N_6684);
or U7551 (N_7551,N_6988,N_6878);
nand U7552 (N_7552,N_6971,N_6595);
or U7553 (N_7553,N_6994,N_6893);
xnor U7554 (N_7554,N_6808,N_6581);
or U7555 (N_7555,N_6739,N_6753);
and U7556 (N_7556,N_6539,N_6650);
or U7557 (N_7557,N_6731,N_7084);
xnor U7558 (N_7558,N_7171,N_6774);
nand U7559 (N_7559,N_6658,N_7095);
nor U7560 (N_7560,N_6647,N_7122);
xor U7561 (N_7561,N_6542,N_6464);
and U7562 (N_7562,N_6453,N_6964);
and U7563 (N_7563,N_6766,N_6463);
xnor U7564 (N_7564,N_7196,N_6989);
nand U7565 (N_7565,N_7056,N_6674);
nor U7566 (N_7566,N_7100,N_6680);
or U7567 (N_7567,N_6528,N_6613);
and U7568 (N_7568,N_6769,N_6978);
nor U7569 (N_7569,N_6561,N_7030);
xnor U7570 (N_7570,N_6459,N_7014);
and U7571 (N_7571,N_6478,N_6724);
nor U7572 (N_7572,N_6411,N_6837);
nor U7573 (N_7573,N_7185,N_6524);
or U7574 (N_7574,N_6776,N_6813);
and U7575 (N_7575,N_6482,N_6483);
and U7576 (N_7576,N_6407,N_7153);
nor U7577 (N_7577,N_6558,N_6760);
xnor U7578 (N_7578,N_7010,N_6940);
nor U7579 (N_7579,N_6985,N_6481);
nand U7580 (N_7580,N_7034,N_6421);
nand U7581 (N_7581,N_6998,N_6409);
or U7582 (N_7582,N_6944,N_6804);
xor U7583 (N_7583,N_6682,N_6514);
or U7584 (N_7584,N_6606,N_7109);
and U7585 (N_7585,N_7197,N_6501);
xnor U7586 (N_7586,N_6961,N_6871);
or U7587 (N_7587,N_7176,N_6860);
nor U7588 (N_7588,N_6695,N_6574);
and U7589 (N_7589,N_6462,N_6881);
and U7590 (N_7590,N_7050,N_7187);
nor U7591 (N_7591,N_6975,N_6798);
or U7592 (N_7592,N_6576,N_6618);
xnor U7593 (N_7593,N_7139,N_6652);
nand U7594 (N_7594,N_6543,N_6821);
or U7595 (N_7595,N_6723,N_6889);
or U7596 (N_7596,N_6757,N_6447);
and U7597 (N_7597,N_6917,N_7057);
or U7598 (N_7598,N_7160,N_6713);
and U7599 (N_7599,N_6679,N_6560);
xor U7600 (N_7600,N_7146,N_7006);
xnor U7601 (N_7601,N_7042,N_6475);
nor U7602 (N_7602,N_7179,N_6543);
and U7603 (N_7603,N_6409,N_7089);
xor U7604 (N_7604,N_7199,N_6917);
nand U7605 (N_7605,N_6504,N_7054);
and U7606 (N_7606,N_7022,N_6626);
nor U7607 (N_7607,N_6740,N_7130);
nand U7608 (N_7608,N_6754,N_6647);
xnor U7609 (N_7609,N_6815,N_6476);
nor U7610 (N_7610,N_7178,N_6508);
or U7611 (N_7611,N_6623,N_6583);
or U7612 (N_7612,N_6994,N_6831);
and U7613 (N_7613,N_7153,N_6783);
or U7614 (N_7614,N_6941,N_6470);
nand U7615 (N_7615,N_6464,N_6475);
nor U7616 (N_7616,N_6631,N_6620);
nor U7617 (N_7617,N_6540,N_7047);
or U7618 (N_7618,N_7094,N_6522);
nand U7619 (N_7619,N_6897,N_7164);
nor U7620 (N_7620,N_6906,N_6636);
or U7621 (N_7621,N_6781,N_6569);
and U7622 (N_7622,N_7166,N_6597);
and U7623 (N_7623,N_6616,N_6638);
xnor U7624 (N_7624,N_6630,N_6828);
nor U7625 (N_7625,N_6552,N_6729);
or U7626 (N_7626,N_6466,N_6446);
nor U7627 (N_7627,N_7141,N_6599);
nand U7628 (N_7628,N_6514,N_7013);
or U7629 (N_7629,N_6959,N_7149);
or U7630 (N_7630,N_6786,N_7190);
xnor U7631 (N_7631,N_7167,N_7099);
and U7632 (N_7632,N_6689,N_6673);
xnor U7633 (N_7633,N_6473,N_6933);
or U7634 (N_7634,N_6539,N_7062);
nor U7635 (N_7635,N_7050,N_6999);
nor U7636 (N_7636,N_7045,N_6537);
xnor U7637 (N_7637,N_6930,N_6402);
xor U7638 (N_7638,N_6970,N_6861);
or U7639 (N_7639,N_7003,N_6844);
and U7640 (N_7640,N_6603,N_6790);
nor U7641 (N_7641,N_6844,N_7050);
nor U7642 (N_7642,N_6728,N_6994);
xnor U7643 (N_7643,N_6788,N_7040);
or U7644 (N_7644,N_7195,N_6627);
nand U7645 (N_7645,N_6625,N_7151);
nand U7646 (N_7646,N_6919,N_6600);
and U7647 (N_7647,N_6869,N_6538);
xnor U7648 (N_7648,N_7198,N_6575);
or U7649 (N_7649,N_6484,N_6916);
xor U7650 (N_7650,N_6881,N_7062);
nor U7651 (N_7651,N_6860,N_7006);
xnor U7652 (N_7652,N_7074,N_6689);
nor U7653 (N_7653,N_6637,N_6572);
nand U7654 (N_7654,N_6634,N_7146);
or U7655 (N_7655,N_6530,N_7045);
nand U7656 (N_7656,N_6421,N_7040);
nor U7657 (N_7657,N_6679,N_7065);
nor U7658 (N_7658,N_6633,N_7040);
nand U7659 (N_7659,N_6505,N_6956);
nor U7660 (N_7660,N_7000,N_6714);
xor U7661 (N_7661,N_6974,N_6570);
nand U7662 (N_7662,N_6913,N_7197);
or U7663 (N_7663,N_6654,N_6698);
and U7664 (N_7664,N_6611,N_6899);
nand U7665 (N_7665,N_6890,N_6957);
and U7666 (N_7666,N_6635,N_7090);
or U7667 (N_7667,N_6466,N_7003);
xnor U7668 (N_7668,N_6890,N_6450);
and U7669 (N_7669,N_6850,N_6430);
xor U7670 (N_7670,N_6755,N_7156);
or U7671 (N_7671,N_6972,N_6773);
nand U7672 (N_7672,N_6853,N_6725);
or U7673 (N_7673,N_6800,N_6714);
or U7674 (N_7674,N_6445,N_6540);
and U7675 (N_7675,N_6461,N_6752);
or U7676 (N_7676,N_6941,N_6596);
or U7677 (N_7677,N_6434,N_6613);
nor U7678 (N_7678,N_7137,N_6935);
and U7679 (N_7679,N_6990,N_7126);
nor U7680 (N_7680,N_6711,N_6548);
nand U7681 (N_7681,N_6765,N_6862);
nor U7682 (N_7682,N_6471,N_7041);
xnor U7683 (N_7683,N_7154,N_6928);
xnor U7684 (N_7684,N_7193,N_6720);
nor U7685 (N_7685,N_6799,N_6961);
nor U7686 (N_7686,N_6444,N_7057);
xor U7687 (N_7687,N_6903,N_7109);
nand U7688 (N_7688,N_6689,N_7107);
xnor U7689 (N_7689,N_6430,N_6406);
xor U7690 (N_7690,N_6414,N_6737);
or U7691 (N_7691,N_6916,N_6539);
and U7692 (N_7692,N_6956,N_7037);
and U7693 (N_7693,N_6904,N_6467);
xor U7694 (N_7694,N_6774,N_6575);
or U7695 (N_7695,N_7116,N_7046);
nor U7696 (N_7696,N_6495,N_6467);
nand U7697 (N_7697,N_6824,N_6464);
or U7698 (N_7698,N_6798,N_6847);
nand U7699 (N_7699,N_6630,N_6854);
nand U7700 (N_7700,N_6718,N_7186);
xnor U7701 (N_7701,N_7170,N_7188);
and U7702 (N_7702,N_6956,N_6845);
or U7703 (N_7703,N_6757,N_7124);
and U7704 (N_7704,N_6480,N_6910);
nor U7705 (N_7705,N_7175,N_7107);
xor U7706 (N_7706,N_6964,N_6703);
nand U7707 (N_7707,N_6436,N_7120);
nand U7708 (N_7708,N_6442,N_7161);
or U7709 (N_7709,N_6739,N_6433);
and U7710 (N_7710,N_6912,N_6838);
or U7711 (N_7711,N_7026,N_6478);
nor U7712 (N_7712,N_6885,N_6658);
or U7713 (N_7713,N_7181,N_7190);
and U7714 (N_7714,N_6586,N_7025);
nor U7715 (N_7715,N_6618,N_6731);
xnor U7716 (N_7716,N_6592,N_6686);
nor U7717 (N_7717,N_6923,N_6571);
nand U7718 (N_7718,N_6839,N_7160);
xnor U7719 (N_7719,N_6688,N_6708);
and U7720 (N_7720,N_6638,N_7114);
and U7721 (N_7721,N_6720,N_6781);
and U7722 (N_7722,N_6708,N_7008);
and U7723 (N_7723,N_6711,N_6896);
and U7724 (N_7724,N_6730,N_6575);
xnor U7725 (N_7725,N_6827,N_6701);
nand U7726 (N_7726,N_6628,N_6458);
nand U7727 (N_7727,N_6646,N_7005);
nand U7728 (N_7728,N_7119,N_6871);
or U7729 (N_7729,N_6681,N_6785);
nand U7730 (N_7730,N_6880,N_6577);
xor U7731 (N_7731,N_6647,N_6636);
nor U7732 (N_7732,N_6655,N_7028);
nor U7733 (N_7733,N_7178,N_6576);
nand U7734 (N_7734,N_6622,N_6541);
or U7735 (N_7735,N_6413,N_6985);
nand U7736 (N_7736,N_7001,N_6761);
nand U7737 (N_7737,N_6997,N_6538);
and U7738 (N_7738,N_6466,N_6798);
or U7739 (N_7739,N_7196,N_6837);
nand U7740 (N_7740,N_7055,N_6820);
or U7741 (N_7741,N_7013,N_6570);
or U7742 (N_7742,N_6661,N_6531);
nand U7743 (N_7743,N_6425,N_6616);
nor U7744 (N_7744,N_6612,N_6546);
or U7745 (N_7745,N_7157,N_6903);
nand U7746 (N_7746,N_7116,N_6433);
nand U7747 (N_7747,N_6767,N_7048);
nand U7748 (N_7748,N_6472,N_7134);
and U7749 (N_7749,N_6602,N_7111);
nand U7750 (N_7750,N_6971,N_6789);
nand U7751 (N_7751,N_6526,N_6813);
nand U7752 (N_7752,N_6603,N_7146);
or U7753 (N_7753,N_6937,N_6437);
nand U7754 (N_7754,N_6472,N_6887);
nand U7755 (N_7755,N_7168,N_6907);
and U7756 (N_7756,N_7196,N_6706);
nand U7757 (N_7757,N_6577,N_7125);
nand U7758 (N_7758,N_6659,N_7047);
nand U7759 (N_7759,N_6766,N_6832);
nor U7760 (N_7760,N_6612,N_6701);
or U7761 (N_7761,N_6512,N_6818);
nand U7762 (N_7762,N_6775,N_6668);
xor U7763 (N_7763,N_6549,N_7184);
nor U7764 (N_7764,N_6405,N_6599);
or U7765 (N_7765,N_6461,N_6660);
nor U7766 (N_7766,N_6645,N_7107);
nor U7767 (N_7767,N_7113,N_6616);
or U7768 (N_7768,N_6655,N_6516);
nand U7769 (N_7769,N_6781,N_6442);
and U7770 (N_7770,N_6977,N_7128);
nor U7771 (N_7771,N_6814,N_7016);
nor U7772 (N_7772,N_7076,N_6691);
xor U7773 (N_7773,N_7090,N_7028);
nand U7774 (N_7774,N_7009,N_6813);
nor U7775 (N_7775,N_6767,N_6621);
or U7776 (N_7776,N_6626,N_7180);
nand U7777 (N_7777,N_6520,N_6427);
and U7778 (N_7778,N_6790,N_6917);
and U7779 (N_7779,N_6517,N_6958);
or U7780 (N_7780,N_6655,N_6745);
xor U7781 (N_7781,N_6490,N_6598);
nor U7782 (N_7782,N_6518,N_7117);
or U7783 (N_7783,N_7021,N_6651);
nor U7784 (N_7784,N_6549,N_6720);
and U7785 (N_7785,N_7161,N_6502);
nand U7786 (N_7786,N_6823,N_6895);
or U7787 (N_7787,N_6520,N_6917);
and U7788 (N_7788,N_7090,N_7082);
xor U7789 (N_7789,N_6658,N_6637);
and U7790 (N_7790,N_6666,N_6404);
xnor U7791 (N_7791,N_6444,N_6794);
nor U7792 (N_7792,N_6677,N_6544);
xnor U7793 (N_7793,N_6640,N_7001);
and U7794 (N_7794,N_6899,N_6745);
nand U7795 (N_7795,N_6787,N_7129);
and U7796 (N_7796,N_6860,N_6508);
nor U7797 (N_7797,N_6709,N_7135);
nand U7798 (N_7798,N_7079,N_6669);
nand U7799 (N_7799,N_6554,N_6854);
nor U7800 (N_7800,N_6711,N_6502);
nand U7801 (N_7801,N_6403,N_6537);
or U7802 (N_7802,N_6456,N_7054);
nor U7803 (N_7803,N_7130,N_6768);
or U7804 (N_7804,N_6653,N_7029);
nand U7805 (N_7805,N_6939,N_6677);
nor U7806 (N_7806,N_6503,N_6939);
and U7807 (N_7807,N_7097,N_6929);
nand U7808 (N_7808,N_7015,N_7163);
or U7809 (N_7809,N_6835,N_7125);
xnor U7810 (N_7810,N_6406,N_6505);
and U7811 (N_7811,N_6820,N_6850);
nor U7812 (N_7812,N_6769,N_6629);
and U7813 (N_7813,N_6862,N_7142);
xnor U7814 (N_7814,N_6668,N_6511);
nor U7815 (N_7815,N_6413,N_6603);
and U7816 (N_7816,N_6709,N_6970);
or U7817 (N_7817,N_6712,N_7058);
nor U7818 (N_7818,N_6546,N_6464);
and U7819 (N_7819,N_6746,N_6804);
or U7820 (N_7820,N_6705,N_6620);
or U7821 (N_7821,N_6711,N_6817);
xnor U7822 (N_7822,N_6881,N_6403);
nand U7823 (N_7823,N_6861,N_6512);
nand U7824 (N_7824,N_7147,N_6908);
and U7825 (N_7825,N_6619,N_6589);
nor U7826 (N_7826,N_6990,N_7009);
and U7827 (N_7827,N_6417,N_6976);
and U7828 (N_7828,N_6940,N_7039);
xnor U7829 (N_7829,N_7166,N_7172);
or U7830 (N_7830,N_7161,N_6800);
or U7831 (N_7831,N_6852,N_6766);
nand U7832 (N_7832,N_6843,N_6623);
or U7833 (N_7833,N_6769,N_6765);
and U7834 (N_7834,N_7000,N_6600);
xor U7835 (N_7835,N_6671,N_7117);
xor U7836 (N_7836,N_6812,N_7029);
and U7837 (N_7837,N_6706,N_6715);
and U7838 (N_7838,N_6413,N_6533);
and U7839 (N_7839,N_7055,N_6419);
xnor U7840 (N_7840,N_6523,N_6417);
xnor U7841 (N_7841,N_6546,N_7175);
and U7842 (N_7842,N_7009,N_6934);
xnor U7843 (N_7843,N_6469,N_6896);
or U7844 (N_7844,N_6625,N_6453);
xor U7845 (N_7845,N_6471,N_7043);
nand U7846 (N_7846,N_6792,N_7050);
nor U7847 (N_7847,N_6703,N_6702);
nor U7848 (N_7848,N_6656,N_6991);
xor U7849 (N_7849,N_6435,N_6508);
or U7850 (N_7850,N_7147,N_6578);
nor U7851 (N_7851,N_6672,N_6540);
nor U7852 (N_7852,N_7147,N_7031);
xnor U7853 (N_7853,N_6641,N_6914);
or U7854 (N_7854,N_6812,N_7149);
nor U7855 (N_7855,N_6858,N_6899);
nor U7856 (N_7856,N_6603,N_6906);
and U7857 (N_7857,N_6744,N_6782);
nand U7858 (N_7858,N_6769,N_6755);
xor U7859 (N_7859,N_6453,N_6950);
xor U7860 (N_7860,N_6586,N_6882);
nor U7861 (N_7861,N_6531,N_6454);
or U7862 (N_7862,N_6995,N_6996);
nand U7863 (N_7863,N_6629,N_6858);
xor U7864 (N_7864,N_6554,N_7185);
nor U7865 (N_7865,N_7027,N_6902);
nor U7866 (N_7866,N_7127,N_6960);
or U7867 (N_7867,N_7089,N_6555);
xnor U7868 (N_7868,N_6901,N_7188);
and U7869 (N_7869,N_6751,N_6736);
nor U7870 (N_7870,N_6613,N_7017);
nand U7871 (N_7871,N_6964,N_6852);
and U7872 (N_7872,N_6435,N_6640);
or U7873 (N_7873,N_6860,N_7057);
and U7874 (N_7874,N_6835,N_7067);
and U7875 (N_7875,N_6910,N_6890);
nand U7876 (N_7876,N_6414,N_7158);
or U7877 (N_7877,N_6931,N_6529);
nor U7878 (N_7878,N_7191,N_6650);
nand U7879 (N_7879,N_6938,N_7153);
or U7880 (N_7880,N_7014,N_6741);
nand U7881 (N_7881,N_6587,N_7076);
and U7882 (N_7882,N_6994,N_6946);
xor U7883 (N_7883,N_6477,N_7153);
xnor U7884 (N_7884,N_6827,N_6978);
and U7885 (N_7885,N_6803,N_6884);
xor U7886 (N_7886,N_6763,N_6898);
or U7887 (N_7887,N_6707,N_7055);
and U7888 (N_7888,N_6686,N_6926);
nor U7889 (N_7889,N_6837,N_7084);
or U7890 (N_7890,N_6738,N_6573);
nor U7891 (N_7891,N_6580,N_6747);
or U7892 (N_7892,N_6843,N_6546);
xor U7893 (N_7893,N_6791,N_6508);
and U7894 (N_7894,N_6682,N_6904);
nand U7895 (N_7895,N_6698,N_6535);
nor U7896 (N_7896,N_6944,N_6659);
xnor U7897 (N_7897,N_6776,N_6755);
or U7898 (N_7898,N_6612,N_6924);
xor U7899 (N_7899,N_6467,N_6526);
or U7900 (N_7900,N_7015,N_6546);
nand U7901 (N_7901,N_6774,N_6425);
nor U7902 (N_7902,N_6568,N_6747);
xnor U7903 (N_7903,N_6925,N_6478);
or U7904 (N_7904,N_6443,N_6656);
or U7905 (N_7905,N_6936,N_6974);
or U7906 (N_7906,N_7088,N_6416);
nand U7907 (N_7907,N_6596,N_6988);
nand U7908 (N_7908,N_6886,N_6708);
nand U7909 (N_7909,N_6778,N_6854);
nand U7910 (N_7910,N_7070,N_7000);
and U7911 (N_7911,N_6849,N_6991);
and U7912 (N_7912,N_6624,N_6647);
xor U7913 (N_7913,N_6500,N_6455);
or U7914 (N_7914,N_6962,N_7062);
xnor U7915 (N_7915,N_6480,N_6835);
and U7916 (N_7916,N_6984,N_6484);
xor U7917 (N_7917,N_7199,N_6629);
nor U7918 (N_7918,N_6402,N_6699);
xor U7919 (N_7919,N_6489,N_6826);
and U7920 (N_7920,N_6891,N_6992);
or U7921 (N_7921,N_6939,N_7038);
nor U7922 (N_7922,N_7067,N_6799);
or U7923 (N_7923,N_6888,N_6936);
and U7924 (N_7924,N_6418,N_7178);
nor U7925 (N_7925,N_6419,N_7032);
nand U7926 (N_7926,N_6596,N_6825);
nor U7927 (N_7927,N_6934,N_7004);
xor U7928 (N_7928,N_7058,N_7087);
nor U7929 (N_7929,N_6907,N_7051);
nor U7930 (N_7930,N_6557,N_6625);
nor U7931 (N_7931,N_7193,N_6464);
xor U7932 (N_7932,N_6783,N_7039);
nand U7933 (N_7933,N_6740,N_6445);
nor U7934 (N_7934,N_6631,N_6589);
nor U7935 (N_7935,N_6884,N_6779);
nor U7936 (N_7936,N_6961,N_6435);
nor U7937 (N_7937,N_6700,N_6951);
nor U7938 (N_7938,N_7095,N_6640);
and U7939 (N_7939,N_6777,N_6736);
nand U7940 (N_7940,N_6557,N_6721);
and U7941 (N_7941,N_7146,N_7120);
nor U7942 (N_7942,N_6605,N_6658);
and U7943 (N_7943,N_6636,N_6970);
xnor U7944 (N_7944,N_6770,N_6909);
and U7945 (N_7945,N_6820,N_6621);
nor U7946 (N_7946,N_6555,N_6834);
nor U7947 (N_7947,N_6919,N_7105);
xor U7948 (N_7948,N_6748,N_6652);
nand U7949 (N_7949,N_6615,N_6472);
nand U7950 (N_7950,N_6447,N_6969);
and U7951 (N_7951,N_6963,N_6996);
nor U7952 (N_7952,N_7011,N_6849);
and U7953 (N_7953,N_7139,N_6859);
nand U7954 (N_7954,N_6915,N_6956);
nor U7955 (N_7955,N_6492,N_6772);
nor U7956 (N_7956,N_7039,N_7131);
nor U7957 (N_7957,N_6545,N_6984);
nor U7958 (N_7958,N_7032,N_6537);
and U7959 (N_7959,N_7174,N_7001);
or U7960 (N_7960,N_7011,N_7139);
or U7961 (N_7961,N_6640,N_6439);
or U7962 (N_7962,N_6720,N_7005);
and U7963 (N_7963,N_6674,N_7026);
nand U7964 (N_7964,N_6405,N_6579);
xor U7965 (N_7965,N_6831,N_6640);
xnor U7966 (N_7966,N_7074,N_6652);
nand U7967 (N_7967,N_7013,N_7008);
or U7968 (N_7968,N_6882,N_6672);
or U7969 (N_7969,N_6858,N_7000);
xnor U7970 (N_7970,N_6555,N_6541);
xnor U7971 (N_7971,N_6553,N_6795);
xnor U7972 (N_7972,N_6447,N_6780);
nor U7973 (N_7973,N_6962,N_7155);
or U7974 (N_7974,N_6876,N_6941);
nand U7975 (N_7975,N_6437,N_6901);
nand U7976 (N_7976,N_6430,N_6550);
nand U7977 (N_7977,N_6583,N_6849);
xor U7978 (N_7978,N_6400,N_7185);
nor U7979 (N_7979,N_7189,N_6931);
nand U7980 (N_7980,N_6617,N_6587);
xnor U7981 (N_7981,N_7032,N_7149);
or U7982 (N_7982,N_6686,N_7128);
xor U7983 (N_7983,N_6874,N_6590);
and U7984 (N_7984,N_6706,N_6990);
and U7985 (N_7985,N_6489,N_6436);
and U7986 (N_7986,N_6561,N_6766);
xnor U7987 (N_7987,N_6873,N_6851);
nor U7988 (N_7988,N_6489,N_7003);
nand U7989 (N_7989,N_6533,N_6480);
xnor U7990 (N_7990,N_7006,N_6917);
xnor U7991 (N_7991,N_6905,N_7158);
nand U7992 (N_7992,N_6571,N_6894);
and U7993 (N_7993,N_6859,N_7131);
nand U7994 (N_7994,N_7075,N_6608);
and U7995 (N_7995,N_6681,N_6818);
and U7996 (N_7996,N_6452,N_7144);
xor U7997 (N_7997,N_7172,N_6920);
nand U7998 (N_7998,N_6540,N_6440);
and U7999 (N_7999,N_6480,N_6948);
nor U8000 (N_8000,N_7485,N_7237);
nor U8001 (N_8001,N_7988,N_7889);
or U8002 (N_8002,N_7217,N_7967);
or U8003 (N_8003,N_7433,N_7783);
xor U8004 (N_8004,N_7868,N_7525);
xor U8005 (N_8005,N_7708,N_7371);
xor U8006 (N_8006,N_7910,N_7798);
xor U8007 (N_8007,N_7509,N_7899);
and U8008 (N_8008,N_7649,N_7903);
nand U8009 (N_8009,N_7363,N_7806);
xnor U8010 (N_8010,N_7373,N_7907);
or U8011 (N_8011,N_7735,N_7892);
and U8012 (N_8012,N_7595,N_7259);
and U8013 (N_8013,N_7420,N_7332);
or U8014 (N_8014,N_7353,N_7906);
xor U8015 (N_8015,N_7502,N_7517);
nand U8016 (N_8016,N_7387,N_7844);
xor U8017 (N_8017,N_7503,N_7667);
nor U8018 (N_8018,N_7864,N_7293);
nor U8019 (N_8019,N_7397,N_7648);
and U8020 (N_8020,N_7820,N_7955);
or U8021 (N_8021,N_7348,N_7867);
nor U8022 (N_8022,N_7638,N_7429);
xnor U8023 (N_8023,N_7566,N_7291);
and U8024 (N_8024,N_7847,N_7247);
nand U8025 (N_8025,N_7966,N_7728);
xnor U8026 (N_8026,N_7315,N_7534);
and U8027 (N_8027,N_7997,N_7584);
or U8028 (N_8028,N_7290,N_7355);
and U8029 (N_8029,N_7942,N_7432);
xor U8030 (N_8030,N_7937,N_7719);
xor U8031 (N_8031,N_7886,N_7632);
and U8032 (N_8032,N_7880,N_7575);
or U8033 (N_8033,N_7925,N_7861);
nand U8034 (N_8034,N_7490,N_7850);
xor U8035 (N_8035,N_7469,N_7318);
nor U8036 (N_8036,N_7896,N_7202);
or U8037 (N_8037,N_7224,N_7830);
nor U8038 (N_8038,N_7483,N_7243);
nand U8039 (N_8039,N_7692,N_7805);
nor U8040 (N_8040,N_7709,N_7857);
and U8041 (N_8041,N_7687,N_7672);
xor U8042 (N_8042,N_7992,N_7265);
or U8043 (N_8043,N_7730,N_7633);
or U8044 (N_8044,N_7496,N_7834);
xor U8045 (N_8045,N_7902,N_7470);
or U8046 (N_8046,N_7507,N_7439);
xor U8047 (N_8047,N_7791,N_7826);
or U8048 (N_8048,N_7929,N_7938);
nand U8049 (N_8049,N_7516,N_7918);
xor U8050 (N_8050,N_7253,N_7334);
and U8051 (N_8051,N_7900,N_7908);
nor U8052 (N_8052,N_7852,N_7924);
xnor U8053 (N_8053,N_7512,N_7477);
and U8054 (N_8054,N_7990,N_7365);
and U8055 (N_8055,N_7456,N_7588);
or U8056 (N_8056,N_7987,N_7273);
and U8057 (N_8057,N_7403,N_7751);
or U8058 (N_8058,N_7645,N_7488);
xnor U8059 (N_8059,N_7859,N_7207);
nand U8060 (N_8060,N_7473,N_7522);
or U8061 (N_8061,N_7214,N_7787);
xor U8062 (N_8062,N_7995,N_7999);
nor U8063 (N_8063,N_7994,N_7402);
nor U8064 (N_8064,N_7206,N_7275);
xor U8065 (N_8065,N_7853,N_7346);
or U8066 (N_8066,N_7416,N_7989);
nand U8067 (N_8067,N_7874,N_7337);
or U8068 (N_8068,N_7628,N_7651);
or U8069 (N_8069,N_7827,N_7372);
xor U8070 (N_8070,N_7492,N_7817);
nand U8071 (N_8071,N_7546,N_7933);
nor U8072 (N_8072,N_7367,N_7710);
or U8073 (N_8073,N_7425,N_7446);
or U8074 (N_8074,N_7779,N_7613);
nand U8075 (N_8075,N_7414,N_7466);
xor U8076 (N_8076,N_7691,N_7845);
nor U8077 (N_8077,N_7210,N_7753);
nor U8078 (N_8078,N_7723,N_7661);
and U8079 (N_8079,N_7335,N_7664);
nand U8080 (N_8080,N_7639,N_7979);
nor U8081 (N_8081,N_7266,N_7921);
nand U8082 (N_8082,N_7982,N_7821);
xnor U8083 (N_8083,N_7922,N_7614);
xor U8084 (N_8084,N_7856,N_7622);
or U8085 (N_8085,N_7686,N_7819);
xnor U8086 (N_8086,N_7352,N_7833);
xor U8087 (N_8087,N_7876,N_7203);
nand U8088 (N_8088,N_7674,N_7306);
nand U8089 (N_8089,N_7458,N_7744);
nor U8090 (N_8090,N_7965,N_7405);
nand U8091 (N_8091,N_7766,N_7611);
nand U8092 (N_8092,N_7777,N_7276);
nand U8093 (N_8093,N_7655,N_7700);
and U8094 (N_8094,N_7765,N_7930);
nand U8095 (N_8095,N_7741,N_7236);
xnor U8096 (N_8096,N_7497,N_7583);
or U8097 (N_8097,N_7288,N_7620);
nand U8098 (N_8098,N_7452,N_7464);
and U8099 (N_8099,N_7643,N_7440);
nor U8100 (N_8100,N_7715,N_7382);
or U8101 (N_8101,N_7493,N_7627);
nand U8102 (N_8102,N_7843,N_7917);
xnor U8103 (N_8103,N_7543,N_7883);
nand U8104 (N_8104,N_7808,N_7280);
nor U8105 (N_8105,N_7569,N_7437);
and U8106 (N_8106,N_7790,N_7298);
nand U8107 (N_8107,N_7364,N_7233);
xnor U8108 (N_8108,N_7736,N_7986);
xor U8109 (N_8109,N_7272,N_7807);
nor U8110 (N_8110,N_7656,N_7615);
and U8111 (N_8111,N_7540,N_7822);
xnor U8112 (N_8112,N_7398,N_7444);
and U8113 (N_8113,N_7369,N_7644);
nor U8114 (N_8114,N_7747,N_7235);
or U8115 (N_8115,N_7685,N_7223);
or U8116 (N_8116,N_7927,N_7300);
and U8117 (N_8117,N_7996,N_7209);
or U8118 (N_8118,N_7720,N_7431);
nand U8119 (N_8119,N_7984,N_7419);
xnor U8120 (N_8120,N_7699,N_7804);
nor U8121 (N_8121,N_7261,N_7901);
nand U8122 (N_8122,N_7796,N_7285);
nand U8123 (N_8123,N_7343,N_7316);
and U8124 (N_8124,N_7558,N_7972);
and U8125 (N_8125,N_7338,N_7506);
nor U8126 (N_8126,N_7637,N_7871);
nor U8127 (N_8127,N_7581,N_7453);
and U8128 (N_8128,N_7200,N_7594);
and U8129 (N_8129,N_7572,N_7676);
nor U8130 (N_8130,N_7683,N_7846);
or U8131 (N_8131,N_7696,N_7279);
and U8132 (N_8132,N_7913,N_7504);
or U8133 (N_8133,N_7375,N_7858);
or U8134 (N_8134,N_7563,N_7376);
xor U8135 (N_8135,N_7287,N_7641);
nand U8136 (N_8136,N_7941,N_7784);
or U8137 (N_8137,N_7342,N_7511);
and U8138 (N_8138,N_7495,N_7600);
or U8139 (N_8139,N_7634,N_7960);
xor U8140 (N_8140,N_7678,N_7267);
nand U8141 (N_8141,N_7976,N_7915);
and U8142 (N_8142,N_7954,N_7435);
nor U8143 (N_8143,N_7604,N_7598);
and U8144 (N_8144,N_7350,N_7961);
xnor U8145 (N_8145,N_7773,N_7561);
xnor U8146 (N_8146,N_7225,N_7680);
and U8147 (N_8147,N_7550,N_7688);
or U8148 (N_8148,N_7697,N_7250);
or U8149 (N_8149,N_7991,N_7256);
nand U8150 (N_8150,N_7893,N_7659);
nand U8151 (N_8151,N_7245,N_7629);
nand U8152 (N_8152,N_7754,N_7229);
nor U8153 (N_8153,N_7312,N_7718);
nor U8154 (N_8154,N_7329,N_7396);
xnor U8155 (N_8155,N_7553,N_7608);
and U8156 (N_8156,N_7792,N_7428);
nor U8157 (N_8157,N_7609,N_7576);
and U8158 (N_8158,N_7411,N_7618);
xor U8159 (N_8159,N_7739,N_7356);
nor U8160 (N_8160,N_7748,N_7932);
nand U8161 (N_8161,N_7542,N_7257);
and U8162 (N_8162,N_7535,N_7457);
nand U8163 (N_8163,N_7760,N_7417);
nor U8164 (N_8164,N_7518,N_7670);
and U8165 (N_8165,N_7508,N_7530);
or U8166 (N_8166,N_7770,N_7460);
nor U8167 (N_8167,N_7339,N_7465);
nor U8168 (N_8168,N_7359,N_7671);
or U8169 (N_8169,N_7263,N_7552);
xnor U8170 (N_8170,N_7646,N_7286);
nor U8171 (N_8171,N_7767,N_7782);
nand U8172 (N_8172,N_7978,N_7675);
nor U8173 (N_8173,N_7776,N_7772);
nand U8174 (N_8174,N_7724,N_7562);
nor U8175 (N_8175,N_7219,N_7379);
or U8176 (N_8176,N_7840,N_7823);
or U8177 (N_8177,N_7653,N_7523);
and U8178 (N_8178,N_7935,N_7564);
nor U8179 (N_8179,N_7836,N_7489);
or U8180 (N_8180,N_7909,N_7851);
xnor U8181 (N_8181,N_7895,N_7325);
xnor U8182 (N_8182,N_7443,N_7570);
nor U8183 (N_8183,N_7809,N_7242);
nand U8184 (N_8184,N_7310,N_7947);
nor U8185 (N_8185,N_7404,N_7392);
nor U8186 (N_8186,N_7317,N_7877);
nand U8187 (N_8187,N_7366,N_7278);
nor U8188 (N_8188,N_7905,N_7409);
or U8189 (N_8189,N_7467,N_7362);
and U8190 (N_8190,N_7212,N_7487);
or U8191 (N_8191,N_7368,N_7571);
nor U8192 (N_8192,N_7215,N_7313);
and U8193 (N_8193,N_7816,N_7590);
xnor U8194 (N_8194,N_7701,N_7946);
and U8195 (N_8195,N_7652,N_7284);
xor U8196 (N_8196,N_7829,N_7585);
nand U8197 (N_8197,N_7221,N_7394);
nor U8198 (N_8198,N_7309,N_7201);
and U8199 (N_8199,N_7408,N_7586);
and U8200 (N_8200,N_7218,N_7998);
nor U8201 (N_8201,N_7271,N_7529);
xnor U8202 (N_8202,N_7788,N_7255);
nand U8203 (N_8203,N_7591,N_7554);
nand U8204 (N_8204,N_7891,N_7450);
nand U8205 (N_8205,N_7746,N_7679);
xor U8206 (N_8206,N_7663,N_7463);
and U8207 (N_8207,N_7204,N_7295);
nand U8208 (N_8208,N_7665,N_7442);
and U8209 (N_8209,N_7757,N_7573);
and U8210 (N_8210,N_7631,N_7380);
or U8211 (N_8211,N_7865,N_7669);
nor U8212 (N_8212,N_7393,N_7526);
and U8213 (N_8213,N_7943,N_7794);
nand U8214 (N_8214,N_7800,N_7835);
nor U8215 (N_8215,N_7422,N_7726);
nand U8216 (N_8216,N_7980,N_7484);
nor U8217 (N_8217,N_7383,N_7541);
nor U8218 (N_8218,N_7389,N_7842);
xor U8219 (N_8219,N_7934,N_7818);
or U8220 (N_8220,N_7789,N_7361);
xor U8221 (N_8221,N_7977,N_7721);
or U8222 (N_8222,N_7601,N_7657);
xor U8223 (N_8223,N_7498,N_7333);
or U8224 (N_8224,N_7412,N_7249);
nor U8225 (N_8225,N_7479,N_7716);
nor U8226 (N_8226,N_7481,N_7547);
nor U8227 (N_8227,N_7349,N_7549);
or U8228 (N_8228,N_7538,N_7722);
and U8229 (N_8229,N_7582,N_7881);
nor U8230 (N_8230,N_7423,N_7769);
nand U8231 (N_8231,N_7238,N_7875);
and U8232 (N_8232,N_7888,N_7258);
xor U8233 (N_8233,N_7574,N_7331);
and U8234 (N_8234,N_7742,N_7587);
or U8235 (N_8235,N_7294,N_7962);
or U8236 (N_8236,N_7662,N_7568);
nand U8237 (N_8237,N_7936,N_7768);
or U8238 (N_8238,N_7737,N_7602);
and U8239 (N_8239,N_7385,N_7514);
nand U8240 (N_8240,N_7551,N_7795);
xor U8241 (N_8241,N_7270,N_7430);
nand U8242 (N_8242,N_7825,N_7959);
or U8243 (N_8243,N_7640,N_7786);
xnor U8244 (N_8244,N_7780,N_7673);
nor U8245 (N_8245,N_7351,N_7923);
and U8246 (N_8246,N_7969,N_7870);
xnor U8247 (N_8247,N_7973,N_7462);
nand U8248 (N_8248,N_7476,N_7642);
nand U8249 (N_8249,N_7545,N_7344);
or U8250 (N_8250,N_7743,N_7559);
xor U8251 (N_8251,N_7911,N_7330);
and U8252 (N_8252,N_7605,N_7328);
nor U8253 (N_8253,N_7964,N_7660);
nor U8254 (N_8254,N_7597,N_7759);
nor U8255 (N_8255,N_7228,N_7580);
nor U8256 (N_8256,N_7555,N_7418);
nor U8257 (N_8257,N_7860,N_7750);
nor U8258 (N_8258,N_7231,N_7734);
xor U8259 (N_8259,N_7413,N_7533);
and U8260 (N_8260,N_7395,N_7515);
nand U8261 (N_8261,N_7578,N_7717);
and U8262 (N_8262,N_7475,N_7706);
nand U8263 (N_8263,N_7619,N_7441);
nand U8264 (N_8264,N_7912,N_7301);
and U8265 (N_8265,N_7323,N_7303);
xnor U8266 (N_8266,N_7707,N_7802);
xnor U8267 (N_8267,N_7289,N_7704);
or U8268 (N_8268,N_7624,N_7702);
nor U8269 (N_8269,N_7854,N_7771);
xnor U8270 (N_8270,N_7478,N_7510);
nand U8271 (N_8271,N_7762,N_7381);
nor U8272 (N_8272,N_7474,N_7849);
or U8273 (N_8273,N_7957,N_7745);
xnor U8274 (N_8274,N_7296,N_7928);
or U8275 (N_8275,N_7885,N_7682);
and U8276 (N_8276,N_7897,N_7341);
and U8277 (N_8277,N_7269,N_7358);
xor U8278 (N_8278,N_7797,N_7761);
nor U8279 (N_8279,N_7548,N_7812);
or U8280 (N_8280,N_7763,N_7695);
nor U8281 (N_8281,N_7519,N_7447);
nor U8282 (N_8282,N_7539,N_7482);
xnor U8283 (N_8283,N_7505,N_7360);
and U8284 (N_8284,N_7322,N_7427);
nand U8285 (N_8285,N_7436,N_7887);
or U8286 (N_8286,N_7244,N_7630);
nor U8287 (N_8287,N_7890,N_7400);
xor U8288 (N_8288,N_7705,N_7406);
and U8289 (N_8289,N_7756,N_7855);
xnor U8290 (N_8290,N_7793,N_7292);
xor U8291 (N_8291,N_7983,N_7274);
xnor U8292 (N_8292,N_7873,N_7951);
and U8293 (N_8293,N_7813,N_7919);
and U8294 (N_8294,N_7544,N_7711);
and U8295 (N_8295,N_7593,N_7448);
or U8296 (N_8296,N_7799,N_7981);
nand U8297 (N_8297,N_7579,N_7304);
nor U8298 (N_8298,N_7810,N_7975);
nand U8299 (N_8299,N_7785,N_7211);
xor U8300 (N_8300,N_7208,N_7811);
nand U8301 (N_8301,N_7326,N_7636);
xor U8302 (N_8302,N_7246,N_7677);
or U8303 (N_8303,N_7626,N_7949);
or U8304 (N_8304,N_7617,N_7282);
nand U8305 (N_8305,N_7970,N_7232);
or U8306 (N_8306,N_7589,N_7898);
xor U8307 (N_8307,N_7621,N_7603);
nor U8308 (N_8308,N_7357,N_7532);
nor U8309 (N_8309,N_7283,N_7388);
and U8310 (N_8310,N_7528,N_7607);
nand U8311 (N_8311,N_7914,N_7950);
xor U8312 (N_8312,N_7264,N_7297);
xnor U8313 (N_8313,N_7449,N_7781);
xor U8314 (N_8314,N_7248,N_7252);
nand U8315 (N_8315,N_7841,N_7832);
and U8316 (N_8316,N_7491,N_7952);
xor U8317 (N_8317,N_7319,N_7714);
or U8318 (N_8318,N_7596,N_7729);
xnor U8319 (N_8319,N_7472,N_7878);
xnor U8320 (N_8320,N_7480,N_7882);
nand U8321 (N_8321,N_7971,N_7299);
xnor U8322 (N_8322,N_7752,N_7262);
or U8323 (N_8323,N_7340,N_7650);
nand U8324 (N_8324,N_7321,N_7486);
or U8325 (N_8325,N_7625,N_7226);
nor U8326 (N_8326,N_7623,N_7426);
xnor U8327 (N_8327,N_7494,N_7205);
xnor U8328 (N_8328,N_7501,N_7524);
nand U8329 (N_8329,N_7945,N_7774);
xnor U8330 (N_8330,N_7500,N_7733);
or U8331 (N_8331,N_7327,N_7520);
nand U8332 (N_8332,N_7985,N_7222);
or U8333 (N_8333,N_7948,N_7521);
nand U8334 (N_8334,N_7916,N_7863);
nor U8335 (N_8335,N_7940,N_7536);
and U8336 (N_8336,N_7926,N_7668);
nor U8337 (N_8337,N_7220,N_7694);
xnor U8338 (N_8338,N_7993,N_7703);
nand U8339 (N_8339,N_7445,N_7241);
or U8340 (N_8340,N_7740,N_7693);
or U8341 (N_8341,N_7527,N_7277);
and U8342 (N_8342,N_7567,N_7531);
and U8343 (N_8343,N_7320,N_7654);
and U8344 (N_8344,N_7599,N_7839);
nor U8345 (N_8345,N_7240,N_7260);
or U8346 (N_8346,N_7213,N_7838);
or U8347 (N_8347,N_7963,N_7537);
and U8348 (N_8348,N_7837,N_7234);
nand U8349 (N_8349,N_7738,N_7370);
and U8350 (N_8350,N_7399,N_7681);
nand U8351 (N_8351,N_7869,N_7302);
nand U8352 (N_8352,N_7421,N_7468);
nand U8353 (N_8353,N_7872,N_7410);
or U8354 (N_8354,N_7311,N_7958);
nand U8355 (N_8355,N_7616,N_7239);
and U8356 (N_8356,N_7968,N_7689);
nand U8357 (N_8357,N_7931,N_7727);
xor U8358 (N_8358,N_7281,N_7658);
xnor U8359 (N_8359,N_7424,N_7386);
or U8360 (N_8360,N_7666,N_7347);
and U8361 (N_8361,N_7251,N_7378);
xnor U8362 (N_8362,N_7815,N_7814);
and U8363 (N_8363,N_7401,N_7953);
and U8364 (N_8364,N_7407,N_7324);
xnor U8365 (N_8365,N_7560,N_7698);
and U8366 (N_8366,N_7713,N_7307);
nand U8367 (N_8367,N_7254,N_7775);
or U8368 (N_8368,N_7939,N_7758);
nor U8369 (N_8369,N_7434,N_7732);
or U8370 (N_8370,N_7755,N_7454);
xnor U8371 (N_8371,N_7904,N_7461);
and U8372 (N_8372,N_7848,N_7824);
nor U8373 (N_8373,N_7314,N_7690);
or U8374 (N_8374,N_7647,N_7894);
xnor U8375 (N_8375,N_7862,N_7712);
nand U8376 (N_8376,N_7556,N_7731);
and U8377 (N_8377,N_7684,N_7956);
xnor U8378 (N_8378,N_7764,N_7384);
and U8379 (N_8379,N_7606,N_7778);
xnor U8380 (N_8380,N_7415,N_7374);
xor U8381 (N_8381,N_7354,N_7471);
and U8382 (N_8382,N_7216,N_7391);
nand U8383 (N_8383,N_7377,N_7612);
and U8384 (N_8384,N_7336,N_7268);
nand U8385 (N_8385,N_7451,N_7944);
or U8386 (N_8386,N_7974,N_7610);
and U8387 (N_8387,N_7879,N_7227);
or U8388 (N_8388,N_7725,N_7749);
nor U8389 (N_8389,N_7308,N_7577);
or U8390 (N_8390,N_7565,N_7513);
and U8391 (N_8391,N_7635,N_7455);
nor U8392 (N_8392,N_7884,N_7866);
xor U8393 (N_8393,N_7801,N_7557);
xor U8394 (N_8394,N_7831,N_7230);
nor U8395 (N_8395,N_7305,N_7592);
xor U8396 (N_8396,N_7345,N_7438);
xor U8397 (N_8397,N_7828,N_7459);
and U8398 (N_8398,N_7499,N_7920);
nor U8399 (N_8399,N_7803,N_7390);
xnor U8400 (N_8400,N_7935,N_7279);
or U8401 (N_8401,N_7831,N_7547);
and U8402 (N_8402,N_7510,N_7589);
xor U8403 (N_8403,N_7736,N_7586);
and U8404 (N_8404,N_7293,N_7695);
xnor U8405 (N_8405,N_7959,N_7910);
nand U8406 (N_8406,N_7293,N_7832);
xor U8407 (N_8407,N_7619,N_7942);
nor U8408 (N_8408,N_7358,N_7990);
and U8409 (N_8409,N_7378,N_7434);
nor U8410 (N_8410,N_7652,N_7610);
and U8411 (N_8411,N_7598,N_7300);
and U8412 (N_8412,N_7244,N_7468);
and U8413 (N_8413,N_7633,N_7723);
and U8414 (N_8414,N_7528,N_7584);
nand U8415 (N_8415,N_7945,N_7212);
and U8416 (N_8416,N_7606,N_7813);
or U8417 (N_8417,N_7891,N_7263);
nand U8418 (N_8418,N_7835,N_7440);
xnor U8419 (N_8419,N_7248,N_7217);
or U8420 (N_8420,N_7825,N_7971);
or U8421 (N_8421,N_7307,N_7247);
or U8422 (N_8422,N_7415,N_7445);
nand U8423 (N_8423,N_7894,N_7342);
xnor U8424 (N_8424,N_7999,N_7689);
xor U8425 (N_8425,N_7324,N_7231);
nand U8426 (N_8426,N_7408,N_7240);
nand U8427 (N_8427,N_7749,N_7614);
xnor U8428 (N_8428,N_7422,N_7501);
xnor U8429 (N_8429,N_7771,N_7845);
xnor U8430 (N_8430,N_7450,N_7423);
nand U8431 (N_8431,N_7767,N_7857);
and U8432 (N_8432,N_7605,N_7692);
nor U8433 (N_8433,N_7441,N_7239);
and U8434 (N_8434,N_7257,N_7869);
nor U8435 (N_8435,N_7654,N_7512);
nand U8436 (N_8436,N_7468,N_7516);
or U8437 (N_8437,N_7785,N_7304);
nand U8438 (N_8438,N_7384,N_7524);
and U8439 (N_8439,N_7716,N_7783);
xnor U8440 (N_8440,N_7801,N_7539);
nand U8441 (N_8441,N_7677,N_7658);
nand U8442 (N_8442,N_7468,N_7472);
nand U8443 (N_8443,N_7302,N_7371);
or U8444 (N_8444,N_7783,N_7292);
nand U8445 (N_8445,N_7785,N_7426);
nor U8446 (N_8446,N_7852,N_7491);
nand U8447 (N_8447,N_7786,N_7773);
xor U8448 (N_8448,N_7998,N_7640);
xnor U8449 (N_8449,N_7823,N_7912);
nand U8450 (N_8450,N_7569,N_7925);
xor U8451 (N_8451,N_7732,N_7814);
xor U8452 (N_8452,N_7972,N_7574);
nor U8453 (N_8453,N_7434,N_7812);
or U8454 (N_8454,N_7626,N_7996);
and U8455 (N_8455,N_7900,N_7858);
or U8456 (N_8456,N_7585,N_7847);
nand U8457 (N_8457,N_7388,N_7370);
nand U8458 (N_8458,N_7915,N_7997);
nor U8459 (N_8459,N_7286,N_7708);
xnor U8460 (N_8460,N_7564,N_7478);
xnor U8461 (N_8461,N_7317,N_7716);
or U8462 (N_8462,N_7615,N_7847);
nand U8463 (N_8463,N_7804,N_7729);
and U8464 (N_8464,N_7537,N_7733);
nand U8465 (N_8465,N_7353,N_7764);
nand U8466 (N_8466,N_7209,N_7952);
xnor U8467 (N_8467,N_7715,N_7608);
xnor U8468 (N_8468,N_7321,N_7335);
nand U8469 (N_8469,N_7560,N_7673);
nor U8470 (N_8470,N_7419,N_7874);
xor U8471 (N_8471,N_7365,N_7718);
or U8472 (N_8472,N_7940,N_7916);
and U8473 (N_8473,N_7363,N_7225);
xor U8474 (N_8474,N_7408,N_7244);
or U8475 (N_8475,N_7911,N_7373);
and U8476 (N_8476,N_7473,N_7663);
or U8477 (N_8477,N_7529,N_7233);
xnor U8478 (N_8478,N_7813,N_7532);
xor U8479 (N_8479,N_7829,N_7269);
nand U8480 (N_8480,N_7734,N_7524);
or U8481 (N_8481,N_7767,N_7975);
xor U8482 (N_8482,N_7791,N_7301);
or U8483 (N_8483,N_7888,N_7560);
or U8484 (N_8484,N_7293,N_7823);
xor U8485 (N_8485,N_7703,N_7930);
or U8486 (N_8486,N_7500,N_7280);
nor U8487 (N_8487,N_7241,N_7796);
nand U8488 (N_8488,N_7241,N_7720);
xnor U8489 (N_8489,N_7386,N_7640);
nor U8490 (N_8490,N_7239,N_7838);
xnor U8491 (N_8491,N_7553,N_7941);
nor U8492 (N_8492,N_7444,N_7485);
xor U8493 (N_8493,N_7520,N_7909);
or U8494 (N_8494,N_7205,N_7747);
or U8495 (N_8495,N_7236,N_7580);
nand U8496 (N_8496,N_7771,N_7976);
nand U8497 (N_8497,N_7891,N_7273);
and U8498 (N_8498,N_7877,N_7709);
or U8499 (N_8499,N_7825,N_7807);
or U8500 (N_8500,N_7203,N_7270);
xor U8501 (N_8501,N_7253,N_7695);
or U8502 (N_8502,N_7456,N_7798);
xor U8503 (N_8503,N_7981,N_7232);
nand U8504 (N_8504,N_7535,N_7869);
nor U8505 (N_8505,N_7883,N_7786);
and U8506 (N_8506,N_7394,N_7203);
nand U8507 (N_8507,N_7651,N_7503);
xor U8508 (N_8508,N_7326,N_7742);
or U8509 (N_8509,N_7850,N_7750);
xor U8510 (N_8510,N_7464,N_7821);
xor U8511 (N_8511,N_7607,N_7884);
nand U8512 (N_8512,N_7900,N_7277);
and U8513 (N_8513,N_7731,N_7410);
or U8514 (N_8514,N_7936,N_7623);
xnor U8515 (N_8515,N_7457,N_7952);
xnor U8516 (N_8516,N_7739,N_7481);
and U8517 (N_8517,N_7472,N_7432);
nand U8518 (N_8518,N_7229,N_7331);
nor U8519 (N_8519,N_7370,N_7380);
and U8520 (N_8520,N_7911,N_7755);
nand U8521 (N_8521,N_7531,N_7700);
xnor U8522 (N_8522,N_7239,N_7945);
nor U8523 (N_8523,N_7369,N_7966);
xor U8524 (N_8524,N_7670,N_7290);
xor U8525 (N_8525,N_7399,N_7669);
nor U8526 (N_8526,N_7629,N_7789);
and U8527 (N_8527,N_7333,N_7946);
xor U8528 (N_8528,N_7243,N_7904);
or U8529 (N_8529,N_7313,N_7547);
xnor U8530 (N_8530,N_7212,N_7617);
nand U8531 (N_8531,N_7403,N_7512);
and U8532 (N_8532,N_7335,N_7424);
xnor U8533 (N_8533,N_7618,N_7451);
and U8534 (N_8534,N_7837,N_7766);
xor U8535 (N_8535,N_7469,N_7731);
or U8536 (N_8536,N_7617,N_7920);
xnor U8537 (N_8537,N_7221,N_7844);
nor U8538 (N_8538,N_7607,N_7665);
xnor U8539 (N_8539,N_7457,N_7417);
nand U8540 (N_8540,N_7551,N_7282);
nand U8541 (N_8541,N_7393,N_7542);
or U8542 (N_8542,N_7968,N_7990);
xor U8543 (N_8543,N_7455,N_7612);
nand U8544 (N_8544,N_7864,N_7532);
and U8545 (N_8545,N_7219,N_7744);
xnor U8546 (N_8546,N_7676,N_7563);
nor U8547 (N_8547,N_7627,N_7375);
xor U8548 (N_8548,N_7589,N_7762);
xor U8549 (N_8549,N_7650,N_7215);
nand U8550 (N_8550,N_7760,N_7806);
or U8551 (N_8551,N_7898,N_7878);
nand U8552 (N_8552,N_7254,N_7724);
xnor U8553 (N_8553,N_7328,N_7260);
nor U8554 (N_8554,N_7909,N_7554);
and U8555 (N_8555,N_7982,N_7895);
nor U8556 (N_8556,N_7647,N_7266);
and U8557 (N_8557,N_7759,N_7265);
and U8558 (N_8558,N_7759,N_7718);
and U8559 (N_8559,N_7401,N_7405);
nor U8560 (N_8560,N_7909,N_7375);
and U8561 (N_8561,N_7321,N_7351);
nor U8562 (N_8562,N_7784,N_7354);
nor U8563 (N_8563,N_7970,N_7360);
and U8564 (N_8564,N_7265,N_7916);
xor U8565 (N_8565,N_7567,N_7564);
or U8566 (N_8566,N_7396,N_7487);
xnor U8567 (N_8567,N_7546,N_7362);
and U8568 (N_8568,N_7353,N_7336);
or U8569 (N_8569,N_7519,N_7645);
or U8570 (N_8570,N_7910,N_7969);
or U8571 (N_8571,N_7514,N_7662);
nor U8572 (N_8572,N_7751,N_7587);
xnor U8573 (N_8573,N_7453,N_7310);
and U8574 (N_8574,N_7848,N_7481);
nor U8575 (N_8575,N_7659,N_7717);
nor U8576 (N_8576,N_7249,N_7586);
xnor U8577 (N_8577,N_7862,N_7938);
or U8578 (N_8578,N_7629,N_7875);
and U8579 (N_8579,N_7942,N_7840);
nor U8580 (N_8580,N_7665,N_7238);
nand U8581 (N_8581,N_7886,N_7905);
or U8582 (N_8582,N_7272,N_7528);
xor U8583 (N_8583,N_7884,N_7799);
and U8584 (N_8584,N_7969,N_7448);
nand U8585 (N_8585,N_7463,N_7373);
and U8586 (N_8586,N_7634,N_7243);
nand U8587 (N_8587,N_7728,N_7274);
xor U8588 (N_8588,N_7866,N_7433);
xor U8589 (N_8589,N_7957,N_7738);
nor U8590 (N_8590,N_7997,N_7862);
xor U8591 (N_8591,N_7350,N_7706);
and U8592 (N_8592,N_7951,N_7376);
or U8593 (N_8593,N_7944,N_7417);
nand U8594 (N_8594,N_7473,N_7783);
or U8595 (N_8595,N_7300,N_7220);
or U8596 (N_8596,N_7868,N_7980);
and U8597 (N_8597,N_7859,N_7517);
and U8598 (N_8598,N_7519,N_7343);
nor U8599 (N_8599,N_7986,N_7550);
xnor U8600 (N_8600,N_7357,N_7726);
nand U8601 (N_8601,N_7800,N_7231);
or U8602 (N_8602,N_7425,N_7466);
and U8603 (N_8603,N_7698,N_7928);
or U8604 (N_8604,N_7208,N_7200);
xnor U8605 (N_8605,N_7417,N_7343);
and U8606 (N_8606,N_7863,N_7514);
xor U8607 (N_8607,N_7878,N_7947);
xor U8608 (N_8608,N_7850,N_7813);
and U8609 (N_8609,N_7248,N_7555);
nand U8610 (N_8610,N_7804,N_7244);
or U8611 (N_8611,N_7700,N_7460);
nand U8612 (N_8612,N_7317,N_7836);
or U8613 (N_8613,N_7734,N_7695);
and U8614 (N_8614,N_7893,N_7288);
and U8615 (N_8615,N_7550,N_7689);
nand U8616 (N_8616,N_7321,N_7484);
nor U8617 (N_8617,N_7645,N_7343);
nor U8618 (N_8618,N_7592,N_7973);
xnor U8619 (N_8619,N_7701,N_7441);
xor U8620 (N_8620,N_7794,N_7566);
nand U8621 (N_8621,N_7716,N_7917);
and U8622 (N_8622,N_7543,N_7260);
xnor U8623 (N_8623,N_7747,N_7547);
and U8624 (N_8624,N_7515,N_7851);
nand U8625 (N_8625,N_7234,N_7826);
or U8626 (N_8626,N_7918,N_7577);
and U8627 (N_8627,N_7338,N_7451);
xor U8628 (N_8628,N_7234,N_7549);
xnor U8629 (N_8629,N_7863,N_7252);
and U8630 (N_8630,N_7943,N_7769);
nand U8631 (N_8631,N_7415,N_7796);
xor U8632 (N_8632,N_7975,N_7328);
xor U8633 (N_8633,N_7405,N_7275);
nand U8634 (N_8634,N_7476,N_7744);
nand U8635 (N_8635,N_7526,N_7771);
xor U8636 (N_8636,N_7948,N_7453);
or U8637 (N_8637,N_7211,N_7710);
xor U8638 (N_8638,N_7401,N_7466);
or U8639 (N_8639,N_7278,N_7379);
or U8640 (N_8640,N_7506,N_7313);
or U8641 (N_8641,N_7560,N_7456);
or U8642 (N_8642,N_7339,N_7442);
or U8643 (N_8643,N_7416,N_7732);
or U8644 (N_8644,N_7412,N_7293);
xor U8645 (N_8645,N_7360,N_7901);
and U8646 (N_8646,N_7292,N_7524);
or U8647 (N_8647,N_7878,N_7528);
nor U8648 (N_8648,N_7695,N_7556);
or U8649 (N_8649,N_7391,N_7851);
nor U8650 (N_8650,N_7999,N_7383);
or U8651 (N_8651,N_7685,N_7658);
nor U8652 (N_8652,N_7652,N_7489);
nor U8653 (N_8653,N_7864,N_7612);
or U8654 (N_8654,N_7801,N_7275);
and U8655 (N_8655,N_7456,N_7616);
or U8656 (N_8656,N_7806,N_7567);
or U8657 (N_8657,N_7215,N_7958);
or U8658 (N_8658,N_7644,N_7529);
nor U8659 (N_8659,N_7388,N_7754);
nand U8660 (N_8660,N_7827,N_7787);
xnor U8661 (N_8661,N_7750,N_7839);
xor U8662 (N_8662,N_7239,N_7712);
nor U8663 (N_8663,N_7778,N_7963);
nor U8664 (N_8664,N_7689,N_7497);
and U8665 (N_8665,N_7939,N_7965);
or U8666 (N_8666,N_7543,N_7499);
or U8667 (N_8667,N_7606,N_7409);
or U8668 (N_8668,N_7894,N_7863);
or U8669 (N_8669,N_7816,N_7380);
xnor U8670 (N_8670,N_7593,N_7655);
nand U8671 (N_8671,N_7827,N_7897);
nor U8672 (N_8672,N_7594,N_7914);
nor U8673 (N_8673,N_7546,N_7419);
and U8674 (N_8674,N_7967,N_7514);
and U8675 (N_8675,N_7587,N_7971);
nand U8676 (N_8676,N_7344,N_7375);
nor U8677 (N_8677,N_7844,N_7962);
xor U8678 (N_8678,N_7456,N_7737);
nor U8679 (N_8679,N_7813,N_7949);
xor U8680 (N_8680,N_7250,N_7327);
nor U8681 (N_8681,N_7641,N_7726);
xor U8682 (N_8682,N_7559,N_7210);
or U8683 (N_8683,N_7646,N_7617);
xor U8684 (N_8684,N_7456,N_7207);
and U8685 (N_8685,N_7634,N_7281);
or U8686 (N_8686,N_7933,N_7457);
and U8687 (N_8687,N_7286,N_7435);
or U8688 (N_8688,N_7975,N_7881);
xor U8689 (N_8689,N_7623,N_7571);
or U8690 (N_8690,N_7678,N_7700);
or U8691 (N_8691,N_7867,N_7692);
nor U8692 (N_8692,N_7646,N_7838);
nand U8693 (N_8693,N_7415,N_7914);
nand U8694 (N_8694,N_7357,N_7756);
or U8695 (N_8695,N_7524,N_7917);
nor U8696 (N_8696,N_7459,N_7554);
nand U8697 (N_8697,N_7775,N_7581);
nor U8698 (N_8698,N_7603,N_7620);
nand U8699 (N_8699,N_7717,N_7950);
xor U8700 (N_8700,N_7805,N_7853);
nor U8701 (N_8701,N_7820,N_7893);
xnor U8702 (N_8702,N_7312,N_7513);
nor U8703 (N_8703,N_7446,N_7842);
xor U8704 (N_8704,N_7446,N_7517);
and U8705 (N_8705,N_7967,N_7461);
nand U8706 (N_8706,N_7321,N_7639);
or U8707 (N_8707,N_7822,N_7632);
or U8708 (N_8708,N_7654,N_7923);
or U8709 (N_8709,N_7717,N_7887);
nand U8710 (N_8710,N_7871,N_7675);
xor U8711 (N_8711,N_7557,N_7603);
xnor U8712 (N_8712,N_7366,N_7450);
nor U8713 (N_8713,N_7888,N_7961);
and U8714 (N_8714,N_7683,N_7596);
nand U8715 (N_8715,N_7444,N_7250);
nor U8716 (N_8716,N_7690,N_7746);
xor U8717 (N_8717,N_7228,N_7992);
nor U8718 (N_8718,N_7451,N_7464);
or U8719 (N_8719,N_7218,N_7707);
and U8720 (N_8720,N_7727,N_7274);
and U8721 (N_8721,N_7258,N_7727);
nand U8722 (N_8722,N_7684,N_7858);
nand U8723 (N_8723,N_7473,N_7384);
xnor U8724 (N_8724,N_7804,N_7458);
and U8725 (N_8725,N_7642,N_7507);
and U8726 (N_8726,N_7270,N_7865);
and U8727 (N_8727,N_7926,N_7605);
and U8728 (N_8728,N_7358,N_7914);
and U8729 (N_8729,N_7687,N_7389);
nor U8730 (N_8730,N_7750,N_7327);
and U8731 (N_8731,N_7300,N_7213);
nor U8732 (N_8732,N_7738,N_7346);
xnor U8733 (N_8733,N_7917,N_7579);
or U8734 (N_8734,N_7986,N_7755);
xnor U8735 (N_8735,N_7717,N_7387);
nor U8736 (N_8736,N_7439,N_7663);
or U8737 (N_8737,N_7603,N_7458);
or U8738 (N_8738,N_7481,N_7401);
xor U8739 (N_8739,N_7515,N_7413);
and U8740 (N_8740,N_7485,N_7539);
and U8741 (N_8741,N_7568,N_7257);
nor U8742 (N_8742,N_7680,N_7568);
or U8743 (N_8743,N_7872,N_7624);
xor U8744 (N_8744,N_7992,N_7851);
or U8745 (N_8745,N_7853,N_7422);
xnor U8746 (N_8746,N_7711,N_7657);
xnor U8747 (N_8747,N_7766,N_7903);
and U8748 (N_8748,N_7659,N_7510);
and U8749 (N_8749,N_7602,N_7210);
xnor U8750 (N_8750,N_7534,N_7543);
nand U8751 (N_8751,N_7890,N_7830);
xnor U8752 (N_8752,N_7398,N_7258);
or U8753 (N_8753,N_7377,N_7473);
or U8754 (N_8754,N_7762,N_7936);
nor U8755 (N_8755,N_7670,N_7316);
and U8756 (N_8756,N_7940,N_7632);
xor U8757 (N_8757,N_7597,N_7335);
nand U8758 (N_8758,N_7609,N_7558);
nand U8759 (N_8759,N_7383,N_7328);
and U8760 (N_8760,N_7976,N_7758);
and U8761 (N_8761,N_7791,N_7706);
nor U8762 (N_8762,N_7526,N_7525);
or U8763 (N_8763,N_7928,N_7207);
xor U8764 (N_8764,N_7422,N_7200);
xnor U8765 (N_8765,N_7213,N_7561);
nor U8766 (N_8766,N_7367,N_7364);
nor U8767 (N_8767,N_7834,N_7482);
and U8768 (N_8768,N_7621,N_7333);
nor U8769 (N_8769,N_7434,N_7852);
nor U8770 (N_8770,N_7333,N_7216);
nand U8771 (N_8771,N_7218,N_7913);
or U8772 (N_8772,N_7770,N_7744);
nor U8773 (N_8773,N_7887,N_7255);
nor U8774 (N_8774,N_7412,N_7479);
or U8775 (N_8775,N_7978,N_7301);
nor U8776 (N_8776,N_7932,N_7741);
nand U8777 (N_8777,N_7871,N_7608);
and U8778 (N_8778,N_7261,N_7871);
and U8779 (N_8779,N_7521,N_7794);
xor U8780 (N_8780,N_7684,N_7521);
nor U8781 (N_8781,N_7634,N_7664);
nor U8782 (N_8782,N_7367,N_7595);
xnor U8783 (N_8783,N_7905,N_7280);
nor U8784 (N_8784,N_7921,N_7340);
nor U8785 (N_8785,N_7698,N_7509);
or U8786 (N_8786,N_7305,N_7438);
and U8787 (N_8787,N_7203,N_7573);
and U8788 (N_8788,N_7442,N_7876);
xor U8789 (N_8789,N_7474,N_7519);
nand U8790 (N_8790,N_7417,N_7702);
or U8791 (N_8791,N_7931,N_7567);
or U8792 (N_8792,N_7722,N_7586);
or U8793 (N_8793,N_7736,N_7980);
xnor U8794 (N_8794,N_7752,N_7288);
or U8795 (N_8795,N_7634,N_7514);
and U8796 (N_8796,N_7938,N_7558);
nor U8797 (N_8797,N_7493,N_7383);
nand U8798 (N_8798,N_7915,N_7201);
nor U8799 (N_8799,N_7571,N_7712);
or U8800 (N_8800,N_8198,N_8486);
or U8801 (N_8801,N_8248,N_8595);
nand U8802 (N_8802,N_8377,N_8205);
or U8803 (N_8803,N_8073,N_8142);
or U8804 (N_8804,N_8481,N_8407);
xnor U8805 (N_8805,N_8523,N_8517);
nand U8806 (N_8806,N_8155,N_8792);
nand U8807 (N_8807,N_8569,N_8176);
nor U8808 (N_8808,N_8615,N_8276);
or U8809 (N_8809,N_8379,N_8398);
and U8810 (N_8810,N_8107,N_8558);
and U8811 (N_8811,N_8571,N_8119);
xor U8812 (N_8812,N_8644,N_8255);
or U8813 (N_8813,N_8663,N_8207);
and U8814 (N_8814,N_8136,N_8752);
xor U8815 (N_8815,N_8202,N_8471);
nor U8816 (N_8816,N_8094,N_8015);
nand U8817 (N_8817,N_8418,N_8568);
nor U8818 (N_8818,N_8223,N_8295);
nor U8819 (N_8819,N_8596,N_8592);
or U8820 (N_8820,N_8635,N_8342);
nand U8821 (N_8821,N_8540,N_8439);
nor U8822 (N_8822,N_8695,N_8472);
nand U8823 (N_8823,N_8030,N_8146);
nor U8824 (N_8824,N_8056,N_8011);
and U8825 (N_8825,N_8326,N_8717);
nand U8826 (N_8826,N_8348,N_8550);
nand U8827 (N_8827,N_8519,N_8704);
xnor U8828 (N_8828,N_8066,N_8389);
nand U8829 (N_8829,N_8562,N_8628);
xnor U8830 (N_8830,N_8288,N_8224);
xor U8831 (N_8831,N_8428,N_8425);
nand U8832 (N_8832,N_8339,N_8547);
nor U8833 (N_8833,N_8747,N_8149);
and U8834 (N_8834,N_8749,N_8676);
or U8835 (N_8835,N_8648,N_8365);
xor U8836 (N_8836,N_8337,N_8275);
nand U8837 (N_8837,N_8419,N_8233);
and U8838 (N_8838,N_8581,N_8078);
or U8839 (N_8839,N_8551,N_8264);
nor U8840 (N_8840,N_8147,N_8725);
and U8841 (N_8841,N_8376,N_8294);
xor U8842 (N_8842,N_8602,N_8456);
and U8843 (N_8843,N_8692,N_8600);
nand U8844 (N_8844,N_8178,N_8089);
nor U8845 (N_8845,N_8382,N_8674);
and U8846 (N_8846,N_8217,N_8664);
xor U8847 (N_8847,N_8196,N_8760);
or U8848 (N_8848,N_8029,N_8772);
or U8849 (N_8849,N_8112,N_8165);
and U8850 (N_8850,N_8062,N_8753);
and U8851 (N_8851,N_8484,N_8733);
xnor U8852 (N_8852,N_8185,N_8302);
or U8853 (N_8853,N_8017,N_8651);
or U8854 (N_8854,N_8361,N_8266);
and U8855 (N_8855,N_8117,N_8021);
nand U8856 (N_8856,N_8312,N_8296);
and U8857 (N_8857,N_8270,N_8222);
and U8858 (N_8858,N_8609,N_8575);
nand U8859 (N_8859,N_8487,N_8622);
nand U8860 (N_8860,N_8114,N_8625);
nor U8861 (N_8861,N_8122,N_8032);
and U8862 (N_8862,N_8755,N_8036);
nand U8863 (N_8863,N_8409,N_8047);
nor U8864 (N_8864,N_8013,N_8197);
or U8865 (N_8865,N_8209,N_8308);
nand U8866 (N_8866,N_8031,N_8284);
or U8867 (N_8867,N_8427,N_8767);
or U8868 (N_8868,N_8229,N_8371);
nand U8869 (N_8869,N_8187,N_8099);
nand U8870 (N_8870,N_8578,N_8335);
or U8871 (N_8871,N_8509,N_8314);
nand U8872 (N_8872,N_8138,N_8152);
and U8873 (N_8873,N_8705,N_8786);
nor U8874 (N_8874,N_8189,N_8057);
nor U8875 (N_8875,N_8506,N_8706);
or U8876 (N_8876,N_8503,N_8763);
nand U8877 (N_8877,N_8433,N_8455);
or U8878 (N_8878,N_8059,N_8492);
nor U8879 (N_8879,N_8203,N_8130);
or U8880 (N_8880,N_8090,N_8160);
or U8881 (N_8881,N_8757,N_8060);
nor U8882 (N_8882,N_8403,N_8590);
nor U8883 (N_8883,N_8265,N_8765);
nor U8884 (N_8884,N_8278,N_8681);
nor U8885 (N_8885,N_8369,N_8247);
nand U8886 (N_8886,N_8037,N_8357);
xor U8887 (N_8887,N_8154,N_8531);
nand U8888 (N_8888,N_8559,N_8680);
or U8889 (N_8889,N_8137,N_8243);
nand U8890 (N_8890,N_8436,N_8024);
or U8891 (N_8891,N_8258,N_8552);
nand U8892 (N_8892,N_8678,N_8544);
or U8893 (N_8893,N_8150,N_8148);
nand U8894 (N_8894,N_8730,N_8360);
nand U8895 (N_8895,N_8659,N_8529);
or U8896 (N_8896,N_8070,N_8754);
and U8897 (N_8897,N_8387,N_8423);
nor U8898 (N_8898,N_8499,N_8785);
nand U8899 (N_8899,N_8109,N_8391);
nor U8900 (N_8900,N_8560,N_8304);
or U8901 (N_8901,N_8452,N_8654);
xnor U8902 (N_8902,N_8536,N_8118);
nand U8903 (N_8903,N_8074,N_8476);
and U8904 (N_8904,N_8333,N_8426);
xnor U8905 (N_8905,N_8175,N_8052);
or U8906 (N_8906,N_8299,N_8097);
xnor U8907 (N_8907,N_8076,N_8077);
nor U8908 (N_8908,N_8632,N_8688);
or U8909 (N_8909,N_8009,N_8171);
xor U8910 (N_8910,N_8035,N_8027);
nor U8911 (N_8911,N_8650,N_8100);
and U8912 (N_8912,N_8158,N_8239);
nor U8913 (N_8913,N_8067,N_8327);
nand U8914 (N_8914,N_8715,N_8180);
nand U8915 (N_8915,N_8631,N_8527);
or U8916 (N_8916,N_8495,N_8385);
nor U8917 (N_8917,N_8534,N_8505);
nor U8918 (N_8918,N_8718,N_8182);
nand U8919 (N_8919,N_8283,N_8338);
and U8920 (N_8920,N_8045,N_8012);
and U8921 (N_8921,N_8043,N_8514);
nor U8922 (N_8922,N_8151,N_8356);
nor U8923 (N_8923,N_8451,N_8634);
nor U8924 (N_8924,N_8216,N_8797);
or U8925 (N_8925,N_8321,N_8474);
and U8926 (N_8926,N_8719,N_8408);
nor U8927 (N_8927,N_8460,N_8344);
nor U8928 (N_8928,N_8723,N_8579);
or U8929 (N_8929,N_8269,N_8424);
nor U8930 (N_8930,N_8777,N_8336);
xor U8931 (N_8931,N_8349,N_8161);
and U8932 (N_8932,N_8058,N_8662);
xor U8933 (N_8933,N_8775,N_8210);
nand U8934 (N_8934,N_8110,N_8002);
nor U8935 (N_8935,N_8140,N_8491);
and U8936 (N_8936,N_8779,N_8623);
nor U8937 (N_8937,N_8159,N_8655);
and U8938 (N_8938,N_8004,N_8298);
nand U8939 (N_8939,N_8000,N_8724);
and U8940 (N_8940,N_8708,N_8322);
or U8941 (N_8941,N_8567,N_8561);
nand U8942 (N_8942,N_8292,N_8199);
nand U8943 (N_8943,N_8186,N_8081);
xnor U8944 (N_8944,N_8006,N_8566);
xor U8945 (N_8945,N_8722,N_8442);
nand U8946 (N_8946,N_8345,N_8141);
or U8947 (N_8947,N_8671,N_8675);
and U8948 (N_8948,N_8039,N_8538);
nor U8949 (N_8949,N_8570,N_8466);
and U8950 (N_8950,N_8286,N_8092);
nand U8951 (N_8951,N_8370,N_8787);
nor U8952 (N_8952,N_8061,N_8438);
xor U8953 (N_8953,N_8670,N_8166);
xnor U8954 (N_8954,N_8605,N_8440);
nor U8955 (N_8955,N_8401,N_8240);
and U8956 (N_8956,N_8454,N_8368);
or U8957 (N_8957,N_8781,N_8591);
nand U8958 (N_8958,N_8657,N_8593);
or U8959 (N_8959,N_8515,N_8016);
xnor U8960 (N_8960,N_8761,N_8383);
or U8961 (N_8961,N_8443,N_8639);
nand U8962 (N_8962,N_8372,N_8684);
nand U8963 (N_8963,N_8019,N_8612);
nand U8964 (N_8964,N_8716,N_8343);
or U8965 (N_8965,N_8301,N_8709);
xor U8966 (N_8966,N_8279,N_8251);
and U8967 (N_8967,N_8572,N_8080);
and U8968 (N_8968,N_8421,N_8018);
xnor U8969 (N_8969,N_8005,N_8588);
or U8970 (N_8970,N_8790,N_8449);
nand U8971 (N_8971,N_8352,N_8771);
xnor U8972 (N_8972,N_8745,N_8250);
or U8973 (N_8973,N_8274,N_8574);
or U8974 (N_8974,N_8145,N_8049);
and U8975 (N_8975,N_8221,N_8316);
or U8976 (N_8976,N_8468,N_8020);
xor U8977 (N_8977,N_8464,N_8597);
nand U8978 (N_8978,N_8524,N_8318);
and U8979 (N_8979,N_8173,N_8402);
nand U8980 (N_8980,N_8620,N_8697);
nor U8981 (N_8981,N_8791,N_8388);
xor U8982 (N_8982,N_8477,N_8798);
nor U8983 (N_8983,N_8710,N_8378);
or U8984 (N_8984,N_8126,N_8297);
and U8985 (N_8985,N_8164,N_8188);
nor U8986 (N_8986,N_8518,N_8415);
and U8987 (N_8987,N_8698,N_8168);
and U8988 (N_8988,N_8516,N_8504);
nor U8989 (N_8989,N_8334,N_8734);
xor U8990 (N_8990,N_8762,N_8702);
nand U8991 (N_8991,N_8317,N_8743);
nand U8992 (N_8992,N_8624,N_8637);
nand U8993 (N_8993,N_8208,N_8267);
nor U8994 (N_8994,N_8381,N_8143);
nor U8995 (N_8995,N_8093,N_8195);
and U8996 (N_8996,N_8375,N_8242);
or U8997 (N_8997,N_8489,N_8774);
and U8998 (N_8998,N_8646,N_8396);
or U8999 (N_8999,N_8124,N_8068);
xnor U9000 (N_9000,N_8627,N_8022);
xnor U9001 (N_9001,N_8236,N_8354);
or U9002 (N_9002,N_8683,N_8545);
nand U9003 (N_9003,N_8135,N_8244);
and U9004 (N_9004,N_8788,N_8323);
xor U9005 (N_9005,N_8127,N_8406);
xor U9006 (N_9006,N_8034,N_8133);
and U9007 (N_9007,N_8621,N_8082);
or U9008 (N_9008,N_8201,N_8497);
xor U9009 (N_9009,N_8025,N_8351);
nand U9010 (N_9010,N_8245,N_8498);
or U9011 (N_9011,N_8102,N_8553);
xor U9012 (N_9012,N_8782,N_8626);
xor U9013 (N_9013,N_8563,N_8399);
nand U9014 (N_9014,N_8768,N_8530);
and U9015 (N_9015,N_8647,N_8618);
and U9016 (N_9016,N_8129,N_8638);
or U9017 (N_9017,N_8330,N_8305);
and U9018 (N_9018,N_8640,N_8448);
and U9019 (N_9019,N_8007,N_8483);
xnor U9020 (N_9020,N_8463,N_8393);
xor U9021 (N_9021,N_8044,N_8508);
and U9022 (N_9022,N_8480,N_8204);
nand U9023 (N_9023,N_8565,N_8268);
nand U9024 (N_9024,N_8307,N_8750);
nor U9025 (N_9025,N_8123,N_8261);
and U9026 (N_9026,N_8384,N_8083);
nor U9027 (N_9027,N_8467,N_8254);
xor U9028 (N_9028,N_8063,N_8072);
nand U9029 (N_9029,N_8218,N_8711);
xor U9030 (N_9030,N_8071,N_8580);
xor U9031 (N_9031,N_8194,N_8610);
nor U9032 (N_9032,N_8457,N_8444);
and U9033 (N_9033,N_8055,N_8096);
and U9034 (N_9034,N_8328,N_8665);
nand U9035 (N_9035,N_8794,N_8598);
or U9036 (N_9036,N_8380,N_8331);
xnor U9037 (N_9037,N_8744,N_8432);
or U9038 (N_9038,N_8796,N_8603);
nand U9039 (N_9039,N_8500,N_8246);
and U9040 (N_9040,N_8053,N_8599);
nor U9041 (N_9041,N_8586,N_8079);
or U9042 (N_9042,N_8450,N_8397);
xnor U9043 (N_9043,N_8652,N_8494);
nand U9044 (N_9044,N_8546,N_8272);
and U9045 (N_9045,N_8513,N_8347);
nor U9046 (N_9046,N_8607,N_8729);
and U9047 (N_9047,N_8736,N_8430);
nand U9048 (N_9048,N_8420,N_8738);
and U9049 (N_9049,N_8488,N_8048);
or U9050 (N_9050,N_8784,N_8253);
and U9051 (N_9051,N_8617,N_8273);
xnor U9052 (N_9052,N_8769,N_8340);
and U9053 (N_9053,N_8277,N_8374);
xnor U9054 (N_9054,N_8630,N_8134);
and U9055 (N_9055,N_8132,N_8179);
nand U9056 (N_9056,N_8104,N_8616);
nor U9057 (N_9057,N_8740,N_8390);
and U9058 (N_9058,N_8511,N_8128);
nand U9059 (N_9059,N_8542,N_8573);
xnor U9060 (N_9060,N_8667,N_8554);
xnor U9061 (N_9061,N_8672,N_8106);
nor U9062 (N_9062,N_8473,N_8543);
nor U9063 (N_9063,N_8645,N_8282);
and U9064 (N_9064,N_8183,N_8643);
and U9065 (N_9065,N_8256,N_8346);
or U9066 (N_9066,N_8341,N_8731);
nand U9067 (N_9067,N_8751,N_8422);
nor U9068 (N_9068,N_8051,N_8789);
and U9069 (N_9069,N_8091,N_8303);
nor U9070 (N_9070,N_8756,N_8167);
nand U9071 (N_9071,N_8703,N_8003);
nor U9072 (N_9072,N_8434,N_8619);
and U9073 (N_9073,N_8319,N_8726);
xnor U9074 (N_9074,N_8174,N_8050);
and U9075 (N_9075,N_8773,N_8577);
and U9076 (N_9076,N_8111,N_8582);
and U9077 (N_9077,N_8230,N_8496);
xor U9078 (N_9078,N_8026,N_8512);
nand U9079 (N_9079,N_8714,N_8776);
or U9080 (N_9080,N_8405,N_8611);
nand U9081 (N_9081,N_8220,N_8746);
nor U9082 (N_9082,N_8228,N_8690);
or U9083 (N_9083,N_8042,N_8701);
and U9084 (N_9084,N_8084,N_8727);
nand U9085 (N_9085,N_8417,N_8686);
nor U9086 (N_9086,N_8362,N_8235);
or U9087 (N_9087,N_8601,N_8105);
or U9088 (N_9088,N_8793,N_8720);
and U9089 (N_9089,N_8411,N_8033);
nor U9090 (N_9090,N_8192,N_8386);
and U9091 (N_9091,N_8555,N_8548);
nor U9092 (N_9092,N_8353,N_8172);
xnor U9093 (N_9093,N_8227,N_8054);
nand U9094 (N_9094,N_8759,N_8713);
or U9095 (N_9095,N_8413,N_8300);
xnor U9096 (N_9096,N_8121,N_8193);
xnor U9097 (N_9097,N_8212,N_8576);
or U9098 (N_9098,N_8085,N_8046);
or U9099 (N_9099,N_8501,N_8162);
xnor U9100 (N_9100,N_8144,N_8666);
xnor U9101 (N_9101,N_8458,N_8075);
and U9102 (N_9102,N_8656,N_8169);
nand U9103 (N_9103,N_8493,N_8758);
or U9104 (N_9104,N_8363,N_8693);
nand U9105 (N_9105,N_8549,N_8157);
and U9106 (N_9106,N_8320,N_8392);
nand U9107 (N_9107,N_8728,N_8677);
or U9108 (N_9108,N_8441,N_8232);
or U9109 (N_9109,N_8641,N_8226);
xnor U9110 (N_9110,N_8533,N_8661);
xnor U9111 (N_9111,N_8289,N_8748);
nand U9112 (N_9112,N_8214,N_8658);
and U9113 (N_9113,N_8490,N_8608);
nor U9114 (N_9114,N_8465,N_8783);
nor U9115 (N_9115,N_8742,N_8732);
nor U9116 (N_9116,N_8170,N_8191);
or U9117 (N_9117,N_8064,N_8311);
nand U9118 (N_9118,N_8556,N_8539);
and U9119 (N_9119,N_8373,N_8329);
or U9120 (N_9120,N_8238,N_8712);
or U9121 (N_9121,N_8478,N_8584);
nor U9122 (N_9122,N_8231,N_8190);
and U9123 (N_9123,N_8234,N_8435);
and U9124 (N_9124,N_8213,N_8799);
nor U9125 (N_9125,N_8285,N_8156);
nand U9126 (N_9126,N_8766,N_8633);
nand U9127 (N_9127,N_8557,N_8290);
nor U9128 (N_9128,N_8001,N_8447);
nand U9129 (N_9129,N_8023,N_8685);
nor U9130 (N_9130,N_8280,N_8525);
nand U9131 (N_9131,N_8679,N_8237);
xnor U9132 (N_9132,N_8115,N_8780);
or U9133 (N_9133,N_8010,N_8737);
nor U9134 (N_9134,N_8367,N_8437);
xnor U9135 (N_9135,N_8585,N_8795);
nand U9136 (N_9136,N_8394,N_8696);
nor U9137 (N_9137,N_8113,N_8535);
xnor U9138 (N_9138,N_8412,N_8520);
or U9139 (N_9139,N_8462,N_8669);
nand U9140 (N_9140,N_8040,N_8532);
xor U9141 (N_9141,N_8332,N_8101);
and U9142 (N_9142,N_8587,N_8673);
xor U9143 (N_9143,N_8778,N_8459);
nor U9144 (N_9144,N_8521,N_8668);
or U9145 (N_9145,N_8008,N_8069);
or U9146 (N_9146,N_8200,N_8163);
xnor U9147 (N_9147,N_8537,N_8694);
or U9148 (N_9148,N_8482,N_8116);
nand U9149 (N_9149,N_8219,N_8522);
nand U9150 (N_9150,N_8502,N_8707);
or U9151 (N_9151,N_8366,N_8038);
nor U9152 (N_9152,N_8541,N_8653);
nor U9153 (N_9153,N_8395,N_8606);
nor U9154 (N_9154,N_8475,N_8260);
and U9155 (N_9155,N_8649,N_8014);
or U9156 (N_9156,N_8125,N_8211);
nand U9157 (N_9157,N_8431,N_8241);
and U9158 (N_9158,N_8699,N_8041);
nor U9159 (N_9159,N_8139,N_8225);
nand U9160 (N_9160,N_8445,N_8291);
nor U9161 (N_9161,N_8741,N_8416);
xor U9162 (N_9162,N_8485,N_8355);
nor U9163 (N_9163,N_8583,N_8770);
or U9164 (N_9164,N_8088,N_8528);
or U9165 (N_9165,N_8410,N_8613);
nand U9166 (N_9166,N_8184,N_8453);
nor U9167 (N_9167,N_8263,N_8594);
nor U9168 (N_9168,N_8086,N_8470);
xor U9169 (N_9169,N_8065,N_8324);
nor U9170 (N_9170,N_8181,N_8564);
or U9171 (N_9171,N_8252,N_8120);
nand U9172 (N_9172,N_8507,N_8469);
and U9173 (N_9173,N_8325,N_8281);
nor U9174 (N_9174,N_8414,N_8510);
nand U9175 (N_9175,N_8177,N_8358);
nand U9176 (N_9176,N_8526,N_8691);
xor U9177 (N_9177,N_8215,N_8604);
or U9178 (N_9178,N_8687,N_8429);
nor U9179 (N_9179,N_8682,N_8310);
and U9180 (N_9180,N_8614,N_8153);
or U9181 (N_9181,N_8271,N_8404);
nand U9182 (N_9182,N_8095,N_8660);
nor U9183 (N_9183,N_8636,N_8359);
nor U9184 (N_9184,N_8309,N_8315);
and U9185 (N_9185,N_8257,N_8293);
xnor U9186 (N_9186,N_8262,N_8313);
xnor U9187 (N_9187,N_8131,N_8479);
and U9188 (N_9188,N_8642,N_8249);
nand U9189 (N_9189,N_8735,N_8629);
or U9190 (N_9190,N_8287,N_8259);
nand U9191 (N_9191,N_8350,N_8446);
xnor U9192 (N_9192,N_8098,N_8400);
nor U9193 (N_9193,N_8739,N_8589);
nor U9194 (N_9194,N_8689,N_8764);
or U9195 (N_9195,N_8721,N_8087);
nand U9196 (N_9196,N_8700,N_8108);
xnor U9197 (N_9197,N_8028,N_8364);
xor U9198 (N_9198,N_8461,N_8306);
nor U9199 (N_9199,N_8206,N_8103);
xor U9200 (N_9200,N_8038,N_8141);
xor U9201 (N_9201,N_8474,N_8083);
xor U9202 (N_9202,N_8678,N_8296);
nand U9203 (N_9203,N_8713,N_8409);
nand U9204 (N_9204,N_8415,N_8318);
nor U9205 (N_9205,N_8499,N_8779);
nand U9206 (N_9206,N_8377,N_8644);
xnor U9207 (N_9207,N_8614,N_8270);
xnor U9208 (N_9208,N_8455,N_8260);
nand U9209 (N_9209,N_8188,N_8482);
or U9210 (N_9210,N_8488,N_8580);
nand U9211 (N_9211,N_8742,N_8738);
and U9212 (N_9212,N_8188,N_8185);
or U9213 (N_9213,N_8299,N_8748);
and U9214 (N_9214,N_8008,N_8095);
or U9215 (N_9215,N_8196,N_8717);
nor U9216 (N_9216,N_8716,N_8267);
xnor U9217 (N_9217,N_8403,N_8467);
or U9218 (N_9218,N_8618,N_8666);
nor U9219 (N_9219,N_8091,N_8035);
xor U9220 (N_9220,N_8322,N_8011);
nand U9221 (N_9221,N_8198,N_8281);
and U9222 (N_9222,N_8616,N_8560);
and U9223 (N_9223,N_8113,N_8626);
nand U9224 (N_9224,N_8262,N_8689);
or U9225 (N_9225,N_8117,N_8711);
and U9226 (N_9226,N_8375,N_8640);
nand U9227 (N_9227,N_8457,N_8072);
or U9228 (N_9228,N_8608,N_8342);
nor U9229 (N_9229,N_8204,N_8189);
xnor U9230 (N_9230,N_8792,N_8514);
xor U9231 (N_9231,N_8347,N_8312);
and U9232 (N_9232,N_8613,N_8166);
or U9233 (N_9233,N_8402,N_8094);
or U9234 (N_9234,N_8262,N_8254);
xnor U9235 (N_9235,N_8350,N_8265);
xor U9236 (N_9236,N_8154,N_8414);
nand U9237 (N_9237,N_8577,N_8764);
and U9238 (N_9238,N_8256,N_8318);
xor U9239 (N_9239,N_8496,N_8102);
and U9240 (N_9240,N_8340,N_8105);
or U9241 (N_9241,N_8178,N_8124);
nand U9242 (N_9242,N_8344,N_8716);
or U9243 (N_9243,N_8111,N_8505);
xor U9244 (N_9244,N_8534,N_8509);
and U9245 (N_9245,N_8437,N_8073);
nand U9246 (N_9246,N_8542,N_8201);
or U9247 (N_9247,N_8252,N_8770);
or U9248 (N_9248,N_8422,N_8202);
or U9249 (N_9249,N_8424,N_8002);
or U9250 (N_9250,N_8257,N_8380);
and U9251 (N_9251,N_8097,N_8435);
nor U9252 (N_9252,N_8228,N_8446);
or U9253 (N_9253,N_8365,N_8777);
nand U9254 (N_9254,N_8705,N_8147);
nor U9255 (N_9255,N_8299,N_8625);
or U9256 (N_9256,N_8485,N_8500);
or U9257 (N_9257,N_8711,N_8732);
and U9258 (N_9258,N_8281,N_8137);
and U9259 (N_9259,N_8201,N_8054);
nor U9260 (N_9260,N_8188,N_8646);
xnor U9261 (N_9261,N_8672,N_8238);
or U9262 (N_9262,N_8139,N_8353);
xnor U9263 (N_9263,N_8111,N_8611);
nor U9264 (N_9264,N_8287,N_8302);
or U9265 (N_9265,N_8732,N_8799);
or U9266 (N_9266,N_8050,N_8170);
xor U9267 (N_9267,N_8543,N_8080);
and U9268 (N_9268,N_8351,N_8246);
xnor U9269 (N_9269,N_8422,N_8046);
or U9270 (N_9270,N_8012,N_8172);
xor U9271 (N_9271,N_8367,N_8760);
nand U9272 (N_9272,N_8010,N_8766);
and U9273 (N_9273,N_8035,N_8405);
nand U9274 (N_9274,N_8689,N_8558);
nand U9275 (N_9275,N_8543,N_8099);
nand U9276 (N_9276,N_8467,N_8670);
or U9277 (N_9277,N_8334,N_8184);
nand U9278 (N_9278,N_8192,N_8476);
or U9279 (N_9279,N_8554,N_8363);
or U9280 (N_9280,N_8110,N_8532);
or U9281 (N_9281,N_8348,N_8138);
or U9282 (N_9282,N_8349,N_8025);
nand U9283 (N_9283,N_8617,N_8133);
nand U9284 (N_9284,N_8727,N_8044);
or U9285 (N_9285,N_8125,N_8464);
nor U9286 (N_9286,N_8737,N_8114);
nand U9287 (N_9287,N_8163,N_8136);
or U9288 (N_9288,N_8054,N_8037);
nand U9289 (N_9289,N_8411,N_8147);
nor U9290 (N_9290,N_8689,N_8125);
nand U9291 (N_9291,N_8489,N_8279);
nand U9292 (N_9292,N_8466,N_8352);
nand U9293 (N_9293,N_8151,N_8058);
nor U9294 (N_9294,N_8746,N_8024);
and U9295 (N_9295,N_8411,N_8193);
and U9296 (N_9296,N_8399,N_8454);
xnor U9297 (N_9297,N_8008,N_8347);
nor U9298 (N_9298,N_8210,N_8764);
xnor U9299 (N_9299,N_8628,N_8106);
and U9300 (N_9300,N_8519,N_8463);
and U9301 (N_9301,N_8245,N_8070);
nor U9302 (N_9302,N_8131,N_8750);
nand U9303 (N_9303,N_8316,N_8378);
xnor U9304 (N_9304,N_8502,N_8630);
nand U9305 (N_9305,N_8476,N_8665);
nor U9306 (N_9306,N_8105,N_8007);
or U9307 (N_9307,N_8563,N_8542);
or U9308 (N_9308,N_8033,N_8642);
nor U9309 (N_9309,N_8178,N_8404);
and U9310 (N_9310,N_8276,N_8733);
nand U9311 (N_9311,N_8218,N_8025);
or U9312 (N_9312,N_8267,N_8288);
xnor U9313 (N_9313,N_8066,N_8515);
and U9314 (N_9314,N_8189,N_8611);
and U9315 (N_9315,N_8358,N_8001);
xor U9316 (N_9316,N_8717,N_8688);
nand U9317 (N_9317,N_8392,N_8163);
or U9318 (N_9318,N_8413,N_8280);
nand U9319 (N_9319,N_8730,N_8004);
nor U9320 (N_9320,N_8006,N_8587);
and U9321 (N_9321,N_8488,N_8316);
nand U9322 (N_9322,N_8003,N_8121);
nor U9323 (N_9323,N_8335,N_8534);
xnor U9324 (N_9324,N_8114,N_8321);
xor U9325 (N_9325,N_8248,N_8122);
or U9326 (N_9326,N_8395,N_8490);
xor U9327 (N_9327,N_8654,N_8308);
and U9328 (N_9328,N_8457,N_8143);
or U9329 (N_9329,N_8439,N_8557);
or U9330 (N_9330,N_8381,N_8657);
nand U9331 (N_9331,N_8163,N_8345);
and U9332 (N_9332,N_8532,N_8588);
nor U9333 (N_9333,N_8728,N_8631);
nor U9334 (N_9334,N_8749,N_8487);
nor U9335 (N_9335,N_8199,N_8046);
and U9336 (N_9336,N_8643,N_8186);
or U9337 (N_9337,N_8197,N_8467);
xor U9338 (N_9338,N_8321,N_8536);
and U9339 (N_9339,N_8620,N_8783);
nor U9340 (N_9340,N_8146,N_8399);
or U9341 (N_9341,N_8383,N_8125);
xor U9342 (N_9342,N_8760,N_8084);
nand U9343 (N_9343,N_8664,N_8568);
or U9344 (N_9344,N_8301,N_8105);
or U9345 (N_9345,N_8241,N_8231);
and U9346 (N_9346,N_8122,N_8253);
and U9347 (N_9347,N_8615,N_8208);
or U9348 (N_9348,N_8655,N_8785);
and U9349 (N_9349,N_8182,N_8419);
nand U9350 (N_9350,N_8389,N_8757);
or U9351 (N_9351,N_8274,N_8358);
and U9352 (N_9352,N_8387,N_8385);
xor U9353 (N_9353,N_8424,N_8020);
xnor U9354 (N_9354,N_8707,N_8376);
xnor U9355 (N_9355,N_8695,N_8175);
nor U9356 (N_9356,N_8365,N_8610);
and U9357 (N_9357,N_8459,N_8445);
or U9358 (N_9358,N_8747,N_8397);
nand U9359 (N_9359,N_8194,N_8263);
xor U9360 (N_9360,N_8255,N_8746);
nand U9361 (N_9361,N_8395,N_8188);
and U9362 (N_9362,N_8579,N_8533);
nand U9363 (N_9363,N_8178,N_8752);
and U9364 (N_9364,N_8448,N_8019);
and U9365 (N_9365,N_8233,N_8301);
xnor U9366 (N_9366,N_8275,N_8241);
or U9367 (N_9367,N_8052,N_8284);
nand U9368 (N_9368,N_8116,N_8144);
nand U9369 (N_9369,N_8053,N_8249);
or U9370 (N_9370,N_8341,N_8291);
or U9371 (N_9371,N_8125,N_8175);
xor U9372 (N_9372,N_8692,N_8205);
nand U9373 (N_9373,N_8522,N_8411);
nor U9374 (N_9374,N_8389,N_8790);
nand U9375 (N_9375,N_8158,N_8767);
and U9376 (N_9376,N_8111,N_8571);
nand U9377 (N_9377,N_8288,N_8285);
and U9378 (N_9378,N_8491,N_8057);
xor U9379 (N_9379,N_8767,N_8530);
xnor U9380 (N_9380,N_8014,N_8239);
nand U9381 (N_9381,N_8550,N_8591);
and U9382 (N_9382,N_8467,N_8444);
or U9383 (N_9383,N_8463,N_8484);
nand U9384 (N_9384,N_8242,N_8116);
nor U9385 (N_9385,N_8795,N_8409);
or U9386 (N_9386,N_8274,N_8009);
or U9387 (N_9387,N_8576,N_8056);
nor U9388 (N_9388,N_8023,N_8455);
nand U9389 (N_9389,N_8660,N_8601);
xnor U9390 (N_9390,N_8699,N_8001);
xnor U9391 (N_9391,N_8025,N_8405);
nand U9392 (N_9392,N_8637,N_8265);
nand U9393 (N_9393,N_8042,N_8373);
nor U9394 (N_9394,N_8235,N_8195);
xor U9395 (N_9395,N_8634,N_8053);
nand U9396 (N_9396,N_8425,N_8199);
nand U9397 (N_9397,N_8127,N_8353);
nand U9398 (N_9398,N_8518,N_8581);
and U9399 (N_9399,N_8143,N_8240);
or U9400 (N_9400,N_8302,N_8662);
nand U9401 (N_9401,N_8315,N_8266);
xor U9402 (N_9402,N_8285,N_8275);
nor U9403 (N_9403,N_8188,N_8469);
xnor U9404 (N_9404,N_8028,N_8189);
nor U9405 (N_9405,N_8594,N_8324);
xnor U9406 (N_9406,N_8356,N_8010);
and U9407 (N_9407,N_8063,N_8414);
or U9408 (N_9408,N_8223,N_8573);
nand U9409 (N_9409,N_8734,N_8446);
xnor U9410 (N_9410,N_8300,N_8132);
nand U9411 (N_9411,N_8529,N_8415);
xnor U9412 (N_9412,N_8639,N_8602);
nor U9413 (N_9413,N_8708,N_8030);
nor U9414 (N_9414,N_8154,N_8159);
xor U9415 (N_9415,N_8296,N_8161);
nor U9416 (N_9416,N_8778,N_8456);
and U9417 (N_9417,N_8440,N_8420);
xnor U9418 (N_9418,N_8500,N_8229);
or U9419 (N_9419,N_8515,N_8443);
xor U9420 (N_9420,N_8111,N_8520);
or U9421 (N_9421,N_8774,N_8147);
or U9422 (N_9422,N_8728,N_8457);
nor U9423 (N_9423,N_8664,N_8374);
nor U9424 (N_9424,N_8112,N_8565);
nor U9425 (N_9425,N_8680,N_8246);
nand U9426 (N_9426,N_8603,N_8023);
nor U9427 (N_9427,N_8297,N_8727);
xor U9428 (N_9428,N_8022,N_8428);
nor U9429 (N_9429,N_8260,N_8106);
xor U9430 (N_9430,N_8281,N_8317);
nor U9431 (N_9431,N_8720,N_8209);
or U9432 (N_9432,N_8249,N_8275);
xnor U9433 (N_9433,N_8715,N_8438);
xnor U9434 (N_9434,N_8559,N_8707);
nand U9435 (N_9435,N_8005,N_8038);
or U9436 (N_9436,N_8556,N_8193);
xor U9437 (N_9437,N_8440,N_8334);
xor U9438 (N_9438,N_8464,N_8161);
xnor U9439 (N_9439,N_8197,N_8570);
xor U9440 (N_9440,N_8327,N_8367);
nor U9441 (N_9441,N_8469,N_8040);
and U9442 (N_9442,N_8605,N_8669);
nor U9443 (N_9443,N_8746,N_8206);
or U9444 (N_9444,N_8243,N_8314);
and U9445 (N_9445,N_8525,N_8570);
or U9446 (N_9446,N_8142,N_8182);
or U9447 (N_9447,N_8488,N_8624);
and U9448 (N_9448,N_8766,N_8738);
or U9449 (N_9449,N_8263,N_8756);
nand U9450 (N_9450,N_8193,N_8543);
and U9451 (N_9451,N_8009,N_8266);
and U9452 (N_9452,N_8686,N_8195);
nand U9453 (N_9453,N_8153,N_8187);
and U9454 (N_9454,N_8125,N_8629);
and U9455 (N_9455,N_8732,N_8008);
xnor U9456 (N_9456,N_8383,N_8007);
xor U9457 (N_9457,N_8213,N_8176);
nand U9458 (N_9458,N_8664,N_8382);
nand U9459 (N_9459,N_8599,N_8439);
nor U9460 (N_9460,N_8446,N_8406);
and U9461 (N_9461,N_8600,N_8790);
nor U9462 (N_9462,N_8081,N_8672);
nand U9463 (N_9463,N_8435,N_8703);
or U9464 (N_9464,N_8080,N_8644);
nand U9465 (N_9465,N_8277,N_8160);
and U9466 (N_9466,N_8549,N_8026);
nand U9467 (N_9467,N_8164,N_8386);
nand U9468 (N_9468,N_8743,N_8026);
and U9469 (N_9469,N_8164,N_8393);
and U9470 (N_9470,N_8674,N_8639);
nand U9471 (N_9471,N_8450,N_8624);
nand U9472 (N_9472,N_8485,N_8371);
xnor U9473 (N_9473,N_8313,N_8132);
nor U9474 (N_9474,N_8435,N_8131);
and U9475 (N_9475,N_8387,N_8740);
or U9476 (N_9476,N_8644,N_8122);
xnor U9477 (N_9477,N_8788,N_8577);
nand U9478 (N_9478,N_8530,N_8079);
xor U9479 (N_9479,N_8550,N_8398);
or U9480 (N_9480,N_8740,N_8777);
nand U9481 (N_9481,N_8373,N_8413);
and U9482 (N_9482,N_8662,N_8660);
or U9483 (N_9483,N_8243,N_8781);
nor U9484 (N_9484,N_8640,N_8042);
or U9485 (N_9485,N_8562,N_8560);
or U9486 (N_9486,N_8768,N_8321);
or U9487 (N_9487,N_8461,N_8571);
xnor U9488 (N_9488,N_8641,N_8556);
nor U9489 (N_9489,N_8123,N_8464);
nor U9490 (N_9490,N_8774,N_8564);
and U9491 (N_9491,N_8312,N_8023);
nand U9492 (N_9492,N_8611,N_8640);
nor U9493 (N_9493,N_8733,N_8234);
or U9494 (N_9494,N_8412,N_8241);
nor U9495 (N_9495,N_8158,N_8075);
or U9496 (N_9496,N_8149,N_8517);
or U9497 (N_9497,N_8551,N_8289);
or U9498 (N_9498,N_8786,N_8418);
nor U9499 (N_9499,N_8436,N_8740);
or U9500 (N_9500,N_8120,N_8038);
nor U9501 (N_9501,N_8192,N_8715);
or U9502 (N_9502,N_8050,N_8435);
or U9503 (N_9503,N_8653,N_8531);
nand U9504 (N_9504,N_8014,N_8269);
and U9505 (N_9505,N_8048,N_8266);
nand U9506 (N_9506,N_8787,N_8382);
nor U9507 (N_9507,N_8708,N_8665);
or U9508 (N_9508,N_8277,N_8327);
nand U9509 (N_9509,N_8031,N_8131);
nor U9510 (N_9510,N_8457,N_8721);
nor U9511 (N_9511,N_8241,N_8398);
and U9512 (N_9512,N_8678,N_8451);
nor U9513 (N_9513,N_8229,N_8218);
xnor U9514 (N_9514,N_8219,N_8300);
xnor U9515 (N_9515,N_8768,N_8133);
xnor U9516 (N_9516,N_8046,N_8659);
nor U9517 (N_9517,N_8213,N_8511);
xor U9518 (N_9518,N_8331,N_8732);
nand U9519 (N_9519,N_8132,N_8713);
nand U9520 (N_9520,N_8755,N_8489);
nor U9521 (N_9521,N_8057,N_8372);
or U9522 (N_9522,N_8585,N_8376);
xor U9523 (N_9523,N_8513,N_8146);
or U9524 (N_9524,N_8472,N_8780);
nor U9525 (N_9525,N_8418,N_8057);
xor U9526 (N_9526,N_8579,N_8274);
and U9527 (N_9527,N_8628,N_8329);
or U9528 (N_9528,N_8116,N_8796);
nor U9529 (N_9529,N_8752,N_8268);
xnor U9530 (N_9530,N_8287,N_8345);
xnor U9531 (N_9531,N_8010,N_8424);
or U9532 (N_9532,N_8169,N_8364);
nor U9533 (N_9533,N_8167,N_8052);
xor U9534 (N_9534,N_8373,N_8122);
and U9535 (N_9535,N_8057,N_8370);
or U9536 (N_9536,N_8158,N_8288);
or U9537 (N_9537,N_8323,N_8438);
or U9538 (N_9538,N_8034,N_8504);
and U9539 (N_9539,N_8061,N_8050);
xor U9540 (N_9540,N_8066,N_8728);
nand U9541 (N_9541,N_8208,N_8720);
nand U9542 (N_9542,N_8143,N_8376);
or U9543 (N_9543,N_8590,N_8685);
nor U9544 (N_9544,N_8496,N_8687);
or U9545 (N_9545,N_8108,N_8777);
nor U9546 (N_9546,N_8650,N_8224);
and U9547 (N_9547,N_8047,N_8255);
nor U9548 (N_9548,N_8597,N_8057);
nor U9549 (N_9549,N_8144,N_8027);
and U9550 (N_9550,N_8651,N_8183);
or U9551 (N_9551,N_8057,N_8391);
or U9552 (N_9552,N_8096,N_8484);
nand U9553 (N_9553,N_8679,N_8245);
and U9554 (N_9554,N_8703,N_8584);
nor U9555 (N_9555,N_8469,N_8356);
and U9556 (N_9556,N_8384,N_8584);
or U9557 (N_9557,N_8502,N_8263);
and U9558 (N_9558,N_8272,N_8537);
xnor U9559 (N_9559,N_8785,N_8231);
nor U9560 (N_9560,N_8136,N_8614);
nand U9561 (N_9561,N_8368,N_8044);
nand U9562 (N_9562,N_8653,N_8650);
or U9563 (N_9563,N_8317,N_8129);
and U9564 (N_9564,N_8511,N_8158);
nand U9565 (N_9565,N_8632,N_8304);
nand U9566 (N_9566,N_8181,N_8719);
nand U9567 (N_9567,N_8172,N_8730);
nand U9568 (N_9568,N_8452,N_8110);
nand U9569 (N_9569,N_8087,N_8283);
or U9570 (N_9570,N_8697,N_8039);
xnor U9571 (N_9571,N_8021,N_8712);
and U9572 (N_9572,N_8704,N_8548);
nand U9573 (N_9573,N_8293,N_8371);
xnor U9574 (N_9574,N_8397,N_8177);
xor U9575 (N_9575,N_8541,N_8432);
nand U9576 (N_9576,N_8532,N_8315);
nor U9577 (N_9577,N_8545,N_8717);
xor U9578 (N_9578,N_8180,N_8116);
and U9579 (N_9579,N_8027,N_8747);
and U9580 (N_9580,N_8749,N_8748);
nor U9581 (N_9581,N_8225,N_8647);
nand U9582 (N_9582,N_8285,N_8284);
or U9583 (N_9583,N_8578,N_8342);
xnor U9584 (N_9584,N_8770,N_8595);
nand U9585 (N_9585,N_8484,N_8143);
and U9586 (N_9586,N_8738,N_8691);
or U9587 (N_9587,N_8373,N_8187);
nand U9588 (N_9588,N_8336,N_8354);
or U9589 (N_9589,N_8304,N_8669);
nor U9590 (N_9590,N_8598,N_8372);
nor U9591 (N_9591,N_8673,N_8448);
and U9592 (N_9592,N_8730,N_8106);
xnor U9593 (N_9593,N_8748,N_8226);
xor U9594 (N_9594,N_8109,N_8550);
xor U9595 (N_9595,N_8347,N_8599);
or U9596 (N_9596,N_8759,N_8385);
xor U9597 (N_9597,N_8368,N_8118);
and U9598 (N_9598,N_8125,N_8050);
nor U9599 (N_9599,N_8667,N_8093);
and U9600 (N_9600,N_9195,N_9024);
nand U9601 (N_9601,N_9181,N_8904);
nand U9602 (N_9602,N_9049,N_9440);
or U9603 (N_9603,N_8802,N_9113);
xor U9604 (N_9604,N_9055,N_9586);
nor U9605 (N_9605,N_9006,N_9079);
xnor U9606 (N_9606,N_9474,N_8987);
nand U9607 (N_9607,N_8846,N_9438);
nand U9608 (N_9608,N_9585,N_8880);
xnor U9609 (N_9609,N_9408,N_8874);
nor U9610 (N_9610,N_9485,N_9383);
nor U9611 (N_9611,N_8868,N_9421);
and U9612 (N_9612,N_9223,N_9483);
nor U9613 (N_9613,N_9159,N_8841);
and U9614 (N_9614,N_9380,N_9269);
nand U9615 (N_9615,N_9236,N_9266);
xnor U9616 (N_9616,N_9022,N_8918);
and U9617 (N_9617,N_9444,N_9522);
or U9618 (N_9618,N_9233,N_9414);
nand U9619 (N_9619,N_9176,N_9561);
nor U9620 (N_9620,N_9240,N_9381);
and U9621 (N_9621,N_9134,N_8915);
and U9622 (N_9622,N_9000,N_9589);
or U9623 (N_9623,N_9241,N_9156);
or U9624 (N_9624,N_8952,N_9477);
nor U9625 (N_9625,N_8875,N_9274);
nor U9626 (N_9626,N_9467,N_9143);
or U9627 (N_9627,N_8825,N_9324);
nor U9628 (N_9628,N_9168,N_8819);
and U9629 (N_9629,N_9307,N_8803);
xnor U9630 (N_9630,N_8873,N_9573);
or U9631 (N_9631,N_9546,N_8964);
or U9632 (N_9632,N_9178,N_9219);
nor U9633 (N_9633,N_9212,N_9460);
or U9634 (N_9634,N_9132,N_8940);
nor U9635 (N_9635,N_9457,N_9061);
and U9636 (N_9636,N_9203,N_9123);
nor U9637 (N_9637,N_9098,N_9217);
and U9638 (N_9638,N_9101,N_9478);
nand U9639 (N_9639,N_9594,N_9391);
nand U9640 (N_9640,N_9596,N_8845);
nand U9641 (N_9641,N_9074,N_9465);
xor U9642 (N_9642,N_8948,N_8833);
xnor U9643 (N_9643,N_9069,N_9202);
and U9644 (N_9644,N_9013,N_8807);
nand U9645 (N_9645,N_9363,N_9025);
and U9646 (N_9646,N_8937,N_9128);
nand U9647 (N_9647,N_8859,N_9067);
nand U9648 (N_9648,N_9503,N_8954);
nand U9649 (N_9649,N_9557,N_9141);
xnor U9650 (N_9650,N_9031,N_8823);
nor U9651 (N_9651,N_8889,N_9336);
or U9652 (N_9652,N_9301,N_9063);
or U9653 (N_9653,N_8929,N_9384);
xnor U9654 (N_9654,N_9375,N_9255);
and U9655 (N_9655,N_9293,N_9590);
xor U9656 (N_9656,N_8913,N_9313);
and U9657 (N_9657,N_9342,N_9286);
nand U9658 (N_9658,N_9220,N_9295);
nand U9659 (N_9659,N_9348,N_9114);
nor U9660 (N_9660,N_9442,N_8884);
nor U9661 (N_9661,N_8977,N_9533);
xnor U9662 (N_9662,N_8998,N_9326);
nand U9663 (N_9663,N_9282,N_9524);
nand U9664 (N_9664,N_9536,N_9158);
xnor U9665 (N_9665,N_9185,N_9062);
nor U9666 (N_9666,N_9012,N_9040);
nor U9667 (N_9667,N_9229,N_9396);
and U9668 (N_9668,N_9280,N_9214);
nor U9669 (N_9669,N_8957,N_9518);
nor U9670 (N_9670,N_9039,N_9463);
xor U9671 (N_9671,N_8848,N_9193);
nor U9672 (N_9672,N_8941,N_8864);
and U9673 (N_9673,N_9058,N_9379);
and U9674 (N_9674,N_9126,N_9435);
and U9675 (N_9675,N_9505,N_8982);
nand U9676 (N_9676,N_9172,N_9002);
nand U9677 (N_9677,N_9528,N_8914);
nor U9678 (N_9678,N_9105,N_9497);
xor U9679 (N_9679,N_9060,N_9455);
nand U9680 (N_9680,N_9535,N_9526);
nand U9681 (N_9681,N_9411,N_8800);
xor U9682 (N_9682,N_8966,N_8903);
nand U9683 (N_9683,N_9323,N_9499);
xnor U9684 (N_9684,N_9345,N_9500);
xnor U9685 (N_9685,N_9088,N_9388);
or U9686 (N_9686,N_9034,N_9166);
nor U9687 (N_9687,N_9433,N_9579);
xor U9688 (N_9688,N_9086,N_9139);
nor U9689 (N_9689,N_8951,N_9028);
nand U9690 (N_9690,N_9510,N_8978);
and U9691 (N_9691,N_9409,N_9205);
and U9692 (N_9692,N_8986,N_9151);
nor U9693 (N_9693,N_8801,N_8894);
and U9694 (N_9694,N_8924,N_9097);
or U9695 (N_9695,N_9210,N_8973);
nand U9696 (N_9696,N_8962,N_9109);
and U9697 (N_9697,N_9155,N_9486);
and U9698 (N_9698,N_9304,N_9213);
and U9699 (N_9699,N_9118,N_9564);
nand U9700 (N_9700,N_8971,N_9093);
and U9701 (N_9701,N_8896,N_9057);
or U9702 (N_9702,N_8900,N_8916);
xor U9703 (N_9703,N_9595,N_9350);
nand U9704 (N_9704,N_9072,N_8806);
nand U9705 (N_9705,N_9417,N_9130);
nor U9706 (N_9706,N_8999,N_9529);
xor U9707 (N_9707,N_8810,N_9360);
xor U9708 (N_9708,N_9198,N_9534);
and U9709 (N_9709,N_9489,N_9145);
nor U9710 (N_9710,N_9111,N_8863);
or U9711 (N_9711,N_9264,N_9581);
nand U9712 (N_9712,N_9027,N_9218);
xor U9713 (N_9713,N_8994,N_9310);
xnor U9714 (N_9714,N_9305,N_8910);
nand U9715 (N_9715,N_9265,N_9466);
nand U9716 (N_9716,N_9085,N_9201);
nor U9717 (N_9717,N_9196,N_9038);
nor U9718 (N_9718,N_8840,N_8947);
and U9719 (N_9719,N_9019,N_9247);
nand U9720 (N_9720,N_9095,N_9144);
nand U9721 (N_9721,N_9279,N_9129);
and U9722 (N_9722,N_9131,N_9285);
and U9723 (N_9723,N_9258,N_9387);
nand U9724 (N_9724,N_8967,N_8821);
nand U9725 (N_9725,N_9583,N_9014);
xor U9726 (N_9726,N_9587,N_9456);
or U9727 (N_9727,N_9330,N_9081);
and U9728 (N_9728,N_9556,N_9221);
xnor U9729 (N_9729,N_9507,N_9385);
xor U9730 (N_9730,N_9402,N_9254);
and U9731 (N_9731,N_9570,N_9325);
nor U9732 (N_9732,N_9354,N_9333);
nor U9733 (N_9733,N_9200,N_9481);
and U9734 (N_9734,N_9356,N_9044);
nand U9735 (N_9735,N_9480,N_8991);
nor U9736 (N_9736,N_9392,N_9576);
xor U9737 (N_9737,N_9394,N_9580);
xnor U9738 (N_9738,N_9395,N_9540);
and U9739 (N_9739,N_9338,N_8939);
nor U9740 (N_9740,N_9412,N_9023);
nand U9741 (N_9741,N_9242,N_9487);
xnor U9742 (N_9742,N_9119,N_9543);
nand U9743 (N_9743,N_9368,N_9152);
and U9744 (N_9744,N_9125,N_9035);
or U9745 (N_9745,N_9506,N_9501);
and U9746 (N_9746,N_8905,N_9386);
and U9747 (N_9747,N_9406,N_8891);
and U9748 (N_9748,N_9239,N_8839);
and U9749 (N_9749,N_8887,N_9413);
xnor U9750 (N_9750,N_9108,N_8876);
and U9751 (N_9751,N_9458,N_9448);
xnor U9752 (N_9752,N_9271,N_9050);
or U9753 (N_9753,N_9186,N_8942);
or U9754 (N_9754,N_9020,N_9558);
xnor U9755 (N_9755,N_9206,N_9592);
xnor U9756 (N_9756,N_9291,N_8861);
xor U9757 (N_9757,N_8844,N_9078);
xor U9758 (N_9758,N_9267,N_8809);
xnor U9759 (N_9759,N_8968,N_9547);
and U9760 (N_9760,N_9127,N_9296);
or U9761 (N_9761,N_9192,N_9041);
nand U9762 (N_9762,N_8981,N_9142);
or U9763 (N_9763,N_8926,N_9364);
or U9764 (N_9764,N_9454,N_9230);
nor U9765 (N_9765,N_9281,N_9495);
or U9766 (N_9766,N_9250,N_8992);
or U9767 (N_9767,N_9490,N_9288);
xnor U9768 (N_9768,N_9297,N_9378);
nand U9769 (N_9769,N_9173,N_8829);
and U9770 (N_9770,N_9115,N_9033);
nor U9771 (N_9771,N_9398,N_9588);
xor U9772 (N_9772,N_9523,N_9316);
nand U9773 (N_9773,N_9312,N_9099);
xnor U9774 (N_9774,N_8933,N_9445);
nor U9775 (N_9775,N_9116,N_9425);
nor U9776 (N_9776,N_9542,N_9393);
or U9777 (N_9777,N_8972,N_9094);
xnor U9778 (N_9778,N_9447,N_9512);
nand U9779 (N_9779,N_8808,N_9479);
xnor U9780 (N_9780,N_9270,N_8858);
nor U9781 (N_9781,N_8883,N_8920);
or U9782 (N_9782,N_9147,N_8925);
and U9783 (N_9783,N_9426,N_9539);
xor U9784 (N_9784,N_9550,N_9459);
nor U9785 (N_9785,N_8826,N_9009);
and U9786 (N_9786,N_9418,N_8974);
nor U9787 (N_9787,N_9369,N_9494);
or U9788 (N_9788,N_9331,N_9177);
xnor U9789 (N_9789,N_8976,N_9311);
or U9790 (N_9790,N_9298,N_8836);
nor U9791 (N_9791,N_9184,N_9578);
xor U9792 (N_9792,N_9308,N_9337);
nand U9793 (N_9793,N_9416,N_9424);
and U9794 (N_9794,N_8958,N_8984);
or U9795 (N_9795,N_9401,N_8907);
or U9796 (N_9796,N_8953,N_9092);
and U9797 (N_9797,N_9183,N_9136);
and U9798 (N_9798,N_9502,N_9294);
nor U9799 (N_9799,N_9260,N_8838);
and U9800 (N_9800,N_9215,N_9243);
nor U9801 (N_9801,N_9498,N_9372);
or U9802 (N_9802,N_9366,N_8908);
xnor U9803 (N_9803,N_8847,N_9005);
xnor U9804 (N_9804,N_8854,N_8862);
and U9805 (N_9805,N_8934,N_8855);
and U9806 (N_9806,N_8969,N_9030);
and U9807 (N_9807,N_9001,N_8816);
and U9808 (N_9808,N_9376,N_9228);
nor U9809 (N_9809,N_9080,N_9190);
xnor U9810 (N_9810,N_9521,N_9249);
nor U9811 (N_9811,N_9231,N_9511);
or U9812 (N_9812,N_8831,N_9537);
and U9813 (N_9813,N_8919,N_9516);
xor U9814 (N_9814,N_9517,N_9509);
nor U9815 (N_9815,N_9315,N_9021);
nor U9816 (N_9816,N_9328,N_9056);
nor U9817 (N_9817,N_9225,N_9572);
nor U9818 (N_9818,N_8830,N_9370);
nor U9819 (N_9819,N_9450,N_9299);
nand U9820 (N_9820,N_9272,N_9224);
nor U9821 (N_9821,N_9591,N_9344);
or U9822 (N_9822,N_9167,N_9397);
and U9823 (N_9823,N_9322,N_9493);
or U9824 (N_9824,N_9046,N_8851);
or U9825 (N_9825,N_9303,N_9248);
and U9826 (N_9826,N_9154,N_9508);
or U9827 (N_9827,N_9026,N_9194);
or U9828 (N_9828,N_9551,N_8818);
nand U9829 (N_9829,N_8866,N_9513);
and U9830 (N_9830,N_9365,N_9153);
nand U9831 (N_9831,N_8956,N_9209);
xor U9832 (N_9832,N_9262,N_9064);
xor U9833 (N_9833,N_9263,N_9289);
xor U9834 (N_9834,N_8997,N_8965);
and U9835 (N_9835,N_9347,N_9472);
or U9836 (N_9836,N_9106,N_9571);
or U9837 (N_9837,N_9133,N_9436);
xnor U9838 (N_9838,N_9016,N_9410);
nor U9839 (N_9839,N_9527,N_9598);
nor U9840 (N_9840,N_8850,N_9355);
nor U9841 (N_9841,N_9584,N_8817);
or U9842 (N_9842,N_9037,N_9562);
xor U9843 (N_9843,N_8882,N_9091);
nor U9844 (N_9844,N_9150,N_9407);
and U9845 (N_9845,N_8945,N_9259);
nand U9846 (N_9846,N_9124,N_9273);
nor U9847 (N_9847,N_9237,N_8881);
xor U9848 (N_9848,N_9138,N_9011);
nor U9849 (N_9849,N_9276,N_8944);
and U9850 (N_9850,N_8814,N_9346);
nand U9851 (N_9851,N_8820,N_9268);
nand U9852 (N_9852,N_8867,N_9162);
nor U9853 (N_9853,N_8988,N_9554);
xnor U9854 (N_9854,N_9373,N_9430);
nand U9855 (N_9855,N_9525,N_9068);
nand U9856 (N_9856,N_9103,N_9319);
nor U9857 (N_9857,N_8897,N_8832);
and U9858 (N_9858,N_9422,N_9340);
xor U9859 (N_9859,N_8901,N_8856);
or U9860 (N_9860,N_8813,N_9100);
xnor U9861 (N_9861,N_8824,N_8950);
nor U9862 (N_9862,N_9565,N_9222);
and U9863 (N_9863,N_9358,N_9469);
and U9864 (N_9864,N_8885,N_9389);
nand U9865 (N_9865,N_9441,N_9188);
xor U9866 (N_9866,N_9290,N_8921);
nor U9867 (N_9867,N_9071,N_9110);
nand U9868 (N_9868,N_9429,N_9275);
and U9869 (N_9869,N_8995,N_9569);
xnor U9870 (N_9870,N_9320,N_9112);
and U9871 (N_9871,N_8980,N_9053);
nor U9872 (N_9872,N_8834,N_9318);
or U9873 (N_9873,N_8928,N_9082);
nand U9874 (N_9874,N_9419,N_9208);
nor U9875 (N_9875,N_8996,N_9334);
and U9876 (N_9876,N_8959,N_8828);
nor U9877 (N_9877,N_9087,N_9059);
and U9878 (N_9878,N_9382,N_9191);
and U9879 (N_9879,N_8892,N_8983);
and U9880 (N_9880,N_9548,N_9399);
and U9881 (N_9881,N_9568,N_9287);
and U9882 (N_9882,N_8890,N_9488);
xnor U9883 (N_9883,N_9361,N_8842);
nor U9884 (N_9884,N_8812,N_9300);
and U9885 (N_9885,N_8877,N_8975);
or U9886 (N_9886,N_9054,N_8849);
nor U9887 (N_9887,N_9452,N_9090);
or U9888 (N_9888,N_9245,N_9470);
nor U9889 (N_9889,N_9453,N_8899);
xnor U9890 (N_9890,N_9427,N_9476);
nor U9891 (N_9891,N_9292,N_9471);
and U9892 (N_9892,N_9560,N_9314);
or U9893 (N_9893,N_8865,N_9149);
xnor U9894 (N_9894,N_9544,N_9434);
xnor U9895 (N_9895,N_9261,N_9165);
and U9896 (N_9896,N_8960,N_9371);
xor U9897 (N_9897,N_9317,N_8804);
nand U9898 (N_9898,N_8938,N_9032);
nand U9899 (N_9899,N_9096,N_8805);
xor U9900 (N_9900,N_9135,N_9335);
and U9901 (N_9901,N_9423,N_9104);
nand U9902 (N_9902,N_9179,N_9042);
and U9903 (N_9903,N_8931,N_8946);
xnor U9904 (N_9904,N_8888,N_9439);
or U9905 (N_9905,N_9070,N_9420);
nor U9906 (N_9906,N_8879,N_9257);
and U9907 (N_9907,N_9309,N_9107);
nor U9908 (N_9908,N_9048,N_9357);
or U9909 (N_9909,N_9514,N_9244);
or U9910 (N_9910,N_9246,N_9226);
nand U9911 (N_9911,N_9353,N_9567);
xnor U9912 (N_9912,N_9204,N_9321);
or U9913 (N_9913,N_9238,N_9004);
or U9914 (N_9914,N_8886,N_8811);
xnor U9915 (N_9915,N_9066,N_9052);
xor U9916 (N_9916,N_9122,N_9446);
and U9917 (N_9917,N_9462,N_9515);
and U9918 (N_9918,N_9146,N_9169);
xnor U9919 (N_9919,N_8930,N_8815);
xnor U9920 (N_9920,N_9157,N_9216);
and U9921 (N_9921,N_9075,N_8963);
xor U9922 (N_9922,N_9349,N_8970);
or U9923 (N_9923,N_9065,N_9390);
xnor U9924 (N_9924,N_9083,N_9161);
nand U9925 (N_9925,N_9302,N_9283);
nand U9926 (N_9926,N_9199,N_8932);
xor U9927 (N_9927,N_9120,N_9415);
and U9928 (N_9928,N_9227,N_9076);
nor U9929 (N_9929,N_9329,N_9464);
xnor U9930 (N_9930,N_9140,N_9545);
nand U9931 (N_9931,N_9180,N_9211);
nand U9932 (N_9932,N_9174,N_9374);
nor U9933 (N_9933,N_8989,N_8902);
nand U9934 (N_9934,N_9148,N_9563);
or U9935 (N_9935,N_9451,N_9284);
nand U9936 (N_9936,N_9182,N_9232);
nor U9937 (N_9937,N_8922,N_9170);
nand U9938 (N_9938,N_9532,N_9377);
and U9939 (N_9939,N_8835,N_9339);
nand U9940 (N_9940,N_9117,N_8852);
and U9941 (N_9941,N_9582,N_9043);
and U9942 (N_9942,N_8990,N_8917);
xor U9943 (N_9943,N_9473,N_8827);
nor U9944 (N_9944,N_9362,N_8911);
xor U9945 (N_9945,N_9504,N_9010);
nor U9946 (N_9946,N_9530,N_8871);
and U9947 (N_9947,N_9553,N_9278);
xor U9948 (N_9948,N_8893,N_9443);
or U9949 (N_9949,N_9359,N_9171);
nand U9950 (N_9950,N_9163,N_9577);
or U9951 (N_9951,N_9256,N_9164);
xor U9952 (N_9952,N_9520,N_8837);
xor U9953 (N_9953,N_9468,N_9251);
and U9954 (N_9954,N_9597,N_9461);
and U9955 (N_9955,N_9253,N_9121);
and U9956 (N_9956,N_8869,N_9538);
xor U9957 (N_9957,N_9332,N_8936);
xor U9958 (N_9958,N_8955,N_9102);
or U9959 (N_9959,N_9015,N_8860);
or U9960 (N_9960,N_9449,N_8878);
xor U9961 (N_9961,N_8906,N_9555);
nand U9962 (N_9962,N_9575,N_9252);
and U9963 (N_9963,N_9566,N_9137);
or U9964 (N_9964,N_9045,N_9492);
nor U9965 (N_9965,N_9482,N_9599);
nand U9966 (N_9966,N_9051,N_9519);
or U9967 (N_9967,N_9047,N_9432);
nor U9968 (N_9968,N_9484,N_8979);
and U9969 (N_9969,N_9491,N_8935);
or U9970 (N_9970,N_9431,N_9404);
nor U9971 (N_9971,N_9559,N_9428);
xnor U9972 (N_9972,N_9175,N_9475);
xnor U9973 (N_9973,N_9029,N_9343);
or U9974 (N_9974,N_9073,N_9306);
and U9975 (N_9975,N_9549,N_8961);
nand U9976 (N_9976,N_9077,N_9234);
nand U9977 (N_9977,N_9018,N_8895);
or U9978 (N_9978,N_8870,N_9541);
or U9979 (N_9979,N_8872,N_9017);
or U9980 (N_9980,N_9403,N_9405);
nor U9981 (N_9981,N_9160,N_8909);
xor U9982 (N_9982,N_9197,N_9574);
xnor U9983 (N_9983,N_9341,N_9207);
nand U9984 (N_9984,N_9352,N_8843);
nand U9985 (N_9985,N_9003,N_9089);
or U9986 (N_9986,N_9008,N_9327);
or U9987 (N_9987,N_8853,N_8912);
and U9988 (N_9988,N_9367,N_9593);
xor U9989 (N_9989,N_9531,N_9400);
xnor U9990 (N_9990,N_9235,N_8993);
and U9991 (N_9991,N_9084,N_8923);
nor U9992 (N_9992,N_9036,N_9496);
and U9993 (N_9993,N_8927,N_9187);
xor U9994 (N_9994,N_9552,N_8822);
or U9995 (N_9995,N_9437,N_8857);
xnor U9996 (N_9996,N_8943,N_8985);
xor U9997 (N_9997,N_8898,N_9007);
nand U9998 (N_9998,N_9351,N_8949);
or U9999 (N_9999,N_9277,N_9189);
and U10000 (N_10000,N_8823,N_8852);
and U10001 (N_10001,N_9263,N_9102);
xnor U10002 (N_10002,N_9528,N_9142);
and U10003 (N_10003,N_9139,N_8957);
or U10004 (N_10004,N_9276,N_9344);
or U10005 (N_10005,N_9019,N_9438);
xnor U10006 (N_10006,N_9036,N_8936);
xor U10007 (N_10007,N_8815,N_9124);
nor U10008 (N_10008,N_9288,N_9240);
xnor U10009 (N_10009,N_9212,N_9543);
nand U10010 (N_10010,N_9318,N_9547);
nand U10011 (N_10011,N_9178,N_8984);
nor U10012 (N_10012,N_9176,N_9356);
or U10013 (N_10013,N_9144,N_8811);
nor U10014 (N_10014,N_9418,N_9504);
and U10015 (N_10015,N_9338,N_9066);
nand U10016 (N_10016,N_9323,N_9195);
nor U10017 (N_10017,N_9294,N_9247);
and U10018 (N_10018,N_9029,N_9529);
and U10019 (N_10019,N_8918,N_8865);
or U10020 (N_10020,N_9277,N_9049);
nor U10021 (N_10021,N_8858,N_9058);
xnor U10022 (N_10022,N_8944,N_9145);
nand U10023 (N_10023,N_9427,N_9278);
nand U10024 (N_10024,N_9020,N_9007);
xnor U10025 (N_10025,N_9303,N_9533);
nor U10026 (N_10026,N_8818,N_8860);
xnor U10027 (N_10027,N_9354,N_9336);
and U10028 (N_10028,N_9104,N_9267);
xnor U10029 (N_10029,N_8876,N_9536);
or U10030 (N_10030,N_9049,N_8871);
or U10031 (N_10031,N_9582,N_9059);
nand U10032 (N_10032,N_8949,N_9074);
xor U10033 (N_10033,N_9410,N_9227);
nand U10034 (N_10034,N_9041,N_8815);
nor U10035 (N_10035,N_9381,N_9376);
nand U10036 (N_10036,N_8883,N_9334);
or U10037 (N_10037,N_9411,N_9371);
xnor U10038 (N_10038,N_8965,N_8854);
nor U10039 (N_10039,N_9032,N_9076);
xor U10040 (N_10040,N_9584,N_8805);
and U10041 (N_10041,N_8894,N_9340);
xor U10042 (N_10042,N_8806,N_9347);
nor U10043 (N_10043,N_9051,N_8906);
xor U10044 (N_10044,N_9135,N_8977);
and U10045 (N_10045,N_9436,N_9377);
xor U10046 (N_10046,N_9310,N_8816);
or U10047 (N_10047,N_8879,N_9329);
nor U10048 (N_10048,N_8955,N_8825);
or U10049 (N_10049,N_8883,N_9301);
xor U10050 (N_10050,N_9176,N_9522);
nor U10051 (N_10051,N_9510,N_9559);
nand U10052 (N_10052,N_9042,N_8804);
xnor U10053 (N_10053,N_8840,N_8948);
and U10054 (N_10054,N_9072,N_8954);
xnor U10055 (N_10055,N_9277,N_9011);
nand U10056 (N_10056,N_8980,N_9112);
nor U10057 (N_10057,N_9330,N_8913);
or U10058 (N_10058,N_9100,N_9281);
xnor U10059 (N_10059,N_9413,N_9587);
and U10060 (N_10060,N_9457,N_9333);
or U10061 (N_10061,N_9040,N_9288);
nand U10062 (N_10062,N_8985,N_9046);
or U10063 (N_10063,N_9503,N_9188);
nand U10064 (N_10064,N_9490,N_9193);
nand U10065 (N_10065,N_9261,N_9565);
or U10066 (N_10066,N_9563,N_9260);
and U10067 (N_10067,N_8814,N_9124);
xor U10068 (N_10068,N_9330,N_9103);
xnor U10069 (N_10069,N_8884,N_9014);
nor U10070 (N_10070,N_9081,N_9055);
nor U10071 (N_10071,N_9223,N_9279);
xor U10072 (N_10072,N_8885,N_8936);
or U10073 (N_10073,N_8882,N_9129);
xor U10074 (N_10074,N_9255,N_9530);
xor U10075 (N_10075,N_8814,N_9405);
nand U10076 (N_10076,N_9411,N_9529);
nand U10077 (N_10077,N_9208,N_9490);
nand U10078 (N_10078,N_9445,N_8840);
and U10079 (N_10079,N_8947,N_9514);
nand U10080 (N_10080,N_8811,N_8914);
or U10081 (N_10081,N_8947,N_9032);
nor U10082 (N_10082,N_9495,N_8814);
nand U10083 (N_10083,N_9070,N_9025);
or U10084 (N_10084,N_9217,N_9240);
or U10085 (N_10085,N_9206,N_9183);
or U10086 (N_10086,N_9216,N_9437);
nor U10087 (N_10087,N_8958,N_9066);
xnor U10088 (N_10088,N_9032,N_9299);
xor U10089 (N_10089,N_9478,N_9215);
nand U10090 (N_10090,N_9112,N_9049);
nor U10091 (N_10091,N_9465,N_9009);
or U10092 (N_10092,N_8837,N_9434);
and U10093 (N_10093,N_9251,N_8889);
nand U10094 (N_10094,N_9017,N_9341);
or U10095 (N_10095,N_9391,N_9432);
and U10096 (N_10096,N_9589,N_9072);
nor U10097 (N_10097,N_8819,N_9299);
nand U10098 (N_10098,N_9454,N_9256);
or U10099 (N_10099,N_9140,N_9241);
or U10100 (N_10100,N_8814,N_9060);
and U10101 (N_10101,N_9075,N_9299);
nand U10102 (N_10102,N_8809,N_8841);
xnor U10103 (N_10103,N_9533,N_9364);
nor U10104 (N_10104,N_8947,N_9407);
and U10105 (N_10105,N_9265,N_8820);
and U10106 (N_10106,N_8822,N_9442);
xnor U10107 (N_10107,N_9551,N_9421);
xor U10108 (N_10108,N_9070,N_9549);
xnor U10109 (N_10109,N_8833,N_8965);
or U10110 (N_10110,N_9079,N_8812);
nand U10111 (N_10111,N_9371,N_9251);
xor U10112 (N_10112,N_9310,N_9243);
nand U10113 (N_10113,N_8987,N_8848);
and U10114 (N_10114,N_8982,N_9234);
and U10115 (N_10115,N_9334,N_9089);
nor U10116 (N_10116,N_8807,N_9571);
or U10117 (N_10117,N_9127,N_9436);
and U10118 (N_10118,N_9599,N_9303);
nand U10119 (N_10119,N_8816,N_8986);
nor U10120 (N_10120,N_8951,N_9306);
and U10121 (N_10121,N_9457,N_9554);
or U10122 (N_10122,N_9044,N_8811);
xor U10123 (N_10123,N_9581,N_9278);
xnor U10124 (N_10124,N_9421,N_9132);
nor U10125 (N_10125,N_8894,N_9116);
and U10126 (N_10126,N_8975,N_8886);
xor U10127 (N_10127,N_9351,N_9050);
nand U10128 (N_10128,N_9517,N_8803);
nand U10129 (N_10129,N_8889,N_9554);
or U10130 (N_10130,N_8843,N_8949);
nand U10131 (N_10131,N_9192,N_8937);
or U10132 (N_10132,N_8838,N_9067);
nand U10133 (N_10133,N_9472,N_8814);
xor U10134 (N_10134,N_8943,N_8989);
or U10135 (N_10135,N_8816,N_8847);
or U10136 (N_10136,N_8983,N_9462);
and U10137 (N_10137,N_9088,N_8897);
xnor U10138 (N_10138,N_9287,N_9132);
or U10139 (N_10139,N_9397,N_8834);
nor U10140 (N_10140,N_9267,N_8936);
or U10141 (N_10141,N_8872,N_9510);
xor U10142 (N_10142,N_8930,N_9444);
nor U10143 (N_10143,N_8856,N_9190);
or U10144 (N_10144,N_9311,N_9576);
nor U10145 (N_10145,N_9489,N_9212);
nor U10146 (N_10146,N_9455,N_9383);
nand U10147 (N_10147,N_9551,N_9113);
nor U10148 (N_10148,N_9501,N_9075);
or U10149 (N_10149,N_9216,N_9247);
or U10150 (N_10150,N_9089,N_9507);
nand U10151 (N_10151,N_9153,N_9577);
nor U10152 (N_10152,N_8865,N_8884);
or U10153 (N_10153,N_8886,N_9491);
nand U10154 (N_10154,N_9092,N_9237);
xor U10155 (N_10155,N_8894,N_9337);
or U10156 (N_10156,N_9451,N_9492);
xor U10157 (N_10157,N_9570,N_9390);
and U10158 (N_10158,N_9346,N_9321);
xor U10159 (N_10159,N_9319,N_8924);
nand U10160 (N_10160,N_8917,N_8902);
nand U10161 (N_10161,N_9169,N_9103);
nand U10162 (N_10162,N_9269,N_9448);
and U10163 (N_10163,N_9576,N_9287);
xor U10164 (N_10164,N_9208,N_9130);
and U10165 (N_10165,N_9452,N_9076);
xnor U10166 (N_10166,N_9540,N_8869);
nand U10167 (N_10167,N_9460,N_9300);
nor U10168 (N_10168,N_9332,N_8867);
and U10169 (N_10169,N_9577,N_9550);
or U10170 (N_10170,N_8986,N_9509);
xor U10171 (N_10171,N_9269,N_9182);
nor U10172 (N_10172,N_9456,N_9075);
and U10173 (N_10173,N_8845,N_9544);
xnor U10174 (N_10174,N_9518,N_8925);
nor U10175 (N_10175,N_9536,N_8807);
nor U10176 (N_10176,N_9290,N_9536);
and U10177 (N_10177,N_9322,N_8835);
nand U10178 (N_10178,N_9192,N_9030);
and U10179 (N_10179,N_8939,N_9211);
or U10180 (N_10180,N_8899,N_8883);
or U10181 (N_10181,N_8982,N_8992);
and U10182 (N_10182,N_9061,N_8917);
nand U10183 (N_10183,N_9445,N_8997);
nand U10184 (N_10184,N_9059,N_9237);
xnor U10185 (N_10185,N_9393,N_9441);
xor U10186 (N_10186,N_8801,N_8910);
and U10187 (N_10187,N_8978,N_9372);
xor U10188 (N_10188,N_8993,N_8954);
and U10189 (N_10189,N_9401,N_9079);
xor U10190 (N_10190,N_9550,N_9088);
or U10191 (N_10191,N_9445,N_9093);
or U10192 (N_10192,N_9295,N_9326);
xor U10193 (N_10193,N_9420,N_9191);
nand U10194 (N_10194,N_9416,N_9293);
and U10195 (N_10195,N_8975,N_9370);
nand U10196 (N_10196,N_8983,N_9071);
xor U10197 (N_10197,N_9080,N_8972);
or U10198 (N_10198,N_9094,N_9145);
and U10199 (N_10199,N_9534,N_9203);
and U10200 (N_10200,N_8871,N_9006);
nor U10201 (N_10201,N_9082,N_9122);
xor U10202 (N_10202,N_8989,N_9405);
or U10203 (N_10203,N_9118,N_8920);
and U10204 (N_10204,N_9175,N_9547);
xor U10205 (N_10205,N_9452,N_8827);
nor U10206 (N_10206,N_9218,N_8836);
nand U10207 (N_10207,N_9207,N_8939);
or U10208 (N_10208,N_9467,N_9367);
xor U10209 (N_10209,N_9422,N_8924);
nor U10210 (N_10210,N_8903,N_8800);
nor U10211 (N_10211,N_9113,N_8945);
nor U10212 (N_10212,N_9393,N_9530);
nand U10213 (N_10213,N_9179,N_9380);
or U10214 (N_10214,N_8966,N_9576);
nand U10215 (N_10215,N_9026,N_8822);
or U10216 (N_10216,N_9187,N_9392);
nand U10217 (N_10217,N_9216,N_9304);
xor U10218 (N_10218,N_9477,N_9051);
nand U10219 (N_10219,N_9465,N_9043);
or U10220 (N_10220,N_9338,N_8807);
or U10221 (N_10221,N_8858,N_9381);
nand U10222 (N_10222,N_8982,N_9551);
and U10223 (N_10223,N_9399,N_8826);
or U10224 (N_10224,N_9468,N_9167);
nor U10225 (N_10225,N_8977,N_9471);
nand U10226 (N_10226,N_9266,N_9390);
xor U10227 (N_10227,N_9049,N_9338);
nor U10228 (N_10228,N_9231,N_9244);
xor U10229 (N_10229,N_9437,N_9122);
or U10230 (N_10230,N_9240,N_9111);
nand U10231 (N_10231,N_9424,N_9331);
and U10232 (N_10232,N_9247,N_8948);
and U10233 (N_10233,N_9437,N_9563);
nand U10234 (N_10234,N_9072,N_9523);
xnor U10235 (N_10235,N_8809,N_9332);
xor U10236 (N_10236,N_8823,N_9098);
nand U10237 (N_10237,N_9128,N_9077);
nand U10238 (N_10238,N_9363,N_9318);
xnor U10239 (N_10239,N_9540,N_9367);
and U10240 (N_10240,N_9483,N_9362);
and U10241 (N_10241,N_9532,N_8811);
and U10242 (N_10242,N_8994,N_8944);
nand U10243 (N_10243,N_9482,N_8875);
nand U10244 (N_10244,N_8851,N_9322);
nand U10245 (N_10245,N_9275,N_9397);
nor U10246 (N_10246,N_9231,N_8909);
nor U10247 (N_10247,N_9519,N_8974);
or U10248 (N_10248,N_9247,N_9505);
xor U10249 (N_10249,N_9529,N_9086);
and U10250 (N_10250,N_9176,N_9428);
and U10251 (N_10251,N_8994,N_8925);
nand U10252 (N_10252,N_9268,N_9571);
xnor U10253 (N_10253,N_9361,N_9596);
and U10254 (N_10254,N_9163,N_9295);
nor U10255 (N_10255,N_9278,N_9347);
or U10256 (N_10256,N_9064,N_8903);
and U10257 (N_10257,N_8843,N_9570);
xnor U10258 (N_10258,N_9047,N_9581);
xnor U10259 (N_10259,N_8985,N_9338);
xnor U10260 (N_10260,N_9482,N_9397);
nand U10261 (N_10261,N_9126,N_9206);
xor U10262 (N_10262,N_8909,N_8933);
nand U10263 (N_10263,N_8869,N_8892);
xnor U10264 (N_10264,N_8978,N_8989);
nand U10265 (N_10265,N_9483,N_9301);
nor U10266 (N_10266,N_9065,N_9371);
and U10267 (N_10267,N_9437,N_9289);
xnor U10268 (N_10268,N_8928,N_8947);
nor U10269 (N_10269,N_8845,N_9495);
nor U10270 (N_10270,N_9490,N_9483);
or U10271 (N_10271,N_9369,N_9394);
or U10272 (N_10272,N_9274,N_8928);
nor U10273 (N_10273,N_9390,N_9351);
or U10274 (N_10274,N_9266,N_9396);
and U10275 (N_10275,N_9564,N_9275);
nor U10276 (N_10276,N_9510,N_9383);
and U10277 (N_10277,N_8808,N_8850);
nor U10278 (N_10278,N_9211,N_9173);
and U10279 (N_10279,N_9016,N_9097);
xor U10280 (N_10280,N_8918,N_9258);
or U10281 (N_10281,N_9014,N_9325);
xor U10282 (N_10282,N_9433,N_8908);
xor U10283 (N_10283,N_8814,N_8848);
nand U10284 (N_10284,N_9467,N_8996);
or U10285 (N_10285,N_9472,N_8982);
xnor U10286 (N_10286,N_9575,N_9249);
nand U10287 (N_10287,N_9057,N_9336);
or U10288 (N_10288,N_9158,N_9265);
and U10289 (N_10289,N_9500,N_9194);
or U10290 (N_10290,N_9257,N_9250);
xor U10291 (N_10291,N_9035,N_8868);
xnor U10292 (N_10292,N_9175,N_9311);
nor U10293 (N_10293,N_8945,N_9463);
or U10294 (N_10294,N_9591,N_9013);
xor U10295 (N_10295,N_9418,N_8844);
nor U10296 (N_10296,N_9300,N_9438);
nor U10297 (N_10297,N_9206,N_9588);
or U10298 (N_10298,N_9220,N_9381);
or U10299 (N_10299,N_9205,N_9512);
xnor U10300 (N_10300,N_9330,N_9188);
and U10301 (N_10301,N_9306,N_9353);
and U10302 (N_10302,N_9362,N_9459);
xnor U10303 (N_10303,N_9206,N_9356);
xor U10304 (N_10304,N_9349,N_9587);
and U10305 (N_10305,N_9187,N_9160);
xnor U10306 (N_10306,N_9320,N_9520);
or U10307 (N_10307,N_8950,N_8852);
or U10308 (N_10308,N_8940,N_8932);
nand U10309 (N_10309,N_9149,N_8862);
or U10310 (N_10310,N_9416,N_9088);
nand U10311 (N_10311,N_9481,N_9490);
xor U10312 (N_10312,N_9108,N_9052);
xnor U10313 (N_10313,N_9379,N_9330);
nor U10314 (N_10314,N_8921,N_9252);
xor U10315 (N_10315,N_9508,N_9312);
nand U10316 (N_10316,N_9259,N_9484);
nand U10317 (N_10317,N_9121,N_9330);
and U10318 (N_10318,N_9083,N_9555);
nand U10319 (N_10319,N_9506,N_9426);
nor U10320 (N_10320,N_9019,N_8842);
xor U10321 (N_10321,N_9378,N_8862);
or U10322 (N_10322,N_9108,N_8963);
and U10323 (N_10323,N_9363,N_9097);
xnor U10324 (N_10324,N_9001,N_9453);
or U10325 (N_10325,N_9223,N_8931);
and U10326 (N_10326,N_9363,N_9163);
or U10327 (N_10327,N_9533,N_9239);
and U10328 (N_10328,N_9370,N_9240);
xor U10329 (N_10329,N_9067,N_8922);
or U10330 (N_10330,N_9182,N_9448);
and U10331 (N_10331,N_9249,N_9029);
and U10332 (N_10332,N_9323,N_9142);
nand U10333 (N_10333,N_9419,N_9181);
xor U10334 (N_10334,N_9304,N_9445);
nand U10335 (N_10335,N_9370,N_9476);
and U10336 (N_10336,N_9151,N_9072);
and U10337 (N_10337,N_8933,N_9246);
nand U10338 (N_10338,N_9487,N_8881);
xnor U10339 (N_10339,N_9389,N_9082);
nand U10340 (N_10340,N_9402,N_9103);
or U10341 (N_10341,N_8915,N_8931);
nor U10342 (N_10342,N_8965,N_8836);
or U10343 (N_10343,N_8873,N_9401);
nor U10344 (N_10344,N_9372,N_9552);
nand U10345 (N_10345,N_9594,N_9531);
nand U10346 (N_10346,N_9553,N_9256);
or U10347 (N_10347,N_9285,N_9340);
nor U10348 (N_10348,N_9438,N_9391);
nor U10349 (N_10349,N_8855,N_9436);
and U10350 (N_10350,N_8865,N_9439);
xor U10351 (N_10351,N_9510,N_9019);
nor U10352 (N_10352,N_9560,N_8931);
or U10353 (N_10353,N_9124,N_9575);
nor U10354 (N_10354,N_9261,N_9327);
xor U10355 (N_10355,N_9270,N_8805);
nand U10356 (N_10356,N_9269,N_9453);
and U10357 (N_10357,N_8954,N_9227);
nand U10358 (N_10358,N_8973,N_9382);
nor U10359 (N_10359,N_9197,N_9428);
nor U10360 (N_10360,N_9597,N_9062);
or U10361 (N_10361,N_8917,N_9230);
nor U10362 (N_10362,N_8889,N_8811);
xnor U10363 (N_10363,N_9275,N_8827);
or U10364 (N_10364,N_9336,N_9158);
xor U10365 (N_10365,N_9220,N_9524);
xor U10366 (N_10366,N_9564,N_9577);
and U10367 (N_10367,N_9258,N_9349);
nand U10368 (N_10368,N_9100,N_9236);
and U10369 (N_10369,N_9075,N_9104);
and U10370 (N_10370,N_9280,N_9215);
nor U10371 (N_10371,N_9195,N_9060);
nor U10372 (N_10372,N_9101,N_9274);
nor U10373 (N_10373,N_9215,N_9577);
xnor U10374 (N_10374,N_9131,N_9127);
nor U10375 (N_10375,N_9156,N_9202);
nor U10376 (N_10376,N_8903,N_9387);
nand U10377 (N_10377,N_9555,N_9198);
and U10378 (N_10378,N_8945,N_9245);
nand U10379 (N_10379,N_8878,N_9446);
and U10380 (N_10380,N_9092,N_9389);
nand U10381 (N_10381,N_9381,N_9577);
and U10382 (N_10382,N_9396,N_9353);
or U10383 (N_10383,N_9225,N_9528);
and U10384 (N_10384,N_9368,N_8994);
xnor U10385 (N_10385,N_9243,N_9096);
and U10386 (N_10386,N_8901,N_8808);
and U10387 (N_10387,N_8917,N_9031);
nor U10388 (N_10388,N_9333,N_8959);
or U10389 (N_10389,N_9006,N_9158);
nor U10390 (N_10390,N_9201,N_9301);
nand U10391 (N_10391,N_9283,N_9522);
or U10392 (N_10392,N_9207,N_9471);
xor U10393 (N_10393,N_9504,N_9598);
or U10394 (N_10394,N_8919,N_8955);
or U10395 (N_10395,N_9592,N_9339);
or U10396 (N_10396,N_9459,N_9246);
xnor U10397 (N_10397,N_8960,N_8816);
xor U10398 (N_10398,N_9145,N_9599);
and U10399 (N_10399,N_8985,N_9443);
and U10400 (N_10400,N_10207,N_10369);
and U10401 (N_10401,N_9767,N_10078);
nor U10402 (N_10402,N_10152,N_9636);
xnor U10403 (N_10403,N_10047,N_10299);
xor U10404 (N_10404,N_9704,N_10263);
or U10405 (N_10405,N_9692,N_10268);
or U10406 (N_10406,N_9856,N_9902);
nor U10407 (N_10407,N_9635,N_10284);
xor U10408 (N_10408,N_9674,N_10051);
nor U10409 (N_10409,N_10352,N_9629);
or U10410 (N_10410,N_10394,N_10059);
and U10411 (N_10411,N_9623,N_10210);
or U10412 (N_10412,N_10069,N_9615);
xor U10413 (N_10413,N_10276,N_9601);
nor U10414 (N_10414,N_10258,N_10092);
or U10415 (N_10415,N_9804,N_10387);
nor U10416 (N_10416,N_10385,N_10338);
or U10417 (N_10417,N_10066,N_9952);
and U10418 (N_10418,N_9651,N_9628);
nor U10419 (N_10419,N_10166,N_10082);
xnor U10420 (N_10420,N_10185,N_10018);
nor U10421 (N_10421,N_10211,N_10359);
or U10422 (N_10422,N_10310,N_10122);
nand U10423 (N_10423,N_9923,N_10247);
nand U10424 (N_10424,N_9865,N_9846);
and U10425 (N_10425,N_10060,N_9777);
nor U10426 (N_10426,N_10164,N_10271);
nand U10427 (N_10427,N_10212,N_10305);
and U10428 (N_10428,N_10302,N_9990);
xnor U10429 (N_10429,N_10091,N_10147);
nor U10430 (N_10430,N_10137,N_10265);
or U10431 (N_10431,N_9673,N_10230);
nand U10432 (N_10432,N_10188,N_9632);
nor U10433 (N_10433,N_9922,N_9737);
nand U10434 (N_10434,N_10264,N_9653);
or U10435 (N_10435,N_9740,N_9835);
and U10436 (N_10436,N_9697,N_10384);
nand U10437 (N_10437,N_9996,N_9717);
nand U10438 (N_10438,N_10100,N_9626);
nor U10439 (N_10439,N_10179,N_9969);
and U10440 (N_10440,N_9751,N_9700);
nor U10441 (N_10441,N_10133,N_10165);
nand U10442 (N_10442,N_9842,N_10195);
nor U10443 (N_10443,N_9761,N_9606);
xnor U10444 (N_10444,N_9621,N_10221);
nand U10445 (N_10445,N_9691,N_10105);
nand U10446 (N_10446,N_9920,N_10234);
and U10447 (N_10447,N_9609,N_10150);
and U10448 (N_10448,N_9983,N_10172);
or U10449 (N_10449,N_9634,N_10000);
nor U10450 (N_10450,N_10358,N_9669);
and U10451 (N_10451,N_10303,N_9799);
nand U10452 (N_10452,N_10058,N_9819);
or U10453 (N_10453,N_9764,N_10161);
and U10454 (N_10454,N_9979,N_10323);
or U10455 (N_10455,N_10329,N_9770);
nand U10456 (N_10456,N_9785,N_10061);
xor U10457 (N_10457,N_9690,N_9695);
xor U10458 (N_10458,N_9872,N_9683);
and U10459 (N_10459,N_10024,N_9627);
or U10460 (N_10460,N_9859,N_10312);
xnor U10461 (N_10461,N_9645,N_10370);
nor U10462 (N_10462,N_9878,N_9736);
nand U10463 (N_10463,N_10139,N_10117);
and U10464 (N_10464,N_9656,N_9986);
or U10465 (N_10465,N_9932,N_10224);
xnor U10466 (N_10466,N_9602,N_9857);
and U10467 (N_10467,N_10344,N_10270);
and U10468 (N_10468,N_10055,N_10392);
xor U10469 (N_10469,N_9714,N_9852);
or U10470 (N_10470,N_10154,N_9929);
or U10471 (N_10471,N_9694,N_9904);
nand U10472 (N_10472,N_9958,N_9985);
nand U10473 (N_10473,N_10374,N_10040);
or U10474 (N_10474,N_10362,N_9892);
nor U10475 (N_10475,N_9721,N_10112);
xnor U10476 (N_10476,N_9912,N_9992);
nor U10477 (N_10477,N_9964,N_9925);
nor U10478 (N_10478,N_9862,N_10007);
nor U10479 (N_10479,N_10277,N_10099);
or U10480 (N_10480,N_9706,N_10238);
nand U10481 (N_10481,N_9988,N_9688);
nor U10482 (N_10482,N_9646,N_9977);
nand U10483 (N_10483,N_10200,N_9625);
xnor U10484 (N_10484,N_9998,N_9843);
or U10485 (N_10485,N_9987,N_9670);
and U10486 (N_10486,N_9924,N_9773);
or U10487 (N_10487,N_9911,N_10118);
and U10488 (N_10488,N_10328,N_10322);
nor U10489 (N_10489,N_9855,N_10288);
nand U10490 (N_10490,N_9624,N_9783);
xnor U10491 (N_10491,N_10022,N_10208);
nand U10492 (N_10492,N_10204,N_10140);
and U10493 (N_10493,N_10318,N_10038);
xor U10494 (N_10494,N_10309,N_9776);
xnor U10495 (N_10495,N_9715,N_9655);
or U10496 (N_10496,N_10054,N_10259);
and U10497 (N_10497,N_9928,N_9800);
or U10498 (N_10498,N_10366,N_9766);
or U10499 (N_10499,N_9847,N_10375);
or U10500 (N_10500,N_9633,N_9798);
xnor U10501 (N_10501,N_10114,N_10155);
and U10502 (N_10502,N_9916,N_9619);
and U10503 (N_10503,N_9890,N_10381);
and U10504 (N_10504,N_9680,N_10176);
xor U10505 (N_10505,N_10135,N_10390);
and U10506 (N_10506,N_9604,N_9891);
xnor U10507 (N_10507,N_10278,N_10044);
nor U10508 (N_10508,N_10115,N_9909);
or U10509 (N_10509,N_9994,N_10039);
nand U10510 (N_10510,N_9757,N_10248);
or U10511 (N_10511,N_9905,N_9951);
and U10512 (N_10512,N_10050,N_10380);
and U10513 (N_10513,N_10102,N_10255);
nor U10514 (N_10514,N_9710,N_9778);
nand U10515 (N_10515,N_9752,N_9617);
xor U10516 (N_10516,N_9818,N_9849);
nand U10517 (N_10517,N_9885,N_9719);
or U10518 (N_10518,N_9803,N_9810);
or U10519 (N_10519,N_10222,N_10081);
xnor U10520 (N_10520,N_10010,N_10218);
nand U10521 (N_10521,N_9889,N_9733);
nor U10522 (N_10522,N_9950,N_9837);
xnor U10523 (N_10523,N_9944,N_10353);
or U10524 (N_10524,N_9967,N_10070);
nor U10525 (N_10525,N_10332,N_9814);
xnor U10526 (N_10526,N_9822,N_10001);
xnor U10527 (N_10527,N_9630,N_10032);
and U10528 (N_10528,N_9833,N_9744);
or U10529 (N_10529,N_9701,N_10151);
and U10530 (N_10530,N_9940,N_9802);
nand U10531 (N_10531,N_10308,N_9899);
and U10532 (N_10532,N_10097,N_10107);
nor U10533 (N_10533,N_10223,N_10254);
or U10534 (N_10534,N_10244,N_9809);
nand U10535 (N_10535,N_9984,N_10233);
or U10536 (N_10536,N_9603,N_9735);
xor U10537 (N_10537,N_10226,N_9795);
xnor U10538 (N_10538,N_10198,N_10042);
nand U10539 (N_10539,N_9935,N_10260);
and U10540 (N_10540,N_9622,N_9848);
or U10541 (N_10541,N_10280,N_10160);
nor U10542 (N_10542,N_10327,N_9726);
nor U10543 (N_10543,N_10023,N_10372);
nor U10544 (N_10544,N_10011,N_9966);
nand U10545 (N_10545,N_10395,N_9637);
and U10546 (N_10546,N_9828,N_10324);
and U10547 (N_10547,N_9768,N_9755);
nand U10548 (N_10548,N_9789,N_10283);
nor U10549 (N_10549,N_10068,N_9941);
and U10550 (N_10550,N_10049,N_10341);
xor U10551 (N_10551,N_9839,N_10232);
and U10552 (N_10552,N_9811,N_9685);
and U10553 (N_10553,N_10124,N_10028);
and U10554 (N_10554,N_10245,N_9732);
and U10555 (N_10555,N_10269,N_9995);
and U10556 (N_10556,N_10216,N_10141);
nand U10557 (N_10557,N_9906,N_9709);
or U10558 (N_10558,N_10377,N_9663);
xnor U10559 (N_10559,N_10062,N_10073);
and U10560 (N_10560,N_10014,N_10237);
and U10561 (N_10561,N_10206,N_10213);
or U10562 (N_10562,N_10174,N_9873);
and U10563 (N_10563,N_10311,N_10340);
or U10564 (N_10564,N_9679,N_10191);
nand U10565 (N_10565,N_9908,N_9711);
and U10566 (N_10566,N_10189,N_10065);
or U10567 (N_10567,N_10257,N_9931);
nor U10568 (N_10568,N_9639,N_10231);
nor U10569 (N_10569,N_9769,N_9649);
and U10570 (N_10570,N_10167,N_9989);
nand U10571 (N_10571,N_9650,N_9863);
nand U10572 (N_10572,N_9827,N_9946);
nor U10573 (N_10573,N_9961,N_9716);
or U10574 (N_10574,N_9771,N_10186);
nand U10575 (N_10575,N_9973,N_10031);
and U10576 (N_10576,N_9641,N_10134);
xor U10577 (N_10577,N_9684,N_9729);
xnor U10578 (N_10578,N_9782,N_9965);
nor U10579 (N_10579,N_9658,N_10330);
nand U10580 (N_10580,N_10389,N_9868);
nand U10581 (N_10581,N_10138,N_10291);
nand U10582 (N_10582,N_9614,N_9661);
nand U10583 (N_10583,N_10052,N_10190);
and U10584 (N_10584,N_9953,N_10080);
xnor U10585 (N_10585,N_9664,N_9871);
xor U10586 (N_10586,N_9841,N_10015);
nand U10587 (N_10587,N_9786,N_9812);
nand U10588 (N_10588,N_9870,N_10398);
and U10589 (N_10589,N_10116,N_10335);
xnor U10590 (N_10590,N_10256,N_10274);
xnor U10591 (N_10591,N_10201,N_9877);
nand U10592 (N_10592,N_9844,N_10184);
and U10593 (N_10593,N_10365,N_9972);
nor U10594 (N_10594,N_10334,N_9753);
or U10595 (N_10595,N_10220,N_10379);
nand U10596 (N_10596,N_9618,N_9763);
nand U10597 (N_10597,N_10246,N_9724);
xor U10598 (N_10598,N_9921,N_10250);
or U10599 (N_10599,N_10316,N_10045);
nand U10600 (N_10600,N_10143,N_10009);
nor U10601 (N_10601,N_9918,N_9762);
nor U10602 (N_10602,N_9886,N_10339);
or U10603 (N_10603,N_10298,N_10388);
and U10604 (N_10604,N_10294,N_9978);
nand U10605 (N_10605,N_10243,N_9853);
nand U10606 (N_10606,N_10202,N_10382);
nor U10607 (N_10607,N_9616,N_10314);
xor U10608 (N_10608,N_9774,N_9743);
xnor U10609 (N_10609,N_10005,N_10085);
and U10610 (N_10610,N_10321,N_10026);
xnor U10611 (N_10611,N_10333,N_10063);
xnor U10612 (N_10612,N_10159,N_9805);
xnor U10613 (N_10613,N_10295,N_10076);
nand U10614 (N_10614,N_10019,N_9725);
nor U10615 (N_10615,N_9980,N_9861);
nand U10616 (N_10616,N_9672,N_10357);
xor U10617 (N_10617,N_10103,N_10229);
or U10618 (N_10618,N_9807,N_10391);
nand U10619 (N_10619,N_10146,N_9657);
xor U10620 (N_10620,N_10214,N_10158);
nand U10621 (N_10621,N_10181,N_9671);
nor U10622 (N_10622,N_10029,N_9917);
or U10623 (N_10623,N_9816,N_10109);
and U10624 (N_10624,N_9832,N_10037);
nand U10625 (N_10625,N_10021,N_9620);
and U10626 (N_10626,N_10219,N_9659);
or U10627 (N_10627,N_10354,N_9647);
xnor U10628 (N_10628,N_10142,N_10048);
or U10629 (N_10629,N_10307,N_9829);
or U10630 (N_10630,N_10197,N_10084);
and U10631 (N_10631,N_9790,N_10378);
or U10632 (N_10632,N_9612,N_9741);
nor U10633 (N_10633,N_10043,N_9954);
xnor U10634 (N_10634,N_10225,N_9875);
and U10635 (N_10635,N_10093,N_9644);
nor U10636 (N_10636,N_10171,N_10349);
xor U10637 (N_10637,N_9727,N_9668);
nand U10638 (N_10638,N_9772,N_9640);
nor U10639 (N_10639,N_9938,N_9815);
and U10640 (N_10640,N_9936,N_10169);
xor U10641 (N_10641,N_10034,N_10035);
nor U10642 (N_10642,N_10033,N_9797);
xor U10643 (N_10643,N_9600,N_10182);
nand U10644 (N_10644,N_10331,N_9792);
nor U10645 (N_10645,N_9826,N_9860);
and U10646 (N_10646,N_9897,N_9817);
or U10647 (N_10647,N_9677,N_10071);
or U10648 (N_10648,N_10083,N_9821);
and U10649 (N_10649,N_10235,N_9718);
xnor U10650 (N_10650,N_9613,N_10347);
and U10651 (N_10651,N_9682,N_9702);
or U10652 (N_10652,N_10096,N_10383);
or U10653 (N_10653,N_10132,N_9887);
nor U10654 (N_10654,N_10285,N_10106);
nor U10655 (N_10655,N_9881,N_10217);
nand U10656 (N_10656,N_10241,N_10317);
and U10657 (N_10657,N_10157,N_10348);
or U10658 (N_10658,N_10129,N_10290);
nand U10659 (N_10659,N_9882,N_9981);
nor U10660 (N_10660,N_9901,N_10006);
xnor U10661 (N_10661,N_9830,N_10337);
xnor U10662 (N_10662,N_9914,N_9907);
or U10663 (N_10663,N_9813,N_9896);
nand U10664 (N_10664,N_9793,N_9993);
or U10665 (N_10665,N_9971,N_9884);
xnor U10666 (N_10666,N_9608,N_9749);
nand U10667 (N_10667,N_10267,N_10304);
nand U10668 (N_10668,N_10002,N_10089);
nand U10669 (N_10669,N_10130,N_10373);
nor U10670 (N_10670,N_9991,N_9708);
and U10671 (N_10671,N_10113,N_9742);
or U10672 (N_10672,N_9693,N_9898);
or U10673 (N_10673,N_10056,N_10004);
or U10674 (N_10674,N_9784,N_10192);
nor U10675 (N_10675,N_9997,N_10396);
nand U10676 (N_10676,N_10281,N_9957);
xor U10677 (N_10677,N_10279,N_9738);
or U10678 (N_10678,N_10363,N_10360);
nor U10679 (N_10679,N_10199,N_10053);
or U10680 (N_10680,N_9903,N_9959);
nand U10681 (N_10681,N_9927,N_9883);
nand U10682 (N_10682,N_10275,N_9960);
and U10683 (N_10683,N_10350,N_9949);
or U10684 (N_10684,N_9939,N_10228);
xnor U10685 (N_10685,N_10123,N_10399);
or U10686 (N_10686,N_9631,N_10016);
nand U10687 (N_10687,N_10205,N_9963);
xnor U10688 (N_10688,N_10397,N_10145);
and U10689 (N_10689,N_9943,N_9945);
or U10690 (N_10690,N_9605,N_10194);
xor U10691 (N_10691,N_10183,N_9610);
nand U10692 (N_10692,N_10193,N_10012);
xor U10693 (N_10693,N_9712,N_9638);
nor U10694 (N_10694,N_9703,N_10110);
and U10695 (N_10695,N_9788,N_10215);
nor U10696 (N_10696,N_9720,N_10036);
xnor U10697 (N_10697,N_10293,N_10090);
and U10698 (N_10698,N_10125,N_10095);
nor U10699 (N_10699,N_10239,N_9643);
and U10700 (N_10700,N_9707,N_9831);
nor U10701 (N_10701,N_9869,N_9806);
and U10702 (N_10702,N_9867,N_9824);
xnor U10703 (N_10703,N_10343,N_10163);
nand U10704 (N_10704,N_10153,N_10162);
xor U10705 (N_10705,N_9746,N_10261);
or U10706 (N_10706,N_10282,N_9760);
nand U10707 (N_10707,N_10272,N_9705);
nor U10708 (N_10708,N_9754,N_10251);
or U10709 (N_10709,N_10175,N_9747);
and U10710 (N_10710,N_9975,N_10030);
nor U10711 (N_10711,N_10273,N_10041);
or U10712 (N_10712,N_10262,N_9675);
xnor U10713 (N_10713,N_9662,N_10227);
xor U10714 (N_10714,N_9956,N_10074);
nor U10715 (N_10715,N_10361,N_9607);
xor U10716 (N_10716,N_9900,N_10098);
xor U10717 (N_10717,N_9825,N_10136);
nor U10718 (N_10718,N_9970,N_10286);
or U10719 (N_10719,N_10156,N_9734);
nor U10720 (N_10720,N_10017,N_9723);
xnor U10721 (N_10721,N_9851,N_9780);
or U10722 (N_10722,N_9687,N_10367);
nor U10723 (N_10723,N_10057,N_10345);
xnor U10724 (N_10724,N_10249,N_10356);
nor U10725 (N_10725,N_9840,N_9808);
xnor U10726 (N_10726,N_10236,N_9934);
nand U10727 (N_10727,N_9836,N_9728);
nand U10728 (N_10728,N_10148,N_10266);
or U10729 (N_10729,N_10300,N_9968);
nand U10730 (N_10730,N_10177,N_10077);
and U10731 (N_10731,N_10368,N_9689);
nand U10732 (N_10732,N_10287,N_10289);
and U10733 (N_10733,N_10170,N_9999);
nor U10734 (N_10734,N_9933,N_10027);
and U10735 (N_10735,N_9748,N_10126);
nor U10736 (N_10736,N_9654,N_10119);
nor U10737 (N_10737,N_9686,N_9820);
nor U10738 (N_10738,N_9866,N_10111);
or U10739 (N_10739,N_9801,N_9779);
nor U10740 (N_10740,N_10313,N_9879);
nand U10741 (N_10741,N_10292,N_9876);
xnor U10742 (N_10742,N_10364,N_9880);
nand U10743 (N_10743,N_9730,N_9915);
nand U10744 (N_10744,N_10240,N_9775);
or U10745 (N_10745,N_10144,N_10376);
nand U10746 (N_10746,N_10242,N_9823);
or U10747 (N_10747,N_9696,N_10088);
and U10748 (N_10748,N_10013,N_9794);
xnor U10749 (N_10749,N_10371,N_10325);
xor U10750 (N_10750,N_10351,N_9948);
xor U10751 (N_10751,N_10319,N_10128);
nand U10752 (N_10752,N_10306,N_10386);
and U10753 (N_10753,N_9791,N_10127);
xor U10754 (N_10754,N_9974,N_9698);
xnor U10755 (N_10755,N_10346,N_9874);
or U10756 (N_10756,N_10149,N_9745);
and U10757 (N_10757,N_9699,N_9681);
and U10758 (N_10758,N_9652,N_9758);
xor U10759 (N_10759,N_10072,N_9731);
nor U10760 (N_10760,N_9864,N_10315);
or U10761 (N_10761,N_9947,N_9642);
and U10762 (N_10762,N_10203,N_9756);
or U10763 (N_10763,N_9787,N_9937);
xor U10764 (N_10764,N_10003,N_9955);
xor U10765 (N_10765,N_9888,N_9942);
nand U10766 (N_10766,N_9660,N_10025);
nor U10767 (N_10767,N_9678,N_9930);
nand U10768 (N_10768,N_10209,N_10008);
nand U10769 (N_10769,N_9781,N_10168);
and U10770 (N_10770,N_10393,N_10320);
nand U10771 (N_10771,N_10252,N_9648);
and U10772 (N_10772,N_10121,N_9611);
or U10773 (N_10773,N_10173,N_10297);
or U10774 (N_10774,N_9796,N_9713);
xor U10775 (N_10775,N_9962,N_9666);
nor U10776 (N_10776,N_9910,N_9919);
and U10777 (N_10777,N_10094,N_9834);
and U10778 (N_10778,N_10131,N_9893);
nand U10779 (N_10779,N_10046,N_10020);
or U10780 (N_10780,N_9854,N_9722);
or U10781 (N_10781,N_9913,N_10326);
or U10782 (N_10782,N_9982,N_10087);
or U10783 (N_10783,N_9926,N_10101);
or U10784 (N_10784,N_10187,N_10108);
nand U10785 (N_10785,N_10075,N_10336);
xor U10786 (N_10786,N_10120,N_9895);
and U10787 (N_10787,N_9845,N_9850);
or U10788 (N_10788,N_9739,N_9976);
nand U10789 (N_10789,N_9759,N_9676);
or U10790 (N_10790,N_10342,N_10064);
nand U10791 (N_10791,N_9765,N_10086);
nand U10792 (N_10792,N_9894,N_10301);
nand U10793 (N_10793,N_10253,N_10180);
xor U10794 (N_10794,N_9838,N_10104);
nand U10795 (N_10795,N_9750,N_9667);
nor U10796 (N_10796,N_10196,N_9665);
or U10797 (N_10797,N_9858,N_10178);
and U10798 (N_10798,N_10296,N_10079);
and U10799 (N_10799,N_10067,N_10355);
xnor U10800 (N_10800,N_9921,N_10375);
xnor U10801 (N_10801,N_9934,N_9957);
nor U10802 (N_10802,N_9847,N_9671);
xor U10803 (N_10803,N_10178,N_9704);
xnor U10804 (N_10804,N_9907,N_9808);
nand U10805 (N_10805,N_10237,N_9804);
or U10806 (N_10806,N_10291,N_9624);
nor U10807 (N_10807,N_10355,N_9744);
nand U10808 (N_10808,N_9760,N_10301);
nand U10809 (N_10809,N_9883,N_9939);
and U10810 (N_10810,N_9841,N_10296);
xor U10811 (N_10811,N_10006,N_9912);
and U10812 (N_10812,N_10191,N_10192);
and U10813 (N_10813,N_9934,N_9674);
nand U10814 (N_10814,N_9764,N_9843);
and U10815 (N_10815,N_10080,N_9660);
or U10816 (N_10816,N_10200,N_9847);
or U10817 (N_10817,N_9702,N_9623);
nor U10818 (N_10818,N_10127,N_10047);
and U10819 (N_10819,N_9784,N_10225);
xor U10820 (N_10820,N_10080,N_10272);
nor U10821 (N_10821,N_9944,N_9806);
nand U10822 (N_10822,N_9605,N_10312);
or U10823 (N_10823,N_10029,N_9933);
and U10824 (N_10824,N_9932,N_10350);
nand U10825 (N_10825,N_9953,N_10366);
xor U10826 (N_10826,N_9940,N_9804);
nand U10827 (N_10827,N_10175,N_10261);
xnor U10828 (N_10828,N_10223,N_9826);
and U10829 (N_10829,N_10197,N_9674);
nand U10830 (N_10830,N_9877,N_10283);
or U10831 (N_10831,N_9716,N_9628);
xnor U10832 (N_10832,N_10394,N_10162);
nor U10833 (N_10833,N_10218,N_10216);
xor U10834 (N_10834,N_10164,N_9678);
or U10835 (N_10835,N_10263,N_10204);
or U10836 (N_10836,N_9950,N_9902);
nor U10837 (N_10837,N_9810,N_10295);
xor U10838 (N_10838,N_9860,N_10191);
and U10839 (N_10839,N_9770,N_10237);
or U10840 (N_10840,N_9606,N_9976);
nor U10841 (N_10841,N_9832,N_10268);
nor U10842 (N_10842,N_10356,N_10131);
or U10843 (N_10843,N_10096,N_9820);
nor U10844 (N_10844,N_10326,N_9606);
and U10845 (N_10845,N_10270,N_10314);
xor U10846 (N_10846,N_10104,N_9650);
nand U10847 (N_10847,N_9671,N_10283);
nor U10848 (N_10848,N_9800,N_9677);
or U10849 (N_10849,N_9790,N_10139);
and U10850 (N_10850,N_9744,N_9809);
xor U10851 (N_10851,N_10155,N_10047);
and U10852 (N_10852,N_9918,N_10271);
nor U10853 (N_10853,N_10104,N_10266);
or U10854 (N_10854,N_10014,N_9777);
nor U10855 (N_10855,N_9933,N_10377);
nand U10856 (N_10856,N_9813,N_10031);
nor U10857 (N_10857,N_10308,N_9902);
nor U10858 (N_10858,N_9972,N_10067);
or U10859 (N_10859,N_10397,N_9871);
and U10860 (N_10860,N_10066,N_9687);
nor U10861 (N_10861,N_10118,N_9638);
nand U10862 (N_10862,N_10299,N_10322);
xnor U10863 (N_10863,N_10293,N_10194);
and U10864 (N_10864,N_9965,N_9939);
nand U10865 (N_10865,N_9728,N_10274);
nand U10866 (N_10866,N_9758,N_9625);
nand U10867 (N_10867,N_9775,N_10083);
nor U10868 (N_10868,N_9718,N_10345);
nor U10869 (N_10869,N_9942,N_10390);
xor U10870 (N_10870,N_9635,N_9889);
nand U10871 (N_10871,N_9881,N_9964);
xnor U10872 (N_10872,N_9725,N_9931);
and U10873 (N_10873,N_9954,N_9653);
nor U10874 (N_10874,N_10154,N_10056);
nand U10875 (N_10875,N_10018,N_10131);
nor U10876 (N_10876,N_9846,N_9793);
or U10877 (N_10877,N_10049,N_10008);
and U10878 (N_10878,N_10082,N_10259);
or U10879 (N_10879,N_9899,N_9992);
or U10880 (N_10880,N_9778,N_9909);
xor U10881 (N_10881,N_10015,N_10308);
nand U10882 (N_10882,N_10356,N_9603);
or U10883 (N_10883,N_9796,N_10344);
and U10884 (N_10884,N_9610,N_10200);
nor U10885 (N_10885,N_10062,N_10329);
xnor U10886 (N_10886,N_10264,N_10242);
xor U10887 (N_10887,N_9619,N_10059);
nor U10888 (N_10888,N_10046,N_10350);
nor U10889 (N_10889,N_10147,N_9832);
xor U10890 (N_10890,N_9727,N_10254);
nand U10891 (N_10891,N_10323,N_9763);
and U10892 (N_10892,N_10341,N_9964);
or U10893 (N_10893,N_10383,N_10020);
or U10894 (N_10894,N_9631,N_9900);
and U10895 (N_10895,N_9712,N_10002);
nand U10896 (N_10896,N_10079,N_10349);
nand U10897 (N_10897,N_9611,N_10340);
or U10898 (N_10898,N_10014,N_9882);
nand U10899 (N_10899,N_9780,N_9827);
nor U10900 (N_10900,N_9849,N_9607);
or U10901 (N_10901,N_10346,N_10087);
nand U10902 (N_10902,N_10139,N_10361);
nor U10903 (N_10903,N_9665,N_9882);
nor U10904 (N_10904,N_10350,N_9641);
and U10905 (N_10905,N_10305,N_10028);
nor U10906 (N_10906,N_10288,N_10197);
or U10907 (N_10907,N_9778,N_9855);
nor U10908 (N_10908,N_9878,N_10388);
nor U10909 (N_10909,N_10280,N_10377);
xnor U10910 (N_10910,N_9685,N_9721);
xnor U10911 (N_10911,N_9923,N_9641);
and U10912 (N_10912,N_10102,N_9750);
and U10913 (N_10913,N_9952,N_10067);
nor U10914 (N_10914,N_9696,N_9756);
and U10915 (N_10915,N_9827,N_10215);
xnor U10916 (N_10916,N_9844,N_10101);
nor U10917 (N_10917,N_10024,N_10184);
and U10918 (N_10918,N_10166,N_10264);
or U10919 (N_10919,N_10322,N_9620);
nand U10920 (N_10920,N_9891,N_9869);
or U10921 (N_10921,N_9758,N_9840);
nand U10922 (N_10922,N_10197,N_10377);
xnor U10923 (N_10923,N_10038,N_9751);
nand U10924 (N_10924,N_10358,N_9627);
and U10925 (N_10925,N_9884,N_10320);
or U10926 (N_10926,N_9950,N_10263);
xnor U10927 (N_10927,N_10150,N_10030);
and U10928 (N_10928,N_10274,N_10353);
and U10929 (N_10929,N_10165,N_9976);
or U10930 (N_10930,N_9935,N_10051);
and U10931 (N_10931,N_9927,N_9677);
or U10932 (N_10932,N_10019,N_10234);
or U10933 (N_10933,N_9743,N_10345);
nand U10934 (N_10934,N_10068,N_10172);
or U10935 (N_10935,N_10168,N_9685);
and U10936 (N_10936,N_10213,N_10096);
xor U10937 (N_10937,N_10370,N_10367);
xnor U10938 (N_10938,N_10123,N_9792);
and U10939 (N_10939,N_10389,N_9823);
nor U10940 (N_10940,N_10105,N_9869);
and U10941 (N_10941,N_9772,N_9841);
or U10942 (N_10942,N_9899,N_10052);
nor U10943 (N_10943,N_10140,N_10215);
nor U10944 (N_10944,N_10365,N_10181);
xor U10945 (N_10945,N_9944,N_9618);
or U10946 (N_10946,N_10254,N_10164);
or U10947 (N_10947,N_10083,N_9726);
xnor U10948 (N_10948,N_10091,N_9778);
nand U10949 (N_10949,N_10320,N_10358);
nor U10950 (N_10950,N_9632,N_9696);
nand U10951 (N_10951,N_10274,N_10118);
or U10952 (N_10952,N_10032,N_9869);
nand U10953 (N_10953,N_9811,N_10327);
xor U10954 (N_10954,N_9630,N_10066);
or U10955 (N_10955,N_10087,N_9760);
xnor U10956 (N_10956,N_9987,N_10249);
nand U10957 (N_10957,N_9724,N_10344);
nor U10958 (N_10958,N_10221,N_10133);
and U10959 (N_10959,N_9831,N_10104);
or U10960 (N_10960,N_9644,N_9967);
or U10961 (N_10961,N_10116,N_10094);
or U10962 (N_10962,N_9713,N_9704);
and U10963 (N_10963,N_10091,N_10044);
and U10964 (N_10964,N_9761,N_10323);
or U10965 (N_10965,N_9671,N_9811);
nand U10966 (N_10966,N_9895,N_9801);
and U10967 (N_10967,N_10280,N_10041);
nand U10968 (N_10968,N_10102,N_10382);
or U10969 (N_10969,N_9618,N_10216);
nor U10970 (N_10970,N_9976,N_10231);
and U10971 (N_10971,N_9791,N_9626);
and U10972 (N_10972,N_10216,N_9743);
nand U10973 (N_10973,N_9886,N_9948);
xnor U10974 (N_10974,N_10058,N_10257);
nand U10975 (N_10975,N_9915,N_9854);
and U10976 (N_10976,N_9621,N_10169);
nand U10977 (N_10977,N_9996,N_9669);
and U10978 (N_10978,N_9715,N_9661);
xnor U10979 (N_10979,N_9875,N_9937);
xnor U10980 (N_10980,N_10381,N_10297);
and U10981 (N_10981,N_10342,N_9761);
or U10982 (N_10982,N_10351,N_10103);
or U10983 (N_10983,N_9778,N_9649);
xor U10984 (N_10984,N_10060,N_9932);
xor U10985 (N_10985,N_10267,N_10041);
xor U10986 (N_10986,N_10182,N_9792);
nand U10987 (N_10987,N_9910,N_10195);
and U10988 (N_10988,N_9664,N_10243);
nand U10989 (N_10989,N_10214,N_10171);
and U10990 (N_10990,N_10323,N_9632);
xor U10991 (N_10991,N_9929,N_9908);
nor U10992 (N_10992,N_9985,N_10236);
and U10993 (N_10993,N_9659,N_10308);
nor U10994 (N_10994,N_9749,N_10123);
nand U10995 (N_10995,N_9630,N_9967);
or U10996 (N_10996,N_9993,N_9977);
xor U10997 (N_10997,N_10236,N_10395);
and U10998 (N_10998,N_9798,N_9912);
nand U10999 (N_10999,N_10372,N_9636);
xnor U11000 (N_11000,N_10129,N_9737);
nand U11001 (N_11001,N_9967,N_10045);
or U11002 (N_11002,N_9965,N_9666);
and U11003 (N_11003,N_9718,N_10304);
nor U11004 (N_11004,N_10180,N_9693);
nor U11005 (N_11005,N_9827,N_9621);
and U11006 (N_11006,N_10123,N_9841);
and U11007 (N_11007,N_10313,N_9910);
and U11008 (N_11008,N_10017,N_10216);
nor U11009 (N_11009,N_9890,N_9744);
and U11010 (N_11010,N_9749,N_10169);
or U11011 (N_11011,N_9747,N_9859);
or U11012 (N_11012,N_9666,N_10032);
and U11013 (N_11013,N_10154,N_9889);
or U11014 (N_11014,N_10118,N_9642);
nor U11015 (N_11015,N_9876,N_10303);
or U11016 (N_11016,N_10101,N_9753);
nor U11017 (N_11017,N_9856,N_10027);
and U11018 (N_11018,N_10309,N_9653);
or U11019 (N_11019,N_10047,N_9767);
and U11020 (N_11020,N_10138,N_9625);
nand U11021 (N_11021,N_9733,N_10039);
nand U11022 (N_11022,N_9763,N_10333);
and U11023 (N_11023,N_10104,N_10267);
and U11024 (N_11024,N_9820,N_10087);
or U11025 (N_11025,N_9748,N_10142);
nor U11026 (N_11026,N_10011,N_10175);
nor U11027 (N_11027,N_10022,N_9633);
xnor U11028 (N_11028,N_10270,N_10068);
or U11029 (N_11029,N_10069,N_9984);
nand U11030 (N_11030,N_10081,N_9735);
and U11031 (N_11031,N_9812,N_10087);
xor U11032 (N_11032,N_10057,N_9669);
or U11033 (N_11033,N_10339,N_10249);
or U11034 (N_11034,N_9715,N_10234);
and U11035 (N_11035,N_9725,N_10269);
xnor U11036 (N_11036,N_9803,N_9624);
or U11037 (N_11037,N_9713,N_10359);
nor U11038 (N_11038,N_10362,N_9629);
nand U11039 (N_11039,N_9641,N_10105);
or U11040 (N_11040,N_9827,N_10369);
xor U11041 (N_11041,N_10305,N_10368);
xnor U11042 (N_11042,N_9953,N_10175);
nand U11043 (N_11043,N_10023,N_10136);
or U11044 (N_11044,N_10012,N_9895);
or U11045 (N_11045,N_10255,N_10342);
and U11046 (N_11046,N_10302,N_9983);
and U11047 (N_11047,N_9875,N_10264);
and U11048 (N_11048,N_10374,N_9767);
nand U11049 (N_11049,N_10124,N_10146);
nor U11050 (N_11050,N_9907,N_10078);
and U11051 (N_11051,N_9805,N_10089);
nor U11052 (N_11052,N_10093,N_10314);
nor U11053 (N_11053,N_9855,N_10123);
nor U11054 (N_11054,N_10269,N_10150);
and U11055 (N_11055,N_10221,N_9892);
xor U11056 (N_11056,N_10146,N_10030);
xnor U11057 (N_11057,N_10019,N_10139);
nand U11058 (N_11058,N_9788,N_10022);
nor U11059 (N_11059,N_9884,N_9769);
or U11060 (N_11060,N_10120,N_9627);
and U11061 (N_11061,N_9974,N_9891);
nand U11062 (N_11062,N_10221,N_9695);
xor U11063 (N_11063,N_9972,N_10330);
nor U11064 (N_11064,N_10184,N_9831);
nor U11065 (N_11065,N_10053,N_9668);
or U11066 (N_11066,N_9800,N_10017);
or U11067 (N_11067,N_10368,N_9706);
and U11068 (N_11068,N_9856,N_10101);
or U11069 (N_11069,N_10338,N_10007);
nand U11070 (N_11070,N_10216,N_10333);
xor U11071 (N_11071,N_10238,N_10312);
or U11072 (N_11072,N_9911,N_10370);
or U11073 (N_11073,N_10250,N_9872);
nand U11074 (N_11074,N_9997,N_9851);
nand U11075 (N_11075,N_10137,N_10224);
or U11076 (N_11076,N_10011,N_9747);
xnor U11077 (N_11077,N_9938,N_9668);
or U11078 (N_11078,N_9961,N_9691);
or U11079 (N_11079,N_10081,N_9648);
nor U11080 (N_11080,N_10376,N_10319);
or U11081 (N_11081,N_10392,N_9779);
or U11082 (N_11082,N_9740,N_10158);
nand U11083 (N_11083,N_9850,N_9810);
or U11084 (N_11084,N_9704,N_9865);
or U11085 (N_11085,N_9889,N_9913);
nor U11086 (N_11086,N_10046,N_9732);
xnor U11087 (N_11087,N_9659,N_10113);
nand U11088 (N_11088,N_10023,N_9937);
and U11089 (N_11089,N_9745,N_9726);
xor U11090 (N_11090,N_9816,N_9765);
or U11091 (N_11091,N_9635,N_9607);
nand U11092 (N_11092,N_9973,N_9844);
nor U11093 (N_11093,N_10245,N_10024);
or U11094 (N_11094,N_9648,N_9655);
nand U11095 (N_11095,N_10009,N_9756);
and U11096 (N_11096,N_9971,N_10173);
xnor U11097 (N_11097,N_10377,N_9830);
nor U11098 (N_11098,N_10217,N_9829);
nor U11099 (N_11099,N_10100,N_10012);
or U11100 (N_11100,N_10070,N_10009);
and U11101 (N_11101,N_10222,N_9696);
nand U11102 (N_11102,N_10222,N_10399);
nand U11103 (N_11103,N_10027,N_9651);
nand U11104 (N_11104,N_9826,N_10364);
and U11105 (N_11105,N_9823,N_9846);
and U11106 (N_11106,N_10176,N_9929);
and U11107 (N_11107,N_10222,N_9705);
nand U11108 (N_11108,N_10178,N_9659);
nand U11109 (N_11109,N_9823,N_9716);
nand U11110 (N_11110,N_9872,N_9818);
nor U11111 (N_11111,N_9639,N_10089);
and U11112 (N_11112,N_10208,N_9995);
or U11113 (N_11113,N_10006,N_9849);
and U11114 (N_11114,N_9735,N_9631);
or U11115 (N_11115,N_10188,N_10015);
nand U11116 (N_11116,N_9653,N_9731);
and U11117 (N_11117,N_10056,N_9853);
nand U11118 (N_11118,N_10364,N_10210);
nand U11119 (N_11119,N_10283,N_10060);
or U11120 (N_11120,N_10127,N_9891);
xnor U11121 (N_11121,N_10389,N_10074);
and U11122 (N_11122,N_10108,N_10054);
and U11123 (N_11123,N_10189,N_10125);
nor U11124 (N_11124,N_10351,N_9855);
or U11125 (N_11125,N_10018,N_10222);
or U11126 (N_11126,N_9983,N_10329);
nor U11127 (N_11127,N_10358,N_9871);
and U11128 (N_11128,N_10000,N_10332);
xnor U11129 (N_11129,N_9644,N_10131);
or U11130 (N_11130,N_9857,N_10154);
nor U11131 (N_11131,N_10054,N_10343);
and U11132 (N_11132,N_9962,N_10257);
nand U11133 (N_11133,N_9756,N_9842);
nor U11134 (N_11134,N_10300,N_10282);
and U11135 (N_11135,N_9672,N_10142);
nor U11136 (N_11136,N_10369,N_9770);
nor U11137 (N_11137,N_10342,N_9710);
xor U11138 (N_11138,N_10365,N_10234);
nor U11139 (N_11139,N_9665,N_9910);
and U11140 (N_11140,N_9641,N_10310);
and U11141 (N_11141,N_10322,N_10027);
nor U11142 (N_11142,N_9617,N_10032);
nand U11143 (N_11143,N_10259,N_10177);
xor U11144 (N_11144,N_9665,N_10088);
xor U11145 (N_11145,N_10286,N_9879);
or U11146 (N_11146,N_10153,N_10218);
xor U11147 (N_11147,N_10084,N_9991);
and U11148 (N_11148,N_9884,N_10220);
xor U11149 (N_11149,N_10091,N_9867);
xor U11150 (N_11150,N_10137,N_9711);
and U11151 (N_11151,N_10165,N_9766);
xor U11152 (N_11152,N_10101,N_9775);
or U11153 (N_11153,N_9690,N_10156);
xor U11154 (N_11154,N_9886,N_10082);
and U11155 (N_11155,N_10366,N_10002);
xnor U11156 (N_11156,N_9981,N_9739);
or U11157 (N_11157,N_9655,N_9716);
nor U11158 (N_11158,N_9693,N_10168);
or U11159 (N_11159,N_9858,N_9914);
nand U11160 (N_11160,N_9752,N_10361);
nor U11161 (N_11161,N_10017,N_9826);
and U11162 (N_11162,N_10050,N_9810);
nand U11163 (N_11163,N_9997,N_10181);
and U11164 (N_11164,N_10247,N_10066);
and U11165 (N_11165,N_9776,N_10390);
and U11166 (N_11166,N_9706,N_9646);
or U11167 (N_11167,N_10059,N_9919);
nor U11168 (N_11168,N_9692,N_10265);
and U11169 (N_11169,N_9914,N_9724);
or U11170 (N_11170,N_10152,N_9836);
nand U11171 (N_11171,N_10152,N_10012);
or U11172 (N_11172,N_9983,N_9889);
or U11173 (N_11173,N_10392,N_9943);
nor U11174 (N_11174,N_9610,N_10249);
or U11175 (N_11175,N_10015,N_9926);
and U11176 (N_11176,N_9767,N_10268);
and U11177 (N_11177,N_9979,N_10112);
nor U11178 (N_11178,N_10295,N_9644);
nor U11179 (N_11179,N_10089,N_10148);
or U11180 (N_11180,N_9927,N_9686);
nand U11181 (N_11181,N_9617,N_10085);
xor U11182 (N_11182,N_10244,N_10373);
or U11183 (N_11183,N_9832,N_10375);
and U11184 (N_11184,N_10274,N_10062);
xnor U11185 (N_11185,N_9961,N_10228);
xor U11186 (N_11186,N_9922,N_10045);
or U11187 (N_11187,N_10263,N_10105);
nor U11188 (N_11188,N_10198,N_10337);
nand U11189 (N_11189,N_10065,N_9738);
or U11190 (N_11190,N_10376,N_10217);
and U11191 (N_11191,N_10103,N_9990);
xnor U11192 (N_11192,N_9694,N_9685);
nand U11193 (N_11193,N_10009,N_10180);
and U11194 (N_11194,N_10342,N_10111);
and U11195 (N_11195,N_10191,N_9836);
xnor U11196 (N_11196,N_9957,N_10376);
nand U11197 (N_11197,N_9864,N_10278);
xor U11198 (N_11198,N_10382,N_9973);
or U11199 (N_11199,N_10005,N_10270);
nand U11200 (N_11200,N_10572,N_11183);
nor U11201 (N_11201,N_11050,N_10683);
and U11202 (N_11202,N_10780,N_10512);
nand U11203 (N_11203,N_10927,N_10619);
nor U11204 (N_11204,N_10941,N_10424);
nor U11205 (N_11205,N_10579,N_11110);
or U11206 (N_11206,N_10756,N_10674);
or U11207 (N_11207,N_10886,N_11017);
nor U11208 (N_11208,N_10670,N_11083);
xor U11209 (N_11209,N_10859,N_10848);
nand U11210 (N_11210,N_10461,N_11026);
nand U11211 (N_11211,N_10812,N_10602);
and U11212 (N_11212,N_10513,N_10934);
nor U11213 (N_11213,N_10928,N_10556);
and U11214 (N_11214,N_10895,N_10853);
and U11215 (N_11215,N_10977,N_10569);
xor U11216 (N_11216,N_10500,N_10457);
xnor U11217 (N_11217,N_10653,N_10975);
xor U11218 (N_11218,N_11071,N_10813);
or U11219 (N_11219,N_10963,N_10548);
nor U11220 (N_11220,N_10559,N_10519);
or U11221 (N_11221,N_11091,N_10531);
and U11222 (N_11222,N_10960,N_10875);
xnor U11223 (N_11223,N_10655,N_10772);
and U11224 (N_11224,N_10452,N_10511);
nor U11225 (N_11225,N_10899,N_10577);
xor U11226 (N_11226,N_10488,N_10789);
xnor U11227 (N_11227,N_10830,N_10405);
nor U11228 (N_11228,N_10465,N_10445);
xnor U11229 (N_11229,N_10764,N_10846);
and U11230 (N_11230,N_10586,N_11192);
nand U11231 (N_11231,N_10735,N_10665);
and U11232 (N_11232,N_10440,N_10643);
xnor U11233 (N_11233,N_10484,N_10404);
xor U11234 (N_11234,N_10797,N_10822);
nor U11235 (N_11235,N_10733,N_10721);
nand U11236 (N_11236,N_11157,N_10673);
nor U11237 (N_11237,N_10959,N_10821);
nand U11238 (N_11238,N_11094,N_10593);
nand U11239 (N_11239,N_10737,N_10738);
nor U11240 (N_11240,N_11182,N_10635);
nor U11241 (N_11241,N_10480,N_11152);
or U11242 (N_11242,N_10468,N_10744);
and U11243 (N_11243,N_10930,N_10545);
nand U11244 (N_11244,N_10757,N_10474);
nand U11245 (N_11245,N_10703,N_10459);
xnor U11246 (N_11246,N_10897,N_10451);
xor U11247 (N_11247,N_11117,N_10564);
nor U11248 (N_11248,N_11007,N_11029);
nand U11249 (N_11249,N_11045,N_11143);
or U11250 (N_11250,N_10419,N_10882);
or U11251 (N_11251,N_10770,N_10801);
or U11252 (N_11252,N_10908,N_10605);
nand U11253 (N_11253,N_10565,N_10932);
nand U11254 (N_11254,N_11019,N_11076);
and U11255 (N_11255,N_10456,N_10496);
nor U11256 (N_11256,N_11008,N_10972);
nand U11257 (N_11257,N_11147,N_11006);
or U11258 (N_11258,N_10811,N_10948);
or U11259 (N_11259,N_10516,N_10621);
and U11260 (N_11260,N_10534,N_10633);
nand U11261 (N_11261,N_10919,N_10486);
nand U11262 (N_11262,N_10539,N_10431);
nand U11263 (N_11263,N_11100,N_10610);
or U11264 (N_11264,N_10755,N_10408);
and U11265 (N_11265,N_10547,N_10438);
nor U11266 (N_11266,N_10667,N_10464);
or U11267 (N_11267,N_11039,N_11175);
xnor U11268 (N_11268,N_11164,N_10551);
nand U11269 (N_11269,N_11186,N_11023);
or U11270 (N_11270,N_11155,N_10971);
nor U11271 (N_11271,N_10810,N_10788);
xnor U11272 (N_11272,N_10428,N_11005);
xor U11273 (N_11273,N_10482,N_10767);
nor U11274 (N_11274,N_10649,N_10689);
xor U11275 (N_11275,N_10728,N_11095);
nand U11276 (N_11276,N_10924,N_11024);
or U11277 (N_11277,N_11139,N_10499);
nand U11278 (N_11278,N_11044,N_10825);
or U11279 (N_11279,N_10759,N_10967);
and U11280 (N_11280,N_10809,N_10422);
xnor U11281 (N_11281,N_11196,N_10437);
nand U11282 (N_11282,N_10656,N_10659);
nand U11283 (N_11283,N_10877,N_10820);
or U11284 (N_11284,N_10563,N_10682);
nand U11285 (N_11285,N_10947,N_10557);
nor U11286 (N_11286,N_10447,N_11031);
nor U11287 (N_11287,N_10760,N_10630);
and U11288 (N_11288,N_10920,N_10916);
nand U11289 (N_11289,N_10640,N_10537);
xnor U11290 (N_11290,N_10543,N_11123);
or U11291 (N_11291,N_10453,N_10961);
nand U11292 (N_11292,N_10792,N_10815);
xnor U11293 (N_11293,N_11114,N_10997);
nand U11294 (N_11294,N_11135,N_10898);
and U11295 (N_11295,N_10976,N_10439);
nor U11296 (N_11296,N_10595,N_11108);
xnor U11297 (N_11297,N_10714,N_10902);
and U11298 (N_11298,N_10742,N_11042);
nor U11299 (N_11299,N_10631,N_10420);
and U11300 (N_11300,N_10858,N_10803);
nand U11301 (N_11301,N_11104,N_10623);
xor U11302 (N_11302,N_10485,N_10890);
nand U11303 (N_11303,N_11122,N_10717);
xnor U11304 (N_11304,N_10910,N_10435);
nand U11305 (N_11305,N_10860,N_11011);
nand U11306 (N_11306,N_10826,N_10805);
or U11307 (N_11307,N_10964,N_10968);
nand U11308 (N_11308,N_10597,N_10831);
or U11309 (N_11309,N_11133,N_11103);
and U11310 (N_11310,N_11158,N_10817);
or U11311 (N_11311,N_10505,N_10974);
xnor U11312 (N_11312,N_10841,N_10998);
and U11313 (N_11313,N_11184,N_11113);
nand U11314 (N_11314,N_10795,N_10926);
xnor U11315 (N_11315,N_10995,N_10679);
nor U11316 (N_11316,N_10704,N_10931);
xnor U11317 (N_11317,N_10582,N_10982);
nand U11318 (N_11318,N_11199,N_10654);
or U11319 (N_11319,N_10617,N_11111);
and U11320 (N_11320,N_11102,N_10680);
nor U11321 (N_11321,N_11025,N_10751);
or U11322 (N_11322,N_10608,N_11087);
nand U11323 (N_11323,N_10601,N_10632);
or U11324 (N_11324,N_11156,N_10802);
xnor U11325 (N_11325,N_11030,N_11150);
nand U11326 (N_11326,N_10940,N_10473);
or U11327 (N_11327,N_10466,N_10449);
xor U11328 (N_11328,N_10868,N_11086);
xor U11329 (N_11329,N_10552,N_10962);
nand U11330 (N_11330,N_10896,N_10829);
and U11331 (N_11331,N_10965,N_11073);
nand U11332 (N_11332,N_10791,N_10423);
and U11333 (N_11333,N_10503,N_10672);
and U11334 (N_11334,N_10695,N_10973);
and U11335 (N_11335,N_10410,N_11062);
nor U11336 (N_11336,N_10720,N_10514);
or U11337 (N_11337,N_10638,N_10685);
nand U11338 (N_11338,N_11079,N_10869);
nor U11339 (N_11339,N_11173,N_10571);
nand U11340 (N_11340,N_11093,N_10598);
or U11341 (N_11341,N_10884,N_10937);
or U11342 (N_11342,N_10528,N_10842);
nor U11343 (N_11343,N_10660,N_10710);
and U11344 (N_11344,N_10736,N_10991);
and U11345 (N_11345,N_11161,N_10994);
or U11346 (N_11346,N_10561,N_10416);
and U11347 (N_11347,N_10690,N_10578);
nand U11348 (N_11348,N_10850,N_11036);
or U11349 (N_11349,N_10828,N_10814);
nor U11350 (N_11350,N_10743,N_10732);
nand U11351 (N_11351,N_11119,N_11098);
or U11352 (N_11352,N_10584,N_11109);
or U11353 (N_11353,N_11193,N_10709);
nor U11354 (N_11354,N_10442,N_10783);
and U11355 (N_11355,N_10527,N_10824);
or U11356 (N_11356,N_10495,N_10705);
xor U11357 (N_11357,N_10723,N_10470);
nor U11358 (N_11358,N_10498,N_11134);
xnor U11359 (N_11359,N_11034,N_11129);
and U11360 (N_11360,N_10872,N_10936);
or U11361 (N_11361,N_11185,N_10980);
or U11362 (N_11362,N_10804,N_10870);
xor U11363 (N_11363,N_10819,N_10574);
or U11364 (N_11364,N_10827,N_11015);
and U11365 (N_11365,N_11027,N_10583);
nand U11366 (N_11366,N_10502,N_10526);
and U11367 (N_11367,N_10581,N_10427);
or U11368 (N_11368,N_11187,N_11021);
xnor U11369 (N_11369,N_11101,N_10530);
nand U11370 (N_11370,N_11174,N_11096);
nor U11371 (N_11371,N_10887,N_10544);
xor U11372 (N_11372,N_10989,N_10818);
nand U11373 (N_11373,N_11099,N_11066);
or U11374 (N_11374,N_10957,N_10587);
xor U11375 (N_11375,N_11009,N_10487);
or U11376 (N_11376,N_10462,N_11142);
xnor U11377 (N_11377,N_10433,N_10712);
nor U11378 (N_11378,N_11162,N_10693);
or U11379 (N_11379,N_10892,N_10769);
nor U11380 (N_11380,N_11120,N_10535);
and U11381 (N_11381,N_11040,N_10532);
xnor U11382 (N_11382,N_10835,N_10648);
nand U11383 (N_11383,N_11057,N_11153);
or U11384 (N_11384,N_11140,N_10677);
nor U11385 (N_11385,N_10634,N_11198);
nand U11386 (N_11386,N_10592,N_10777);
or U11387 (N_11387,N_11128,N_11177);
nor U11388 (N_11388,N_10430,N_10836);
and U11389 (N_11389,N_10701,N_10686);
or U11390 (N_11390,N_11061,N_11178);
nor U11391 (N_11391,N_10722,N_10696);
and U11392 (N_11392,N_10663,N_10506);
xnor U11393 (N_11393,N_10412,N_10774);
nor U11394 (N_11394,N_10874,N_10807);
and U11395 (N_11395,N_11126,N_10675);
or U11396 (N_11396,N_11059,N_10477);
xor U11397 (N_11397,N_10808,N_10984);
or U11398 (N_11398,N_10901,N_10851);
nor U11399 (N_11399,N_10861,N_10881);
xor U11400 (N_11400,N_10585,N_10854);
or U11401 (N_11401,N_11176,N_10713);
xnor U11402 (N_11402,N_10981,N_10407);
nand U11403 (N_11403,N_10450,N_10411);
nor U11404 (N_11404,N_11188,N_11127);
and U11405 (N_11405,N_10469,N_10522);
xor U11406 (N_11406,N_10515,N_10951);
and U11407 (N_11407,N_10642,N_10700);
and U11408 (N_11408,N_10894,N_10871);
xor U11409 (N_11409,N_10730,N_10922);
and U11410 (N_11410,N_10956,N_10766);
and U11411 (N_11411,N_11166,N_10843);
nand U11412 (N_11412,N_10490,N_10970);
nand U11413 (N_11413,N_10987,N_10501);
xor U11414 (N_11414,N_10504,N_11072);
nand U11415 (N_11415,N_10876,N_10523);
and U11416 (N_11416,N_11179,N_10454);
or U11417 (N_11417,N_11180,N_11171);
or U11418 (N_11418,N_10923,N_10400);
nand U11419 (N_11419,N_10553,N_10988);
or U11420 (N_11420,N_11085,N_10839);
nand U11421 (N_11421,N_11190,N_11130);
xnor U11422 (N_11422,N_10911,N_10691);
or U11423 (N_11423,N_10570,N_10865);
or U11424 (N_11424,N_11075,N_10857);
and U11425 (N_11425,N_10460,N_10576);
nand U11426 (N_11426,N_10588,N_11001);
or U11427 (N_11427,N_10758,N_11089);
nor U11428 (N_11428,N_10731,N_10879);
nor U11429 (N_11429,N_10845,N_10999);
or U11430 (N_11430,N_11052,N_10517);
nor U11431 (N_11431,N_10694,N_10699);
xnor U11432 (N_11432,N_10942,N_10671);
or U11433 (N_11433,N_10580,N_10426);
and U11434 (N_11434,N_11049,N_11090);
nor U11435 (N_11435,N_11149,N_11078);
and U11436 (N_11436,N_10607,N_10939);
or U11437 (N_11437,N_11022,N_10955);
xnor U11438 (N_11438,N_10418,N_10775);
and U11439 (N_11439,N_11004,N_10429);
nor U11440 (N_11440,N_10609,N_10915);
nand U11441 (N_11441,N_10668,N_10873);
nor U11442 (N_11442,N_10885,N_11195);
and U11443 (N_11443,N_10778,N_10935);
xnor U11444 (N_11444,N_10866,N_10856);
nor U11445 (N_11445,N_10837,N_10944);
and U11446 (N_11446,N_10785,N_10929);
or U11447 (N_11447,N_10888,N_10855);
or U11448 (N_11448,N_10542,N_10520);
xor U11449 (N_11449,N_10666,N_10463);
nor U11450 (N_11450,N_10616,N_10840);
nor U11451 (N_11451,N_11154,N_10844);
nor U11452 (N_11452,N_10953,N_10799);
xor U11453 (N_11453,N_10753,N_11016);
nand U11454 (N_11454,N_10421,N_10492);
xor U11455 (N_11455,N_10471,N_11028);
nor U11456 (N_11456,N_10952,N_10906);
or U11457 (N_11457,N_11146,N_10455);
or U11458 (N_11458,N_10446,N_10697);
nor U11459 (N_11459,N_10626,N_11170);
and U11460 (N_11460,N_10636,N_10741);
nor U11461 (N_11461,N_10750,N_10567);
nor U11462 (N_11462,N_11063,N_11084);
or U11463 (N_11463,N_10917,N_11197);
xor U11464 (N_11464,N_11013,N_10590);
or U11465 (N_11465,N_10692,N_10533);
and U11466 (N_11466,N_10637,N_11065);
and U11467 (N_11467,N_10776,N_10681);
or U11468 (N_11468,N_10414,N_10734);
xnor U11469 (N_11469,N_10483,N_10779);
or U11470 (N_11470,N_10624,N_10688);
xnor U11471 (N_11471,N_11000,N_10669);
nor U11472 (N_11472,N_10508,N_10925);
and U11473 (N_11473,N_10641,N_10740);
nand U11474 (N_11474,N_11132,N_10432);
xnor U11475 (N_11475,N_10611,N_10706);
or U11476 (N_11476,N_11080,N_10990);
and U11477 (N_11477,N_11136,N_10662);
nand U11478 (N_11478,N_10747,N_10782);
or U11479 (N_11479,N_10707,N_10847);
xnor U11480 (N_11480,N_11070,N_10794);
nand U11481 (N_11481,N_10625,N_10762);
and U11482 (N_11482,N_10541,N_10415);
xnor U11483 (N_11483,N_10644,N_10497);
nand U11484 (N_11484,N_10784,N_10752);
nand U11485 (N_11485,N_10443,N_10768);
xnor U11486 (N_11486,N_10949,N_10684);
nand U11487 (N_11487,N_10651,N_10676);
nor U11488 (N_11488,N_10748,N_10629);
nor U11489 (N_11489,N_10979,N_11032);
or U11490 (N_11490,N_10467,N_10652);
or U11491 (N_11491,N_11163,N_10945);
nand U11492 (N_11492,N_11038,N_10773);
or U11493 (N_11493,N_10554,N_10664);
nand U11494 (N_11494,N_11003,N_10893);
nor U11495 (N_11495,N_10904,N_11067);
nor U11496 (N_11496,N_10606,N_11053);
nor U11497 (N_11497,N_10509,N_10614);
and U11498 (N_11498,N_10800,N_10798);
xnor U11499 (N_11499,N_10568,N_11068);
or U11500 (N_11500,N_11125,N_11033);
nand U11501 (N_11501,N_10479,N_10627);
xnor U11502 (N_11502,N_10529,N_11082);
nor U11503 (N_11503,N_10823,N_11159);
or U11504 (N_11504,N_10838,N_10604);
xor U11505 (N_11505,N_11112,N_11048);
nor U11506 (N_11506,N_10986,N_11077);
nand U11507 (N_11507,N_11035,N_10903);
nand U11508 (N_11508,N_10746,N_10536);
xor U11509 (N_11509,N_10596,N_10978);
and U11510 (N_11510,N_10719,N_11131);
nand U11511 (N_11511,N_10754,N_11124);
or U11512 (N_11512,N_10862,N_10954);
xor U11513 (N_11513,N_10992,N_10763);
nor U11514 (N_11514,N_11144,N_11115);
and U11515 (N_11515,N_10540,N_10786);
nand U11516 (N_11516,N_10781,N_11056);
nand U11517 (N_11517,N_10489,N_11055);
nand U11518 (N_11518,N_11064,N_10761);
xor U11519 (N_11519,N_10806,N_10555);
xor U11520 (N_11520,N_11116,N_11141);
nand U11521 (N_11521,N_10969,N_10434);
and U11522 (N_11522,N_10646,N_10628);
nand U11523 (N_11523,N_11088,N_10613);
nor U11524 (N_11524,N_10771,N_11181);
and U11525 (N_11525,N_11041,N_10448);
or U11526 (N_11526,N_10863,N_10510);
or U11527 (N_11527,N_10864,N_10562);
and U11528 (N_11528,N_10612,N_10657);
xnor U11529 (N_11529,N_11194,N_10725);
xnor U11530 (N_11530,N_11145,N_10639);
nor U11531 (N_11531,N_10406,N_10711);
and U11532 (N_11532,N_11169,N_10594);
and U11533 (N_11533,N_10417,N_11121);
and U11534 (N_11534,N_10524,N_10933);
nor U11535 (N_11535,N_10891,N_10475);
or U11536 (N_11536,N_10834,N_11172);
nor U11537 (N_11537,N_10918,N_10726);
or U11538 (N_11538,N_10441,N_11107);
and U11539 (N_11539,N_10718,N_10600);
nand U11540 (N_11540,N_10790,N_10476);
nor U11541 (N_11541,N_10745,N_10938);
xor U11542 (N_11542,N_10494,N_10481);
and U11543 (N_11543,N_10425,N_11189);
nand U11544 (N_11544,N_10615,N_10907);
nand U11545 (N_11545,N_10793,N_10702);
nand U11546 (N_11546,N_10724,N_10727);
and U11547 (N_11547,N_10716,N_11037);
nor U11548 (N_11548,N_10566,N_11191);
nand U11549 (N_11549,N_10983,N_11010);
nor U11550 (N_11550,N_10889,N_11137);
xnor U11551 (N_11551,N_11018,N_11014);
nand U11552 (N_11552,N_10436,N_10589);
nor U11553 (N_11553,N_10645,N_11051);
xor U11554 (N_11554,N_10966,N_10913);
xnor U11555 (N_11555,N_10787,N_10958);
xor U11556 (N_11556,N_10914,N_10573);
and U11557 (N_11557,N_10912,N_10715);
and U11558 (N_11558,N_10849,N_10878);
and U11559 (N_11559,N_10900,N_11097);
and U11560 (N_11560,N_10402,N_10993);
xor U11561 (N_11561,N_10729,N_10796);
nor U11562 (N_11562,N_10921,N_10525);
nor U11563 (N_11563,N_11043,N_10620);
and U11564 (N_11564,N_11012,N_11138);
xnor U11565 (N_11565,N_11106,N_10618);
xor U11566 (N_11566,N_10658,N_10943);
nor U11567 (N_11567,N_10950,N_10996);
nor U11568 (N_11568,N_11105,N_11047);
and U11569 (N_11569,N_10599,N_10401);
nand U11570 (N_11570,N_11081,N_10905);
nor U11571 (N_11571,N_11167,N_10852);
xnor U11572 (N_11572,N_11020,N_10946);
nand U11573 (N_11573,N_11118,N_10521);
xor U11574 (N_11574,N_11060,N_10493);
nand U11575 (N_11575,N_10546,N_10409);
or U11576 (N_11576,N_11058,N_10749);
and U11577 (N_11577,N_10647,N_10765);
and U11578 (N_11578,N_11002,N_10867);
nor U11579 (N_11579,N_10833,N_11168);
nor U11580 (N_11580,N_10413,N_10603);
nand U11581 (N_11581,N_11069,N_10708);
and U11582 (N_11582,N_10650,N_10549);
or U11583 (N_11583,N_10560,N_10444);
or U11584 (N_11584,N_10678,N_10883);
nor U11585 (N_11585,N_10403,N_10816);
xor U11586 (N_11586,N_10538,N_10518);
xnor U11587 (N_11587,N_10507,N_10458);
xor U11588 (N_11588,N_10739,N_11046);
nand U11589 (N_11589,N_10880,N_10575);
nor U11590 (N_11590,N_10661,N_10491);
nor U11591 (N_11591,N_11054,N_11074);
or U11592 (N_11592,N_10558,N_11092);
nor U11593 (N_11593,N_10698,N_10622);
nand U11594 (N_11594,N_11160,N_10591);
nor U11595 (N_11595,N_10478,N_10985);
nor U11596 (N_11596,N_10687,N_11148);
xor U11597 (N_11597,N_10832,N_11151);
xor U11598 (N_11598,N_10550,N_10472);
and U11599 (N_11599,N_10909,N_11165);
nand U11600 (N_11600,N_10733,N_10955);
xnor U11601 (N_11601,N_10727,N_10983);
nand U11602 (N_11602,N_10494,N_10706);
or U11603 (N_11603,N_10593,N_10671);
and U11604 (N_11604,N_11017,N_10807);
nor U11605 (N_11605,N_10890,N_10957);
nand U11606 (N_11606,N_11012,N_10811);
nand U11607 (N_11607,N_11160,N_11127);
or U11608 (N_11608,N_10829,N_10995);
xor U11609 (N_11609,N_10663,N_10548);
and U11610 (N_11610,N_10582,N_10616);
and U11611 (N_11611,N_10509,N_11175);
and U11612 (N_11612,N_10690,N_11160);
or U11613 (N_11613,N_10718,N_10744);
nor U11614 (N_11614,N_10716,N_10811);
nor U11615 (N_11615,N_11187,N_10957);
nand U11616 (N_11616,N_10420,N_10586);
and U11617 (N_11617,N_11130,N_10520);
nand U11618 (N_11618,N_11153,N_10800);
and U11619 (N_11619,N_10968,N_10547);
and U11620 (N_11620,N_11092,N_11060);
nor U11621 (N_11621,N_11100,N_10775);
or U11622 (N_11622,N_10621,N_10640);
nand U11623 (N_11623,N_10565,N_10676);
nand U11624 (N_11624,N_10582,N_10467);
nor U11625 (N_11625,N_11158,N_10639);
and U11626 (N_11626,N_10954,N_10757);
and U11627 (N_11627,N_11096,N_10445);
or U11628 (N_11628,N_10407,N_10841);
xnor U11629 (N_11629,N_10836,N_11003);
or U11630 (N_11630,N_10608,N_10815);
nor U11631 (N_11631,N_10746,N_10552);
xor U11632 (N_11632,N_10901,N_10678);
and U11633 (N_11633,N_10450,N_10567);
nand U11634 (N_11634,N_10653,N_10998);
or U11635 (N_11635,N_10877,N_10499);
nand U11636 (N_11636,N_10825,N_10945);
and U11637 (N_11637,N_10455,N_10622);
xor U11638 (N_11638,N_10823,N_10552);
xor U11639 (N_11639,N_11110,N_10448);
nor U11640 (N_11640,N_10490,N_11013);
or U11641 (N_11641,N_10462,N_11025);
xnor U11642 (N_11642,N_11081,N_10993);
xnor U11643 (N_11643,N_11193,N_11046);
xnor U11644 (N_11644,N_10939,N_11162);
nor U11645 (N_11645,N_10942,N_10931);
xor U11646 (N_11646,N_11036,N_10460);
nor U11647 (N_11647,N_10544,N_11049);
and U11648 (N_11648,N_10568,N_11166);
nand U11649 (N_11649,N_10435,N_11025);
nor U11650 (N_11650,N_10657,N_11017);
nand U11651 (N_11651,N_11038,N_10792);
nor U11652 (N_11652,N_10982,N_10646);
nand U11653 (N_11653,N_10908,N_10817);
and U11654 (N_11654,N_11166,N_10642);
nand U11655 (N_11655,N_10619,N_10845);
nor U11656 (N_11656,N_10422,N_10945);
or U11657 (N_11657,N_10425,N_10940);
nor U11658 (N_11658,N_10948,N_10856);
and U11659 (N_11659,N_10582,N_10676);
or U11660 (N_11660,N_10680,N_11162);
nand U11661 (N_11661,N_11168,N_11010);
xnor U11662 (N_11662,N_10909,N_10974);
nor U11663 (N_11663,N_10723,N_10536);
and U11664 (N_11664,N_10975,N_10707);
or U11665 (N_11665,N_10405,N_10531);
nor U11666 (N_11666,N_10692,N_10626);
or U11667 (N_11667,N_10890,N_10459);
and U11668 (N_11668,N_10793,N_10692);
and U11669 (N_11669,N_10829,N_10425);
or U11670 (N_11670,N_10668,N_10473);
nor U11671 (N_11671,N_11157,N_10969);
or U11672 (N_11672,N_11071,N_11085);
xor U11673 (N_11673,N_10646,N_10639);
and U11674 (N_11674,N_11118,N_11101);
xnor U11675 (N_11675,N_10660,N_10609);
xnor U11676 (N_11676,N_10869,N_10845);
nor U11677 (N_11677,N_10482,N_10443);
or U11678 (N_11678,N_10982,N_10502);
and U11679 (N_11679,N_10484,N_10642);
nor U11680 (N_11680,N_10509,N_10504);
xnor U11681 (N_11681,N_10438,N_10520);
nand U11682 (N_11682,N_10724,N_10599);
and U11683 (N_11683,N_10927,N_10565);
or U11684 (N_11684,N_10555,N_10974);
nor U11685 (N_11685,N_11111,N_11085);
and U11686 (N_11686,N_11121,N_10874);
and U11687 (N_11687,N_10650,N_10959);
or U11688 (N_11688,N_10570,N_10886);
xnor U11689 (N_11689,N_10806,N_11101);
nor U11690 (N_11690,N_10796,N_10609);
nor U11691 (N_11691,N_10800,N_10606);
or U11692 (N_11692,N_10657,N_10818);
nand U11693 (N_11693,N_10666,N_10926);
nand U11694 (N_11694,N_10935,N_10771);
nand U11695 (N_11695,N_10984,N_11038);
or U11696 (N_11696,N_10958,N_10986);
nor U11697 (N_11697,N_11028,N_10989);
or U11698 (N_11698,N_10441,N_10414);
xor U11699 (N_11699,N_10740,N_11044);
nand U11700 (N_11700,N_10454,N_10581);
xor U11701 (N_11701,N_10500,N_10999);
and U11702 (N_11702,N_11194,N_11094);
nand U11703 (N_11703,N_10511,N_11155);
nor U11704 (N_11704,N_11093,N_10666);
nand U11705 (N_11705,N_11037,N_10853);
nor U11706 (N_11706,N_10492,N_10413);
or U11707 (N_11707,N_10966,N_10897);
nor U11708 (N_11708,N_10732,N_10769);
and U11709 (N_11709,N_10674,N_10660);
xnor U11710 (N_11710,N_10853,N_11020);
or U11711 (N_11711,N_10855,N_10619);
nand U11712 (N_11712,N_11083,N_10611);
xnor U11713 (N_11713,N_10536,N_10808);
nand U11714 (N_11714,N_10858,N_11020);
xor U11715 (N_11715,N_10569,N_11118);
nor U11716 (N_11716,N_10421,N_10803);
and U11717 (N_11717,N_10633,N_10904);
xor U11718 (N_11718,N_10996,N_10400);
or U11719 (N_11719,N_10617,N_10589);
xor U11720 (N_11720,N_11095,N_10612);
and U11721 (N_11721,N_10600,N_10763);
nand U11722 (N_11722,N_11130,N_11030);
or U11723 (N_11723,N_11098,N_10722);
nor U11724 (N_11724,N_10765,N_10916);
nor U11725 (N_11725,N_10856,N_10715);
nor U11726 (N_11726,N_11014,N_10561);
nand U11727 (N_11727,N_10715,N_10708);
or U11728 (N_11728,N_10475,N_10929);
and U11729 (N_11729,N_10563,N_10820);
nor U11730 (N_11730,N_10742,N_10649);
or U11731 (N_11731,N_10731,N_10434);
or U11732 (N_11732,N_10888,N_10623);
nor U11733 (N_11733,N_10498,N_10529);
nand U11734 (N_11734,N_10772,N_10708);
or U11735 (N_11735,N_10457,N_10467);
nand U11736 (N_11736,N_10761,N_10706);
nor U11737 (N_11737,N_10566,N_10567);
nand U11738 (N_11738,N_10769,N_11015);
and U11739 (N_11739,N_10421,N_11070);
and U11740 (N_11740,N_10655,N_10565);
nor U11741 (N_11741,N_10744,N_10502);
xor U11742 (N_11742,N_10928,N_10830);
and U11743 (N_11743,N_10543,N_11093);
xor U11744 (N_11744,N_10512,N_11012);
and U11745 (N_11745,N_10917,N_11028);
nor U11746 (N_11746,N_11143,N_11015);
and U11747 (N_11747,N_10605,N_10884);
and U11748 (N_11748,N_11136,N_10775);
xor U11749 (N_11749,N_10605,N_10816);
nand U11750 (N_11750,N_10840,N_10845);
and U11751 (N_11751,N_10633,N_10632);
and U11752 (N_11752,N_10613,N_10910);
nor U11753 (N_11753,N_10651,N_10892);
nor U11754 (N_11754,N_10801,N_10526);
xor U11755 (N_11755,N_10460,N_10943);
nor U11756 (N_11756,N_11117,N_10786);
and U11757 (N_11757,N_11097,N_10941);
or U11758 (N_11758,N_10696,N_11088);
nand U11759 (N_11759,N_10676,N_10835);
nor U11760 (N_11760,N_10857,N_10781);
nor U11761 (N_11761,N_10838,N_10958);
xnor U11762 (N_11762,N_11050,N_10537);
and U11763 (N_11763,N_11056,N_11176);
and U11764 (N_11764,N_10630,N_10884);
nor U11765 (N_11765,N_10901,N_10976);
or U11766 (N_11766,N_10854,N_10693);
xnor U11767 (N_11767,N_10907,N_10725);
xnor U11768 (N_11768,N_10887,N_10447);
xor U11769 (N_11769,N_10654,N_10728);
and U11770 (N_11770,N_10952,N_10770);
nand U11771 (N_11771,N_11154,N_11002);
xor U11772 (N_11772,N_10427,N_11019);
and U11773 (N_11773,N_10954,N_10435);
nand U11774 (N_11774,N_10785,N_11082);
and U11775 (N_11775,N_10696,N_10752);
and U11776 (N_11776,N_10554,N_10537);
nor U11777 (N_11777,N_10742,N_10752);
nand U11778 (N_11778,N_10600,N_10965);
xor U11779 (N_11779,N_10999,N_11141);
and U11780 (N_11780,N_10758,N_10627);
nand U11781 (N_11781,N_10971,N_10960);
or U11782 (N_11782,N_10849,N_10755);
or U11783 (N_11783,N_11140,N_10648);
nor U11784 (N_11784,N_10798,N_10841);
and U11785 (N_11785,N_10522,N_10823);
or U11786 (N_11786,N_10947,N_10831);
and U11787 (N_11787,N_10965,N_10468);
or U11788 (N_11788,N_11030,N_10604);
and U11789 (N_11789,N_10924,N_11145);
nor U11790 (N_11790,N_10979,N_10936);
nand U11791 (N_11791,N_10510,N_10989);
nand U11792 (N_11792,N_10704,N_11104);
xor U11793 (N_11793,N_11010,N_11112);
or U11794 (N_11794,N_10768,N_11092);
and U11795 (N_11795,N_10403,N_10834);
or U11796 (N_11796,N_10719,N_10989);
nor U11797 (N_11797,N_10665,N_10840);
and U11798 (N_11798,N_10639,N_10935);
or U11799 (N_11799,N_10842,N_11085);
nand U11800 (N_11800,N_10581,N_10647);
or U11801 (N_11801,N_10790,N_10766);
and U11802 (N_11802,N_10769,N_10983);
or U11803 (N_11803,N_10586,N_11016);
xnor U11804 (N_11804,N_11166,N_11036);
nor U11805 (N_11805,N_10630,N_11071);
nand U11806 (N_11806,N_10969,N_10573);
nand U11807 (N_11807,N_10926,N_11034);
nor U11808 (N_11808,N_10401,N_11037);
or U11809 (N_11809,N_10906,N_10511);
nor U11810 (N_11810,N_10436,N_10692);
nor U11811 (N_11811,N_10827,N_11160);
xnor U11812 (N_11812,N_10770,N_10680);
xor U11813 (N_11813,N_11011,N_10945);
nor U11814 (N_11814,N_10811,N_10574);
nor U11815 (N_11815,N_10952,N_10635);
xor U11816 (N_11816,N_10785,N_10673);
nor U11817 (N_11817,N_10506,N_10616);
nand U11818 (N_11818,N_10792,N_10406);
xnor U11819 (N_11819,N_10732,N_10576);
nand U11820 (N_11820,N_10991,N_11084);
or U11821 (N_11821,N_10443,N_10845);
nand U11822 (N_11822,N_10879,N_11140);
nand U11823 (N_11823,N_10749,N_10475);
nand U11824 (N_11824,N_10451,N_10638);
xor U11825 (N_11825,N_11026,N_10901);
xor U11826 (N_11826,N_10719,N_10713);
or U11827 (N_11827,N_10718,N_11137);
or U11828 (N_11828,N_10836,N_10716);
xnor U11829 (N_11829,N_10541,N_10796);
xnor U11830 (N_11830,N_10961,N_10412);
and U11831 (N_11831,N_10682,N_10649);
nand U11832 (N_11832,N_10459,N_11104);
and U11833 (N_11833,N_10508,N_11193);
or U11834 (N_11834,N_10567,N_10440);
nand U11835 (N_11835,N_10746,N_11082);
and U11836 (N_11836,N_11029,N_10703);
nand U11837 (N_11837,N_11178,N_10708);
nand U11838 (N_11838,N_10808,N_10845);
or U11839 (N_11839,N_11056,N_10420);
nand U11840 (N_11840,N_11132,N_10598);
and U11841 (N_11841,N_10531,N_10814);
nand U11842 (N_11842,N_10487,N_10832);
xnor U11843 (N_11843,N_11105,N_10685);
and U11844 (N_11844,N_11198,N_10577);
xnor U11845 (N_11845,N_10900,N_11000);
or U11846 (N_11846,N_10517,N_10773);
nor U11847 (N_11847,N_10745,N_10770);
nor U11848 (N_11848,N_10790,N_10603);
xnor U11849 (N_11849,N_10742,N_10610);
or U11850 (N_11850,N_10960,N_11147);
or U11851 (N_11851,N_10776,N_10664);
nor U11852 (N_11852,N_10823,N_10672);
and U11853 (N_11853,N_11002,N_10593);
xnor U11854 (N_11854,N_10785,N_10619);
nor U11855 (N_11855,N_10697,N_10601);
and U11856 (N_11856,N_10862,N_11105);
or U11857 (N_11857,N_10655,N_10610);
nand U11858 (N_11858,N_10654,N_10488);
nor U11859 (N_11859,N_11149,N_11163);
nor U11860 (N_11860,N_10812,N_11052);
nor U11861 (N_11861,N_10511,N_10740);
nor U11862 (N_11862,N_10644,N_10890);
and U11863 (N_11863,N_10492,N_10737);
nand U11864 (N_11864,N_10608,N_10917);
and U11865 (N_11865,N_10913,N_10592);
or U11866 (N_11866,N_11198,N_10557);
or U11867 (N_11867,N_10969,N_11043);
or U11868 (N_11868,N_10827,N_10580);
and U11869 (N_11869,N_10977,N_10494);
or U11870 (N_11870,N_10968,N_10808);
nand U11871 (N_11871,N_10435,N_11175);
or U11872 (N_11872,N_10510,N_10944);
or U11873 (N_11873,N_10416,N_10572);
and U11874 (N_11874,N_10508,N_10900);
and U11875 (N_11875,N_10872,N_10515);
xnor U11876 (N_11876,N_11192,N_10964);
and U11877 (N_11877,N_10482,N_11145);
and U11878 (N_11878,N_10939,N_10969);
and U11879 (N_11879,N_10430,N_11016);
nor U11880 (N_11880,N_11156,N_11185);
xor U11881 (N_11881,N_10852,N_10610);
nor U11882 (N_11882,N_10818,N_10549);
nor U11883 (N_11883,N_10556,N_11095);
and U11884 (N_11884,N_10415,N_10709);
nor U11885 (N_11885,N_11126,N_10689);
nor U11886 (N_11886,N_10718,N_10667);
nand U11887 (N_11887,N_10956,N_10774);
xnor U11888 (N_11888,N_10642,N_10968);
nor U11889 (N_11889,N_11098,N_11143);
or U11890 (N_11890,N_10587,N_11130);
or U11891 (N_11891,N_11109,N_10560);
nor U11892 (N_11892,N_10975,N_10461);
nand U11893 (N_11893,N_10508,N_11095);
and U11894 (N_11894,N_10490,N_10462);
and U11895 (N_11895,N_11115,N_10429);
nor U11896 (N_11896,N_11084,N_10617);
and U11897 (N_11897,N_10448,N_10818);
or U11898 (N_11898,N_10827,N_10421);
or U11899 (N_11899,N_11102,N_11172);
and U11900 (N_11900,N_10501,N_10557);
nor U11901 (N_11901,N_10941,N_10659);
nand U11902 (N_11902,N_10847,N_10682);
xor U11903 (N_11903,N_10889,N_10472);
or U11904 (N_11904,N_10475,N_10615);
nand U11905 (N_11905,N_10594,N_10616);
xor U11906 (N_11906,N_10915,N_10799);
or U11907 (N_11907,N_10619,N_10757);
and U11908 (N_11908,N_10674,N_10699);
xnor U11909 (N_11909,N_11184,N_10894);
xor U11910 (N_11910,N_10411,N_10444);
nor U11911 (N_11911,N_11113,N_10712);
xnor U11912 (N_11912,N_10584,N_10700);
and U11913 (N_11913,N_10529,N_11062);
xor U11914 (N_11914,N_10980,N_10429);
and U11915 (N_11915,N_10879,N_10629);
or U11916 (N_11916,N_10816,N_11062);
and U11917 (N_11917,N_10554,N_10808);
nor U11918 (N_11918,N_10502,N_10606);
nor U11919 (N_11919,N_11093,N_11128);
nor U11920 (N_11920,N_11100,N_11019);
nand U11921 (N_11921,N_10571,N_10680);
or U11922 (N_11922,N_10401,N_10667);
nand U11923 (N_11923,N_10810,N_10434);
nand U11924 (N_11924,N_10824,N_10638);
and U11925 (N_11925,N_10633,N_10782);
and U11926 (N_11926,N_11124,N_11185);
nor U11927 (N_11927,N_11120,N_10422);
or U11928 (N_11928,N_10677,N_11160);
and U11929 (N_11929,N_10625,N_10490);
nor U11930 (N_11930,N_10421,N_11043);
nand U11931 (N_11931,N_10749,N_10496);
or U11932 (N_11932,N_11071,N_11180);
xnor U11933 (N_11933,N_10824,N_10971);
and U11934 (N_11934,N_10404,N_10900);
and U11935 (N_11935,N_10565,N_11026);
and U11936 (N_11936,N_11172,N_10829);
nor U11937 (N_11937,N_11007,N_11005);
or U11938 (N_11938,N_10604,N_11048);
and U11939 (N_11939,N_10403,N_10738);
xor U11940 (N_11940,N_10738,N_10714);
and U11941 (N_11941,N_10875,N_10835);
nand U11942 (N_11942,N_11165,N_10954);
nor U11943 (N_11943,N_10866,N_10790);
nor U11944 (N_11944,N_10943,N_10942);
and U11945 (N_11945,N_11122,N_10785);
or U11946 (N_11946,N_10703,N_11167);
nand U11947 (N_11947,N_10456,N_10676);
and U11948 (N_11948,N_11022,N_10792);
xnor U11949 (N_11949,N_11101,N_11175);
nor U11950 (N_11950,N_11172,N_10935);
nand U11951 (N_11951,N_10783,N_10732);
nand U11952 (N_11952,N_11127,N_10595);
and U11953 (N_11953,N_10999,N_10651);
and U11954 (N_11954,N_10642,N_11130);
nand U11955 (N_11955,N_10564,N_10741);
and U11956 (N_11956,N_10670,N_10911);
xnor U11957 (N_11957,N_10797,N_10773);
xnor U11958 (N_11958,N_10516,N_11093);
or U11959 (N_11959,N_10433,N_10577);
nor U11960 (N_11960,N_10749,N_10808);
and U11961 (N_11961,N_11153,N_10481);
and U11962 (N_11962,N_10856,N_10592);
and U11963 (N_11963,N_11182,N_10497);
nand U11964 (N_11964,N_10802,N_10421);
nor U11965 (N_11965,N_11079,N_10463);
nor U11966 (N_11966,N_10542,N_11105);
nor U11967 (N_11967,N_11044,N_10781);
xor U11968 (N_11968,N_10963,N_10685);
nor U11969 (N_11969,N_10662,N_10530);
and U11970 (N_11970,N_11014,N_10781);
nand U11971 (N_11971,N_10428,N_10469);
nor U11972 (N_11972,N_10695,N_10710);
xnor U11973 (N_11973,N_10939,N_10469);
nand U11974 (N_11974,N_10667,N_11186);
or U11975 (N_11975,N_10688,N_11091);
nand U11976 (N_11976,N_10790,N_11096);
or U11977 (N_11977,N_10867,N_10498);
or U11978 (N_11978,N_10816,N_11094);
nand U11979 (N_11979,N_11037,N_10702);
and U11980 (N_11980,N_10863,N_10911);
and U11981 (N_11981,N_10583,N_10405);
xor U11982 (N_11982,N_11046,N_10622);
and U11983 (N_11983,N_10514,N_11131);
or U11984 (N_11984,N_10872,N_10774);
nor U11985 (N_11985,N_10518,N_11098);
xnor U11986 (N_11986,N_10583,N_10654);
nor U11987 (N_11987,N_10634,N_10716);
or U11988 (N_11988,N_11089,N_10657);
and U11989 (N_11989,N_10845,N_11018);
or U11990 (N_11990,N_10506,N_10788);
xor U11991 (N_11991,N_10664,N_10668);
xor U11992 (N_11992,N_10506,N_11071);
nor U11993 (N_11993,N_10417,N_10497);
xnor U11994 (N_11994,N_10538,N_10555);
or U11995 (N_11995,N_10544,N_11007);
xnor U11996 (N_11996,N_10680,N_11002);
nor U11997 (N_11997,N_10522,N_10943);
nor U11998 (N_11998,N_10661,N_10748);
nor U11999 (N_11999,N_10945,N_10513);
nor U12000 (N_12000,N_11575,N_11925);
or U12001 (N_12001,N_11871,N_11222);
nand U12002 (N_12002,N_11943,N_11322);
and U12003 (N_12003,N_11376,N_11874);
nand U12004 (N_12004,N_11541,N_11588);
xor U12005 (N_12005,N_11423,N_11641);
and U12006 (N_12006,N_11658,N_11794);
nand U12007 (N_12007,N_11891,N_11256);
nand U12008 (N_12008,N_11321,N_11500);
and U12009 (N_12009,N_11275,N_11628);
xor U12010 (N_12010,N_11517,N_11862);
nor U12011 (N_12011,N_11563,N_11251);
and U12012 (N_12012,N_11604,N_11753);
or U12013 (N_12013,N_11977,N_11512);
and U12014 (N_12014,N_11411,N_11360);
and U12015 (N_12015,N_11260,N_11238);
nor U12016 (N_12016,N_11418,N_11413);
xor U12017 (N_12017,N_11684,N_11945);
nor U12018 (N_12018,N_11282,N_11240);
nand U12019 (N_12019,N_11813,N_11744);
nand U12020 (N_12020,N_11546,N_11781);
nand U12021 (N_12021,N_11552,N_11537);
or U12022 (N_12022,N_11897,N_11242);
or U12023 (N_12023,N_11284,N_11732);
nand U12024 (N_12024,N_11345,N_11485);
and U12025 (N_12025,N_11911,N_11585);
or U12026 (N_12026,N_11634,N_11728);
xnor U12027 (N_12027,N_11498,N_11851);
xor U12028 (N_12028,N_11442,N_11958);
xnor U12029 (N_12029,N_11907,N_11329);
or U12030 (N_12030,N_11361,N_11347);
or U12031 (N_12031,N_11384,N_11599);
nand U12032 (N_12032,N_11814,N_11557);
xnor U12033 (N_12033,N_11355,N_11730);
or U12034 (N_12034,N_11327,N_11392);
or U12035 (N_12035,N_11457,N_11333);
nand U12036 (N_12036,N_11829,N_11265);
and U12037 (N_12037,N_11961,N_11858);
xnor U12038 (N_12038,N_11424,N_11673);
or U12039 (N_12039,N_11473,N_11499);
nor U12040 (N_12040,N_11957,N_11481);
nor U12041 (N_12041,N_11932,N_11854);
nand U12042 (N_12042,N_11562,N_11551);
and U12043 (N_12043,N_11336,N_11865);
nor U12044 (N_12044,N_11723,N_11901);
nor U12045 (N_12045,N_11886,N_11852);
nor U12046 (N_12046,N_11351,N_11773);
xor U12047 (N_12047,N_11403,N_11530);
nand U12048 (N_12048,N_11808,N_11236);
and U12049 (N_12049,N_11683,N_11954);
or U12050 (N_12050,N_11691,N_11234);
nand U12051 (N_12051,N_11332,N_11227);
nor U12052 (N_12052,N_11246,N_11210);
nor U12053 (N_12053,N_11678,N_11428);
nor U12054 (N_12054,N_11608,N_11710);
nor U12055 (N_12055,N_11453,N_11690);
xnor U12056 (N_12056,N_11339,N_11845);
and U12057 (N_12057,N_11340,N_11848);
nor U12058 (N_12058,N_11324,N_11381);
nor U12059 (N_12059,N_11908,N_11778);
nor U12060 (N_12060,N_11786,N_11878);
nor U12061 (N_12061,N_11522,N_11746);
or U12062 (N_12062,N_11822,N_11731);
nor U12063 (N_12063,N_11930,N_11790);
and U12064 (N_12064,N_11859,N_11715);
and U12065 (N_12065,N_11801,N_11688);
nor U12066 (N_12066,N_11479,N_11497);
nor U12067 (N_12067,N_11545,N_11695);
xor U12068 (N_12068,N_11326,N_11910);
or U12069 (N_12069,N_11916,N_11669);
nand U12070 (N_12070,N_11573,N_11652);
and U12071 (N_12071,N_11748,N_11456);
and U12072 (N_12072,N_11547,N_11212);
and U12073 (N_12073,N_11255,N_11229);
nor U12074 (N_12074,N_11763,N_11582);
nand U12075 (N_12075,N_11576,N_11887);
or U12076 (N_12076,N_11389,N_11452);
or U12077 (N_12077,N_11965,N_11760);
xor U12078 (N_12078,N_11200,N_11316);
nand U12079 (N_12079,N_11263,N_11992);
xnor U12080 (N_12080,N_11410,N_11572);
nand U12081 (N_12081,N_11523,N_11761);
xor U12082 (N_12082,N_11692,N_11806);
or U12083 (N_12083,N_11350,N_11579);
xor U12084 (N_12084,N_11767,N_11698);
xnor U12085 (N_12085,N_11649,N_11672);
nand U12086 (N_12086,N_11906,N_11627);
xor U12087 (N_12087,N_11631,N_11221);
or U12088 (N_12088,N_11402,N_11883);
xnor U12089 (N_12089,N_11226,N_11618);
xor U12090 (N_12090,N_11740,N_11733);
xnor U12091 (N_12091,N_11616,N_11869);
or U12092 (N_12092,N_11510,N_11567);
and U12093 (N_12093,N_11568,N_11338);
or U12094 (N_12094,N_11521,N_11527);
xor U12095 (N_12095,N_11759,N_11849);
or U12096 (N_12096,N_11755,N_11460);
and U12097 (N_12097,N_11602,N_11972);
nand U12098 (N_12098,N_11622,N_11232);
nor U12099 (N_12099,N_11475,N_11917);
and U12100 (N_12100,N_11580,N_11953);
nor U12101 (N_12101,N_11950,N_11589);
or U12102 (N_12102,N_11668,N_11860);
xnor U12103 (N_12103,N_11720,N_11973);
nand U12104 (N_12104,N_11613,N_11268);
xnor U12105 (N_12105,N_11518,N_11877);
nand U12106 (N_12106,N_11896,N_11762);
or U12107 (N_12107,N_11736,N_11843);
nor U12108 (N_12108,N_11554,N_11290);
nand U12109 (N_12109,N_11375,N_11704);
and U12110 (N_12110,N_11959,N_11379);
nand U12111 (N_12111,N_11409,N_11368);
nor U12112 (N_12112,N_11323,N_11768);
and U12113 (N_12113,N_11819,N_11994);
and U12114 (N_12114,N_11454,N_11466);
nor U12115 (N_12115,N_11624,N_11991);
or U12116 (N_12116,N_11880,N_11661);
nor U12117 (N_12117,N_11921,N_11207);
and U12118 (N_12118,N_11348,N_11919);
nand U12119 (N_12119,N_11528,N_11488);
xor U12120 (N_12120,N_11821,N_11370);
xnor U12121 (N_12121,N_11941,N_11560);
nand U12122 (N_12122,N_11396,N_11279);
xor U12123 (N_12123,N_11591,N_11940);
nor U12124 (N_12124,N_11675,N_11224);
or U12125 (N_12125,N_11446,N_11873);
nor U12126 (N_12126,N_11920,N_11553);
and U12127 (N_12127,N_11706,N_11543);
nand U12128 (N_12128,N_11436,N_11470);
nand U12129 (N_12129,N_11237,N_11833);
or U12130 (N_12130,N_11904,N_11367);
or U12131 (N_12131,N_11798,N_11532);
xor U12132 (N_12132,N_11511,N_11539);
nand U12133 (N_12133,N_11495,N_11654);
or U12134 (N_12134,N_11603,N_11832);
or U12135 (N_12135,N_11931,N_11807);
xor U12136 (N_12136,N_11600,N_11742);
nor U12137 (N_12137,N_11827,N_11407);
nand U12138 (N_12138,N_11391,N_11266);
or U12139 (N_12139,N_11489,N_11853);
and U12140 (N_12140,N_11635,N_11369);
nand U12141 (N_12141,N_11985,N_11846);
and U12142 (N_12142,N_11870,N_11964);
and U12143 (N_12143,N_11830,N_11923);
nor U12144 (N_12144,N_11534,N_11325);
nor U12145 (N_12145,N_11824,N_11749);
and U12146 (N_12146,N_11671,N_11271);
nand U12147 (N_12147,N_11484,N_11211);
nand U12148 (N_12148,N_11726,N_11660);
and U12149 (N_12149,N_11487,N_11254);
nor U12150 (N_12150,N_11431,N_11995);
and U12151 (N_12151,N_11443,N_11533);
xnor U12152 (N_12152,N_11346,N_11955);
and U12153 (N_12153,N_11948,N_11772);
xnor U12154 (N_12154,N_11802,N_11913);
and U12155 (N_12155,N_11927,N_11300);
xnor U12156 (N_12156,N_11997,N_11598);
and U12157 (N_12157,N_11937,N_11774);
nand U12158 (N_12158,N_11963,N_11835);
nor U12159 (N_12159,N_11610,N_11272);
xor U12160 (N_12160,N_11525,N_11253);
nand U12161 (N_12161,N_11235,N_11636);
and U12162 (N_12162,N_11217,N_11981);
nand U12163 (N_12163,N_11366,N_11952);
or U12164 (N_12164,N_11751,N_11612);
xnor U12165 (N_12165,N_11344,N_11799);
nand U12166 (N_12166,N_11826,N_11583);
or U12167 (N_12167,N_11885,N_11960);
and U12168 (N_12168,N_11993,N_11294);
nor U12169 (N_12169,N_11241,N_11875);
or U12170 (N_12170,N_11922,N_11390);
and U12171 (N_12171,N_11445,N_11216);
nand U12172 (N_12172,N_11299,N_11313);
nand U12173 (N_12173,N_11974,N_11422);
nor U12174 (N_12174,N_11914,N_11483);
nand U12175 (N_12175,N_11501,N_11421);
nand U12176 (N_12176,N_11334,N_11397);
xnor U12177 (N_12177,N_11291,N_11597);
and U12178 (N_12178,N_11727,N_11219);
or U12179 (N_12179,N_11924,N_11987);
or U12180 (N_12180,N_11839,N_11476);
nor U12181 (N_12181,N_11292,N_11743);
xnor U12182 (N_12182,N_11879,N_11319);
nor U12183 (N_12183,N_11680,N_11811);
nand U12184 (N_12184,N_11784,N_11298);
xnor U12185 (N_12185,N_11218,N_11270);
or U12186 (N_12186,N_11225,N_11855);
and U12187 (N_12187,N_11592,N_11293);
xor U12188 (N_12188,N_11406,N_11872);
nor U12189 (N_12189,N_11892,N_11739);
or U12190 (N_12190,N_11505,N_11335);
nand U12191 (N_12191,N_11363,N_11408);
nor U12192 (N_12192,N_11273,N_11594);
nor U12193 (N_12193,N_11777,N_11388);
or U12194 (N_12194,N_11864,N_11629);
xor U12195 (N_12195,N_11644,N_11330);
or U12196 (N_12196,N_11971,N_11352);
and U12197 (N_12197,N_11435,N_11465);
nor U12198 (N_12198,N_11988,N_11549);
xor U12199 (N_12199,N_11249,N_11311);
nand U12200 (N_12200,N_11689,N_11535);
nor U12201 (N_12201,N_11354,N_11520);
nor U12202 (N_12202,N_11626,N_11439);
nor U12203 (N_12203,N_11861,N_11477);
and U12204 (N_12204,N_11474,N_11513);
nand U12205 (N_12205,N_11666,N_11949);
or U12206 (N_12206,N_11449,N_11213);
and U12207 (N_12207,N_11968,N_11427);
and U12208 (N_12208,N_11378,N_11606);
and U12209 (N_12209,N_11239,N_11425);
or U12210 (N_12210,N_11788,N_11502);
xnor U12211 (N_12211,N_11288,N_11942);
or U12212 (N_12212,N_11747,N_11737);
or U12213 (N_12213,N_11850,N_11555);
nand U12214 (N_12214,N_11933,N_11304);
nand U12215 (N_12215,N_11642,N_11946);
xnor U12216 (N_12216,N_11693,N_11586);
nor U12217 (N_12217,N_11486,N_11277);
or U12218 (N_12218,N_11362,N_11373);
xor U12219 (N_12219,N_11699,N_11882);
nand U12220 (N_12220,N_11662,N_11729);
xnor U12221 (N_12221,N_11419,N_11638);
and U12222 (N_12222,N_11711,N_11531);
xnor U12223 (N_12223,N_11385,N_11414);
or U12224 (N_12224,N_11214,N_11577);
and U12225 (N_12225,N_11667,N_11783);
or U12226 (N_12226,N_11463,N_11984);
xnor U12227 (N_12227,N_11838,N_11769);
and U12228 (N_12228,N_11983,N_11401);
nor U12229 (N_12229,N_11703,N_11353);
xnor U12230 (N_12230,N_11472,N_11990);
xnor U12231 (N_12231,N_11503,N_11825);
or U12232 (N_12232,N_11317,N_11526);
nand U12233 (N_12233,N_11979,N_11630);
or U12234 (N_12234,N_11494,N_11364);
and U12235 (N_12235,N_11301,N_11653);
nor U12236 (N_12236,N_11434,N_11970);
nor U12237 (N_12237,N_11278,N_11394);
nand U12238 (N_12238,N_11305,N_11556);
and U12239 (N_12239,N_11840,N_11371);
xnor U12240 (N_12240,N_11309,N_11621);
xnor U12241 (N_12241,N_11269,N_11912);
nand U12242 (N_12242,N_11247,N_11696);
and U12243 (N_12243,N_11674,N_11561);
xnor U12244 (N_12244,N_11285,N_11252);
nor U12245 (N_12245,N_11876,N_11818);
xor U12246 (N_12246,N_11303,N_11685);
and U12247 (N_12247,N_11209,N_11752);
xnor U12248 (N_12248,N_11890,N_11437);
nand U12249 (N_12249,N_11857,N_11766);
or U12250 (N_12250,N_11365,N_11220);
or U12251 (N_12251,N_11318,N_11776);
xnor U12252 (N_12252,N_11721,N_11697);
or U12253 (N_12253,N_11947,N_11228);
and U12254 (N_12254,N_11800,N_11357);
nand U12255 (N_12255,N_11262,N_11999);
or U12256 (N_12256,N_11380,N_11450);
and U12257 (N_12257,N_11462,N_11529);
or U12258 (N_12258,N_11754,N_11996);
and U12259 (N_12259,N_11312,N_11468);
or U12260 (N_12260,N_11287,N_11797);
xor U12261 (N_12261,N_11758,N_11645);
nand U12262 (N_12262,N_11491,N_11633);
and U12263 (N_12263,N_11934,N_11565);
nand U12264 (N_12264,N_11519,N_11359);
nor U12265 (N_12265,N_11926,N_11719);
and U12266 (N_12266,N_11815,N_11718);
and U12267 (N_12267,N_11918,N_11458);
nor U12268 (N_12268,N_11596,N_11429);
nand U12269 (N_12269,N_11650,N_11928);
or U12270 (N_12270,N_11208,N_11416);
and U12271 (N_12271,N_11461,N_11998);
and U12272 (N_12272,N_11202,N_11889);
nor U12273 (N_12273,N_11420,N_11374);
nor U12274 (N_12274,N_11888,N_11791);
nor U12275 (N_12275,N_11898,N_11250);
and U12276 (N_12276,N_11459,N_11686);
and U12277 (N_12277,N_11708,N_11276);
or U12278 (N_12278,N_11976,N_11595);
or U12279 (N_12279,N_11866,N_11516);
xor U12280 (N_12280,N_11405,N_11283);
nand U12281 (N_12281,N_11863,N_11734);
and U12282 (N_12282,N_11601,N_11515);
nor U12283 (N_12283,N_11245,N_11386);
nor U12284 (N_12284,N_11570,N_11643);
or U12285 (N_12285,N_11625,N_11393);
nor U12286 (N_12286,N_11793,N_11493);
nor U12287 (N_12287,N_11823,N_11639);
or U12288 (N_12288,N_11544,N_11709);
xor U12289 (N_12289,N_11975,N_11756);
nor U12290 (N_12290,N_11356,N_11647);
or U12291 (N_12291,N_11935,N_11509);
xor U12292 (N_12292,N_11905,N_11700);
nand U12293 (N_12293,N_11310,N_11441);
nand U12294 (N_12294,N_11584,N_11302);
xor U12295 (N_12295,N_11349,N_11296);
xnor U12296 (N_12296,N_11713,N_11426);
and U12297 (N_12297,N_11430,N_11295);
nand U12298 (N_12298,N_11478,N_11682);
nand U12299 (N_12299,N_11681,N_11615);
xor U12300 (N_12300,N_11902,N_11632);
nand U12301 (N_12301,N_11780,N_11536);
nand U12302 (N_12302,N_11508,N_11956);
xnor U12303 (N_12303,N_11764,N_11550);
nand U12304 (N_12304,N_11231,N_11480);
or U12305 (N_12305,N_11938,N_11842);
and U12306 (N_12306,N_11448,N_11915);
or U12307 (N_12307,N_11646,N_11257);
nor U12308 (N_12308,N_11724,N_11506);
nor U12309 (N_12309,N_11440,N_11805);
or U12310 (N_12310,N_11881,N_11617);
nand U12311 (N_12311,N_11548,N_11640);
nor U12312 (N_12312,N_11722,N_11571);
nor U12313 (N_12313,N_11651,N_11782);
nand U12314 (N_12314,N_11372,N_11274);
and U12315 (N_12315,N_11201,N_11656);
xor U12316 (N_12316,N_11337,N_11929);
or U12317 (N_12317,N_11540,N_11796);
nor U12318 (N_12318,N_11387,N_11750);
or U12319 (N_12319,N_11578,N_11687);
nand U12320 (N_12320,N_11308,N_11659);
xnor U12321 (N_12321,N_11267,N_11204);
nor U12322 (N_12322,N_11614,N_11205);
nor U12323 (N_12323,N_11433,N_11469);
nand U12324 (N_12324,N_11705,N_11900);
nand U12325 (N_12325,N_11820,N_11451);
nor U12326 (N_12326,N_11670,N_11320);
nand U12327 (N_12327,N_11828,N_11894);
and U12328 (N_12328,N_11607,N_11939);
nand U12329 (N_12329,N_11447,N_11261);
nand U12330 (N_12330,N_11609,N_11590);
nand U12331 (N_12331,N_11694,N_11215);
nand U12332 (N_12332,N_11741,N_11831);
and U12333 (N_12333,N_11779,N_11738);
nand U12334 (N_12334,N_11812,N_11909);
or U12335 (N_12335,N_11417,N_11792);
xor U12336 (N_12336,N_11559,N_11398);
nand U12337 (N_12337,N_11714,N_11593);
and U12338 (N_12338,N_11514,N_11258);
nand U12339 (N_12339,N_11903,N_11248);
nor U12340 (N_12340,N_11712,N_11837);
or U12341 (N_12341,N_11306,N_11785);
nor U12342 (N_12342,N_11230,N_11765);
xnor U12343 (N_12343,N_11243,N_11982);
xor U12344 (N_12344,N_11455,N_11969);
or U12345 (N_12345,N_11847,N_11412);
nand U12346 (N_12346,N_11771,N_11504);
xnor U12347 (N_12347,N_11564,N_11444);
or U12348 (N_12348,N_11395,N_11404);
and U12349 (N_12349,N_11735,N_11507);
nor U12350 (N_12350,N_11936,N_11657);
nor U12351 (N_12351,N_11438,N_11676);
or U12352 (N_12352,N_11620,N_11524);
nor U12353 (N_12353,N_11895,N_11868);
and U12354 (N_12354,N_11377,N_11400);
nand U12355 (N_12355,N_11605,N_11566);
nand U12356 (N_12356,N_11611,N_11745);
nand U12357 (N_12357,N_11358,N_11331);
or U12358 (N_12358,N_11623,N_11538);
nand U12359 (N_12359,N_11314,N_11966);
xor U12360 (N_12360,N_11775,N_11619);
nor U12361 (N_12361,N_11482,N_11884);
or U12362 (N_12362,N_11962,N_11637);
nor U12363 (N_12363,N_11259,N_11834);
nor U12364 (N_12364,N_11716,N_11856);
nor U12365 (N_12365,N_11496,N_11289);
nand U12366 (N_12366,N_11967,N_11893);
or U12367 (N_12367,N_11809,N_11280);
nand U12368 (N_12368,N_11297,N_11817);
or U12369 (N_12369,N_11844,N_11542);
and U12370 (N_12370,N_11899,N_11803);
and U12371 (N_12371,N_11665,N_11789);
and U12372 (N_12372,N_11342,N_11343);
or U12373 (N_12373,N_11281,N_11663);
nor U12374 (N_12374,N_11307,N_11980);
or U12375 (N_12375,N_11770,N_11867);
and U12376 (N_12376,N_11492,N_11223);
xnor U12377 (N_12377,N_11702,N_11558);
and U12378 (N_12378,N_11810,N_11490);
xor U12379 (N_12379,N_11233,N_11382);
xnor U12380 (N_12380,N_11836,N_11315);
or U12381 (N_12381,N_11383,N_11757);
or U12382 (N_12382,N_11203,N_11951);
nor U12383 (N_12383,N_11664,N_11816);
and U12384 (N_12384,N_11679,N_11328);
nor U12385 (N_12385,N_11989,N_11655);
and U12386 (N_12386,N_11415,N_11587);
xor U12387 (N_12387,N_11581,N_11286);
or U12388 (N_12388,N_11707,N_11341);
nand U12389 (N_12389,N_11795,N_11944);
and U12390 (N_12390,N_11978,N_11574);
and U12391 (N_12391,N_11569,N_11264);
and U12392 (N_12392,N_11244,N_11717);
and U12393 (N_12393,N_11432,N_11841);
or U12394 (N_12394,N_11986,N_11464);
xor U12395 (N_12395,N_11787,N_11701);
xnor U12396 (N_12396,N_11467,N_11677);
xnor U12397 (N_12397,N_11471,N_11648);
nor U12398 (N_12398,N_11206,N_11399);
or U12399 (N_12399,N_11804,N_11725);
xnor U12400 (N_12400,N_11267,N_11576);
or U12401 (N_12401,N_11208,N_11888);
or U12402 (N_12402,N_11909,N_11375);
nand U12403 (N_12403,N_11464,N_11468);
nor U12404 (N_12404,N_11670,N_11647);
and U12405 (N_12405,N_11531,N_11395);
nand U12406 (N_12406,N_11312,N_11842);
xnor U12407 (N_12407,N_11901,N_11323);
nor U12408 (N_12408,N_11361,N_11517);
or U12409 (N_12409,N_11366,N_11387);
or U12410 (N_12410,N_11845,N_11574);
nand U12411 (N_12411,N_11453,N_11488);
or U12412 (N_12412,N_11995,N_11363);
nor U12413 (N_12413,N_11615,N_11787);
nor U12414 (N_12414,N_11986,N_11379);
and U12415 (N_12415,N_11778,N_11712);
and U12416 (N_12416,N_11323,N_11365);
and U12417 (N_12417,N_11931,N_11906);
nor U12418 (N_12418,N_11569,N_11878);
or U12419 (N_12419,N_11296,N_11373);
nor U12420 (N_12420,N_11535,N_11605);
and U12421 (N_12421,N_11711,N_11360);
xnor U12422 (N_12422,N_11745,N_11468);
nor U12423 (N_12423,N_11552,N_11767);
nor U12424 (N_12424,N_11567,N_11625);
and U12425 (N_12425,N_11245,N_11470);
or U12426 (N_12426,N_11313,N_11922);
or U12427 (N_12427,N_11369,N_11548);
nor U12428 (N_12428,N_11497,N_11867);
or U12429 (N_12429,N_11555,N_11711);
xor U12430 (N_12430,N_11711,N_11318);
and U12431 (N_12431,N_11693,N_11990);
nand U12432 (N_12432,N_11508,N_11255);
nor U12433 (N_12433,N_11938,N_11280);
and U12434 (N_12434,N_11790,N_11774);
xnor U12435 (N_12435,N_11319,N_11762);
and U12436 (N_12436,N_11936,N_11489);
xor U12437 (N_12437,N_11791,N_11251);
and U12438 (N_12438,N_11938,N_11779);
nand U12439 (N_12439,N_11488,N_11351);
xnor U12440 (N_12440,N_11804,N_11337);
xnor U12441 (N_12441,N_11780,N_11301);
xor U12442 (N_12442,N_11492,N_11865);
or U12443 (N_12443,N_11429,N_11468);
and U12444 (N_12444,N_11721,N_11380);
or U12445 (N_12445,N_11332,N_11859);
xnor U12446 (N_12446,N_11217,N_11245);
nor U12447 (N_12447,N_11230,N_11323);
and U12448 (N_12448,N_11670,N_11449);
nand U12449 (N_12449,N_11812,N_11597);
xnor U12450 (N_12450,N_11703,N_11679);
nand U12451 (N_12451,N_11797,N_11648);
nor U12452 (N_12452,N_11425,N_11579);
nor U12453 (N_12453,N_11495,N_11581);
or U12454 (N_12454,N_11328,N_11785);
or U12455 (N_12455,N_11386,N_11609);
or U12456 (N_12456,N_11904,N_11499);
or U12457 (N_12457,N_11795,N_11971);
xnor U12458 (N_12458,N_11479,N_11586);
nand U12459 (N_12459,N_11354,N_11799);
xnor U12460 (N_12460,N_11788,N_11515);
nor U12461 (N_12461,N_11948,N_11411);
nand U12462 (N_12462,N_11619,N_11714);
xnor U12463 (N_12463,N_11371,N_11462);
xnor U12464 (N_12464,N_11925,N_11453);
nand U12465 (N_12465,N_11731,N_11871);
and U12466 (N_12466,N_11829,N_11686);
xnor U12467 (N_12467,N_11490,N_11967);
or U12468 (N_12468,N_11905,N_11291);
xnor U12469 (N_12469,N_11314,N_11635);
xor U12470 (N_12470,N_11974,N_11939);
nor U12471 (N_12471,N_11373,N_11234);
and U12472 (N_12472,N_11215,N_11227);
xnor U12473 (N_12473,N_11716,N_11620);
or U12474 (N_12474,N_11858,N_11352);
xor U12475 (N_12475,N_11903,N_11961);
nor U12476 (N_12476,N_11741,N_11657);
nand U12477 (N_12477,N_11253,N_11735);
xnor U12478 (N_12478,N_11230,N_11341);
xor U12479 (N_12479,N_11206,N_11268);
and U12480 (N_12480,N_11461,N_11415);
nand U12481 (N_12481,N_11913,N_11536);
nor U12482 (N_12482,N_11426,N_11756);
nor U12483 (N_12483,N_11780,N_11788);
nand U12484 (N_12484,N_11599,N_11410);
xor U12485 (N_12485,N_11717,N_11692);
nor U12486 (N_12486,N_11444,N_11368);
and U12487 (N_12487,N_11802,N_11381);
xnor U12488 (N_12488,N_11443,N_11491);
nor U12489 (N_12489,N_11917,N_11581);
and U12490 (N_12490,N_11238,N_11728);
xor U12491 (N_12491,N_11899,N_11972);
or U12492 (N_12492,N_11575,N_11596);
nor U12493 (N_12493,N_11521,N_11382);
or U12494 (N_12494,N_11320,N_11501);
nor U12495 (N_12495,N_11710,N_11737);
nand U12496 (N_12496,N_11645,N_11801);
and U12497 (N_12497,N_11587,N_11405);
nand U12498 (N_12498,N_11621,N_11438);
and U12499 (N_12499,N_11916,N_11638);
or U12500 (N_12500,N_11399,N_11410);
or U12501 (N_12501,N_11546,N_11516);
nand U12502 (N_12502,N_11869,N_11658);
and U12503 (N_12503,N_11934,N_11548);
nand U12504 (N_12504,N_11575,N_11230);
or U12505 (N_12505,N_11981,N_11572);
or U12506 (N_12506,N_11725,N_11443);
or U12507 (N_12507,N_11586,N_11461);
and U12508 (N_12508,N_11450,N_11429);
nand U12509 (N_12509,N_11405,N_11499);
nor U12510 (N_12510,N_11252,N_11693);
nor U12511 (N_12511,N_11838,N_11657);
or U12512 (N_12512,N_11714,N_11748);
xor U12513 (N_12513,N_11939,N_11469);
nand U12514 (N_12514,N_11287,N_11897);
nor U12515 (N_12515,N_11265,N_11600);
and U12516 (N_12516,N_11699,N_11282);
or U12517 (N_12517,N_11947,N_11603);
nor U12518 (N_12518,N_11684,N_11539);
nor U12519 (N_12519,N_11715,N_11852);
or U12520 (N_12520,N_11211,N_11382);
nor U12521 (N_12521,N_11747,N_11293);
nor U12522 (N_12522,N_11576,N_11622);
xnor U12523 (N_12523,N_11626,N_11924);
or U12524 (N_12524,N_11553,N_11386);
xnor U12525 (N_12525,N_11874,N_11206);
nor U12526 (N_12526,N_11753,N_11944);
and U12527 (N_12527,N_11521,N_11315);
xor U12528 (N_12528,N_11365,N_11281);
xnor U12529 (N_12529,N_11295,N_11901);
nand U12530 (N_12530,N_11846,N_11645);
and U12531 (N_12531,N_11388,N_11256);
nor U12532 (N_12532,N_11253,N_11715);
nor U12533 (N_12533,N_11956,N_11278);
xor U12534 (N_12534,N_11792,N_11874);
or U12535 (N_12535,N_11543,N_11878);
xnor U12536 (N_12536,N_11411,N_11545);
nand U12537 (N_12537,N_11560,N_11398);
or U12538 (N_12538,N_11252,N_11679);
xor U12539 (N_12539,N_11671,N_11976);
nor U12540 (N_12540,N_11898,N_11469);
and U12541 (N_12541,N_11660,N_11419);
xnor U12542 (N_12542,N_11317,N_11550);
xnor U12543 (N_12543,N_11636,N_11901);
nor U12544 (N_12544,N_11538,N_11795);
xnor U12545 (N_12545,N_11918,N_11849);
nand U12546 (N_12546,N_11840,N_11249);
or U12547 (N_12547,N_11279,N_11438);
and U12548 (N_12548,N_11747,N_11477);
xnor U12549 (N_12549,N_11403,N_11665);
nand U12550 (N_12550,N_11328,N_11885);
nand U12551 (N_12551,N_11690,N_11252);
nor U12552 (N_12552,N_11608,N_11330);
and U12553 (N_12553,N_11653,N_11374);
nand U12554 (N_12554,N_11562,N_11383);
nand U12555 (N_12555,N_11660,N_11839);
and U12556 (N_12556,N_11434,N_11948);
and U12557 (N_12557,N_11760,N_11456);
and U12558 (N_12558,N_11285,N_11659);
nor U12559 (N_12559,N_11453,N_11978);
nor U12560 (N_12560,N_11882,N_11388);
nor U12561 (N_12561,N_11741,N_11344);
or U12562 (N_12562,N_11327,N_11469);
nor U12563 (N_12563,N_11355,N_11993);
and U12564 (N_12564,N_11624,N_11839);
and U12565 (N_12565,N_11653,N_11496);
and U12566 (N_12566,N_11706,N_11675);
nor U12567 (N_12567,N_11665,N_11387);
and U12568 (N_12568,N_11222,N_11402);
and U12569 (N_12569,N_11827,N_11480);
or U12570 (N_12570,N_11865,N_11741);
nand U12571 (N_12571,N_11982,N_11393);
or U12572 (N_12572,N_11900,N_11870);
nor U12573 (N_12573,N_11334,N_11283);
or U12574 (N_12574,N_11838,N_11987);
nand U12575 (N_12575,N_11962,N_11544);
nor U12576 (N_12576,N_11515,N_11340);
or U12577 (N_12577,N_11310,N_11947);
or U12578 (N_12578,N_11708,N_11342);
or U12579 (N_12579,N_11790,N_11725);
nor U12580 (N_12580,N_11334,N_11883);
or U12581 (N_12581,N_11554,N_11816);
nand U12582 (N_12582,N_11208,N_11916);
nand U12583 (N_12583,N_11628,N_11448);
nor U12584 (N_12584,N_11590,N_11982);
nand U12585 (N_12585,N_11915,N_11631);
and U12586 (N_12586,N_11820,N_11316);
nor U12587 (N_12587,N_11390,N_11952);
nor U12588 (N_12588,N_11253,N_11239);
or U12589 (N_12589,N_11698,N_11291);
nor U12590 (N_12590,N_11958,N_11702);
or U12591 (N_12591,N_11605,N_11444);
xor U12592 (N_12592,N_11662,N_11796);
and U12593 (N_12593,N_11300,N_11503);
or U12594 (N_12594,N_11383,N_11874);
or U12595 (N_12595,N_11645,N_11536);
nand U12596 (N_12596,N_11349,N_11375);
nor U12597 (N_12597,N_11748,N_11572);
or U12598 (N_12598,N_11274,N_11499);
nor U12599 (N_12599,N_11655,N_11994);
and U12600 (N_12600,N_11930,N_11917);
and U12601 (N_12601,N_11723,N_11867);
nor U12602 (N_12602,N_11306,N_11711);
xor U12603 (N_12603,N_11201,N_11945);
or U12604 (N_12604,N_11282,N_11569);
and U12605 (N_12605,N_11483,N_11666);
xnor U12606 (N_12606,N_11384,N_11589);
xnor U12607 (N_12607,N_11686,N_11484);
nor U12608 (N_12608,N_11822,N_11770);
nand U12609 (N_12609,N_11644,N_11721);
nor U12610 (N_12610,N_11235,N_11800);
nand U12611 (N_12611,N_11407,N_11432);
and U12612 (N_12612,N_11307,N_11200);
nand U12613 (N_12613,N_11213,N_11991);
nand U12614 (N_12614,N_11548,N_11354);
and U12615 (N_12615,N_11777,N_11405);
or U12616 (N_12616,N_11306,N_11965);
nor U12617 (N_12617,N_11591,N_11525);
nor U12618 (N_12618,N_11724,N_11967);
nand U12619 (N_12619,N_11242,N_11453);
xor U12620 (N_12620,N_11376,N_11263);
xor U12621 (N_12621,N_11729,N_11554);
and U12622 (N_12622,N_11281,N_11425);
nand U12623 (N_12623,N_11353,N_11648);
xnor U12624 (N_12624,N_11253,N_11309);
nand U12625 (N_12625,N_11892,N_11697);
nand U12626 (N_12626,N_11743,N_11794);
or U12627 (N_12627,N_11560,N_11916);
xor U12628 (N_12628,N_11666,N_11535);
xnor U12629 (N_12629,N_11844,N_11357);
and U12630 (N_12630,N_11404,N_11514);
xnor U12631 (N_12631,N_11976,N_11444);
or U12632 (N_12632,N_11214,N_11371);
nand U12633 (N_12633,N_11526,N_11306);
nor U12634 (N_12634,N_11343,N_11877);
xor U12635 (N_12635,N_11569,N_11884);
xnor U12636 (N_12636,N_11794,N_11252);
xor U12637 (N_12637,N_11282,N_11363);
nand U12638 (N_12638,N_11955,N_11800);
xnor U12639 (N_12639,N_11814,N_11309);
nor U12640 (N_12640,N_11752,N_11874);
xnor U12641 (N_12641,N_11548,N_11941);
or U12642 (N_12642,N_11942,N_11248);
xnor U12643 (N_12643,N_11756,N_11965);
and U12644 (N_12644,N_11231,N_11842);
nand U12645 (N_12645,N_11581,N_11767);
xor U12646 (N_12646,N_11505,N_11739);
or U12647 (N_12647,N_11754,N_11451);
xnor U12648 (N_12648,N_11668,N_11993);
and U12649 (N_12649,N_11721,N_11627);
nor U12650 (N_12650,N_11997,N_11355);
or U12651 (N_12651,N_11494,N_11318);
nand U12652 (N_12652,N_11675,N_11969);
xnor U12653 (N_12653,N_11343,N_11674);
xnor U12654 (N_12654,N_11478,N_11486);
nand U12655 (N_12655,N_11458,N_11408);
xnor U12656 (N_12656,N_11435,N_11268);
and U12657 (N_12657,N_11788,N_11857);
and U12658 (N_12658,N_11554,N_11362);
and U12659 (N_12659,N_11226,N_11685);
nor U12660 (N_12660,N_11556,N_11716);
and U12661 (N_12661,N_11733,N_11261);
nand U12662 (N_12662,N_11879,N_11217);
nor U12663 (N_12663,N_11814,N_11217);
nor U12664 (N_12664,N_11853,N_11694);
or U12665 (N_12665,N_11305,N_11554);
xor U12666 (N_12666,N_11448,N_11655);
and U12667 (N_12667,N_11682,N_11234);
xnor U12668 (N_12668,N_11783,N_11466);
nand U12669 (N_12669,N_11369,N_11738);
or U12670 (N_12670,N_11856,N_11303);
xor U12671 (N_12671,N_11591,N_11551);
nor U12672 (N_12672,N_11911,N_11311);
nor U12673 (N_12673,N_11621,N_11524);
xnor U12674 (N_12674,N_11881,N_11328);
and U12675 (N_12675,N_11424,N_11860);
and U12676 (N_12676,N_11457,N_11739);
or U12677 (N_12677,N_11663,N_11651);
xor U12678 (N_12678,N_11420,N_11614);
nand U12679 (N_12679,N_11972,N_11444);
nor U12680 (N_12680,N_11949,N_11204);
nor U12681 (N_12681,N_11820,N_11661);
or U12682 (N_12682,N_11688,N_11299);
nand U12683 (N_12683,N_11908,N_11462);
nor U12684 (N_12684,N_11687,N_11431);
xor U12685 (N_12685,N_11942,N_11810);
and U12686 (N_12686,N_11762,N_11293);
nor U12687 (N_12687,N_11204,N_11604);
and U12688 (N_12688,N_11714,N_11844);
nand U12689 (N_12689,N_11255,N_11845);
nor U12690 (N_12690,N_11228,N_11273);
nor U12691 (N_12691,N_11356,N_11309);
and U12692 (N_12692,N_11988,N_11589);
xor U12693 (N_12693,N_11514,N_11739);
or U12694 (N_12694,N_11375,N_11389);
nor U12695 (N_12695,N_11945,N_11654);
and U12696 (N_12696,N_11660,N_11398);
and U12697 (N_12697,N_11492,N_11939);
and U12698 (N_12698,N_11649,N_11610);
xnor U12699 (N_12699,N_11279,N_11818);
and U12700 (N_12700,N_11259,N_11983);
and U12701 (N_12701,N_11258,N_11480);
and U12702 (N_12702,N_11395,N_11837);
and U12703 (N_12703,N_11202,N_11260);
nor U12704 (N_12704,N_11732,N_11270);
or U12705 (N_12705,N_11573,N_11499);
xor U12706 (N_12706,N_11765,N_11399);
or U12707 (N_12707,N_11906,N_11997);
nand U12708 (N_12708,N_11838,N_11884);
or U12709 (N_12709,N_11448,N_11484);
xnor U12710 (N_12710,N_11305,N_11714);
nand U12711 (N_12711,N_11530,N_11370);
and U12712 (N_12712,N_11295,N_11477);
nand U12713 (N_12713,N_11743,N_11937);
nand U12714 (N_12714,N_11522,N_11959);
and U12715 (N_12715,N_11891,N_11611);
nand U12716 (N_12716,N_11230,N_11864);
and U12717 (N_12717,N_11984,N_11971);
nor U12718 (N_12718,N_11408,N_11561);
or U12719 (N_12719,N_11790,N_11390);
or U12720 (N_12720,N_11941,N_11623);
xnor U12721 (N_12721,N_11991,N_11569);
xnor U12722 (N_12722,N_11277,N_11570);
xnor U12723 (N_12723,N_11249,N_11752);
nor U12724 (N_12724,N_11417,N_11899);
nor U12725 (N_12725,N_11405,N_11458);
and U12726 (N_12726,N_11873,N_11453);
or U12727 (N_12727,N_11238,N_11883);
or U12728 (N_12728,N_11372,N_11777);
and U12729 (N_12729,N_11883,N_11311);
xor U12730 (N_12730,N_11371,N_11616);
and U12731 (N_12731,N_11587,N_11955);
nor U12732 (N_12732,N_11759,N_11239);
and U12733 (N_12733,N_11634,N_11726);
xor U12734 (N_12734,N_11634,N_11626);
xnor U12735 (N_12735,N_11579,N_11916);
xor U12736 (N_12736,N_11993,N_11301);
and U12737 (N_12737,N_11270,N_11831);
nand U12738 (N_12738,N_11895,N_11624);
xor U12739 (N_12739,N_11548,N_11607);
xor U12740 (N_12740,N_11363,N_11603);
nor U12741 (N_12741,N_11275,N_11216);
nand U12742 (N_12742,N_11308,N_11676);
nand U12743 (N_12743,N_11446,N_11831);
or U12744 (N_12744,N_11229,N_11673);
and U12745 (N_12745,N_11972,N_11378);
nand U12746 (N_12746,N_11703,N_11429);
xor U12747 (N_12747,N_11897,N_11636);
and U12748 (N_12748,N_11698,N_11226);
nand U12749 (N_12749,N_11316,N_11558);
and U12750 (N_12750,N_11971,N_11219);
xnor U12751 (N_12751,N_11850,N_11622);
and U12752 (N_12752,N_11386,N_11673);
nor U12753 (N_12753,N_11319,N_11398);
or U12754 (N_12754,N_11759,N_11735);
xnor U12755 (N_12755,N_11432,N_11304);
or U12756 (N_12756,N_11824,N_11278);
or U12757 (N_12757,N_11359,N_11941);
xor U12758 (N_12758,N_11717,N_11508);
or U12759 (N_12759,N_11436,N_11528);
or U12760 (N_12760,N_11790,N_11491);
nor U12761 (N_12761,N_11655,N_11920);
nand U12762 (N_12762,N_11904,N_11682);
nand U12763 (N_12763,N_11876,N_11912);
nor U12764 (N_12764,N_11902,N_11829);
and U12765 (N_12765,N_11353,N_11699);
xor U12766 (N_12766,N_11788,N_11734);
nor U12767 (N_12767,N_11992,N_11869);
or U12768 (N_12768,N_11546,N_11609);
xor U12769 (N_12769,N_11276,N_11879);
xor U12770 (N_12770,N_11331,N_11900);
and U12771 (N_12771,N_11726,N_11620);
and U12772 (N_12772,N_11919,N_11875);
nand U12773 (N_12773,N_11947,N_11706);
and U12774 (N_12774,N_11989,N_11904);
or U12775 (N_12775,N_11587,N_11363);
nor U12776 (N_12776,N_11936,N_11552);
nor U12777 (N_12777,N_11368,N_11870);
nor U12778 (N_12778,N_11202,N_11737);
or U12779 (N_12779,N_11427,N_11844);
and U12780 (N_12780,N_11582,N_11459);
or U12781 (N_12781,N_11604,N_11551);
or U12782 (N_12782,N_11870,N_11604);
xor U12783 (N_12783,N_11860,N_11523);
xor U12784 (N_12784,N_11854,N_11271);
nand U12785 (N_12785,N_11865,N_11740);
xor U12786 (N_12786,N_11523,N_11800);
xnor U12787 (N_12787,N_11608,N_11859);
or U12788 (N_12788,N_11617,N_11292);
nor U12789 (N_12789,N_11280,N_11805);
nor U12790 (N_12790,N_11492,N_11266);
nand U12791 (N_12791,N_11269,N_11947);
and U12792 (N_12792,N_11699,N_11328);
and U12793 (N_12793,N_11556,N_11507);
or U12794 (N_12794,N_11399,N_11831);
nor U12795 (N_12795,N_11758,N_11757);
or U12796 (N_12796,N_11772,N_11893);
nor U12797 (N_12797,N_11581,N_11819);
or U12798 (N_12798,N_11264,N_11891);
nand U12799 (N_12799,N_11355,N_11413);
xor U12800 (N_12800,N_12327,N_12483);
or U12801 (N_12801,N_12496,N_12727);
nor U12802 (N_12802,N_12619,N_12288);
xor U12803 (N_12803,N_12768,N_12644);
or U12804 (N_12804,N_12588,N_12354);
and U12805 (N_12805,N_12450,N_12543);
nand U12806 (N_12806,N_12023,N_12088);
and U12807 (N_12807,N_12604,N_12099);
and U12808 (N_12808,N_12469,N_12117);
nand U12809 (N_12809,N_12784,N_12539);
and U12810 (N_12810,N_12172,N_12092);
xor U12811 (N_12811,N_12057,N_12187);
or U12812 (N_12812,N_12050,N_12038);
nand U12813 (N_12813,N_12674,N_12150);
nand U12814 (N_12814,N_12458,N_12005);
nand U12815 (N_12815,N_12586,N_12340);
or U12816 (N_12816,N_12369,N_12140);
nand U12817 (N_12817,N_12781,N_12213);
xnor U12818 (N_12818,N_12090,N_12170);
or U12819 (N_12819,N_12773,N_12281);
and U12820 (N_12820,N_12589,N_12331);
and U12821 (N_12821,N_12221,N_12168);
or U12822 (N_12822,N_12356,N_12471);
nor U12823 (N_12823,N_12617,N_12308);
nor U12824 (N_12824,N_12279,N_12511);
and U12825 (N_12825,N_12384,N_12366);
nand U12826 (N_12826,N_12008,N_12510);
xor U12827 (N_12827,N_12111,N_12525);
and U12828 (N_12828,N_12612,N_12519);
nor U12829 (N_12829,N_12045,N_12782);
nor U12830 (N_12830,N_12318,N_12553);
and U12831 (N_12831,N_12767,N_12635);
xor U12832 (N_12832,N_12376,N_12724);
and U12833 (N_12833,N_12418,N_12737);
or U12834 (N_12834,N_12098,N_12192);
or U12835 (N_12835,N_12438,N_12058);
nor U12836 (N_12836,N_12078,N_12443);
nor U12837 (N_12837,N_12248,N_12252);
nor U12838 (N_12838,N_12176,N_12738);
xnor U12839 (N_12839,N_12052,N_12367);
and U12840 (N_12840,N_12199,N_12591);
nor U12841 (N_12841,N_12363,N_12417);
xor U12842 (N_12842,N_12527,N_12601);
nand U12843 (N_12843,N_12555,N_12382);
nor U12844 (N_12844,N_12643,N_12787);
and U12845 (N_12845,N_12600,N_12693);
and U12846 (N_12846,N_12607,N_12731);
nor U12847 (N_12847,N_12069,N_12408);
nand U12848 (N_12848,N_12200,N_12236);
nor U12849 (N_12849,N_12720,N_12013);
nor U12850 (N_12850,N_12122,N_12173);
or U12851 (N_12851,N_12270,N_12735);
nand U12852 (N_12852,N_12549,N_12572);
and U12853 (N_12853,N_12665,N_12491);
nand U12854 (N_12854,N_12663,N_12733);
and U12855 (N_12855,N_12700,N_12383);
or U12856 (N_12856,N_12155,N_12680);
or U12857 (N_12857,N_12159,N_12753);
nor U12858 (N_12858,N_12602,N_12289);
xnor U12859 (N_12859,N_12285,N_12436);
nor U12860 (N_12860,N_12029,N_12701);
or U12861 (N_12861,N_12178,N_12158);
or U12862 (N_12862,N_12467,N_12464);
nor U12863 (N_12863,N_12267,N_12495);
xor U12864 (N_12864,N_12147,N_12330);
xnor U12865 (N_12865,N_12097,N_12191);
nor U12866 (N_12866,N_12007,N_12286);
nand U12867 (N_12867,N_12235,N_12666);
nand U12868 (N_12868,N_12163,N_12296);
xnor U12869 (N_12869,N_12262,N_12444);
and U12870 (N_12870,N_12370,N_12004);
nor U12871 (N_12871,N_12009,N_12681);
and U12872 (N_12872,N_12247,N_12695);
nand U12873 (N_12873,N_12125,N_12403);
or U12874 (N_12874,N_12217,N_12710);
nand U12875 (N_12875,N_12068,N_12110);
nand U12876 (N_12876,N_12489,N_12410);
nand U12877 (N_12877,N_12258,N_12368);
or U12878 (N_12878,N_12031,N_12709);
and U12879 (N_12879,N_12646,N_12578);
nand U12880 (N_12880,N_12307,N_12184);
or U12881 (N_12881,N_12290,N_12630);
or U12882 (N_12882,N_12425,N_12636);
or U12883 (N_12883,N_12295,N_12722);
nand U12884 (N_12884,N_12419,N_12703);
or U12885 (N_12885,N_12723,N_12545);
nand U12886 (N_12886,N_12439,N_12357);
nor U12887 (N_12887,N_12713,N_12512);
nor U12888 (N_12888,N_12675,N_12291);
or U12889 (N_12889,N_12528,N_12162);
or U12890 (N_12890,N_12317,N_12338);
and U12891 (N_12891,N_12181,N_12596);
or U12892 (N_12892,N_12476,N_12309);
or U12893 (N_12893,N_12791,N_12079);
nor U12894 (N_12894,N_12256,N_12441);
and U12895 (N_12895,N_12505,N_12668);
or U12896 (N_12896,N_12345,N_12397);
nor U12897 (N_12897,N_12466,N_12740);
or U12898 (N_12898,N_12673,N_12141);
xor U12899 (N_12899,N_12287,N_12603);
xnor U12900 (N_12900,N_12440,N_12581);
and U12901 (N_12901,N_12284,N_12412);
nor U12902 (N_12902,N_12540,N_12796);
xor U12903 (N_12903,N_12560,N_12435);
nor U12904 (N_12904,N_12224,N_12255);
and U12905 (N_12905,N_12576,N_12210);
nand U12906 (N_12906,N_12660,N_12592);
or U12907 (N_12907,N_12715,N_12716);
xor U12908 (N_12908,N_12315,N_12361);
and U12909 (N_12909,N_12018,N_12563);
or U12910 (N_12910,N_12334,N_12485);
and U12911 (N_12911,N_12022,N_12532);
nor U12912 (N_12912,N_12146,N_12303);
xnor U12913 (N_12913,N_12772,N_12550);
and U12914 (N_12914,N_12725,N_12011);
nor U12915 (N_12915,N_12034,N_12437);
nor U12916 (N_12916,N_12794,N_12647);
and U12917 (N_12917,N_12396,N_12142);
nand U12918 (N_12918,N_12554,N_12135);
and U12919 (N_12919,N_12153,N_12786);
or U12920 (N_12920,N_12131,N_12475);
and U12921 (N_12921,N_12112,N_12770);
nor U12922 (N_12922,N_12442,N_12492);
xnor U12923 (N_12923,N_12537,N_12652);
nand U12924 (N_12924,N_12204,N_12292);
or U12925 (N_12925,N_12661,N_12413);
xnor U12926 (N_12926,N_12712,N_12745);
and U12927 (N_12927,N_12728,N_12667);
and U12928 (N_12928,N_12348,N_12730);
nor U12929 (N_12929,N_12502,N_12465);
xor U12930 (N_12930,N_12708,N_12126);
nand U12931 (N_12931,N_12228,N_12503);
or U12932 (N_12932,N_12683,N_12324);
and U12933 (N_12933,N_12169,N_12624);
xnor U12934 (N_12934,N_12477,N_12254);
or U12935 (N_12935,N_12275,N_12257);
nand U12936 (N_12936,N_12342,N_12676);
and U12937 (N_12937,N_12721,N_12684);
xor U12938 (N_12938,N_12616,N_12096);
nor U12939 (N_12939,N_12016,N_12197);
and U12940 (N_12940,N_12598,N_12774);
xor U12941 (N_12941,N_12574,N_12251);
xor U12942 (N_12942,N_12139,N_12468);
or U12943 (N_12943,N_12748,N_12570);
nand U12944 (N_12944,N_12121,N_12427);
nand U12945 (N_12945,N_12755,N_12487);
or U12946 (N_12946,N_12167,N_12148);
nor U12947 (N_12947,N_12628,N_12185);
xor U12948 (N_12948,N_12564,N_12350);
and U12949 (N_12949,N_12638,N_12229);
and U12950 (N_12950,N_12205,N_12717);
xnor U12951 (N_12951,N_12025,N_12634);
and U12952 (N_12952,N_12779,N_12156);
xor U12953 (N_12953,N_12060,N_12494);
or U12954 (N_12954,N_12249,N_12653);
and U12955 (N_12955,N_12014,N_12758);
nor U12956 (N_12956,N_12546,N_12416);
nor U12957 (N_12957,N_12694,N_12788);
or U12958 (N_12958,N_12411,N_12744);
xor U12959 (N_12959,N_12565,N_12119);
xnor U12960 (N_12960,N_12201,N_12035);
nor U12961 (N_12961,N_12750,N_12455);
xnor U12962 (N_12962,N_12107,N_12032);
nand U12963 (N_12963,N_12103,N_12319);
or U12964 (N_12964,N_12343,N_12682);
xnor U12965 (N_12965,N_12568,N_12529);
xnor U12966 (N_12966,N_12102,N_12658);
nor U12967 (N_12967,N_12518,N_12585);
nor U12968 (N_12968,N_12329,N_12771);
or U12969 (N_12969,N_12394,N_12209);
nor U12970 (N_12970,N_12669,N_12797);
nand U12971 (N_12971,N_12552,N_12390);
or U12972 (N_12972,N_12792,N_12633);
and U12973 (N_12973,N_12595,N_12691);
and U12974 (N_12974,N_12049,N_12759);
nand U12975 (N_12975,N_12061,N_12372);
nor U12976 (N_12976,N_12451,N_12705);
xor U12977 (N_12977,N_12645,N_12375);
xor U12978 (N_12978,N_12180,N_12493);
nand U12979 (N_12979,N_12130,N_12692);
xnor U12980 (N_12980,N_12323,N_12063);
or U12981 (N_12981,N_12697,N_12349);
and U12982 (N_12982,N_12777,N_12017);
xnor U12983 (N_12983,N_12182,N_12196);
xnor U12984 (N_12984,N_12120,N_12672);
nor U12985 (N_12985,N_12763,N_12274);
or U12986 (N_12986,N_12015,N_12039);
nor U12987 (N_12987,N_12339,N_12073);
xnor U12988 (N_12988,N_12202,N_12127);
xor U12989 (N_12989,N_12143,N_12082);
nand U12990 (N_12990,N_12152,N_12314);
nand U12991 (N_12991,N_12402,N_12044);
and U12992 (N_12992,N_12230,N_12104);
nor U12993 (N_12993,N_12608,N_12632);
or U12994 (N_12994,N_12190,N_12640);
nand U12995 (N_12995,N_12071,N_12136);
xor U12996 (N_12996,N_12655,N_12749);
and U12997 (N_12997,N_12567,N_12028);
nand U12998 (N_12998,N_12040,N_12116);
and U12999 (N_12999,N_12515,N_12409);
nand U13000 (N_13000,N_12359,N_12268);
nand U13001 (N_13001,N_12179,N_12580);
and U13002 (N_13002,N_12571,N_12304);
or U13003 (N_13003,N_12757,N_12206);
nand U13004 (N_13004,N_12093,N_12431);
nand U13005 (N_13005,N_12726,N_12462);
nand U13006 (N_13006,N_12280,N_12743);
nand U13007 (N_13007,N_12649,N_12795);
nand U13008 (N_13008,N_12569,N_12393);
xnor U13009 (N_13009,N_12461,N_12799);
nand U13010 (N_13010,N_12002,N_12548);
or U13011 (N_13011,N_12301,N_12651);
xnor U13012 (N_13012,N_12445,N_12610);
xnor U13013 (N_13013,N_12074,N_12095);
xor U13014 (N_13014,N_12566,N_12706);
and U13015 (N_13015,N_12526,N_12648);
or U13016 (N_13016,N_12488,N_12584);
nor U13017 (N_13017,N_12059,N_12123);
xor U13018 (N_13018,N_12227,N_12457);
and U13019 (N_13019,N_12046,N_12144);
xnor U13020 (N_13020,N_12283,N_12497);
nor U13021 (N_13021,N_12133,N_12037);
nand U13022 (N_13022,N_12358,N_12747);
and U13023 (N_13023,N_12702,N_12341);
or U13024 (N_13024,N_12704,N_12534);
and U13025 (N_13025,N_12310,N_12083);
nor U13026 (N_13026,N_12042,N_12535);
nor U13027 (N_13027,N_12094,N_12305);
or U13028 (N_13028,N_12793,N_12003);
nand U13029 (N_13029,N_12513,N_12657);
nor U13030 (N_13030,N_12531,N_12398);
xor U13031 (N_13031,N_12212,N_12400);
or U13032 (N_13032,N_12211,N_12664);
or U13033 (N_13033,N_12226,N_12689);
nor U13034 (N_13034,N_12353,N_12484);
nand U13035 (N_13035,N_12686,N_12481);
or U13036 (N_13036,N_12377,N_12208);
xnor U13037 (N_13037,N_12010,N_12798);
xnor U13038 (N_13038,N_12091,N_12420);
and U13039 (N_13039,N_12193,N_12240);
nor U13040 (N_13040,N_12297,N_12105);
nor U13041 (N_13041,N_12764,N_12429);
and U13042 (N_13042,N_12177,N_12790);
xnor U13043 (N_13043,N_12500,N_12081);
or U13044 (N_13044,N_12473,N_12277);
and U13045 (N_13045,N_12355,N_12312);
xnor U13046 (N_13046,N_12752,N_12401);
nand U13047 (N_13047,N_12734,N_12785);
xor U13048 (N_13048,N_12611,N_12276);
nand U13049 (N_13049,N_12609,N_12084);
nor U13050 (N_13050,N_12106,N_12222);
or U13051 (N_13051,N_12459,N_12250);
or U13052 (N_13052,N_12021,N_12207);
nor U13053 (N_13053,N_12020,N_12536);
or U13054 (N_13054,N_12129,N_12298);
nor U13055 (N_13055,N_12587,N_12508);
nor U13056 (N_13056,N_12605,N_12718);
nor U13057 (N_13057,N_12762,N_12072);
and U13058 (N_13058,N_12080,N_12335);
nor U13059 (N_13059,N_12599,N_12621);
nand U13060 (N_13060,N_12360,N_12165);
nand U13061 (N_13061,N_12577,N_12428);
nor U13062 (N_13062,N_12538,N_12326);
and U13063 (N_13063,N_12062,N_12769);
and U13064 (N_13064,N_12421,N_12741);
nor U13065 (N_13065,N_12556,N_12195);
xnor U13066 (N_13066,N_12659,N_12504);
and U13067 (N_13067,N_12688,N_12478);
and U13068 (N_13068,N_12597,N_12313);
nand U13069 (N_13069,N_12365,N_12265);
xnor U13070 (N_13070,N_12378,N_12479);
or U13071 (N_13071,N_12637,N_12460);
nor U13072 (N_13072,N_12043,N_12364);
xor U13073 (N_13073,N_12087,N_12362);
nor U13074 (N_13074,N_12189,N_12244);
and U13075 (N_13075,N_12124,N_12373);
nand U13076 (N_13076,N_12732,N_12754);
nor U13077 (N_13077,N_12054,N_12399);
and U13078 (N_13078,N_12593,N_12171);
nand U13079 (N_13079,N_12294,N_12328);
xor U13080 (N_13080,N_12100,N_12542);
nor U13081 (N_13081,N_12070,N_12241);
nand U13082 (N_13082,N_12690,N_12499);
nand U13083 (N_13083,N_12547,N_12389);
and U13084 (N_13084,N_12064,N_12371);
nor U13085 (N_13085,N_12203,N_12077);
or U13086 (N_13086,N_12789,N_12641);
or U13087 (N_13087,N_12223,N_12259);
nor U13088 (N_13088,N_12742,N_12490);
or U13089 (N_13089,N_12387,N_12344);
and U13090 (N_13090,N_12385,N_12557);
or U13091 (N_13091,N_12001,N_12594);
and U13092 (N_13092,N_12024,N_12656);
xnor U13093 (N_13093,N_12134,N_12678);
xor U13094 (N_13094,N_12260,N_12216);
xnor U13095 (N_13095,N_12448,N_12245);
nor U13096 (N_13096,N_12562,N_12685);
nor U13097 (N_13097,N_12422,N_12426);
nand U13098 (N_13098,N_12622,N_12474);
xnor U13099 (N_13099,N_12756,N_12320);
xor U13100 (N_13100,N_12639,N_12388);
nor U13101 (N_13101,N_12533,N_12101);
nor U13102 (N_13102,N_12631,N_12414);
nand U13103 (N_13103,N_12620,N_12423);
or U13104 (N_13104,N_12530,N_12233);
xor U13105 (N_13105,N_12115,N_12671);
or U13106 (N_13106,N_12332,N_12379);
nor U13107 (N_13107,N_12606,N_12128);
and U13108 (N_13108,N_12114,N_12108);
nor U13109 (N_13109,N_12424,N_12157);
or U13110 (N_13110,N_12246,N_12337);
or U13111 (N_13111,N_12273,N_12579);
xor U13112 (N_13112,N_12415,N_12000);
or U13113 (N_13113,N_12027,N_12736);
nand U13114 (N_13114,N_12089,N_12166);
or U13115 (N_13115,N_12696,N_12778);
xnor U13116 (N_13116,N_12719,N_12521);
and U13117 (N_13117,N_12149,N_12541);
nand U13118 (N_13118,N_12293,N_12454);
nor U13119 (N_13119,N_12041,N_12558);
nand U13120 (N_13120,N_12306,N_12266);
nor U13121 (N_13121,N_12780,N_12272);
nor U13122 (N_13122,N_12514,N_12160);
or U13123 (N_13123,N_12463,N_12615);
nor U13124 (N_13124,N_12407,N_12761);
xor U13125 (N_13125,N_12739,N_12218);
nand U13126 (N_13126,N_12381,N_12056);
xnor U13127 (N_13127,N_12447,N_12670);
or U13128 (N_13128,N_12507,N_12237);
or U13129 (N_13129,N_12405,N_12012);
or U13130 (N_13130,N_12629,N_12433);
nand U13131 (N_13131,N_12452,N_12524);
and U13132 (N_13132,N_12006,N_12300);
nor U13133 (N_13133,N_12234,N_12188);
nor U13134 (N_13134,N_12776,N_12746);
xor U13135 (N_13135,N_12480,N_12582);
nand U13136 (N_13136,N_12783,N_12198);
nor U13137 (N_13137,N_12765,N_12194);
nor U13138 (N_13138,N_12085,N_12699);
nor U13139 (N_13139,N_12517,N_12453);
nor U13140 (N_13140,N_12642,N_12374);
and U13141 (N_13141,N_12430,N_12161);
and U13142 (N_13142,N_12271,N_12316);
and U13143 (N_13143,N_12775,N_12751);
nor U13144 (N_13144,N_12264,N_12714);
and U13145 (N_13145,N_12109,N_12076);
xor U13146 (N_13146,N_12623,N_12446);
nor U13147 (N_13147,N_12520,N_12498);
and U13148 (N_13148,N_12154,N_12030);
and U13149 (N_13149,N_12352,N_12231);
nand U13150 (N_13150,N_12174,N_12687);
nor U13151 (N_13151,N_12346,N_12075);
nor U13152 (N_13152,N_12066,N_12132);
or U13153 (N_13153,N_12501,N_12321);
and U13154 (N_13154,N_12729,N_12626);
or U13155 (N_13155,N_12573,N_12559);
xor U13156 (N_13156,N_12164,N_12048);
and U13157 (N_13157,N_12766,N_12220);
and U13158 (N_13158,N_12386,N_12033);
nand U13159 (N_13159,N_12261,N_12138);
or U13160 (N_13160,N_12711,N_12065);
and U13161 (N_13161,N_12239,N_12051);
and U13162 (N_13162,N_12186,N_12036);
nor U13163 (N_13163,N_12395,N_12137);
xnor U13164 (N_13164,N_12055,N_12561);
xnor U13165 (N_13165,N_12232,N_12456);
or U13166 (N_13166,N_12575,N_12242);
nand U13167 (N_13167,N_12047,N_12053);
or U13168 (N_13168,N_12432,N_12067);
nor U13169 (N_13169,N_12322,N_12225);
or U13170 (N_13170,N_12392,N_12613);
nor U13171 (N_13171,N_12391,N_12472);
and U13172 (N_13172,N_12299,N_12614);
or U13173 (N_13173,N_12311,N_12679);
nand U13174 (N_13174,N_12650,N_12509);
and U13175 (N_13175,N_12618,N_12677);
and U13176 (N_13176,N_12625,N_12151);
and U13177 (N_13177,N_12183,N_12175);
nand U13178 (N_13178,N_12551,N_12760);
or U13179 (N_13179,N_12238,N_12333);
and U13180 (N_13180,N_12406,N_12253);
and U13181 (N_13181,N_12026,N_12282);
nor U13182 (N_13182,N_12544,N_12434);
nor U13183 (N_13183,N_12118,N_12351);
nor U13184 (N_13184,N_12019,N_12523);
nor U13185 (N_13185,N_12269,N_12219);
or U13186 (N_13186,N_12662,N_12380);
and U13187 (N_13187,N_12449,N_12243);
nand U13188 (N_13188,N_12482,N_12698);
and U13189 (N_13189,N_12086,N_12336);
nor U13190 (N_13190,N_12486,N_12583);
or U13191 (N_13191,N_12263,N_12516);
nor U13192 (N_13192,N_12707,N_12470);
and U13193 (N_13193,N_12404,N_12522);
and U13194 (N_13194,N_12278,N_12654);
and U13195 (N_13195,N_12627,N_12145);
xnor U13196 (N_13196,N_12506,N_12113);
xnor U13197 (N_13197,N_12325,N_12590);
and U13198 (N_13198,N_12347,N_12214);
and U13199 (N_13199,N_12302,N_12215);
and U13200 (N_13200,N_12639,N_12313);
nor U13201 (N_13201,N_12189,N_12210);
or U13202 (N_13202,N_12671,N_12460);
nor U13203 (N_13203,N_12444,N_12371);
and U13204 (N_13204,N_12793,N_12752);
nor U13205 (N_13205,N_12691,N_12766);
or U13206 (N_13206,N_12272,N_12497);
nand U13207 (N_13207,N_12772,N_12137);
and U13208 (N_13208,N_12274,N_12593);
nor U13209 (N_13209,N_12480,N_12578);
nor U13210 (N_13210,N_12197,N_12061);
nor U13211 (N_13211,N_12196,N_12407);
nand U13212 (N_13212,N_12129,N_12706);
and U13213 (N_13213,N_12610,N_12249);
nand U13214 (N_13214,N_12412,N_12121);
and U13215 (N_13215,N_12206,N_12398);
xnor U13216 (N_13216,N_12199,N_12727);
nor U13217 (N_13217,N_12792,N_12442);
and U13218 (N_13218,N_12457,N_12226);
nor U13219 (N_13219,N_12565,N_12695);
xnor U13220 (N_13220,N_12728,N_12796);
and U13221 (N_13221,N_12455,N_12260);
or U13222 (N_13222,N_12694,N_12307);
xor U13223 (N_13223,N_12766,N_12416);
nand U13224 (N_13224,N_12035,N_12147);
or U13225 (N_13225,N_12228,N_12649);
and U13226 (N_13226,N_12326,N_12579);
xnor U13227 (N_13227,N_12502,N_12739);
xor U13228 (N_13228,N_12772,N_12787);
nor U13229 (N_13229,N_12515,N_12544);
xor U13230 (N_13230,N_12409,N_12735);
or U13231 (N_13231,N_12075,N_12331);
nand U13232 (N_13232,N_12768,N_12568);
nand U13233 (N_13233,N_12728,N_12357);
or U13234 (N_13234,N_12770,N_12798);
and U13235 (N_13235,N_12785,N_12398);
nor U13236 (N_13236,N_12337,N_12701);
xor U13237 (N_13237,N_12054,N_12333);
xnor U13238 (N_13238,N_12588,N_12242);
and U13239 (N_13239,N_12197,N_12183);
xor U13240 (N_13240,N_12220,N_12671);
or U13241 (N_13241,N_12696,N_12398);
nand U13242 (N_13242,N_12255,N_12597);
xor U13243 (N_13243,N_12123,N_12797);
xor U13244 (N_13244,N_12738,N_12484);
nand U13245 (N_13245,N_12053,N_12493);
nand U13246 (N_13246,N_12473,N_12098);
xnor U13247 (N_13247,N_12104,N_12435);
or U13248 (N_13248,N_12395,N_12497);
and U13249 (N_13249,N_12772,N_12588);
and U13250 (N_13250,N_12133,N_12209);
and U13251 (N_13251,N_12737,N_12633);
nor U13252 (N_13252,N_12122,N_12655);
and U13253 (N_13253,N_12078,N_12492);
nand U13254 (N_13254,N_12136,N_12534);
xnor U13255 (N_13255,N_12052,N_12313);
nand U13256 (N_13256,N_12092,N_12589);
or U13257 (N_13257,N_12433,N_12357);
xor U13258 (N_13258,N_12379,N_12502);
nor U13259 (N_13259,N_12323,N_12019);
nand U13260 (N_13260,N_12668,N_12313);
xor U13261 (N_13261,N_12456,N_12580);
xnor U13262 (N_13262,N_12085,N_12335);
xor U13263 (N_13263,N_12464,N_12630);
and U13264 (N_13264,N_12106,N_12480);
and U13265 (N_13265,N_12109,N_12088);
xnor U13266 (N_13266,N_12016,N_12587);
nand U13267 (N_13267,N_12022,N_12036);
nand U13268 (N_13268,N_12239,N_12664);
xnor U13269 (N_13269,N_12718,N_12499);
xor U13270 (N_13270,N_12478,N_12056);
xnor U13271 (N_13271,N_12724,N_12134);
and U13272 (N_13272,N_12116,N_12599);
nor U13273 (N_13273,N_12722,N_12088);
and U13274 (N_13274,N_12331,N_12203);
nor U13275 (N_13275,N_12718,N_12525);
nand U13276 (N_13276,N_12462,N_12322);
nor U13277 (N_13277,N_12663,N_12734);
nand U13278 (N_13278,N_12227,N_12507);
and U13279 (N_13279,N_12494,N_12217);
xnor U13280 (N_13280,N_12560,N_12463);
and U13281 (N_13281,N_12335,N_12653);
and U13282 (N_13282,N_12196,N_12431);
nor U13283 (N_13283,N_12632,N_12579);
or U13284 (N_13284,N_12268,N_12698);
nand U13285 (N_13285,N_12708,N_12620);
or U13286 (N_13286,N_12281,N_12400);
and U13287 (N_13287,N_12687,N_12105);
xor U13288 (N_13288,N_12533,N_12539);
nand U13289 (N_13289,N_12465,N_12067);
nor U13290 (N_13290,N_12662,N_12603);
or U13291 (N_13291,N_12479,N_12179);
nand U13292 (N_13292,N_12076,N_12377);
xor U13293 (N_13293,N_12546,N_12290);
and U13294 (N_13294,N_12088,N_12724);
nand U13295 (N_13295,N_12114,N_12237);
or U13296 (N_13296,N_12259,N_12609);
or U13297 (N_13297,N_12713,N_12724);
nor U13298 (N_13298,N_12345,N_12420);
or U13299 (N_13299,N_12735,N_12681);
or U13300 (N_13300,N_12036,N_12241);
nand U13301 (N_13301,N_12296,N_12166);
or U13302 (N_13302,N_12207,N_12512);
xnor U13303 (N_13303,N_12349,N_12362);
and U13304 (N_13304,N_12233,N_12239);
nor U13305 (N_13305,N_12242,N_12634);
nor U13306 (N_13306,N_12232,N_12497);
and U13307 (N_13307,N_12752,N_12402);
or U13308 (N_13308,N_12729,N_12688);
or U13309 (N_13309,N_12560,N_12563);
nand U13310 (N_13310,N_12748,N_12616);
and U13311 (N_13311,N_12322,N_12543);
xor U13312 (N_13312,N_12032,N_12555);
xor U13313 (N_13313,N_12713,N_12166);
nor U13314 (N_13314,N_12376,N_12440);
and U13315 (N_13315,N_12663,N_12478);
nand U13316 (N_13316,N_12002,N_12397);
nor U13317 (N_13317,N_12510,N_12481);
nand U13318 (N_13318,N_12689,N_12113);
and U13319 (N_13319,N_12289,N_12604);
nand U13320 (N_13320,N_12298,N_12677);
and U13321 (N_13321,N_12792,N_12588);
or U13322 (N_13322,N_12557,N_12295);
xnor U13323 (N_13323,N_12216,N_12222);
or U13324 (N_13324,N_12392,N_12029);
xnor U13325 (N_13325,N_12272,N_12094);
nand U13326 (N_13326,N_12405,N_12018);
nor U13327 (N_13327,N_12558,N_12127);
xnor U13328 (N_13328,N_12775,N_12546);
and U13329 (N_13329,N_12181,N_12100);
and U13330 (N_13330,N_12674,N_12066);
and U13331 (N_13331,N_12056,N_12131);
or U13332 (N_13332,N_12416,N_12380);
nand U13333 (N_13333,N_12398,N_12642);
xor U13334 (N_13334,N_12016,N_12270);
nand U13335 (N_13335,N_12072,N_12459);
nor U13336 (N_13336,N_12449,N_12083);
xor U13337 (N_13337,N_12303,N_12782);
and U13338 (N_13338,N_12139,N_12005);
nor U13339 (N_13339,N_12127,N_12471);
nand U13340 (N_13340,N_12165,N_12586);
and U13341 (N_13341,N_12125,N_12565);
or U13342 (N_13342,N_12257,N_12304);
xnor U13343 (N_13343,N_12075,N_12482);
and U13344 (N_13344,N_12261,N_12224);
or U13345 (N_13345,N_12662,N_12114);
xor U13346 (N_13346,N_12658,N_12605);
xor U13347 (N_13347,N_12690,N_12739);
nor U13348 (N_13348,N_12784,N_12031);
and U13349 (N_13349,N_12467,N_12010);
or U13350 (N_13350,N_12481,N_12068);
xor U13351 (N_13351,N_12250,N_12446);
nand U13352 (N_13352,N_12745,N_12552);
xnor U13353 (N_13353,N_12215,N_12233);
nand U13354 (N_13354,N_12001,N_12097);
nand U13355 (N_13355,N_12594,N_12362);
xnor U13356 (N_13356,N_12359,N_12339);
and U13357 (N_13357,N_12125,N_12453);
or U13358 (N_13358,N_12570,N_12301);
and U13359 (N_13359,N_12226,N_12339);
or U13360 (N_13360,N_12514,N_12494);
or U13361 (N_13361,N_12239,N_12591);
nand U13362 (N_13362,N_12161,N_12527);
nand U13363 (N_13363,N_12722,N_12729);
nor U13364 (N_13364,N_12655,N_12154);
nand U13365 (N_13365,N_12317,N_12577);
nand U13366 (N_13366,N_12691,N_12217);
nor U13367 (N_13367,N_12577,N_12397);
nor U13368 (N_13368,N_12687,N_12319);
or U13369 (N_13369,N_12345,N_12753);
or U13370 (N_13370,N_12606,N_12205);
nor U13371 (N_13371,N_12607,N_12734);
or U13372 (N_13372,N_12789,N_12153);
nand U13373 (N_13373,N_12650,N_12287);
xnor U13374 (N_13374,N_12115,N_12087);
nand U13375 (N_13375,N_12703,N_12293);
nor U13376 (N_13376,N_12095,N_12337);
xor U13377 (N_13377,N_12429,N_12066);
or U13378 (N_13378,N_12450,N_12208);
nand U13379 (N_13379,N_12324,N_12589);
or U13380 (N_13380,N_12614,N_12050);
nand U13381 (N_13381,N_12717,N_12381);
nor U13382 (N_13382,N_12278,N_12361);
nand U13383 (N_13383,N_12523,N_12673);
xor U13384 (N_13384,N_12156,N_12457);
nor U13385 (N_13385,N_12373,N_12796);
nor U13386 (N_13386,N_12776,N_12458);
xnor U13387 (N_13387,N_12549,N_12399);
and U13388 (N_13388,N_12643,N_12394);
xnor U13389 (N_13389,N_12155,N_12379);
nor U13390 (N_13390,N_12304,N_12466);
nor U13391 (N_13391,N_12266,N_12113);
nor U13392 (N_13392,N_12534,N_12106);
or U13393 (N_13393,N_12524,N_12208);
xnor U13394 (N_13394,N_12678,N_12742);
nor U13395 (N_13395,N_12422,N_12765);
xnor U13396 (N_13396,N_12673,N_12152);
nand U13397 (N_13397,N_12010,N_12542);
nand U13398 (N_13398,N_12652,N_12416);
and U13399 (N_13399,N_12203,N_12138);
or U13400 (N_13400,N_12054,N_12142);
xor U13401 (N_13401,N_12490,N_12214);
xnor U13402 (N_13402,N_12411,N_12741);
and U13403 (N_13403,N_12383,N_12362);
nor U13404 (N_13404,N_12586,N_12445);
nand U13405 (N_13405,N_12405,N_12261);
nand U13406 (N_13406,N_12662,N_12607);
nor U13407 (N_13407,N_12744,N_12509);
and U13408 (N_13408,N_12030,N_12106);
nand U13409 (N_13409,N_12643,N_12346);
and U13410 (N_13410,N_12181,N_12474);
nor U13411 (N_13411,N_12440,N_12727);
nand U13412 (N_13412,N_12103,N_12794);
xnor U13413 (N_13413,N_12715,N_12662);
or U13414 (N_13414,N_12182,N_12078);
or U13415 (N_13415,N_12632,N_12006);
or U13416 (N_13416,N_12521,N_12343);
or U13417 (N_13417,N_12096,N_12225);
xor U13418 (N_13418,N_12027,N_12090);
xor U13419 (N_13419,N_12440,N_12009);
or U13420 (N_13420,N_12184,N_12447);
nand U13421 (N_13421,N_12443,N_12106);
xnor U13422 (N_13422,N_12474,N_12363);
nor U13423 (N_13423,N_12540,N_12383);
xor U13424 (N_13424,N_12398,N_12759);
xor U13425 (N_13425,N_12389,N_12116);
and U13426 (N_13426,N_12582,N_12178);
or U13427 (N_13427,N_12663,N_12466);
nor U13428 (N_13428,N_12597,N_12586);
or U13429 (N_13429,N_12735,N_12315);
and U13430 (N_13430,N_12455,N_12051);
and U13431 (N_13431,N_12073,N_12299);
nor U13432 (N_13432,N_12178,N_12703);
nand U13433 (N_13433,N_12415,N_12351);
nor U13434 (N_13434,N_12421,N_12066);
nor U13435 (N_13435,N_12759,N_12196);
and U13436 (N_13436,N_12497,N_12171);
xor U13437 (N_13437,N_12375,N_12755);
or U13438 (N_13438,N_12122,N_12613);
nand U13439 (N_13439,N_12071,N_12210);
or U13440 (N_13440,N_12309,N_12397);
nor U13441 (N_13441,N_12751,N_12100);
and U13442 (N_13442,N_12219,N_12632);
and U13443 (N_13443,N_12054,N_12563);
nor U13444 (N_13444,N_12356,N_12037);
nand U13445 (N_13445,N_12096,N_12142);
or U13446 (N_13446,N_12196,N_12329);
xor U13447 (N_13447,N_12020,N_12522);
and U13448 (N_13448,N_12786,N_12544);
and U13449 (N_13449,N_12449,N_12700);
xor U13450 (N_13450,N_12764,N_12586);
xnor U13451 (N_13451,N_12347,N_12357);
and U13452 (N_13452,N_12250,N_12430);
nor U13453 (N_13453,N_12020,N_12500);
nand U13454 (N_13454,N_12539,N_12025);
nor U13455 (N_13455,N_12388,N_12460);
nand U13456 (N_13456,N_12226,N_12202);
and U13457 (N_13457,N_12205,N_12044);
and U13458 (N_13458,N_12563,N_12280);
nor U13459 (N_13459,N_12425,N_12569);
and U13460 (N_13460,N_12038,N_12088);
and U13461 (N_13461,N_12764,N_12111);
or U13462 (N_13462,N_12392,N_12650);
nand U13463 (N_13463,N_12211,N_12483);
nor U13464 (N_13464,N_12432,N_12026);
nor U13465 (N_13465,N_12310,N_12427);
xor U13466 (N_13466,N_12448,N_12077);
nand U13467 (N_13467,N_12621,N_12103);
nor U13468 (N_13468,N_12041,N_12183);
xnor U13469 (N_13469,N_12693,N_12200);
nor U13470 (N_13470,N_12218,N_12448);
and U13471 (N_13471,N_12672,N_12009);
nand U13472 (N_13472,N_12798,N_12291);
or U13473 (N_13473,N_12361,N_12212);
or U13474 (N_13474,N_12041,N_12047);
nor U13475 (N_13475,N_12121,N_12654);
nand U13476 (N_13476,N_12782,N_12302);
xor U13477 (N_13477,N_12643,N_12755);
nand U13478 (N_13478,N_12384,N_12161);
or U13479 (N_13479,N_12653,N_12776);
nand U13480 (N_13480,N_12308,N_12656);
nor U13481 (N_13481,N_12770,N_12387);
nand U13482 (N_13482,N_12299,N_12678);
or U13483 (N_13483,N_12284,N_12036);
nor U13484 (N_13484,N_12008,N_12720);
nand U13485 (N_13485,N_12333,N_12084);
nor U13486 (N_13486,N_12514,N_12082);
or U13487 (N_13487,N_12004,N_12447);
xor U13488 (N_13488,N_12108,N_12707);
nand U13489 (N_13489,N_12750,N_12530);
nor U13490 (N_13490,N_12434,N_12472);
xor U13491 (N_13491,N_12328,N_12160);
nand U13492 (N_13492,N_12410,N_12150);
or U13493 (N_13493,N_12408,N_12499);
xor U13494 (N_13494,N_12526,N_12035);
nand U13495 (N_13495,N_12515,N_12498);
or U13496 (N_13496,N_12663,N_12120);
or U13497 (N_13497,N_12259,N_12551);
and U13498 (N_13498,N_12378,N_12030);
and U13499 (N_13499,N_12343,N_12029);
and U13500 (N_13500,N_12180,N_12457);
and U13501 (N_13501,N_12272,N_12147);
nand U13502 (N_13502,N_12695,N_12230);
nand U13503 (N_13503,N_12733,N_12432);
or U13504 (N_13504,N_12711,N_12027);
nor U13505 (N_13505,N_12190,N_12531);
or U13506 (N_13506,N_12075,N_12303);
xor U13507 (N_13507,N_12264,N_12249);
and U13508 (N_13508,N_12499,N_12733);
xnor U13509 (N_13509,N_12201,N_12099);
nand U13510 (N_13510,N_12499,N_12563);
or U13511 (N_13511,N_12769,N_12617);
and U13512 (N_13512,N_12691,N_12728);
and U13513 (N_13513,N_12466,N_12513);
xor U13514 (N_13514,N_12323,N_12481);
and U13515 (N_13515,N_12155,N_12533);
nand U13516 (N_13516,N_12650,N_12205);
xor U13517 (N_13517,N_12265,N_12549);
nor U13518 (N_13518,N_12477,N_12226);
nand U13519 (N_13519,N_12198,N_12563);
xor U13520 (N_13520,N_12602,N_12379);
xnor U13521 (N_13521,N_12711,N_12419);
xnor U13522 (N_13522,N_12391,N_12480);
nand U13523 (N_13523,N_12375,N_12799);
nand U13524 (N_13524,N_12741,N_12727);
nor U13525 (N_13525,N_12277,N_12017);
and U13526 (N_13526,N_12535,N_12163);
xnor U13527 (N_13527,N_12319,N_12100);
nor U13528 (N_13528,N_12556,N_12457);
nand U13529 (N_13529,N_12615,N_12554);
or U13530 (N_13530,N_12120,N_12714);
xor U13531 (N_13531,N_12182,N_12084);
nor U13532 (N_13532,N_12796,N_12494);
xnor U13533 (N_13533,N_12724,N_12082);
or U13534 (N_13534,N_12286,N_12700);
nor U13535 (N_13535,N_12175,N_12687);
and U13536 (N_13536,N_12486,N_12792);
nand U13537 (N_13537,N_12297,N_12773);
nand U13538 (N_13538,N_12433,N_12571);
and U13539 (N_13539,N_12764,N_12542);
nand U13540 (N_13540,N_12694,N_12439);
or U13541 (N_13541,N_12174,N_12320);
nand U13542 (N_13542,N_12579,N_12208);
xor U13543 (N_13543,N_12243,N_12133);
xnor U13544 (N_13544,N_12506,N_12038);
or U13545 (N_13545,N_12672,N_12741);
nor U13546 (N_13546,N_12589,N_12595);
nand U13547 (N_13547,N_12293,N_12212);
nor U13548 (N_13548,N_12197,N_12028);
xor U13549 (N_13549,N_12590,N_12611);
nand U13550 (N_13550,N_12656,N_12118);
xnor U13551 (N_13551,N_12112,N_12066);
nor U13552 (N_13552,N_12165,N_12674);
or U13553 (N_13553,N_12779,N_12001);
and U13554 (N_13554,N_12625,N_12158);
nand U13555 (N_13555,N_12728,N_12217);
or U13556 (N_13556,N_12345,N_12353);
and U13557 (N_13557,N_12581,N_12217);
nand U13558 (N_13558,N_12002,N_12040);
nor U13559 (N_13559,N_12758,N_12591);
and U13560 (N_13560,N_12319,N_12141);
xnor U13561 (N_13561,N_12408,N_12450);
or U13562 (N_13562,N_12612,N_12703);
or U13563 (N_13563,N_12647,N_12371);
and U13564 (N_13564,N_12285,N_12126);
nand U13565 (N_13565,N_12166,N_12591);
nand U13566 (N_13566,N_12702,N_12680);
xor U13567 (N_13567,N_12260,N_12255);
or U13568 (N_13568,N_12341,N_12503);
and U13569 (N_13569,N_12246,N_12320);
nand U13570 (N_13570,N_12438,N_12414);
nand U13571 (N_13571,N_12023,N_12760);
nor U13572 (N_13572,N_12331,N_12299);
nor U13573 (N_13573,N_12389,N_12641);
and U13574 (N_13574,N_12782,N_12546);
and U13575 (N_13575,N_12175,N_12711);
xor U13576 (N_13576,N_12643,N_12059);
and U13577 (N_13577,N_12190,N_12441);
nand U13578 (N_13578,N_12468,N_12496);
or U13579 (N_13579,N_12368,N_12440);
nor U13580 (N_13580,N_12650,N_12625);
or U13581 (N_13581,N_12099,N_12290);
xnor U13582 (N_13582,N_12245,N_12041);
xnor U13583 (N_13583,N_12157,N_12574);
nor U13584 (N_13584,N_12227,N_12407);
nand U13585 (N_13585,N_12784,N_12730);
nor U13586 (N_13586,N_12241,N_12522);
and U13587 (N_13587,N_12478,N_12516);
xnor U13588 (N_13588,N_12117,N_12680);
xor U13589 (N_13589,N_12556,N_12078);
and U13590 (N_13590,N_12391,N_12453);
and U13591 (N_13591,N_12334,N_12647);
xor U13592 (N_13592,N_12398,N_12386);
xnor U13593 (N_13593,N_12490,N_12110);
or U13594 (N_13594,N_12720,N_12090);
xor U13595 (N_13595,N_12349,N_12463);
nor U13596 (N_13596,N_12120,N_12248);
xor U13597 (N_13597,N_12120,N_12351);
xor U13598 (N_13598,N_12144,N_12006);
xor U13599 (N_13599,N_12040,N_12226);
nand U13600 (N_13600,N_13153,N_12901);
and U13601 (N_13601,N_12878,N_13003);
nand U13602 (N_13602,N_12936,N_13392);
xor U13603 (N_13603,N_13370,N_13404);
and U13604 (N_13604,N_12986,N_12910);
or U13605 (N_13605,N_13063,N_13120);
or U13606 (N_13606,N_12985,N_13199);
nor U13607 (N_13607,N_12871,N_13538);
xor U13608 (N_13608,N_13462,N_13200);
nand U13609 (N_13609,N_13517,N_12854);
xnor U13610 (N_13610,N_13220,N_12867);
or U13611 (N_13611,N_13324,N_12995);
nand U13612 (N_13612,N_13189,N_13436);
nand U13613 (N_13613,N_13505,N_13539);
nor U13614 (N_13614,N_13323,N_13276);
nand U13615 (N_13615,N_12969,N_13218);
nor U13616 (N_13616,N_12888,N_12813);
nand U13617 (N_13617,N_13183,N_13130);
or U13618 (N_13618,N_13408,N_12821);
nand U13619 (N_13619,N_13359,N_12832);
nor U13620 (N_13620,N_13108,N_12992);
or U13621 (N_13621,N_13221,N_13033);
xnor U13622 (N_13622,N_13504,N_12946);
and U13623 (N_13623,N_13048,N_13080);
nand U13624 (N_13624,N_13417,N_13001);
and U13625 (N_13625,N_13149,N_13371);
nor U13626 (N_13626,N_13467,N_13393);
or U13627 (N_13627,N_12926,N_13527);
or U13628 (N_13628,N_13055,N_13262);
nand U13629 (N_13629,N_13259,N_13077);
or U13630 (N_13630,N_13439,N_13308);
and U13631 (N_13631,N_13296,N_12998);
nand U13632 (N_13632,N_13512,N_13552);
nor U13633 (N_13633,N_13550,N_13249);
or U13634 (N_13634,N_13481,N_13314);
xnor U13635 (N_13635,N_13514,N_12864);
and U13636 (N_13636,N_13352,N_13533);
and U13637 (N_13637,N_13047,N_13483);
nor U13638 (N_13638,N_13415,N_12925);
xnor U13639 (N_13639,N_13398,N_13434);
and U13640 (N_13640,N_13469,N_13253);
and U13641 (N_13641,N_13555,N_13528);
nor U13642 (N_13642,N_12912,N_12918);
or U13643 (N_13643,N_12982,N_13433);
nor U13644 (N_13644,N_13111,N_13362);
and U13645 (N_13645,N_12853,N_13360);
and U13646 (N_13646,N_12991,N_13516);
nor U13647 (N_13647,N_13566,N_12805);
or U13648 (N_13648,N_13597,N_13133);
nand U13649 (N_13649,N_13228,N_13124);
xnor U13650 (N_13650,N_13287,N_13313);
nand U13651 (N_13651,N_13395,N_12807);
and U13652 (N_13652,N_13400,N_13087);
xnor U13653 (N_13653,N_12863,N_13160);
xnor U13654 (N_13654,N_12810,N_13523);
xnor U13655 (N_13655,N_13045,N_12856);
nor U13656 (N_13656,N_13180,N_12876);
nor U13657 (N_13657,N_13424,N_13591);
nand U13658 (N_13658,N_13092,N_13416);
and U13659 (N_13659,N_13449,N_13034);
nand U13660 (N_13660,N_13099,N_13163);
and U13661 (N_13661,N_12922,N_13302);
xnor U13662 (N_13662,N_12808,N_13530);
nor U13663 (N_13663,N_13260,N_13268);
nor U13664 (N_13664,N_13537,N_13458);
or U13665 (N_13665,N_13140,N_12989);
xor U13666 (N_13666,N_13511,N_13237);
and U13667 (N_13667,N_12839,N_12978);
nor U13668 (N_13668,N_13225,N_13201);
nor U13669 (N_13669,N_13212,N_13447);
and U13670 (N_13670,N_13122,N_13044);
nand U13671 (N_13671,N_12824,N_13599);
nand U13672 (N_13672,N_13049,N_13454);
xor U13673 (N_13673,N_12851,N_13182);
or U13674 (N_13674,N_13448,N_13509);
and U13675 (N_13675,N_13148,N_12885);
xor U13676 (N_13676,N_13236,N_13430);
nor U13677 (N_13677,N_13510,N_13191);
nor U13678 (N_13678,N_13508,N_13244);
xnor U13679 (N_13679,N_13580,N_12972);
nand U13680 (N_13680,N_13194,N_13506);
and U13681 (N_13681,N_12939,N_13355);
nor U13682 (N_13682,N_13142,N_13356);
nor U13683 (N_13683,N_13275,N_13305);
xnor U13684 (N_13684,N_13184,N_13116);
nor U13685 (N_13685,N_13471,N_12980);
and U13686 (N_13686,N_13094,N_13382);
and U13687 (N_13687,N_13503,N_13522);
nand U13688 (N_13688,N_13050,N_13345);
xor U13689 (N_13689,N_12861,N_13226);
or U13690 (N_13690,N_13559,N_12836);
and U13691 (N_13691,N_12932,N_12844);
nand U13692 (N_13692,N_13132,N_13227);
and U13693 (N_13693,N_13389,N_13329);
nand U13694 (N_13694,N_12873,N_13304);
nand U13695 (N_13695,N_13307,N_13038);
xor U13696 (N_13696,N_12865,N_13072);
or U13697 (N_13697,N_13411,N_13586);
and U13698 (N_13698,N_13068,N_13394);
and U13699 (N_13699,N_13401,N_13119);
nand U13700 (N_13700,N_13257,N_13380);
xnor U13701 (N_13701,N_13577,N_13455);
or U13702 (N_13702,N_13117,N_13565);
nand U13703 (N_13703,N_13294,N_12881);
nor U13704 (N_13704,N_13171,N_13057);
or U13705 (N_13705,N_13123,N_13542);
xor U13706 (N_13706,N_12815,N_13583);
and U13707 (N_13707,N_13562,N_13278);
nor U13708 (N_13708,N_13595,N_12875);
xor U13709 (N_13709,N_13106,N_13131);
and U13710 (N_13710,N_13279,N_13554);
xnor U13711 (N_13711,N_12957,N_12891);
nand U13712 (N_13712,N_13485,N_13426);
and U13713 (N_13713,N_13283,N_13342);
xor U13714 (N_13714,N_12840,N_13281);
or U13715 (N_13715,N_13385,N_13206);
and U13716 (N_13716,N_12850,N_13435);
or U13717 (N_13717,N_12977,N_13147);
xor U13718 (N_13718,N_13176,N_12830);
and U13719 (N_13719,N_13026,N_13493);
nand U13720 (N_13720,N_12937,N_13575);
nand U13721 (N_13721,N_13407,N_13128);
xor U13722 (N_13722,N_13386,N_12883);
or U13723 (N_13723,N_12874,N_12971);
nor U13724 (N_13724,N_13245,N_12921);
and U13725 (N_13725,N_13029,N_12984);
nor U13726 (N_13726,N_13334,N_12803);
nor U13727 (N_13727,N_13513,N_13306);
nand U13728 (N_13728,N_12823,N_13497);
nor U13729 (N_13729,N_13388,N_13053);
or U13730 (N_13730,N_12812,N_13054);
nor U13731 (N_13731,N_13520,N_13070);
and U13732 (N_13732,N_13097,N_12819);
xor U13733 (N_13733,N_13582,N_13335);
nor U13734 (N_13734,N_12827,N_13596);
xor U13735 (N_13735,N_12806,N_12965);
or U13736 (N_13736,N_12904,N_13250);
or U13737 (N_13737,N_12898,N_13195);
xnor U13738 (N_13738,N_13446,N_13476);
or U13739 (N_13739,N_13223,N_13325);
nand U13740 (N_13740,N_13548,N_13420);
and U13741 (N_13741,N_13322,N_13020);
nor U13742 (N_13742,N_13137,N_13000);
and U13743 (N_13743,N_13367,N_13037);
xnor U13744 (N_13744,N_12930,N_13112);
or U13745 (N_13745,N_13368,N_13079);
and U13746 (N_13746,N_12954,N_13081);
nand U13747 (N_13747,N_12802,N_13246);
nor U13748 (N_13748,N_13238,N_13406);
nand U13749 (N_13749,N_13272,N_13046);
or U13750 (N_13750,N_13491,N_13129);
nand U13751 (N_13751,N_13529,N_12983);
nand U13752 (N_13752,N_12988,N_13061);
xor U13753 (N_13753,N_13492,N_13031);
or U13754 (N_13754,N_13351,N_13211);
nand U13755 (N_13755,N_13310,N_13499);
and U13756 (N_13756,N_13549,N_13006);
nor U13757 (N_13757,N_12981,N_13175);
nand U13758 (N_13758,N_13480,N_13387);
nor U13759 (N_13759,N_13316,N_13340);
and U13760 (N_13760,N_13421,N_12947);
nor U13761 (N_13761,N_12869,N_13210);
nor U13762 (N_13762,N_12826,N_12835);
and U13763 (N_13763,N_12825,N_13576);
or U13764 (N_13764,N_13282,N_13203);
xor U13765 (N_13765,N_12811,N_12968);
or U13766 (N_13766,N_13377,N_13546);
nor U13767 (N_13767,N_13273,N_13572);
nand U13768 (N_13768,N_13564,N_12848);
or U13769 (N_13769,N_12841,N_13265);
or U13770 (N_13770,N_13178,N_13291);
nor U13771 (N_13771,N_13069,N_13012);
or U13772 (N_13772,N_13311,N_12817);
nor U13773 (N_13773,N_13254,N_12996);
or U13774 (N_13774,N_12934,N_13010);
or U13775 (N_13775,N_13016,N_13127);
or U13776 (N_13776,N_13321,N_13412);
or U13777 (N_13777,N_13285,N_13219);
nor U13778 (N_13778,N_12914,N_13557);
nor U13779 (N_13779,N_13234,N_12993);
or U13780 (N_13780,N_12858,N_12956);
and U13781 (N_13781,N_13150,N_12919);
nor U13782 (N_13782,N_13159,N_13269);
nand U13783 (N_13783,N_13292,N_12820);
or U13784 (N_13784,N_12927,N_13437);
and U13785 (N_13785,N_13284,N_12990);
and U13786 (N_13786,N_13074,N_13478);
or U13787 (N_13787,N_13466,N_13186);
nor U13788 (N_13788,N_13109,N_13135);
and U13789 (N_13789,N_13428,N_13333);
or U13790 (N_13790,N_12952,N_13544);
and U13791 (N_13791,N_12870,N_12890);
or U13792 (N_13792,N_13134,N_12879);
or U13793 (N_13793,N_13330,N_13312);
nand U13794 (N_13794,N_12907,N_12857);
nand U13795 (N_13795,N_12942,N_12951);
or U13796 (N_13796,N_13543,N_13354);
or U13797 (N_13797,N_13332,N_13463);
nor U13798 (N_13798,N_13299,N_13479);
or U13799 (N_13799,N_13241,N_13578);
nand U13800 (N_13800,N_13464,N_13381);
and U13801 (N_13801,N_13264,N_13300);
nand U13802 (N_13802,N_12855,N_13532);
and U13803 (N_13803,N_13235,N_13270);
nand U13804 (N_13804,N_13453,N_13598);
nand U13805 (N_13805,N_13521,N_13052);
nor U13806 (N_13806,N_12877,N_13041);
xor U13807 (N_13807,N_12905,N_13427);
and U13808 (N_13808,N_12868,N_13418);
xor U13809 (N_13809,N_13442,N_13013);
xor U13810 (N_13810,N_13303,N_13076);
nor U13811 (N_13811,N_13484,N_12962);
and U13812 (N_13812,N_13067,N_13040);
xor U13813 (N_13813,N_13208,N_13460);
xnor U13814 (N_13814,N_13438,N_13202);
nor U13815 (N_13815,N_13440,N_13198);
nand U13816 (N_13816,N_13118,N_13290);
nand U13817 (N_13817,N_12953,N_13229);
nor U13818 (N_13818,N_13473,N_13405);
xnor U13819 (N_13819,N_13414,N_12909);
nand U13820 (N_13820,N_13422,N_13197);
and U13821 (N_13821,N_13457,N_12899);
or U13822 (N_13822,N_12960,N_13581);
xnor U13823 (N_13823,N_13167,N_13196);
nor U13824 (N_13824,N_13343,N_13173);
nand U13825 (N_13825,N_13373,N_13369);
or U13826 (N_13826,N_13376,N_13255);
or U13827 (N_13827,N_12964,N_13363);
xnor U13828 (N_13828,N_13256,N_13139);
nand U13829 (N_13829,N_12994,N_13289);
nand U13830 (N_13830,N_13589,N_13162);
and U13831 (N_13831,N_12958,N_13177);
xnor U13832 (N_13832,N_13166,N_13535);
or U13833 (N_13833,N_12882,N_13588);
xnor U13834 (N_13834,N_13341,N_12892);
nor U13835 (N_13835,N_13561,N_13372);
nand U13836 (N_13836,N_13531,N_12893);
and U13837 (N_13837,N_12970,N_13030);
xor U13838 (N_13838,N_13494,N_13207);
xnor U13839 (N_13839,N_12945,N_13353);
nor U13840 (N_13840,N_13168,N_12902);
nand U13841 (N_13841,N_12804,N_12997);
and U13842 (N_13842,N_13429,N_12928);
or U13843 (N_13843,N_13592,N_13169);
xnor U13844 (N_13844,N_13024,N_13214);
and U13845 (N_13845,N_13425,N_13399);
or U13846 (N_13846,N_13089,N_12959);
or U13847 (N_13847,N_13443,N_13298);
nor U13848 (N_13848,N_13570,N_13271);
and U13849 (N_13849,N_13495,N_13059);
nor U13850 (N_13850,N_13025,N_13375);
or U13851 (N_13851,N_13023,N_13115);
xnor U13852 (N_13852,N_13242,N_13027);
nor U13853 (N_13853,N_13568,N_13105);
nand U13854 (N_13854,N_13103,N_13174);
nor U13855 (N_13855,N_13482,N_12859);
xnor U13856 (N_13856,N_13361,N_13192);
and U13857 (N_13857,N_13378,N_13459);
xor U13858 (N_13858,N_13213,N_13232);
or U13859 (N_13859,N_13519,N_13594);
and U13860 (N_13860,N_13066,N_13144);
nor U13861 (N_13861,N_13295,N_12963);
xnor U13862 (N_13862,N_13204,N_13315);
nand U13863 (N_13863,N_12849,N_13179);
and U13864 (N_13864,N_13500,N_13102);
nand U13865 (N_13865,N_12895,N_13409);
nand U13866 (N_13866,N_13158,N_13110);
xor U13867 (N_13867,N_13121,N_13217);
or U13868 (N_13868,N_12852,N_13558);
and U13869 (N_13869,N_13216,N_13515);
or U13870 (N_13870,N_13338,N_13317);
and U13871 (N_13871,N_12897,N_13233);
nor U13872 (N_13872,N_13157,N_13441);
xnor U13873 (N_13873,N_12974,N_13266);
and U13874 (N_13874,N_13193,N_13078);
xor U13875 (N_13875,N_12911,N_12886);
or U13876 (N_13876,N_13563,N_13185);
nand U13877 (N_13877,N_13337,N_13161);
xor U13878 (N_13878,N_13018,N_13374);
and U13879 (N_13879,N_12924,N_12846);
and U13880 (N_13880,N_13101,N_13518);
nand U13881 (N_13881,N_13569,N_13277);
nor U13882 (N_13882,N_13344,N_13536);
nor U13883 (N_13883,N_13205,N_13496);
nor U13884 (N_13884,N_13571,N_13093);
nand U13885 (N_13885,N_12929,N_13239);
or U13886 (N_13886,N_13021,N_13560);
xor U13887 (N_13887,N_13541,N_13498);
nand U13888 (N_13888,N_12833,N_13347);
nand U13889 (N_13889,N_13320,N_12941);
or U13890 (N_13890,N_13318,N_13545);
nor U13891 (N_13891,N_13587,N_13240);
and U13892 (N_13892,N_12917,N_13286);
xnor U13893 (N_13893,N_12976,N_12860);
or U13894 (N_13894,N_12940,N_12862);
and U13895 (N_13895,N_12814,N_13231);
nand U13896 (N_13896,N_13082,N_13274);
nand U13897 (N_13897,N_13465,N_13098);
nand U13898 (N_13898,N_13301,N_13293);
xor U13899 (N_13899,N_12935,N_13502);
and U13900 (N_13900,N_13141,N_13501);
and U13901 (N_13901,N_13083,N_13489);
or U13902 (N_13902,N_13019,N_12908);
xnor U13903 (N_13903,N_13075,N_13009);
xnor U13904 (N_13904,N_12801,N_13507);
nand U13905 (N_13905,N_13267,N_13252);
xor U13906 (N_13906,N_13579,N_13151);
nor U13907 (N_13907,N_13574,N_13104);
or U13908 (N_13908,N_12923,N_13039);
xor U13909 (N_13909,N_13590,N_12900);
nand U13910 (N_13910,N_12979,N_12966);
nor U13911 (N_13911,N_13002,N_12818);
and U13912 (N_13912,N_13410,N_13247);
and U13913 (N_13913,N_13136,N_12938);
or U13914 (N_13914,N_13475,N_13451);
xor U13915 (N_13915,N_13084,N_13470);
xnor U13916 (N_13916,N_13477,N_13015);
or U13917 (N_13917,N_13524,N_13060);
nor U13918 (N_13918,N_13043,N_13042);
and U13919 (N_13919,N_13125,N_13065);
xnor U13920 (N_13920,N_13357,N_12828);
xor U13921 (N_13921,N_13585,N_13114);
nor U13922 (N_13922,N_12915,N_13190);
nor U13923 (N_13923,N_12884,N_13486);
and U13924 (N_13924,N_12943,N_13403);
and U13925 (N_13925,N_13062,N_13379);
and U13926 (N_13926,N_13014,N_13222);
nand U13927 (N_13927,N_13445,N_12916);
or U13928 (N_13928,N_13251,N_13090);
xnor U13929 (N_13929,N_13584,N_13051);
nor U13930 (N_13930,N_13525,N_13056);
and U13931 (N_13931,N_13096,N_13573);
and U13932 (N_13932,N_12838,N_13336);
nand U13933 (N_13933,N_13547,N_13113);
nand U13934 (N_13934,N_13172,N_13526);
nand U13935 (N_13935,N_13358,N_13071);
nand U13936 (N_13936,N_13472,N_12896);
and U13937 (N_13937,N_12920,N_12894);
and U13938 (N_13938,N_13085,N_12950);
xnor U13939 (N_13939,N_12800,N_12831);
and U13940 (N_13940,N_13450,N_13263);
and U13941 (N_13941,N_13488,N_13396);
and U13942 (N_13942,N_13346,N_12975);
nor U13943 (N_13943,N_13164,N_12843);
nor U13944 (N_13944,N_13468,N_12967);
nand U13945 (N_13945,N_13419,N_13143);
or U13946 (N_13946,N_13339,N_13230);
and U13947 (N_13947,N_13154,N_12866);
xnor U13948 (N_13948,N_12809,N_13064);
and U13949 (N_13949,N_12847,N_13261);
and U13950 (N_13950,N_13364,N_13553);
and U13951 (N_13951,N_13391,N_13397);
and U13952 (N_13952,N_13224,N_13008);
or U13953 (N_13953,N_13155,N_13138);
and U13954 (N_13954,N_13534,N_12987);
or U13955 (N_13955,N_13551,N_13086);
and U13956 (N_13956,N_13297,N_13209);
xor U13957 (N_13957,N_13366,N_13593);
and U13958 (N_13958,N_12948,N_13348);
and U13959 (N_13959,N_13073,N_13431);
xor U13960 (N_13960,N_13091,N_13017);
or U13961 (N_13961,N_13309,N_13452);
nor U13962 (N_13962,N_12906,N_13187);
xnor U13963 (N_13963,N_13100,N_13258);
or U13964 (N_13964,N_13058,N_12955);
and U13965 (N_13965,N_13402,N_12973);
and U13966 (N_13966,N_13487,N_13145);
and U13967 (N_13967,N_13107,N_13028);
xor U13968 (N_13968,N_13215,N_13461);
nand U13969 (N_13969,N_12903,N_12944);
or U13970 (N_13970,N_13011,N_12872);
nor U13971 (N_13971,N_13004,N_13349);
and U13972 (N_13972,N_13088,N_12961);
or U13973 (N_13973,N_12829,N_13567);
xor U13974 (N_13974,N_13319,N_12845);
xor U13975 (N_13975,N_13383,N_13350);
and U13976 (N_13976,N_13146,N_13288);
and U13977 (N_13977,N_12931,N_13007);
xor U13978 (N_13978,N_12933,N_12887);
nand U13979 (N_13979,N_13331,N_12842);
nand U13980 (N_13980,N_13390,N_13126);
nor U13981 (N_13981,N_13413,N_13540);
nand U13982 (N_13982,N_13035,N_13556);
xor U13983 (N_13983,N_12837,N_13326);
nand U13984 (N_13984,N_12880,N_13328);
nor U13985 (N_13985,N_13152,N_13384);
and U13986 (N_13986,N_13474,N_12816);
or U13987 (N_13987,N_13432,N_13423);
xnor U13988 (N_13988,N_12822,N_13032);
nor U13989 (N_13989,N_13036,N_12913);
or U13990 (N_13990,N_13490,N_13170);
or U13991 (N_13991,N_13365,N_13444);
or U13992 (N_13992,N_13005,N_13248);
nand U13993 (N_13993,N_13165,N_13280);
nor U13994 (N_13994,N_13456,N_12834);
nor U13995 (N_13995,N_13327,N_13181);
nor U13996 (N_13996,N_13156,N_13243);
or U13997 (N_13997,N_13022,N_12949);
xor U13998 (N_13998,N_12889,N_13188);
and U13999 (N_13999,N_13095,N_12999);
xor U14000 (N_14000,N_13495,N_13448);
nor U14001 (N_14001,N_13400,N_12962);
nor U14002 (N_14002,N_13063,N_13556);
nor U14003 (N_14003,N_13550,N_12815);
xor U14004 (N_14004,N_13515,N_13598);
nand U14005 (N_14005,N_13438,N_12865);
nand U14006 (N_14006,N_13019,N_13429);
nand U14007 (N_14007,N_13513,N_13301);
or U14008 (N_14008,N_13147,N_13138);
nand U14009 (N_14009,N_13070,N_13590);
or U14010 (N_14010,N_12874,N_12922);
xor U14011 (N_14011,N_13234,N_13013);
xor U14012 (N_14012,N_13367,N_12917);
and U14013 (N_14013,N_12846,N_13171);
or U14014 (N_14014,N_12902,N_13281);
and U14015 (N_14015,N_13345,N_13035);
nor U14016 (N_14016,N_13420,N_13035);
xor U14017 (N_14017,N_13019,N_12900);
and U14018 (N_14018,N_12887,N_13523);
nand U14019 (N_14019,N_12923,N_13179);
nor U14020 (N_14020,N_13392,N_13440);
or U14021 (N_14021,N_12831,N_13473);
nor U14022 (N_14022,N_13548,N_12984);
or U14023 (N_14023,N_13098,N_13410);
nor U14024 (N_14024,N_13345,N_12840);
nor U14025 (N_14025,N_13545,N_13353);
nand U14026 (N_14026,N_13517,N_13238);
nand U14027 (N_14027,N_13510,N_12970);
or U14028 (N_14028,N_13446,N_12983);
and U14029 (N_14029,N_13576,N_13249);
and U14030 (N_14030,N_13533,N_13356);
xnor U14031 (N_14031,N_13304,N_13257);
nand U14032 (N_14032,N_12934,N_13103);
and U14033 (N_14033,N_12817,N_13057);
xor U14034 (N_14034,N_13260,N_13148);
nor U14035 (N_14035,N_13448,N_13541);
or U14036 (N_14036,N_13097,N_12967);
nand U14037 (N_14037,N_13270,N_12921);
and U14038 (N_14038,N_13272,N_13182);
or U14039 (N_14039,N_13016,N_13042);
and U14040 (N_14040,N_12938,N_12957);
or U14041 (N_14041,N_12977,N_13578);
and U14042 (N_14042,N_12854,N_13497);
and U14043 (N_14043,N_13386,N_13012);
nor U14044 (N_14044,N_13303,N_13097);
nor U14045 (N_14045,N_13090,N_13195);
or U14046 (N_14046,N_12903,N_12929);
and U14047 (N_14047,N_13180,N_13112);
or U14048 (N_14048,N_13350,N_13541);
xor U14049 (N_14049,N_13538,N_13596);
and U14050 (N_14050,N_13116,N_13574);
xnor U14051 (N_14051,N_13297,N_13414);
and U14052 (N_14052,N_12978,N_12927);
xnor U14053 (N_14053,N_13095,N_12983);
nand U14054 (N_14054,N_13114,N_12870);
nor U14055 (N_14055,N_12816,N_13248);
and U14056 (N_14056,N_13240,N_13287);
or U14057 (N_14057,N_13036,N_12954);
and U14058 (N_14058,N_13331,N_12815);
nand U14059 (N_14059,N_13519,N_12891);
xnor U14060 (N_14060,N_13123,N_13032);
and U14061 (N_14061,N_13082,N_13581);
nand U14062 (N_14062,N_13118,N_13230);
nor U14063 (N_14063,N_13055,N_13502);
xor U14064 (N_14064,N_12887,N_12941);
xor U14065 (N_14065,N_13372,N_13029);
or U14066 (N_14066,N_13430,N_13012);
xor U14067 (N_14067,N_12982,N_13117);
and U14068 (N_14068,N_12830,N_12810);
nor U14069 (N_14069,N_13390,N_13428);
or U14070 (N_14070,N_13012,N_12925);
and U14071 (N_14071,N_13389,N_13068);
nand U14072 (N_14072,N_13058,N_13490);
nand U14073 (N_14073,N_13010,N_13279);
xnor U14074 (N_14074,N_13228,N_12970);
nor U14075 (N_14075,N_13208,N_13173);
xnor U14076 (N_14076,N_12826,N_13135);
or U14077 (N_14077,N_13085,N_13136);
or U14078 (N_14078,N_13088,N_13538);
xnor U14079 (N_14079,N_13403,N_13110);
and U14080 (N_14080,N_13561,N_12920);
and U14081 (N_14081,N_12963,N_13212);
xor U14082 (N_14082,N_13513,N_12801);
or U14083 (N_14083,N_13333,N_13309);
xnor U14084 (N_14084,N_13456,N_13511);
xnor U14085 (N_14085,N_13544,N_13584);
xor U14086 (N_14086,N_13547,N_12957);
nor U14087 (N_14087,N_13167,N_12958);
or U14088 (N_14088,N_13134,N_13294);
and U14089 (N_14089,N_13091,N_13282);
or U14090 (N_14090,N_13307,N_12914);
nand U14091 (N_14091,N_12849,N_13080);
nand U14092 (N_14092,N_13588,N_13503);
nor U14093 (N_14093,N_13427,N_13416);
nand U14094 (N_14094,N_12992,N_13398);
nor U14095 (N_14095,N_13354,N_13189);
nand U14096 (N_14096,N_13006,N_13061);
and U14097 (N_14097,N_13299,N_12847);
nor U14098 (N_14098,N_13104,N_13477);
xor U14099 (N_14099,N_12865,N_12928);
xor U14100 (N_14100,N_13282,N_13332);
nand U14101 (N_14101,N_13213,N_13342);
xor U14102 (N_14102,N_13041,N_13112);
or U14103 (N_14103,N_13125,N_13329);
xnor U14104 (N_14104,N_13011,N_13551);
or U14105 (N_14105,N_13325,N_13504);
and U14106 (N_14106,N_12877,N_13266);
nor U14107 (N_14107,N_12845,N_13588);
or U14108 (N_14108,N_13500,N_13019);
xor U14109 (N_14109,N_13542,N_12942);
or U14110 (N_14110,N_13201,N_12879);
or U14111 (N_14111,N_12853,N_13569);
nand U14112 (N_14112,N_13149,N_13289);
and U14113 (N_14113,N_13521,N_13407);
nor U14114 (N_14114,N_13175,N_13173);
or U14115 (N_14115,N_12895,N_12898);
nor U14116 (N_14116,N_12865,N_12827);
nand U14117 (N_14117,N_12853,N_13033);
nand U14118 (N_14118,N_12883,N_13485);
xor U14119 (N_14119,N_12837,N_13083);
nand U14120 (N_14120,N_13519,N_13288);
or U14121 (N_14121,N_12818,N_13534);
xnor U14122 (N_14122,N_13494,N_13060);
xor U14123 (N_14123,N_13394,N_12850);
xor U14124 (N_14124,N_12923,N_13563);
xnor U14125 (N_14125,N_13334,N_12820);
nor U14126 (N_14126,N_12881,N_13347);
or U14127 (N_14127,N_13054,N_12905);
or U14128 (N_14128,N_13102,N_12952);
nand U14129 (N_14129,N_12855,N_13231);
nand U14130 (N_14130,N_13356,N_13060);
nor U14131 (N_14131,N_13017,N_13368);
xnor U14132 (N_14132,N_12844,N_13067);
xor U14133 (N_14133,N_12932,N_13044);
xor U14134 (N_14134,N_13325,N_13505);
or U14135 (N_14135,N_13443,N_13472);
or U14136 (N_14136,N_12890,N_13123);
and U14137 (N_14137,N_12970,N_12861);
and U14138 (N_14138,N_12895,N_12994);
nand U14139 (N_14139,N_13064,N_13498);
nor U14140 (N_14140,N_13568,N_13049);
or U14141 (N_14141,N_13346,N_13199);
nand U14142 (N_14142,N_13048,N_13159);
nand U14143 (N_14143,N_13424,N_13105);
and U14144 (N_14144,N_13369,N_13442);
nor U14145 (N_14145,N_13251,N_13555);
nand U14146 (N_14146,N_13189,N_13371);
and U14147 (N_14147,N_13197,N_13346);
and U14148 (N_14148,N_13078,N_13337);
nor U14149 (N_14149,N_13308,N_13376);
and U14150 (N_14150,N_13125,N_12849);
nand U14151 (N_14151,N_13068,N_13172);
or U14152 (N_14152,N_13190,N_13493);
nand U14153 (N_14153,N_13093,N_13389);
and U14154 (N_14154,N_13000,N_13581);
nor U14155 (N_14155,N_12957,N_13026);
or U14156 (N_14156,N_13348,N_13068);
nand U14157 (N_14157,N_13120,N_13562);
xnor U14158 (N_14158,N_13361,N_13041);
xnor U14159 (N_14159,N_13023,N_13139);
nor U14160 (N_14160,N_13372,N_13348);
and U14161 (N_14161,N_13306,N_13437);
and U14162 (N_14162,N_13202,N_13087);
and U14163 (N_14163,N_13037,N_13503);
nor U14164 (N_14164,N_13182,N_13090);
nand U14165 (N_14165,N_12860,N_12843);
or U14166 (N_14166,N_13346,N_13116);
nor U14167 (N_14167,N_13144,N_13535);
nand U14168 (N_14168,N_13578,N_13478);
or U14169 (N_14169,N_12954,N_12986);
xnor U14170 (N_14170,N_13235,N_13378);
or U14171 (N_14171,N_13090,N_13073);
and U14172 (N_14172,N_12963,N_13147);
xnor U14173 (N_14173,N_12960,N_13251);
nand U14174 (N_14174,N_13164,N_13381);
xor U14175 (N_14175,N_13521,N_12868);
and U14176 (N_14176,N_12969,N_12816);
nand U14177 (N_14177,N_12829,N_12868);
and U14178 (N_14178,N_12973,N_13584);
and U14179 (N_14179,N_13595,N_13088);
nor U14180 (N_14180,N_12847,N_13281);
or U14181 (N_14181,N_13476,N_13336);
and U14182 (N_14182,N_13475,N_13213);
xnor U14183 (N_14183,N_13265,N_13070);
xor U14184 (N_14184,N_13467,N_13395);
nor U14185 (N_14185,N_12962,N_13493);
nand U14186 (N_14186,N_13470,N_13124);
and U14187 (N_14187,N_12984,N_12916);
nor U14188 (N_14188,N_13046,N_13526);
or U14189 (N_14189,N_13253,N_13413);
nand U14190 (N_14190,N_13102,N_13465);
nand U14191 (N_14191,N_13026,N_13176);
or U14192 (N_14192,N_12873,N_13444);
and U14193 (N_14193,N_13389,N_13308);
and U14194 (N_14194,N_12971,N_13172);
xor U14195 (N_14195,N_13095,N_13449);
nor U14196 (N_14196,N_12851,N_13109);
nand U14197 (N_14197,N_13079,N_13019);
nand U14198 (N_14198,N_13179,N_13580);
nand U14199 (N_14199,N_13087,N_12960);
nor U14200 (N_14200,N_12821,N_13279);
and U14201 (N_14201,N_13053,N_13158);
and U14202 (N_14202,N_13043,N_12857);
nand U14203 (N_14203,N_13498,N_12947);
and U14204 (N_14204,N_13353,N_12967);
xor U14205 (N_14205,N_13516,N_12980);
or U14206 (N_14206,N_13547,N_13157);
and U14207 (N_14207,N_12942,N_13129);
nor U14208 (N_14208,N_13128,N_13372);
and U14209 (N_14209,N_13221,N_13500);
and U14210 (N_14210,N_13138,N_13353);
or U14211 (N_14211,N_12923,N_13154);
xnor U14212 (N_14212,N_13168,N_13158);
nand U14213 (N_14213,N_12854,N_13463);
xor U14214 (N_14214,N_13276,N_12971);
nand U14215 (N_14215,N_12829,N_13012);
or U14216 (N_14216,N_13163,N_13247);
or U14217 (N_14217,N_13549,N_13552);
and U14218 (N_14218,N_13446,N_13248);
nor U14219 (N_14219,N_13526,N_13164);
nand U14220 (N_14220,N_13345,N_13445);
or U14221 (N_14221,N_13352,N_13242);
xnor U14222 (N_14222,N_13241,N_12957);
or U14223 (N_14223,N_13453,N_13493);
nand U14224 (N_14224,N_12831,N_13042);
nor U14225 (N_14225,N_13084,N_13403);
xnor U14226 (N_14226,N_13222,N_13426);
and U14227 (N_14227,N_13497,N_13333);
nor U14228 (N_14228,N_13369,N_13339);
nand U14229 (N_14229,N_13001,N_13322);
and U14230 (N_14230,N_13014,N_12974);
xor U14231 (N_14231,N_13455,N_12919);
or U14232 (N_14232,N_13005,N_13386);
and U14233 (N_14233,N_12801,N_12899);
nor U14234 (N_14234,N_13034,N_12948);
and U14235 (N_14235,N_13313,N_13479);
and U14236 (N_14236,N_13066,N_13342);
nand U14237 (N_14237,N_13027,N_12855);
xnor U14238 (N_14238,N_13076,N_12839);
and U14239 (N_14239,N_13363,N_13462);
nor U14240 (N_14240,N_13300,N_12831);
or U14241 (N_14241,N_13327,N_12981);
or U14242 (N_14242,N_13149,N_12971);
and U14243 (N_14243,N_13529,N_12995);
xnor U14244 (N_14244,N_13123,N_12938);
nand U14245 (N_14245,N_13399,N_13046);
or U14246 (N_14246,N_13119,N_12832);
nor U14247 (N_14247,N_13492,N_12812);
nor U14248 (N_14248,N_13508,N_12859);
nand U14249 (N_14249,N_13228,N_12956);
nand U14250 (N_14250,N_13043,N_13511);
nor U14251 (N_14251,N_13570,N_13462);
nor U14252 (N_14252,N_12847,N_12895);
and U14253 (N_14253,N_13406,N_12859);
xor U14254 (N_14254,N_12872,N_13017);
xor U14255 (N_14255,N_13041,N_13271);
xor U14256 (N_14256,N_12856,N_13513);
or U14257 (N_14257,N_13108,N_13094);
nor U14258 (N_14258,N_13187,N_13552);
nor U14259 (N_14259,N_12915,N_12850);
nand U14260 (N_14260,N_12892,N_13536);
xor U14261 (N_14261,N_12982,N_13525);
and U14262 (N_14262,N_13050,N_13290);
nor U14263 (N_14263,N_13034,N_13356);
or U14264 (N_14264,N_13320,N_13597);
or U14265 (N_14265,N_12930,N_12841);
or U14266 (N_14266,N_13058,N_13471);
nand U14267 (N_14267,N_13185,N_12927);
xor U14268 (N_14268,N_13538,N_13576);
and U14269 (N_14269,N_13556,N_13061);
xor U14270 (N_14270,N_13500,N_13264);
and U14271 (N_14271,N_12810,N_13288);
and U14272 (N_14272,N_13349,N_13453);
nor U14273 (N_14273,N_13516,N_13038);
nor U14274 (N_14274,N_12874,N_12945);
or U14275 (N_14275,N_13262,N_13047);
and U14276 (N_14276,N_13164,N_13537);
nand U14277 (N_14277,N_13128,N_12931);
nand U14278 (N_14278,N_12883,N_13197);
xnor U14279 (N_14279,N_13400,N_13170);
nand U14280 (N_14280,N_13228,N_13444);
xnor U14281 (N_14281,N_13217,N_13231);
nor U14282 (N_14282,N_12890,N_12982);
and U14283 (N_14283,N_13475,N_13365);
or U14284 (N_14284,N_13540,N_13171);
xnor U14285 (N_14285,N_12931,N_13570);
or U14286 (N_14286,N_12814,N_13208);
xor U14287 (N_14287,N_13005,N_13160);
or U14288 (N_14288,N_13060,N_13192);
nand U14289 (N_14289,N_13563,N_13414);
xor U14290 (N_14290,N_13265,N_13326);
and U14291 (N_14291,N_13364,N_13128);
nand U14292 (N_14292,N_13121,N_13027);
nor U14293 (N_14293,N_13067,N_12986);
and U14294 (N_14294,N_13545,N_13524);
nor U14295 (N_14295,N_13311,N_12984);
xnor U14296 (N_14296,N_13473,N_13384);
and U14297 (N_14297,N_13137,N_13262);
or U14298 (N_14298,N_13094,N_13420);
or U14299 (N_14299,N_13203,N_12871);
nor U14300 (N_14300,N_12921,N_12940);
nor U14301 (N_14301,N_13136,N_13270);
xor U14302 (N_14302,N_12810,N_13418);
nand U14303 (N_14303,N_13513,N_13596);
xor U14304 (N_14304,N_13050,N_13143);
xnor U14305 (N_14305,N_13507,N_12825);
nand U14306 (N_14306,N_13352,N_13132);
nand U14307 (N_14307,N_13527,N_13287);
xor U14308 (N_14308,N_13578,N_13098);
and U14309 (N_14309,N_13410,N_12950);
nand U14310 (N_14310,N_13290,N_13115);
or U14311 (N_14311,N_13360,N_13146);
nand U14312 (N_14312,N_13290,N_13447);
nor U14313 (N_14313,N_12973,N_12933);
nor U14314 (N_14314,N_13585,N_13253);
nand U14315 (N_14315,N_13332,N_12848);
xnor U14316 (N_14316,N_12927,N_12901);
xnor U14317 (N_14317,N_12867,N_13183);
and U14318 (N_14318,N_13040,N_12933);
nor U14319 (N_14319,N_12978,N_12996);
xnor U14320 (N_14320,N_12857,N_13444);
nor U14321 (N_14321,N_13438,N_13571);
nand U14322 (N_14322,N_12863,N_13455);
and U14323 (N_14323,N_13352,N_13267);
and U14324 (N_14324,N_13092,N_12915);
or U14325 (N_14325,N_13475,N_13427);
nand U14326 (N_14326,N_13579,N_13306);
nand U14327 (N_14327,N_13318,N_13373);
nand U14328 (N_14328,N_13145,N_12924);
nor U14329 (N_14329,N_13531,N_13156);
and U14330 (N_14330,N_13013,N_13575);
xnor U14331 (N_14331,N_13315,N_13376);
and U14332 (N_14332,N_13497,N_13437);
nor U14333 (N_14333,N_13012,N_13218);
and U14334 (N_14334,N_13557,N_12908);
xor U14335 (N_14335,N_13032,N_13356);
xor U14336 (N_14336,N_13243,N_12878);
nand U14337 (N_14337,N_13115,N_13080);
and U14338 (N_14338,N_13464,N_13156);
xnor U14339 (N_14339,N_13052,N_12979);
or U14340 (N_14340,N_12818,N_13306);
nor U14341 (N_14341,N_13534,N_13284);
nand U14342 (N_14342,N_12896,N_12834);
or U14343 (N_14343,N_12825,N_13016);
xor U14344 (N_14344,N_13441,N_13351);
nand U14345 (N_14345,N_13409,N_12851);
xor U14346 (N_14346,N_13599,N_12924);
nand U14347 (N_14347,N_13160,N_13228);
and U14348 (N_14348,N_13111,N_13206);
and U14349 (N_14349,N_13247,N_13115);
xnor U14350 (N_14350,N_13041,N_12844);
and U14351 (N_14351,N_13197,N_13149);
nand U14352 (N_14352,N_13122,N_13185);
nand U14353 (N_14353,N_13391,N_13243);
nand U14354 (N_14354,N_12823,N_12934);
nand U14355 (N_14355,N_13489,N_13418);
nand U14356 (N_14356,N_13329,N_13450);
xor U14357 (N_14357,N_13472,N_13263);
or U14358 (N_14358,N_12836,N_12938);
nand U14359 (N_14359,N_12842,N_13162);
or U14360 (N_14360,N_13503,N_13017);
nor U14361 (N_14361,N_12937,N_12936);
or U14362 (N_14362,N_12949,N_13482);
xnor U14363 (N_14363,N_12983,N_13197);
and U14364 (N_14364,N_13116,N_12977);
and U14365 (N_14365,N_13565,N_13556);
and U14366 (N_14366,N_12842,N_13497);
xnor U14367 (N_14367,N_12976,N_12967);
nor U14368 (N_14368,N_13140,N_12922);
nand U14369 (N_14369,N_12939,N_13318);
or U14370 (N_14370,N_13122,N_12917);
nand U14371 (N_14371,N_12986,N_12848);
nand U14372 (N_14372,N_12904,N_12915);
and U14373 (N_14373,N_13352,N_13193);
or U14374 (N_14374,N_13538,N_13054);
nor U14375 (N_14375,N_13333,N_13118);
or U14376 (N_14376,N_13496,N_13018);
nand U14377 (N_14377,N_13565,N_13245);
and U14378 (N_14378,N_13427,N_12947);
or U14379 (N_14379,N_13098,N_13012);
or U14380 (N_14380,N_13102,N_13248);
xor U14381 (N_14381,N_13504,N_12902);
and U14382 (N_14382,N_13197,N_13122);
nand U14383 (N_14383,N_13585,N_13279);
nor U14384 (N_14384,N_13407,N_13396);
nand U14385 (N_14385,N_13105,N_12859);
or U14386 (N_14386,N_13592,N_12882);
nor U14387 (N_14387,N_13235,N_13598);
nand U14388 (N_14388,N_13387,N_13473);
xor U14389 (N_14389,N_13590,N_12915);
xor U14390 (N_14390,N_13246,N_13300);
and U14391 (N_14391,N_13384,N_13439);
and U14392 (N_14392,N_12945,N_12950);
and U14393 (N_14393,N_13403,N_13044);
nor U14394 (N_14394,N_13140,N_13266);
nor U14395 (N_14395,N_13117,N_12959);
nand U14396 (N_14396,N_13484,N_12808);
xor U14397 (N_14397,N_13513,N_13016);
or U14398 (N_14398,N_13046,N_12846);
nand U14399 (N_14399,N_13350,N_12851);
or U14400 (N_14400,N_14017,N_14398);
or U14401 (N_14401,N_14271,N_14021);
or U14402 (N_14402,N_14259,N_13813);
xor U14403 (N_14403,N_14365,N_13919);
nand U14404 (N_14404,N_14393,N_13737);
or U14405 (N_14405,N_14343,N_13778);
nor U14406 (N_14406,N_14205,N_13655);
and U14407 (N_14407,N_13618,N_13612);
nor U14408 (N_14408,N_13985,N_13939);
xnor U14409 (N_14409,N_14008,N_13722);
nand U14410 (N_14410,N_14378,N_14221);
xnor U14411 (N_14411,N_13614,N_13971);
nor U14412 (N_14412,N_13706,N_14219);
and U14413 (N_14413,N_14064,N_13607);
nand U14414 (N_14414,N_14048,N_13780);
or U14415 (N_14415,N_13853,N_13872);
nand U14416 (N_14416,N_14287,N_14023);
or U14417 (N_14417,N_13633,N_13981);
xor U14418 (N_14418,N_13752,N_13852);
xor U14419 (N_14419,N_13608,N_13837);
or U14420 (N_14420,N_14012,N_14309);
nand U14421 (N_14421,N_13673,N_13721);
and U14422 (N_14422,N_14199,N_13745);
and U14423 (N_14423,N_14188,N_13874);
xnor U14424 (N_14424,N_14191,N_14030);
or U14425 (N_14425,N_14097,N_13738);
and U14426 (N_14426,N_13811,N_14034);
nand U14427 (N_14427,N_13651,N_13848);
xor U14428 (N_14428,N_13807,N_13905);
or U14429 (N_14429,N_13687,N_13834);
or U14430 (N_14430,N_13949,N_14356);
or U14431 (N_14431,N_13674,N_14290);
or U14432 (N_14432,N_13683,N_14032);
or U14433 (N_14433,N_13652,N_14068);
and U14434 (N_14434,N_13767,N_14374);
and U14435 (N_14435,N_13793,N_13820);
and U14436 (N_14436,N_13978,N_13856);
xnor U14437 (N_14437,N_14136,N_13615);
or U14438 (N_14438,N_14235,N_14078);
xnor U14439 (N_14439,N_13804,N_13634);
or U14440 (N_14440,N_13987,N_14169);
xor U14441 (N_14441,N_14013,N_13774);
and U14442 (N_14442,N_14019,N_13705);
nor U14443 (N_14443,N_13649,N_13851);
or U14444 (N_14444,N_13864,N_13660);
or U14445 (N_14445,N_13876,N_13995);
nor U14446 (N_14446,N_13912,N_13697);
and U14447 (N_14447,N_13845,N_13766);
or U14448 (N_14448,N_13830,N_14260);
and U14449 (N_14449,N_13894,N_14011);
or U14450 (N_14450,N_14211,N_14389);
xnor U14451 (N_14451,N_14330,N_14256);
xor U14452 (N_14452,N_14142,N_14088);
or U14453 (N_14453,N_14296,N_14237);
xor U14454 (N_14454,N_13688,N_14214);
nor U14455 (N_14455,N_13938,N_13935);
xor U14456 (N_14456,N_13893,N_13801);
nand U14457 (N_14457,N_13784,N_14137);
or U14458 (N_14458,N_13960,N_13689);
nor U14459 (N_14459,N_14104,N_13986);
nand U14460 (N_14460,N_14186,N_13887);
and U14461 (N_14461,N_14195,N_13881);
xnor U14462 (N_14462,N_14268,N_14046);
and U14463 (N_14463,N_14129,N_14122);
xor U14464 (N_14464,N_14361,N_13694);
nor U14465 (N_14465,N_14298,N_13976);
nand U14466 (N_14466,N_14266,N_14117);
and U14467 (N_14467,N_14248,N_13730);
or U14468 (N_14468,N_13891,N_13998);
nand U14469 (N_14469,N_13809,N_13913);
or U14470 (N_14470,N_13901,N_14255);
nand U14471 (N_14471,N_13825,N_13627);
and U14472 (N_14472,N_13942,N_13654);
xor U14473 (N_14473,N_13923,N_14141);
nor U14474 (N_14474,N_13719,N_14193);
xnor U14475 (N_14475,N_13950,N_14348);
nand U14476 (N_14476,N_14166,N_13656);
xnor U14477 (N_14477,N_14293,N_13924);
or U14478 (N_14478,N_14077,N_14208);
or U14479 (N_14479,N_13623,N_14106);
xnor U14480 (N_14480,N_13857,N_14110);
nand U14481 (N_14481,N_14331,N_13645);
and U14482 (N_14482,N_14156,N_14158);
nand U14483 (N_14483,N_13729,N_13639);
xor U14484 (N_14484,N_13782,N_14038);
xnor U14485 (N_14485,N_14375,N_14070);
or U14486 (N_14486,N_13962,N_14215);
nor U14487 (N_14487,N_13812,N_13704);
xnor U14488 (N_14488,N_13658,N_13613);
and U14489 (N_14489,N_13797,N_14212);
or U14490 (N_14490,N_13882,N_13828);
xnor U14491 (N_14491,N_14316,N_13750);
nand U14492 (N_14492,N_13790,N_13824);
xnor U14493 (N_14493,N_14347,N_14171);
and U14494 (N_14494,N_14152,N_14052);
nor U14495 (N_14495,N_13833,N_13988);
and U14496 (N_14496,N_14140,N_13967);
nor U14497 (N_14497,N_14261,N_13779);
xnor U14498 (N_14498,N_13787,N_14100);
and U14499 (N_14499,N_13999,N_14204);
or U14500 (N_14500,N_13647,N_14194);
and U14501 (N_14501,N_13764,N_14089);
xor U14502 (N_14502,N_13865,N_13631);
and U14503 (N_14503,N_13823,N_14105);
nor U14504 (N_14504,N_13661,N_14118);
and U14505 (N_14505,N_13819,N_13756);
nor U14506 (N_14506,N_14396,N_13928);
nor U14507 (N_14507,N_13948,N_13895);
nand U14508 (N_14508,N_13871,N_14377);
nor U14509 (N_14509,N_14123,N_13943);
nor U14510 (N_14510,N_13711,N_13922);
or U14511 (N_14511,N_14138,N_14222);
xnor U14512 (N_14512,N_14345,N_13696);
or U14513 (N_14513,N_13671,N_14190);
or U14514 (N_14514,N_14380,N_13902);
nand U14515 (N_14515,N_14056,N_13684);
nor U14516 (N_14516,N_14210,N_13690);
and U14517 (N_14517,N_13692,N_13907);
xor U14518 (N_14518,N_13878,N_14133);
nor U14519 (N_14519,N_13936,N_13873);
nor U14520 (N_14520,N_13941,N_14251);
and U14521 (N_14521,N_14167,N_14341);
nand U14522 (N_14522,N_13736,N_14144);
or U14523 (N_14523,N_14311,N_14340);
nor U14524 (N_14524,N_13831,N_13972);
xor U14525 (N_14525,N_13786,N_13979);
or U14526 (N_14526,N_14326,N_14111);
nor U14527 (N_14527,N_14279,N_13817);
and U14528 (N_14528,N_14099,N_14312);
nand U14529 (N_14529,N_13897,N_14310);
nor U14530 (N_14530,N_13744,N_13751);
nand U14531 (N_14531,N_13847,N_13947);
nand U14532 (N_14532,N_13632,N_14264);
or U14533 (N_14533,N_14177,N_14130);
or U14534 (N_14534,N_14163,N_14346);
xnor U14535 (N_14535,N_14172,N_13885);
or U14536 (N_14536,N_14007,N_14323);
and U14537 (N_14537,N_14024,N_13727);
or U14538 (N_14538,N_13970,N_13753);
nor U14539 (N_14539,N_14390,N_14004);
and U14540 (N_14540,N_13803,N_14357);
or U14541 (N_14541,N_14228,N_13641);
or U14542 (N_14542,N_13934,N_14081);
nand U14543 (N_14543,N_13760,N_13701);
nor U14544 (N_14544,N_14209,N_13716);
xnor U14545 (N_14545,N_13642,N_13796);
xnor U14546 (N_14546,N_13965,N_14155);
nand U14547 (N_14547,N_14076,N_13816);
and U14548 (N_14548,N_14329,N_14313);
nand U14549 (N_14549,N_14233,N_13795);
and U14550 (N_14550,N_14270,N_14206);
nor U14551 (N_14551,N_14262,N_13932);
nor U14552 (N_14552,N_14381,N_14098);
xor U14553 (N_14553,N_13788,N_13822);
xnor U14554 (N_14554,N_13982,N_14213);
xor U14555 (N_14555,N_14382,N_14027);
nor U14556 (N_14556,N_13867,N_14086);
or U14557 (N_14557,N_13815,N_13945);
or U14558 (N_14558,N_14053,N_13669);
or U14559 (N_14559,N_13791,N_13648);
nor U14560 (N_14560,N_14291,N_14128);
xor U14561 (N_14561,N_13703,N_13685);
and U14562 (N_14562,N_13731,N_13638);
nand U14563 (N_14563,N_13846,N_13636);
nand U14564 (N_14564,N_14041,N_14322);
and U14565 (N_14565,N_13611,N_14159);
or U14566 (N_14566,N_14305,N_14354);
xor U14567 (N_14567,N_13713,N_14288);
nor U14568 (N_14568,N_14238,N_13785);
nor U14569 (N_14569,N_14282,N_14232);
nor U14570 (N_14570,N_14239,N_14303);
nor U14571 (N_14571,N_13914,N_13653);
nand U14572 (N_14572,N_13850,N_14134);
nor U14573 (N_14573,N_13918,N_14314);
and U14574 (N_14574,N_14332,N_13672);
or U14575 (N_14575,N_14164,N_14360);
nor U14576 (N_14576,N_13821,N_13747);
nor U14577 (N_14577,N_14327,N_13622);
nand U14578 (N_14578,N_14185,N_14014);
xor U14579 (N_14579,N_14094,N_14263);
xor U14580 (N_14580,N_14015,N_14132);
or U14581 (N_14581,N_13870,N_13646);
and U14582 (N_14582,N_14154,N_14127);
nor U14583 (N_14583,N_14049,N_13798);
nand U14584 (N_14584,N_13783,N_13915);
xnor U14585 (N_14585,N_14247,N_14043);
xor U14586 (N_14586,N_14297,N_14395);
xnor U14587 (N_14587,N_14145,N_14028);
xor U14588 (N_14588,N_13663,N_13955);
and U14589 (N_14589,N_13808,N_14174);
and U14590 (N_14590,N_14058,N_14003);
nor U14591 (N_14591,N_14267,N_14253);
nand U14592 (N_14592,N_14246,N_14265);
xnor U14593 (N_14593,N_13889,N_14350);
nand U14594 (N_14594,N_14005,N_14121);
or U14595 (N_14595,N_14168,N_13617);
or U14596 (N_14596,N_13640,N_13933);
and U14597 (N_14597,N_13680,N_14236);
nand U14598 (N_14598,N_14179,N_14045);
nor U14599 (N_14599,N_13792,N_13643);
nand U14600 (N_14600,N_13794,N_14391);
and U14601 (N_14601,N_13910,N_13678);
xor U14602 (N_14602,N_14103,N_13603);
nor U14603 (N_14603,N_13973,N_14230);
xnor U14604 (N_14604,N_14201,N_14119);
or U14605 (N_14605,N_14299,N_14384);
or U14606 (N_14606,N_13710,N_13699);
nand U14607 (N_14607,N_14368,N_14304);
nand U14608 (N_14608,N_14072,N_14320);
and U14609 (N_14609,N_14328,N_14301);
nand U14610 (N_14610,N_14318,N_14302);
or U14611 (N_14611,N_14025,N_14223);
or U14612 (N_14612,N_14274,N_14370);
and U14613 (N_14613,N_13954,N_13700);
or U14614 (N_14614,N_14338,N_14170);
xnor U14615 (N_14615,N_14009,N_13802);
xnor U14616 (N_14616,N_14160,N_14020);
nor U14617 (N_14617,N_13810,N_13869);
nor U14618 (N_14618,N_14225,N_13602);
xor U14619 (N_14619,N_14231,N_13707);
nor U14620 (N_14620,N_13725,N_13620);
nand U14621 (N_14621,N_13728,N_14092);
and U14622 (N_14622,N_14241,N_14216);
or U14623 (N_14623,N_14367,N_13994);
nand U14624 (N_14624,N_13827,N_14275);
or U14625 (N_14625,N_14385,N_14042);
xor U14626 (N_14626,N_14153,N_13667);
nor U14627 (N_14627,N_13968,N_13606);
xnor U14628 (N_14628,N_14061,N_14065);
or U14629 (N_14629,N_14372,N_13904);
xnor U14630 (N_14630,N_13920,N_14278);
and U14631 (N_14631,N_13600,N_14383);
xor U14632 (N_14632,N_13621,N_13739);
and U14633 (N_14633,N_13957,N_13628);
and U14634 (N_14634,N_13890,N_14001);
nand U14635 (N_14635,N_14373,N_14234);
and U14636 (N_14636,N_14150,N_14161);
or U14637 (N_14637,N_13844,N_13676);
or U14638 (N_14638,N_14087,N_13925);
nor U14639 (N_14639,N_13984,N_13983);
and U14640 (N_14640,N_14376,N_13691);
xor U14641 (N_14641,N_14349,N_13836);
nand U14642 (N_14642,N_13605,N_13855);
nor U14643 (N_14643,N_13734,N_13757);
or U14644 (N_14644,N_14369,N_14120);
nand U14645 (N_14645,N_14067,N_14273);
or U14646 (N_14646,N_13826,N_14074);
nand U14647 (N_14647,N_13718,N_14245);
and U14648 (N_14648,N_14090,N_13805);
nand U14649 (N_14649,N_13749,N_13959);
nor U14650 (N_14650,N_13859,N_13761);
xor U14651 (N_14651,N_13880,N_14192);
and U14652 (N_14652,N_13843,N_13863);
xnor U14653 (N_14653,N_14362,N_14392);
and U14654 (N_14654,N_13624,N_13709);
xnor U14655 (N_14655,N_13698,N_13755);
nor U14656 (N_14656,N_14397,N_13635);
nand U14657 (N_14657,N_13682,N_13686);
nand U14658 (N_14658,N_14022,N_13974);
nor U14659 (N_14659,N_13679,N_14276);
xnor U14660 (N_14660,N_13835,N_13849);
or U14661 (N_14661,N_13861,N_13909);
nand U14662 (N_14662,N_13659,N_14180);
or U14663 (N_14663,N_13921,N_13969);
and U14664 (N_14664,N_14342,N_14358);
xnor U14665 (N_14665,N_14029,N_14040);
nand U14666 (N_14666,N_14036,N_14151);
and U14667 (N_14667,N_13715,N_14295);
or U14668 (N_14668,N_13989,N_14084);
nand U14669 (N_14669,N_14173,N_14224);
and U14670 (N_14670,N_13630,N_14114);
xor U14671 (N_14671,N_14254,N_13650);
xnor U14672 (N_14672,N_13818,N_13931);
xor U14673 (N_14673,N_14016,N_13806);
nand U14674 (N_14674,N_14006,N_14187);
xor U14675 (N_14675,N_14083,N_14039);
or U14676 (N_14676,N_13769,N_14198);
and U14677 (N_14677,N_14344,N_14336);
and U14678 (N_14678,N_13875,N_13892);
nand U14679 (N_14679,N_14227,N_13926);
or U14680 (N_14680,N_14044,N_14289);
and U14681 (N_14681,N_14252,N_14181);
xnor U14682 (N_14682,N_13996,N_13733);
nand U14683 (N_14683,N_14010,N_13712);
nand U14684 (N_14684,N_14306,N_13868);
nand U14685 (N_14685,N_14351,N_14143);
nand U14686 (N_14686,N_14307,N_14242);
and U14687 (N_14687,N_13992,N_13666);
xor U14688 (N_14688,N_13740,N_13765);
nor U14689 (N_14689,N_13681,N_13772);
or U14690 (N_14690,N_14147,N_13977);
xnor U14691 (N_14691,N_14363,N_14281);
nor U14692 (N_14692,N_13637,N_13644);
or U14693 (N_14693,N_14283,N_14178);
or U14694 (N_14694,N_14324,N_13886);
xor U14695 (N_14695,N_13832,N_14207);
xnor U14696 (N_14696,N_13610,N_13723);
nand U14697 (N_14697,N_14280,N_14217);
and U14698 (N_14698,N_14047,N_14146);
nand U14699 (N_14699,N_14162,N_13741);
nor U14700 (N_14700,N_13937,N_13768);
or U14701 (N_14701,N_14286,N_14321);
xnor U14702 (N_14702,N_13693,N_14243);
nand U14703 (N_14703,N_13775,N_13664);
nor U14704 (N_14704,N_13946,N_14124);
nor U14705 (N_14705,N_14037,N_14317);
nor U14706 (N_14706,N_13883,N_14300);
nand U14707 (N_14707,N_14157,N_13838);
or U14708 (N_14708,N_14277,N_13702);
nor U14709 (N_14709,N_14131,N_14229);
nand U14710 (N_14710,N_13980,N_13776);
nand U14711 (N_14711,N_13990,N_13899);
nand U14712 (N_14712,N_13748,N_14220);
xnor U14713 (N_14713,N_13668,N_13911);
xor U14714 (N_14714,N_14200,N_14308);
nand U14715 (N_14715,N_13720,N_13917);
nand U14716 (N_14716,N_13814,N_13900);
nor U14717 (N_14717,N_14226,N_14294);
nand U14718 (N_14718,N_14082,N_14135);
nand U14719 (N_14719,N_13742,N_14059);
and U14720 (N_14720,N_13754,N_14080);
nor U14721 (N_14721,N_13609,N_14399);
and U14722 (N_14722,N_13670,N_13665);
and U14723 (N_14723,N_14366,N_14189);
or U14724 (N_14724,N_14050,N_13717);
or U14725 (N_14725,N_13927,N_13625);
nand U14726 (N_14726,N_14108,N_13963);
xnor U14727 (N_14727,N_14292,N_13898);
nor U14728 (N_14728,N_13732,N_13888);
and U14729 (N_14729,N_14379,N_13916);
or U14730 (N_14730,N_13662,N_13604);
or U14731 (N_14731,N_14148,N_14066);
and U14732 (N_14732,N_14257,N_13773);
nor U14733 (N_14733,N_14394,N_13997);
nand U14734 (N_14734,N_14250,N_13964);
nor U14735 (N_14735,N_13726,N_14352);
or U14736 (N_14736,N_13896,N_14102);
or U14737 (N_14737,N_14109,N_14096);
or U14738 (N_14738,N_13746,N_13619);
xor U14739 (N_14739,N_14116,N_14057);
and U14740 (N_14740,N_13966,N_14079);
xor U14741 (N_14741,N_14202,N_13944);
and U14742 (N_14742,N_14033,N_14240);
nand U14743 (N_14743,N_14337,N_14272);
nand U14744 (N_14744,N_14165,N_14218);
or U14745 (N_14745,N_13929,N_14364);
nor U14746 (N_14746,N_13858,N_14075);
nand U14747 (N_14747,N_13903,N_14000);
nor U14748 (N_14748,N_13657,N_14184);
or U14749 (N_14749,N_14051,N_13762);
or U14750 (N_14750,N_13677,N_14018);
xnor U14751 (N_14751,N_14149,N_14060);
and U14752 (N_14752,N_14055,N_13629);
or U14753 (N_14753,N_13626,N_13777);
xor U14754 (N_14754,N_13884,N_14071);
nand U14755 (N_14755,N_14333,N_14285);
nor U14756 (N_14756,N_13735,N_14063);
xnor U14757 (N_14757,N_13759,N_13839);
or U14758 (N_14758,N_14269,N_14319);
or U14759 (N_14759,N_14339,N_14371);
nand U14760 (N_14760,N_14054,N_13952);
nand U14761 (N_14761,N_13616,N_13877);
and U14762 (N_14762,N_14115,N_13789);
nor U14763 (N_14763,N_14093,N_14026);
nor U14764 (N_14764,N_13714,N_14196);
nand U14765 (N_14765,N_14176,N_14388);
nor U14766 (N_14766,N_13708,N_14258);
nor U14767 (N_14767,N_13771,N_14113);
nor U14768 (N_14768,N_14035,N_14073);
nor U14769 (N_14769,N_13993,N_13763);
nand U14770 (N_14770,N_14284,N_13866);
nand U14771 (N_14771,N_13842,N_13695);
nand U14772 (N_14772,N_13743,N_14139);
nor U14773 (N_14773,N_13930,N_13840);
or U14774 (N_14774,N_13800,N_13908);
xor U14775 (N_14775,N_14062,N_13953);
nand U14776 (N_14776,N_13879,N_14107);
nor U14777 (N_14777,N_14125,N_13906);
and U14778 (N_14778,N_14387,N_13862);
and U14779 (N_14779,N_13991,N_13956);
nor U14780 (N_14780,N_14353,N_14203);
nor U14781 (N_14781,N_14069,N_13770);
and U14782 (N_14782,N_14325,N_14126);
xor U14783 (N_14783,N_13675,N_14355);
and U14784 (N_14784,N_14315,N_13940);
or U14785 (N_14785,N_14112,N_14183);
or U14786 (N_14786,N_14359,N_14085);
nand U14787 (N_14787,N_14335,N_13975);
nor U14788 (N_14788,N_13601,N_13951);
or U14789 (N_14789,N_13841,N_14101);
and U14790 (N_14790,N_13758,N_13724);
and U14791 (N_14791,N_13860,N_14334);
and U14792 (N_14792,N_14175,N_14002);
or U14793 (N_14793,N_14249,N_14091);
or U14794 (N_14794,N_13961,N_14095);
xnor U14795 (N_14795,N_14244,N_14182);
and U14796 (N_14796,N_14386,N_13781);
nand U14797 (N_14797,N_13799,N_13829);
or U14798 (N_14798,N_14197,N_13854);
nor U14799 (N_14799,N_14031,N_13958);
and U14800 (N_14800,N_14287,N_14215);
or U14801 (N_14801,N_13927,N_13894);
or U14802 (N_14802,N_13911,N_13914);
or U14803 (N_14803,N_14294,N_14195);
nor U14804 (N_14804,N_13869,N_13750);
nand U14805 (N_14805,N_14284,N_13809);
xnor U14806 (N_14806,N_13705,N_14368);
or U14807 (N_14807,N_14081,N_13831);
and U14808 (N_14808,N_13818,N_14221);
and U14809 (N_14809,N_14019,N_13691);
or U14810 (N_14810,N_13696,N_14307);
or U14811 (N_14811,N_13718,N_14307);
or U14812 (N_14812,N_14173,N_13799);
or U14813 (N_14813,N_13768,N_14278);
nor U14814 (N_14814,N_14226,N_14151);
or U14815 (N_14815,N_13879,N_13720);
or U14816 (N_14816,N_13645,N_13709);
or U14817 (N_14817,N_14231,N_13909);
and U14818 (N_14818,N_14111,N_14342);
and U14819 (N_14819,N_14253,N_14236);
xor U14820 (N_14820,N_14173,N_14076);
or U14821 (N_14821,N_13792,N_13978);
nand U14822 (N_14822,N_13981,N_13704);
and U14823 (N_14823,N_14327,N_14371);
or U14824 (N_14824,N_14025,N_14136);
and U14825 (N_14825,N_14199,N_14019);
xnor U14826 (N_14826,N_13971,N_14384);
or U14827 (N_14827,N_13686,N_13999);
nand U14828 (N_14828,N_13879,N_13826);
nand U14829 (N_14829,N_14214,N_13794);
nor U14830 (N_14830,N_14390,N_13802);
and U14831 (N_14831,N_13643,N_13958);
and U14832 (N_14832,N_13866,N_14269);
nor U14833 (N_14833,N_14166,N_13626);
and U14834 (N_14834,N_14296,N_14073);
nor U14835 (N_14835,N_13836,N_13905);
nor U14836 (N_14836,N_13663,N_13886);
and U14837 (N_14837,N_14183,N_13941);
nand U14838 (N_14838,N_14285,N_13642);
xnor U14839 (N_14839,N_13810,N_14051);
nand U14840 (N_14840,N_14065,N_14384);
or U14841 (N_14841,N_13999,N_14051);
or U14842 (N_14842,N_14252,N_13779);
nor U14843 (N_14843,N_13615,N_13745);
nand U14844 (N_14844,N_13837,N_14310);
nor U14845 (N_14845,N_14085,N_14160);
or U14846 (N_14846,N_13886,N_13902);
xor U14847 (N_14847,N_13632,N_14308);
nor U14848 (N_14848,N_13744,N_13816);
nor U14849 (N_14849,N_13961,N_14129);
nor U14850 (N_14850,N_14155,N_13791);
and U14851 (N_14851,N_13718,N_14298);
and U14852 (N_14852,N_13813,N_13997);
or U14853 (N_14853,N_13602,N_13923);
and U14854 (N_14854,N_13890,N_14031);
xor U14855 (N_14855,N_13786,N_13650);
nor U14856 (N_14856,N_14296,N_13905);
xor U14857 (N_14857,N_14303,N_14199);
and U14858 (N_14858,N_14069,N_13989);
and U14859 (N_14859,N_13985,N_14327);
xor U14860 (N_14860,N_14272,N_14304);
nor U14861 (N_14861,N_14364,N_13691);
and U14862 (N_14862,N_14396,N_14134);
xor U14863 (N_14863,N_13623,N_14321);
nand U14864 (N_14864,N_13904,N_14091);
xor U14865 (N_14865,N_14116,N_13850);
nor U14866 (N_14866,N_14308,N_13963);
or U14867 (N_14867,N_13604,N_14216);
and U14868 (N_14868,N_13763,N_14367);
nor U14869 (N_14869,N_13705,N_14191);
nor U14870 (N_14870,N_13979,N_13656);
nor U14871 (N_14871,N_14066,N_14237);
nor U14872 (N_14872,N_13768,N_13853);
nand U14873 (N_14873,N_13675,N_13966);
or U14874 (N_14874,N_13677,N_13845);
or U14875 (N_14875,N_14253,N_14200);
and U14876 (N_14876,N_14338,N_14015);
and U14877 (N_14877,N_14229,N_14039);
and U14878 (N_14878,N_14215,N_13604);
and U14879 (N_14879,N_13881,N_13965);
or U14880 (N_14880,N_13914,N_13728);
and U14881 (N_14881,N_14331,N_13759);
or U14882 (N_14882,N_14096,N_13758);
or U14883 (N_14883,N_14069,N_13973);
and U14884 (N_14884,N_13865,N_13656);
or U14885 (N_14885,N_13928,N_13835);
and U14886 (N_14886,N_13963,N_14055);
xnor U14887 (N_14887,N_13738,N_14042);
nor U14888 (N_14888,N_14237,N_13850);
and U14889 (N_14889,N_13788,N_13818);
and U14890 (N_14890,N_13801,N_13678);
or U14891 (N_14891,N_14019,N_13785);
and U14892 (N_14892,N_13826,N_14359);
nand U14893 (N_14893,N_13661,N_14152);
nand U14894 (N_14894,N_13986,N_14034);
xor U14895 (N_14895,N_13816,N_14070);
or U14896 (N_14896,N_14195,N_14172);
and U14897 (N_14897,N_13610,N_14013);
nand U14898 (N_14898,N_13703,N_14296);
nand U14899 (N_14899,N_13683,N_14383);
nor U14900 (N_14900,N_13900,N_13943);
or U14901 (N_14901,N_14023,N_14286);
and U14902 (N_14902,N_13814,N_13844);
xor U14903 (N_14903,N_14303,N_14162);
nand U14904 (N_14904,N_14284,N_13738);
or U14905 (N_14905,N_13897,N_14304);
nand U14906 (N_14906,N_13953,N_14083);
nand U14907 (N_14907,N_14258,N_14166);
nor U14908 (N_14908,N_14365,N_13701);
nand U14909 (N_14909,N_13986,N_14225);
and U14910 (N_14910,N_14247,N_14120);
or U14911 (N_14911,N_13659,N_13925);
nand U14912 (N_14912,N_13738,N_14265);
or U14913 (N_14913,N_13914,N_13622);
nor U14914 (N_14914,N_14340,N_14366);
or U14915 (N_14915,N_14360,N_13622);
or U14916 (N_14916,N_14360,N_14350);
xor U14917 (N_14917,N_14110,N_13786);
nor U14918 (N_14918,N_14194,N_13777);
and U14919 (N_14919,N_14101,N_13853);
xnor U14920 (N_14920,N_14175,N_13781);
and U14921 (N_14921,N_13697,N_14144);
or U14922 (N_14922,N_14310,N_13708);
nand U14923 (N_14923,N_14182,N_13766);
and U14924 (N_14924,N_13630,N_13900);
nand U14925 (N_14925,N_13945,N_13717);
nand U14926 (N_14926,N_13824,N_13691);
nor U14927 (N_14927,N_13816,N_14177);
xor U14928 (N_14928,N_14116,N_14244);
or U14929 (N_14929,N_14256,N_14144);
nor U14930 (N_14930,N_14387,N_14224);
nor U14931 (N_14931,N_13827,N_13781);
xnor U14932 (N_14932,N_13975,N_13820);
and U14933 (N_14933,N_14291,N_13745);
nor U14934 (N_14934,N_13639,N_13604);
nand U14935 (N_14935,N_14164,N_13673);
xor U14936 (N_14936,N_14094,N_13659);
xnor U14937 (N_14937,N_13692,N_14068);
xor U14938 (N_14938,N_14235,N_13809);
nand U14939 (N_14939,N_14317,N_13623);
xnor U14940 (N_14940,N_13837,N_14069);
and U14941 (N_14941,N_14083,N_14381);
nor U14942 (N_14942,N_14000,N_14224);
and U14943 (N_14943,N_13940,N_14145);
or U14944 (N_14944,N_14273,N_14340);
xor U14945 (N_14945,N_14270,N_14181);
or U14946 (N_14946,N_14289,N_13915);
nor U14947 (N_14947,N_13847,N_14210);
or U14948 (N_14948,N_14155,N_14170);
nand U14949 (N_14949,N_14178,N_13632);
xnor U14950 (N_14950,N_13749,N_14126);
or U14951 (N_14951,N_13744,N_13768);
or U14952 (N_14952,N_14155,N_14103);
nand U14953 (N_14953,N_14263,N_14322);
nand U14954 (N_14954,N_14289,N_13709);
xnor U14955 (N_14955,N_14273,N_14177);
nand U14956 (N_14956,N_14086,N_13827);
and U14957 (N_14957,N_13699,N_14298);
xnor U14958 (N_14958,N_13974,N_13972);
or U14959 (N_14959,N_14168,N_14024);
and U14960 (N_14960,N_13878,N_14067);
nand U14961 (N_14961,N_14334,N_14065);
nor U14962 (N_14962,N_14216,N_13719);
nor U14963 (N_14963,N_14207,N_14381);
and U14964 (N_14964,N_14256,N_13766);
nor U14965 (N_14965,N_13703,N_13958);
and U14966 (N_14966,N_14157,N_14064);
and U14967 (N_14967,N_13842,N_14161);
xnor U14968 (N_14968,N_13691,N_14035);
xor U14969 (N_14969,N_14203,N_14090);
xor U14970 (N_14970,N_14313,N_13864);
xnor U14971 (N_14971,N_14316,N_14068);
xor U14972 (N_14972,N_13709,N_14242);
nand U14973 (N_14973,N_14093,N_13898);
and U14974 (N_14974,N_14359,N_14068);
and U14975 (N_14975,N_14301,N_13971);
and U14976 (N_14976,N_14112,N_13751);
nor U14977 (N_14977,N_13780,N_13872);
nand U14978 (N_14978,N_13936,N_13734);
xnor U14979 (N_14979,N_14133,N_13954);
and U14980 (N_14980,N_14154,N_14104);
or U14981 (N_14981,N_14007,N_13705);
xnor U14982 (N_14982,N_14055,N_13721);
xnor U14983 (N_14983,N_13790,N_13812);
or U14984 (N_14984,N_13916,N_13640);
xnor U14985 (N_14985,N_14176,N_14133);
or U14986 (N_14986,N_13875,N_13831);
and U14987 (N_14987,N_13623,N_14207);
xnor U14988 (N_14988,N_14398,N_13853);
and U14989 (N_14989,N_13881,N_14272);
and U14990 (N_14990,N_14306,N_13975);
nand U14991 (N_14991,N_13970,N_14230);
nand U14992 (N_14992,N_14344,N_14328);
and U14993 (N_14993,N_13959,N_14198);
or U14994 (N_14994,N_13920,N_13858);
nor U14995 (N_14995,N_13648,N_14358);
xor U14996 (N_14996,N_14269,N_14244);
and U14997 (N_14997,N_14242,N_14363);
or U14998 (N_14998,N_14094,N_14173);
nand U14999 (N_14999,N_13966,N_14291);
nand U15000 (N_15000,N_14278,N_13666);
nor U15001 (N_15001,N_14057,N_13976);
nor U15002 (N_15002,N_13899,N_13838);
nor U15003 (N_15003,N_14166,N_14377);
and U15004 (N_15004,N_13607,N_14275);
xnor U15005 (N_15005,N_14203,N_14028);
xor U15006 (N_15006,N_14015,N_13857);
or U15007 (N_15007,N_13630,N_13708);
nand U15008 (N_15008,N_14353,N_14265);
and U15009 (N_15009,N_14163,N_14372);
and U15010 (N_15010,N_13942,N_13768);
nor U15011 (N_15011,N_14018,N_14317);
or U15012 (N_15012,N_13948,N_13949);
nand U15013 (N_15013,N_14399,N_13845);
or U15014 (N_15014,N_14054,N_13695);
xnor U15015 (N_15015,N_13728,N_14246);
or U15016 (N_15016,N_14030,N_14219);
xor U15017 (N_15017,N_13746,N_14395);
nor U15018 (N_15018,N_13842,N_14275);
and U15019 (N_15019,N_13921,N_13832);
nor U15020 (N_15020,N_13680,N_14213);
and U15021 (N_15021,N_14268,N_13782);
or U15022 (N_15022,N_13894,N_14036);
xnor U15023 (N_15023,N_14375,N_13888);
nand U15024 (N_15024,N_14360,N_13606);
nand U15025 (N_15025,N_14126,N_13998);
and U15026 (N_15026,N_13781,N_13899);
xnor U15027 (N_15027,N_14103,N_13892);
nand U15028 (N_15028,N_13957,N_14250);
nand U15029 (N_15029,N_13682,N_14385);
and U15030 (N_15030,N_13918,N_13831);
nand U15031 (N_15031,N_13604,N_13619);
or U15032 (N_15032,N_14240,N_13894);
nand U15033 (N_15033,N_13686,N_14104);
nand U15034 (N_15034,N_13862,N_13642);
or U15035 (N_15035,N_14042,N_13890);
and U15036 (N_15036,N_13703,N_13925);
or U15037 (N_15037,N_14382,N_14294);
nor U15038 (N_15038,N_14122,N_14282);
or U15039 (N_15039,N_13608,N_13648);
or U15040 (N_15040,N_13899,N_14015);
xnor U15041 (N_15041,N_13842,N_13615);
nand U15042 (N_15042,N_13691,N_13625);
nand U15043 (N_15043,N_13639,N_14159);
nand U15044 (N_15044,N_14388,N_14232);
and U15045 (N_15045,N_14063,N_13876);
and U15046 (N_15046,N_14007,N_13890);
nor U15047 (N_15047,N_14122,N_14054);
nor U15048 (N_15048,N_13629,N_13659);
nor U15049 (N_15049,N_13667,N_14260);
nand U15050 (N_15050,N_14220,N_14287);
or U15051 (N_15051,N_13633,N_14294);
nor U15052 (N_15052,N_13747,N_13819);
nand U15053 (N_15053,N_13871,N_14175);
and U15054 (N_15054,N_13796,N_14092);
and U15055 (N_15055,N_14229,N_13950);
nor U15056 (N_15056,N_14296,N_14340);
nor U15057 (N_15057,N_14017,N_14220);
nand U15058 (N_15058,N_13843,N_13673);
or U15059 (N_15059,N_14044,N_13850);
nand U15060 (N_15060,N_14368,N_14027);
nand U15061 (N_15061,N_14144,N_13732);
xor U15062 (N_15062,N_13903,N_14110);
or U15063 (N_15063,N_13919,N_14121);
nor U15064 (N_15064,N_13813,N_14383);
nand U15065 (N_15065,N_13798,N_13843);
and U15066 (N_15066,N_13661,N_14145);
nor U15067 (N_15067,N_13975,N_13885);
and U15068 (N_15068,N_14207,N_13610);
and U15069 (N_15069,N_14390,N_13950);
xor U15070 (N_15070,N_13895,N_14164);
and U15071 (N_15071,N_13653,N_14042);
and U15072 (N_15072,N_13868,N_13663);
xnor U15073 (N_15073,N_13948,N_14005);
and U15074 (N_15074,N_13824,N_14394);
and U15075 (N_15075,N_13681,N_14294);
xnor U15076 (N_15076,N_14005,N_13913);
or U15077 (N_15077,N_13790,N_13643);
nand U15078 (N_15078,N_14323,N_13785);
xor U15079 (N_15079,N_13648,N_14327);
and U15080 (N_15080,N_13802,N_13859);
and U15081 (N_15081,N_14335,N_14019);
nor U15082 (N_15082,N_13809,N_13739);
nand U15083 (N_15083,N_14267,N_13693);
xnor U15084 (N_15084,N_13799,N_13839);
or U15085 (N_15085,N_13939,N_13707);
and U15086 (N_15086,N_14016,N_13653);
nor U15087 (N_15087,N_13726,N_14139);
and U15088 (N_15088,N_13975,N_13768);
nor U15089 (N_15089,N_14004,N_13689);
and U15090 (N_15090,N_13639,N_13891);
nand U15091 (N_15091,N_13637,N_13624);
and U15092 (N_15092,N_14038,N_13983);
xor U15093 (N_15093,N_13743,N_13753);
nor U15094 (N_15094,N_14094,N_13950);
nor U15095 (N_15095,N_13847,N_13756);
or U15096 (N_15096,N_14093,N_14303);
xor U15097 (N_15097,N_13612,N_14049);
xor U15098 (N_15098,N_13860,N_13898);
or U15099 (N_15099,N_13991,N_13797);
xnor U15100 (N_15100,N_14357,N_13726);
and U15101 (N_15101,N_13917,N_14102);
nand U15102 (N_15102,N_14065,N_14104);
xor U15103 (N_15103,N_13681,N_13684);
nor U15104 (N_15104,N_14200,N_13868);
and U15105 (N_15105,N_13899,N_13628);
or U15106 (N_15106,N_13946,N_13883);
and U15107 (N_15107,N_13953,N_13702);
nand U15108 (N_15108,N_13748,N_13784);
nor U15109 (N_15109,N_13949,N_14383);
or U15110 (N_15110,N_14382,N_14357);
nand U15111 (N_15111,N_13715,N_14043);
nor U15112 (N_15112,N_13864,N_14364);
nand U15113 (N_15113,N_13796,N_13704);
or U15114 (N_15114,N_13846,N_13723);
nand U15115 (N_15115,N_13909,N_14127);
nand U15116 (N_15116,N_13828,N_14358);
and U15117 (N_15117,N_13893,N_13937);
nor U15118 (N_15118,N_14196,N_13725);
or U15119 (N_15119,N_13931,N_13862);
nand U15120 (N_15120,N_13702,N_13698);
nand U15121 (N_15121,N_13625,N_14069);
nand U15122 (N_15122,N_14332,N_13652);
nor U15123 (N_15123,N_13649,N_14307);
and U15124 (N_15124,N_14335,N_14064);
nand U15125 (N_15125,N_14135,N_13981);
nor U15126 (N_15126,N_14021,N_13857);
xnor U15127 (N_15127,N_13816,N_14147);
nor U15128 (N_15128,N_13986,N_14136);
nand U15129 (N_15129,N_13880,N_13827);
nor U15130 (N_15130,N_13925,N_13878);
and U15131 (N_15131,N_13774,N_13942);
xor U15132 (N_15132,N_13991,N_13724);
nor U15133 (N_15133,N_14100,N_14345);
xor U15134 (N_15134,N_14046,N_13823);
and U15135 (N_15135,N_14367,N_13928);
nand U15136 (N_15136,N_14073,N_14229);
nand U15137 (N_15137,N_14257,N_14068);
or U15138 (N_15138,N_13714,N_14275);
nor U15139 (N_15139,N_14055,N_13923);
nand U15140 (N_15140,N_13995,N_14273);
xnor U15141 (N_15141,N_13604,N_14180);
xor U15142 (N_15142,N_14287,N_14295);
nand U15143 (N_15143,N_13641,N_13910);
xor U15144 (N_15144,N_13651,N_14396);
nor U15145 (N_15145,N_14164,N_14048);
nand U15146 (N_15146,N_13864,N_13819);
xor U15147 (N_15147,N_13863,N_14250);
nor U15148 (N_15148,N_13750,N_14219);
xnor U15149 (N_15149,N_14056,N_14383);
and U15150 (N_15150,N_14339,N_14071);
nand U15151 (N_15151,N_13982,N_13857);
or U15152 (N_15152,N_14352,N_13690);
or U15153 (N_15153,N_13939,N_13716);
and U15154 (N_15154,N_14247,N_14157);
nand U15155 (N_15155,N_14340,N_13949);
xnor U15156 (N_15156,N_14057,N_14036);
nor U15157 (N_15157,N_13649,N_14214);
nor U15158 (N_15158,N_14393,N_14348);
nand U15159 (N_15159,N_14277,N_14374);
nor U15160 (N_15160,N_13682,N_14023);
xnor U15161 (N_15161,N_14356,N_13813);
nor U15162 (N_15162,N_14020,N_13721);
xnor U15163 (N_15163,N_14146,N_13621);
and U15164 (N_15164,N_14010,N_14023);
and U15165 (N_15165,N_14073,N_13681);
nor U15166 (N_15166,N_13752,N_13801);
and U15167 (N_15167,N_14398,N_14087);
nor U15168 (N_15168,N_14015,N_14079);
and U15169 (N_15169,N_14101,N_14171);
nor U15170 (N_15170,N_14147,N_13705);
and U15171 (N_15171,N_14177,N_13738);
nor U15172 (N_15172,N_13643,N_14317);
and U15173 (N_15173,N_13681,N_14321);
and U15174 (N_15174,N_13943,N_14026);
nand U15175 (N_15175,N_13752,N_14306);
nor U15176 (N_15176,N_14391,N_13642);
or U15177 (N_15177,N_13610,N_14214);
nand U15178 (N_15178,N_14000,N_13917);
and U15179 (N_15179,N_13617,N_13740);
or U15180 (N_15180,N_13622,N_13638);
nand U15181 (N_15181,N_14124,N_14049);
nand U15182 (N_15182,N_14201,N_14223);
or U15183 (N_15183,N_14096,N_14258);
or U15184 (N_15184,N_13726,N_14011);
nor U15185 (N_15185,N_13636,N_14383);
and U15186 (N_15186,N_14035,N_13645);
nand U15187 (N_15187,N_14165,N_13686);
or U15188 (N_15188,N_14196,N_14114);
and U15189 (N_15189,N_14156,N_13814);
nand U15190 (N_15190,N_13865,N_14199);
and U15191 (N_15191,N_13997,N_13954);
nor U15192 (N_15192,N_14297,N_14163);
nand U15193 (N_15193,N_14000,N_13784);
and U15194 (N_15194,N_14206,N_14215);
and U15195 (N_15195,N_14399,N_14218);
nand U15196 (N_15196,N_14230,N_14109);
or U15197 (N_15197,N_14276,N_13672);
nand U15198 (N_15198,N_13787,N_13775);
nor U15199 (N_15199,N_13974,N_14118);
and U15200 (N_15200,N_14811,N_15074);
xor U15201 (N_15201,N_15021,N_14826);
nand U15202 (N_15202,N_14901,N_15137);
and U15203 (N_15203,N_14499,N_14790);
and U15204 (N_15204,N_14498,N_15175);
xnor U15205 (N_15205,N_14484,N_14475);
xor U15206 (N_15206,N_15095,N_14794);
xnor U15207 (N_15207,N_14633,N_14796);
and U15208 (N_15208,N_15163,N_14709);
nand U15209 (N_15209,N_15155,N_14688);
nand U15210 (N_15210,N_15084,N_15096);
nor U15211 (N_15211,N_14403,N_14741);
nor U15212 (N_15212,N_14420,N_14686);
nand U15213 (N_15213,N_14559,N_14402);
nor U15214 (N_15214,N_15143,N_14889);
nor U15215 (N_15215,N_14431,N_15154);
nand U15216 (N_15216,N_14508,N_14707);
and U15217 (N_15217,N_14531,N_15146);
xor U15218 (N_15218,N_15159,N_14757);
and U15219 (N_15219,N_14868,N_14933);
or U15220 (N_15220,N_14733,N_14478);
nor U15221 (N_15221,N_14834,N_14614);
xnor U15222 (N_15222,N_14501,N_15189);
xor U15223 (N_15223,N_14777,N_14831);
nand U15224 (N_15224,N_15157,N_14791);
and U15225 (N_15225,N_14685,N_14620);
xnor U15226 (N_15226,N_14763,N_14819);
and U15227 (N_15227,N_15044,N_14795);
nand U15228 (N_15228,N_14609,N_14929);
nor U15229 (N_15229,N_15029,N_14829);
or U15230 (N_15230,N_14601,N_15142);
nor U15231 (N_15231,N_15153,N_15134);
and U15232 (N_15232,N_14896,N_14443);
xor U15233 (N_15233,N_14664,N_14532);
and U15234 (N_15234,N_14881,N_14982);
or U15235 (N_15235,N_14586,N_15080);
and U15236 (N_15236,N_14738,N_15123);
nand U15237 (N_15237,N_14674,N_14976);
nor U15238 (N_15238,N_14936,N_14770);
nand U15239 (N_15239,N_14666,N_15145);
xnor U15240 (N_15240,N_14765,N_14618);
nand U15241 (N_15241,N_14466,N_15152);
nor U15242 (N_15242,N_14463,N_15090);
or U15243 (N_15243,N_14673,N_14862);
xor U15244 (N_15244,N_14989,N_14556);
nor U15245 (N_15245,N_14818,N_15129);
nor U15246 (N_15246,N_15094,N_14458);
or U15247 (N_15247,N_14595,N_14997);
or U15248 (N_15248,N_15144,N_14840);
nor U15249 (N_15249,N_15151,N_15100);
or U15250 (N_15250,N_14900,N_15086);
and U15251 (N_15251,N_15050,N_15078);
or U15252 (N_15252,N_15024,N_14596);
xor U15253 (N_15253,N_15106,N_14668);
and U15254 (N_15254,N_14932,N_14805);
and U15255 (N_15255,N_15149,N_14477);
and U15256 (N_15256,N_14870,N_14564);
nand U15257 (N_15257,N_15131,N_14812);
xnor U15258 (N_15258,N_14766,N_14636);
nor U15259 (N_15259,N_14429,N_15199);
xor U15260 (N_15260,N_14621,N_15121);
nor U15261 (N_15261,N_14942,N_14582);
and U15262 (N_15262,N_14680,N_15102);
xnor U15263 (N_15263,N_15048,N_15170);
and U15264 (N_15264,N_14504,N_14612);
xnor U15265 (N_15265,N_14563,N_14585);
nand U15266 (N_15266,N_15103,N_14937);
or U15267 (N_15267,N_14972,N_14503);
and U15268 (N_15268,N_15197,N_14474);
and U15269 (N_15269,N_14873,N_14592);
nor U15270 (N_15270,N_14914,N_14682);
and U15271 (N_15271,N_14720,N_15133);
nor U15272 (N_15272,N_14439,N_14782);
and U15273 (N_15273,N_14607,N_14441);
or U15274 (N_15274,N_15196,N_15191);
xor U15275 (N_15275,N_14800,N_14945);
and U15276 (N_15276,N_14877,N_14671);
and U15277 (N_15277,N_14574,N_14412);
and U15278 (N_15278,N_15188,N_14657);
xor U15279 (N_15279,N_14573,N_14539);
nor U15280 (N_15280,N_14602,N_14645);
xor U15281 (N_15281,N_14507,N_15171);
nor U15282 (N_15282,N_14572,N_14658);
xor U15283 (N_15283,N_15039,N_14428);
xnor U15284 (N_15284,N_14605,N_14462);
nand U15285 (N_15285,N_14995,N_14405);
xor U15286 (N_15286,N_15006,N_14784);
and U15287 (N_15287,N_14486,N_14561);
or U15288 (N_15288,N_14404,N_14825);
nand U15289 (N_15289,N_14670,N_14489);
nand U15290 (N_15290,N_14957,N_14437);
nor U15291 (N_15291,N_15122,N_14640);
xor U15292 (N_15292,N_14922,N_14724);
or U15293 (N_15293,N_14919,N_14654);
xnor U15294 (N_15294,N_14599,N_14655);
and U15295 (N_15295,N_14481,N_14844);
nand U15296 (N_15296,N_14760,N_14952);
nor U15297 (N_15297,N_14701,N_14464);
and U15298 (N_15298,N_14468,N_15003);
nor U15299 (N_15299,N_14704,N_14822);
nor U15300 (N_15300,N_14597,N_14820);
or U15301 (N_15301,N_14759,N_14912);
xor U15302 (N_15302,N_14438,N_14642);
nand U15303 (N_15303,N_14648,N_15043);
xnor U15304 (N_15304,N_14669,N_15194);
nand U15305 (N_15305,N_14465,N_15112);
or U15306 (N_15306,N_14581,N_14742);
xnor U15307 (N_15307,N_14743,N_14702);
xnor U15308 (N_15308,N_15088,N_14547);
nand U15309 (N_15309,N_14440,N_14970);
xnor U15310 (N_15310,N_14899,N_14697);
or U15311 (N_15311,N_14600,N_14778);
and U15312 (N_15312,N_14786,N_15184);
xor U15313 (N_15313,N_15054,N_14793);
nand U15314 (N_15314,N_15045,N_14689);
or U15315 (N_15315,N_14783,N_14435);
xnor U15316 (N_15316,N_14538,N_14959);
nor U15317 (N_15317,N_14421,N_14413);
or U15318 (N_15318,N_14522,N_14543);
nor U15319 (N_15319,N_15014,N_14677);
and U15320 (N_15320,N_14603,N_14551);
or U15321 (N_15321,N_14434,N_14731);
nand U15322 (N_15322,N_14994,N_14857);
nor U15323 (N_15323,N_14576,N_15178);
nor U15324 (N_15324,N_14888,N_15023);
and U15325 (N_15325,N_14517,N_14588);
nand U15326 (N_15326,N_14898,N_14909);
xnor U15327 (N_15327,N_14913,N_14905);
nor U15328 (N_15328,N_15051,N_14789);
nor U15329 (N_15329,N_14652,N_14734);
nor U15330 (N_15330,N_14717,N_14848);
xor U15331 (N_15331,N_14852,N_14509);
and U15332 (N_15332,N_14983,N_15119);
and U15333 (N_15333,N_14892,N_14529);
nand U15334 (N_15334,N_14758,N_14448);
nor U15335 (N_15335,N_14647,N_14549);
xor U15336 (N_15336,N_14955,N_14562);
and U15337 (N_15337,N_15047,N_15064);
xor U15338 (N_15338,N_14611,N_14527);
nor U15339 (N_15339,N_14617,N_14569);
nand U15340 (N_15340,N_14984,N_14842);
nand U15341 (N_15341,N_14943,N_15139);
and U15342 (N_15342,N_14502,N_14737);
nor U15343 (N_15343,N_14537,N_14662);
nand U15344 (N_15344,N_15030,N_14453);
and U15345 (N_15345,N_14941,N_14423);
xnor U15346 (N_15346,N_14926,N_14823);
nand U15347 (N_15347,N_14452,N_14485);
xor U15348 (N_15348,N_15111,N_14968);
nor U15349 (N_15349,N_14946,N_14807);
xor U15350 (N_15350,N_14653,N_14418);
and U15351 (N_15351,N_15010,N_14623);
xnor U15352 (N_15352,N_14885,N_14882);
or U15353 (N_15353,N_14513,N_14860);
xnor U15354 (N_15354,N_14838,N_14841);
and U15355 (N_15355,N_14866,N_14634);
nor U15356 (N_15356,N_14749,N_14487);
nor U15357 (N_15357,N_14444,N_14753);
xor U15358 (N_15358,N_14449,N_14571);
nand U15359 (N_15359,N_14663,N_14471);
nand U15360 (N_15360,N_14739,N_15173);
xor U15361 (N_15361,N_14925,N_14960);
or U15362 (N_15362,N_14523,N_15069);
and U15363 (N_15363,N_14804,N_14643);
xor U15364 (N_15364,N_15049,N_14545);
nor U15365 (N_15365,N_14872,N_14850);
nor U15366 (N_15366,N_14988,N_14698);
xor U15367 (N_15367,N_14797,N_14803);
nor U15368 (N_15368,N_14917,N_15098);
nor U15369 (N_15369,N_14775,N_14986);
nor U15370 (N_15370,N_14718,N_14506);
xnor U15371 (N_15371,N_14525,N_15198);
nand U15372 (N_15372,N_15038,N_15002);
xor U15373 (N_15373,N_15081,N_14521);
nand U15374 (N_15374,N_14526,N_15185);
nand U15375 (N_15375,N_14419,N_14990);
and U15376 (N_15376,N_14962,N_14833);
nor U15377 (N_15377,N_14726,N_15034);
nand U15378 (N_15378,N_14802,N_14921);
nor U15379 (N_15379,N_15075,N_14625);
or U15380 (N_15380,N_14678,N_14846);
nor U15381 (N_15381,N_14514,N_14713);
or U15382 (N_15382,N_15042,N_14771);
nor U15383 (N_15383,N_15190,N_15031);
and U15384 (N_15384,N_14637,N_14849);
or U15385 (N_15385,N_14510,N_14540);
and U15386 (N_15386,N_14656,N_14616);
xnor U15387 (N_15387,N_14948,N_14967);
and U15388 (N_15388,N_14815,N_15033);
nor U15389 (N_15389,N_14944,N_14954);
xnor U15390 (N_15390,N_14975,N_14740);
nand U15391 (N_15391,N_14542,N_14461);
nor U15392 (N_15392,N_14512,N_14401);
and U15393 (N_15393,N_14426,N_15057);
nand U15394 (N_15394,N_14493,N_14861);
and U15395 (N_15395,N_14978,N_14703);
and U15396 (N_15396,N_15169,N_14830);
nor U15397 (N_15397,N_15053,N_14411);
nor U15398 (N_15398,N_14554,N_14548);
nand U15399 (N_15399,N_14934,N_15135);
and U15400 (N_15400,N_15176,N_15126);
nand U15401 (N_15401,N_14971,N_14446);
or U15402 (N_15402,N_14858,N_14949);
and U15403 (N_15403,N_14706,N_14774);
xnor U15404 (N_15404,N_14495,N_15093);
and U15405 (N_15405,N_15182,N_15109);
nor U15406 (N_15406,N_14692,N_15150);
xnor U15407 (N_15407,N_14956,N_14496);
or U15408 (N_15408,N_14469,N_14751);
xnor U15409 (N_15409,N_14890,N_15046);
xor U15410 (N_15410,N_14998,N_14627);
or U15411 (N_15411,N_14589,N_14644);
xnor U15412 (N_15412,N_14999,N_14750);
or U15413 (N_15413,N_15160,N_14483);
nor U15414 (N_15414,N_15183,N_14817);
nand U15415 (N_15415,N_14828,N_14708);
nor U15416 (N_15416,N_15092,N_14565);
nor U15417 (N_15417,N_14410,N_14746);
nor U15418 (N_15418,N_14785,N_14553);
and U15419 (N_15419,N_14631,N_14808);
nand U15420 (N_15420,N_15013,N_15124);
xor U15421 (N_15421,N_14409,N_14604);
and U15422 (N_15422,N_15132,N_14966);
nand U15423 (N_15423,N_14725,N_14855);
xor U15424 (N_15424,N_14460,N_14594);
and U15425 (N_15425,N_15179,N_14883);
or U15426 (N_15426,N_15138,N_14583);
nor U15427 (N_15427,N_14768,N_15097);
and U15428 (N_15428,N_14824,N_14691);
xnor U15429 (N_15429,N_14615,N_14608);
and U15430 (N_15430,N_14492,N_15165);
xor U15431 (N_15431,N_14871,N_14963);
xnor U15432 (N_15432,N_14406,N_14884);
and U15433 (N_15433,N_14488,N_14683);
xnor U15434 (N_15434,N_14414,N_14927);
and U15435 (N_15435,N_14518,N_14696);
nor U15436 (N_15436,N_14788,N_14752);
and U15437 (N_15437,N_15022,N_14544);
and U15438 (N_15438,N_15099,N_14856);
and U15439 (N_15439,N_14575,N_14675);
nor U15440 (N_15440,N_14442,N_15065);
xnor U15441 (N_15441,N_14735,N_15187);
nor U15442 (N_15442,N_14425,N_14814);
nand U15443 (N_15443,N_14451,N_15161);
or U15444 (N_15444,N_15177,N_14570);
and U15445 (N_15445,N_14695,N_15073);
nor U15446 (N_15446,N_15041,N_14969);
nand U15447 (N_15447,N_15027,N_14646);
nor U15448 (N_15448,N_14580,N_15089);
xor U15449 (N_15449,N_14520,N_14613);
and U15450 (N_15450,N_14908,N_15125);
or U15451 (N_15451,N_14938,N_14920);
or U15452 (N_15452,N_14756,N_14910);
xnor U15453 (N_15453,N_14979,N_14953);
nor U15454 (N_15454,N_14904,N_14710);
and U15455 (N_15455,N_14832,N_15077);
or U15456 (N_15456,N_15001,N_14447);
or U15457 (N_15457,N_14864,N_15181);
or U15458 (N_15458,N_15108,N_14558);
nor U15459 (N_15459,N_14931,N_14454);
and U15460 (N_15460,N_14649,N_14996);
or U15461 (N_15461,N_14799,N_14810);
nor U15462 (N_15462,N_14773,N_14473);
or U15463 (N_15463,N_15068,N_14874);
or U15464 (N_15464,N_15082,N_15004);
nor U15465 (N_15465,N_14991,N_15059);
nor U15466 (N_15466,N_15066,N_14672);
xor U15467 (N_15467,N_14534,N_14598);
xnor U15468 (N_15468,N_15018,N_14456);
nor U15469 (N_15469,N_14835,N_14781);
and U15470 (N_15470,N_14610,N_14433);
nand U15471 (N_15471,N_15117,N_14516);
and U15472 (N_15472,N_14745,N_14470);
nor U15473 (N_15473,N_15020,N_14711);
nor U15474 (N_15474,N_15110,N_14619);
nand U15475 (N_15475,N_14515,N_14755);
and U15476 (N_15476,N_15067,N_15072);
and U15477 (N_15477,N_14584,N_14935);
xor U15478 (N_15478,N_15147,N_14965);
xnor U15479 (N_15479,N_15140,N_14903);
nand U15480 (N_15480,N_14816,N_14568);
or U15481 (N_15481,N_15167,N_14730);
xor U15482 (N_15482,N_15158,N_14630);
nor U15483 (N_15483,N_14762,N_14587);
and U15484 (N_15484,N_14827,N_14843);
nor U15485 (N_15485,N_14736,N_14641);
nor U15486 (N_15486,N_14906,N_15087);
nand U15487 (N_15487,N_15083,N_14930);
nand U15488 (N_15488,N_14550,N_15012);
nor U15489 (N_15489,N_14459,N_15141);
xnor U15490 (N_15490,N_14891,N_15172);
nor U15491 (N_15491,N_14727,N_14407);
nand U15492 (N_15492,N_15168,N_14776);
xnor U15493 (N_15493,N_14639,N_14536);
nor U15494 (N_15494,N_14422,N_15127);
and U15495 (N_15495,N_15104,N_15008);
or U15496 (N_15496,N_14552,N_14651);
nand U15497 (N_15497,N_14687,N_14923);
and U15498 (N_15498,N_14867,N_15101);
or U15499 (N_15499,N_14894,N_14676);
or U15500 (N_15500,N_14974,N_14836);
xor U15501 (N_15501,N_15015,N_14809);
nand U15502 (N_15502,N_14940,N_14694);
nand U15503 (N_15503,N_15061,N_14787);
and U15504 (N_15504,N_14902,N_14699);
xnor U15505 (N_15505,N_14723,N_15091);
nor U15506 (N_15506,N_14457,N_15017);
nand U15507 (N_15507,N_14764,N_15156);
nand U15508 (N_15508,N_15019,N_14907);
nand U15509 (N_15509,N_14721,N_14432);
or U15510 (N_15510,N_15076,N_15186);
nand U15511 (N_15511,N_15195,N_14528);
xor U15512 (N_15512,N_14916,N_15040);
and U15513 (N_15513,N_14450,N_14780);
nor U15514 (N_15514,N_14590,N_15037);
or U15515 (N_15515,N_14436,N_15136);
or U15516 (N_15516,N_14557,N_14494);
or U15517 (N_15517,N_15192,N_14579);
or U15518 (N_15518,N_14497,N_14744);
xnor U15519 (N_15519,N_14977,N_14684);
nor U15520 (N_15520,N_14924,N_14500);
and U15521 (N_15521,N_14415,N_14491);
or U15522 (N_15522,N_14801,N_14511);
xor U15523 (N_15523,N_14530,N_14593);
nand U15524 (N_15524,N_14918,N_15032);
xnor U15525 (N_15525,N_14728,N_14661);
nand U15526 (N_15526,N_14524,N_15116);
or U15527 (N_15527,N_14679,N_14626);
nor U15528 (N_15528,N_15120,N_14869);
or U15529 (N_15529,N_15009,N_14719);
nor U15530 (N_15530,N_14577,N_15063);
xnor U15531 (N_15531,N_14981,N_14839);
and U15532 (N_15532,N_14408,N_15005);
nand U15533 (N_15533,N_14772,N_14876);
xnor U15534 (N_15534,N_14992,N_15174);
xnor U15535 (N_15535,N_14535,N_14417);
and U15536 (N_15536,N_14400,N_14628);
or U15537 (N_15537,N_14427,N_14928);
nand U15538 (N_15538,N_14445,N_14961);
nand U15539 (N_15539,N_14947,N_14851);
or U15540 (N_15540,N_15056,N_15052);
nand U15541 (N_15541,N_14754,N_14690);
xor U15542 (N_15542,N_15007,N_15000);
nand U15543 (N_15543,N_15011,N_15055);
nor U15544 (N_15544,N_14886,N_14560);
nand U15545 (N_15545,N_14813,N_14939);
xor U15546 (N_15546,N_14566,N_14424);
and U15547 (N_15547,N_14878,N_14490);
nor U15548 (N_15548,N_15036,N_14430);
xnor U15549 (N_15549,N_14769,N_14865);
xnor U15550 (N_15550,N_14480,N_15058);
or U15551 (N_15551,N_14629,N_14806);
xnor U15552 (N_15552,N_14519,N_14951);
nor U15553 (N_15553,N_14779,N_14650);
xnor U15554 (N_15554,N_15035,N_14712);
nand U15555 (N_15555,N_14845,N_14681);
nor U15556 (N_15556,N_14897,N_14467);
nor U15557 (N_15557,N_15128,N_14748);
nor U15558 (N_15558,N_14455,N_15115);
and U15559 (N_15559,N_14847,N_14732);
xnor U15560 (N_15560,N_14798,N_14638);
xnor U15561 (N_15561,N_15164,N_15026);
nor U15562 (N_15562,N_14911,N_15114);
xor U15563 (N_15563,N_14714,N_15107);
nor U15564 (N_15564,N_14591,N_14985);
nand U15565 (N_15565,N_15060,N_14567);
nand U15566 (N_15566,N_14722,N_15070);
or U15567 (N_15567,N_14482,N_14700);
nand U15568 (N_15568,N_14622,N_14505);
nor U15569 (N_15569,N_14705,N_14837);
and U15570 (N_15570,N_15118,N_14767);
or U15571 (N_15571,N_14476,N_15016);
nand U15572 (N_15572,N_14555,N_14624);
or U15573 (N_15573,N_15162,N_14761);
and U15574 (N_15574,N_14606,N_15079);
or U15575 (N_15575,N_15113,N_14667);
xnor U15576 (N_15576,N_14853,N_15180);
nand U15577 (N_15577,N_15166,N_14747);
nand U15578 (N_15578,N_14980,N_14541);
and U15579 (N_15579,N_14821,N_15071);
or U15580 (N_15580,N_14863,N_14533);
or U15581 (N_15581,N_14546,N_14693);
nor U15582 (N_15582,N_14854,N_15062);
xor U15583 (N_15583,N_14950,N_15028);
nor U15584 (N_15584,N_15085,N_14973);
and U15585 (N_15585,N_14578,N_14895);
xnor U15586 (N_15586,N_14879,N_14716);
nand U15587 (N_15587,N_14635,N_14964);
xor U15588 (N_15588,N_14958,N_15148);
nand U15589 (N_15589,N_14416,N_14893);
nor U15590 (N_15590,N_14915,N_14479);
and U15591 (N_15591,N_14887,N_14792);
xnor U15592 (N_15592,N_14715,N_14472);
and U15593 (N_15593,N_14729,N_15193);
and U15594 (N_15594,N_15130,N_14665);
or U15595 (N_15595,N_15105,N_14993);
nor U15596 (N_15596,N_14987,N_14660);
or U15597 (N_15597,N_15025,N_14659);
nand U15598 (N_15598,N_14875,N_14880);
xor U15599 (N_15599,N_14859,N_14632);
xnor U15600 (N_15600,N_14687,N_14430);
nand U15601 (N_15601,N_14826,N_14659);
or U15602 (N_15602,N_15155,N_14933);
nand U15603 (N_15603,N_14880,N_14653);
and U15604 (N_15604,N_14658,N_14884);
and U15605 (N_15605,N_14672,N_14553);
or U15606 (N_15606,N_14601,N_14745);
xor U15607 (N_15607,N_14419,N_14517);
xor U15608 (N_15608,N_14519,N_14697);
nand U15609 (N_15609,N_15086,N_14683);
or U15610 (N_15610,N_14870,N_14800);
nand U15611 (N_15611,N_14700,N_15068);
and U15612 (N_15612,N_14479,N_15059);
nor U15613 (N_15613,N_14925,N_14709);
and U15614 (N_15614,N_14723,N_14895);
nand U15615 (N_15615,N_15037,N_14487);
xnor U15616 (N_15616,N_15172,N_14767);
or U15617 (N_15617,N_14812,N_14909);
xnor U15618 (N_15618,N_14921,N_15071);
or U15619 (N_15619,N_14846,N_15064);
nor U15620 (N_15620,N_14499,N_15019);
nand U15621 (N_15621,N_15108,N_14569);
xor U15622 (N_15622,N_14851,N_14756);
nor U15623 (N_15623,N_14718,N_14942);
and U15624 (N_15624,N_14980,N_14969);
or U15625 (N_15625,N_14541,N_14483);
nand U15626 (N_15626,N_14910,N_14858);
nand U15627 (N_15627,N_14775,N_15014);
and U15628 (N_15628,N_15009,N_14771);
or U15629 (N_15629,N_15033,N_15046);
or U15630 (N_15630,N_14788,N_14453);
and U15631 (N_15631,N_14856,N_14560);
and U15632 (N_15632,N_14628,N_14972);
nand U15633 (N_15633,N_15048,N_14538);
nor U15634 (N_15634,N_15035,N_14713);
and U15635 (N_15635,N_14460,N_14439);
nand U15636 (N_15636,N_15053,N_15106);
nand U15637 (N_15637,N_15105,N_14865);
or U15638 (N_15638,N_15141,N_15078);
nor U15639 (N_15639,N_14782,N_14742);
and U15640 (N_15640,N_14622,N_14479);
nor U15641 (N_15641,N_14533,N_14920);
and U15642 (N_15642,N_14405,N_15162);
and U15643 (N_15643,N_14962,N_15032);
xor U15644 (N_15644,N_14907,N_15116);
nand U15645 (N_15645,N_14748,N_14650);
nor U15646 (N_15646,N_15126,N_15081);
or U15647 (N_15647,N_14432,N_15016);
nand U15648 (N_15648,N_14440,N_14607);
nor U15649 (N_15649,N_15143,N_14576);
and U15650 (N_15650,N_14938,N_14478);
xnor U15651 (N_15651,N_14768,N_14570);
nor U15652 (N_15652,N_14765,N_14430);
and U15653 (N_15653,N_14587,N_14418);
nand U15654 (N_15654,N_15007,N_14833);
nor U15655 (N_15655,N_14495,N_14407);
xor U15656 (N_15656,N_14799,N_15100);
nand U15657 (N_15657,N_14659,N_14853);
xor U15658 (N_15658,N_14940,N_15150);
nor U15659 (N_15659,N_14416,N_14606);
and U15660 (N_15660,N_14593,N_14985);
and U15661 (N_15661,N_14707,N_14557);
nand U15662 (N_15662,N_14500,N_14769);
nor U15663 (N_15663,N_15143,N_14748);
xnor U15664 (N_15664,N_14997,N_14920);
or U15665 (N_15665,N_14623,N_15030);
or U15666 (N_15666,N_14805,N_15006);
or U15667 (N_15667,N_15030,N_15061);
xnor U15668 (N_15668,N_14883,N_15167);
and U15669 (N_15669,N_14406,N_14958);
or U15670 (N_15670,N_14424,N_14849);
xnor U15671 (N_15671,N_14779,N_14530);
and U15672 (N_15672,N_14409,N_14563);
nor U15673 (N_15673,N_15154,N_14501);
and U15674 (N_15674,N_14670,N_14962);
xnor U15675 (N_15675,N_14484,N_14469);
nand U15676 (N_15676,N_14591,N_14742);
nand U15677 (N_15677,N_14990,N_15102);
and U15678 (N_15678,N_14604,N_14951);
nand U15679 (N_15679,N_15007,N_15002);
nand U15680 (N_15680,N_14688,N_14979);
xor U15681 (N_15681,N_14891,N_15194);
xnor U15682 (N_15682,N_14696,N_15164);
or U15683 (N_15683,N_14588,N_14551);
or U15684 (N_15684,N_14462,N_15031);
and U15685 (N_15685,N_14712,N_14762);
and U15686 (N_15686,N_15072,N_14440);
nand U15687 (N_15687,N_14985,N_14423);
nand U15688 (N_15688,N_15188,N_14540);
nand U15689 (N_15689,N_14732,N_14619);
or U15690 (N_15690,N_14422,N_14821);
and U15691 (N_15691,N_14634,N_14937);
xor U15692 (N_15692,N_14748,N_14775);
nor U15693 (N_15693,N_14535,N_14822);
or U15694 (N_15694,N_14792,N_14937);
or U15695 (N_15695,N_14684,N_14429);
nor U15696 (N_15696,N_14564,N_14413);
and U15697 (N_15697,N_14956,N_14490);
or U15698 (N_15698,N_14930,N_15072);
and U15699 (N_15699,N_15176,N_14498);
and U15700 (N_15700,N_15089,N_14789);
nand U15701 (N_15701,N_14791,N_14556);
and U15702 (N_15702,N_14969,N_14591);
nand U15703 (N_15703,N_14854,N_15097);
xor U15704 (N_15704,N_15042,N_14621);
nor U15705 (N_15705,N_14467,N_14493);
or U15706 (N_15706,N_14666,N_14969);
or U15707 (N_15707,N_15136,N_15062);
nand U15708 (N_15708,N_14514,N_15081);
xor U15709 (N_15709,N_14450,N_14884);
and U15710 (N_15710,N_14788,N_14815);
nand U15711 (N_15711,N_14928,N_14676);
or U15712 (N_15712,N_14855,N_15097);
nand U15713 (N_15713,N_14742,N_14564);
or U15714 (N_15714,N_14748,N_14958);
nand U15715 (N_15715,N_15127,N_14919);
and U15716 (N_15716,N_15169,N_15163);
nor U15717 (N_15717,N_15042,N_14778);
nand U15718 (N_15718,N_14422,N_14818);
xnor U15719 (N_15719,N_14507,N_14658);
nand U15720 (N_15720,N_15007,N_15084);
nand U15721 (N_15721,N_14578,N_15026);
xor U15722 (N_15722,N_14857,N_15115);
or U15723 (N_15723,N_15185,N_15085);
xnor U15724 (N_15724,N_14442,N_14518);
nor U15725 (N_15725,N_14451,N_14593);
nand U15726 (N_15726,N_14968,N_14662);
and U15727 (N_15727,N_15133,N_14668);
and U15728 (N_15728,N_15134,N_14939);
xnor U15729 (N_15729,N_14495,N_14519);
or U15730 (N_15730,N_14410,N_14475);
and U15731 (N_15731,N_14686,N_14666);
nor U15732 (N_15732,N_14414,N_15069);
nor U15733 (N_15733,N_14984,N_15103);
or U15734 (N_15734,N_14949,N_14580);
nand U15735 (N_15735,N_14658,N_15131);
nor U15736 (N_15736,N_14667,N_14986);
or U15737 (N_15737,N_14624,N_14852);
nand U15738 (N_15738,N_14857,N_14674);
or U15739 (N_15739,N_14964,N_14883);
nor U15740 (N_15740,N_14569,N_14497);
nor U15741 (N_15741,N_14587,N_14781);
nor U15742 (N_15742,N_15003,N_14655);
or U15743 (N_15743,N_14554,N_15105);
or U15744 (N_15744,N_14892,N_14742);
and U15745 (N_15745,N_15196,N_14867);
xor U15746 (N_15746,N_14445,N_15105);
nand U15747 (N_15747,N_14652,N_14547);
or U15748 (N_15748,N_14667,N_15139);
and U15749 (N_15749,N_15145,N_14658);
nand U15750 (N_15750,N_14885,N_14927);
nand U15751 (N_15751,N_14418,N_14484);
nand U15752 (N_15752,N_14864,N_15030);
xnor U15753 (N_15753,N_14901,N_14803);
xnor U15754 (N_15754,N_14741,N_15123);
and U15755 (N_15755,N_14729,N_14771);
and U15756 (N_15756,N_15152,N_14947);
nand U15757 (N_15757,N_14925,N_14589);
nor U15758 (N_15758,N_14683,N_15198);
and U15759 (N_15759,N_14496,N_14546);
nor U15760 (N_15760,N_14799,N_14853);
and U15761 (N_15761,N_15022,N_15070);
and U15762 (N_15762,N_14607,N_14433);
or U15763 (N_15763,N_15127,N_15096);
nand U15764 (N_15764,N_14575,N_15006);
nand U15765 (N_15765,N_14538,N_14463);
nand U15766 (N_15766,N_14608,N_14966);
xnor U15767 (N_15767,N_15028,N_14615);
xor U15768 (N_15768,N_14863,N_14853);
or U15769 (N_15769,N_14563,N_15136);
nor U15770 (N_15770,N_14897,N_14969);
nor U15771 (N_15771,N_14709,N_14622);
and U15772 (N_15772,N_14758,N_14498);
xnor U15773 (N_15773,N_14817,N_14529);
and U15774 (N_15774,N_14687,N_14897);
xor U15775 (N_15775,N_14489,N_14789);
nand U15776 (N_15776,N_15196,N_14703);
or U15777 (N_15777,N_15109,N_14466);
xnor U15778 (N_15778,N_14671,N_14849);
nand U15779 (N_15779,N_14451,N_15188);
or U15780 (N_15780,N_14677,N_14626);
xor U15781 (N_15781,N_15190,N_15010);
or U15782 (N_15782,N_14471,N_14445);
nor U15783 (N_15783,N_14438,N_14708);
nor U15784 (N_15784,N_14772,N_14505);
and U15785 (N_15785,N_14507,N_14790);
or U15786 (N_15786,N_14540,N_14715);
nor U15787 (N_15787,N_15079,N_14981);
nand U15788 (N_15788,N_14545,N_14460);
xnor U15789 (N_15789,N_15180,N_14457);
nor U15790 (N_15790,N_15164,N_14888);
xnor U15791 (N_15791,N_14648,N_14517);
and U15792 (N_15792,N_14907,N_14962);
or U15793 (N_15793,N_14803,N_14995);
nor U15794 (N_15794,N_15075,N_14472);
xnor U15795 (N_15795,N_15184,N_14873);
nand U15796 (N_15796,N_14442,N_14926);
xnor U15797 (N_15797,N_14943,N_14790);
xor U15798 (N_15798,N_14919,N_15028);
nand U15799 (N_15799,N_14636,N_14768);
or U15800 (N_15800,N_15152,N_14439);
nand U15801 (N_15801,N_14984,N_15162);
nor U15802 (N_15802,N_14597,N_14504);
nor U15803 (N_15803,N_14651,N_14564);
nand U15804 (N_15804,N_14594,N_15189);
and U15805 (N_15805,N_14619,N_14875);
or U15806 (N_15806,N_15075,N_14887);
or U15807 (N_15807,N_14628,N_14474);
nor U15808 (N_15808,N_14420,N_15012);
or U15809 (N_15809,N_14854,N_15195);
or U15810 (N_15810,N_15104,N_14405);
xnor U15811 (N_15811,N_14865,N_14405);
xnor U15812 (N_15812,N_15180,N_14723);
xor U15813 (N_15813,N_14893,N_14491);
xnor U15814 (N_15814,N_14710,N_14520);
and U15815 (N_15815,N_14542,N_15035);
and U15816 (N_15816,N_14914,N_14918);
nand U15817 (N_15817,N_14488,N_15170);
or U15818 (N_15818,N_15174,N_15093);
nand U15819 (N_15819,N_14463,N_14706);
xnor U15820 (N_15820,N_14431,N_14902);
and U15821 (N_15821,N_14950,N_15049);
nor U15822 (N_15822,N_14599,N_14555);
and U15823 (N_15823,N_14555,N_14967);
or U15824 (N_15824,N_14963,N_14644);
or U15825 (N_15825,N_14756,N_15027);
nand U15826 (N_15826,N_14681,N_14496);
xor U15827 (N_15827,N_14575,N_14999);
or U15828 (N_15828,N_14468,N_14759);
xor U15829 (N_15829,N_15007,N_14664);
xor U15830 (N_15830,N_14944,N_14994);
or U15831 (N_15831,N_14641,N_14694);
nor U15832 (N_15832,N_15083,N_14411);
xor U15833 (N_15833,N_14816,N_14636);
nand U15834 (N_15834,N_14569,N_14605);
or U15835 (N_15835,N_14440,N_15141);
nand U15836 (N_15836,N_14799,N_14552);
or U15837 (N_15837,N_15071,N_14749);
nor U15838 (N_15838,N_14514,N_14889);
xnor U15839 (N_15839,N_14733,N_14582);
or U15840 (N_15840,N_14901,N_14946);
xnor U15841 (N_15841,N_14986,N_14594);
nand U15842 (N_15842,N_14662,N_14819);
nor U15843 (N_15843,N_14875,N_14506);
xor U15844 (N_15844,N_14954,N_14507);
xnor U15845 (N_15845,N_15103,N_14777);
and U15846 (N_15846,N_14631,N_15077);
nand U15847 (N_15847,N_15169,N_14904);
and U15848 (N_15848,N_14807,N_15161);
or U15849 (N_15849,N_14429,N_14633);
xor U15850 (N_15850,N_14569,N_15187);
nor U15851 (N_15851,N_14596,N_15048);
nor U15852 (N_15852,N_15059,N_14740);
or U15853 (N_15853,N_14779,N_14748);
and U15854 (N_15854,N_14713,N_15052);
and U15855 (N_15855,N_15168,N_14692);
and U15856 (N_15856,N_14505,N_14483);
and U15857 (N_15857,N_15026,N_14577);
or U15858 (N_15858,N_15077,N_14914);
or U15859 (N_15859,N_14443,N_15137);
nor U15860 (N_15860,N_14656,N_14760);
nor U15861 (N_15861,N_15064,N_15142);
or U15862 (N_15862,N_14932,N_14585);
nand U15863 (N_15863,N_15096,N_15124);
nand U15864 (N_15864,N_14458,N_14677);
nand U15865 (N_15865,N_14547,N_14818);
nor U15866 (N_15866,N_14452,N_14932);
and U15867 (N_15867,N_14871,N_15059);
xnor U15868 (N_15868,N_15190,N_14819);
xor U15869 (N_15869,N_15095,N_15114);
xor U15870 (N_15870,N_14549,N_15195);
or U15871 (N_15871,N_14494,N_14456);
nand U15872 (N_15872,N_14902,N_14770);
nor U15873 (N_15873,N_14680,N_14442);
nor U15874 (N_15874,N_14668,N_15018);
nor U15875 (N_15875,N_14405,N_14462);
and U15876 (N_15876,N_14693,N_15100);
nand U15877 (N_15877,N_14845,N_14599);
or U15878 (N_15878,N_14771,N_14520);
and U15879 (N_15879,N_14529,N_14813);
or U15880 (N_15880,N_14449,N_15185);
or U15881 (N_15881,N_14806,N_14857);
xnor U15882 (N_15882,N_15159,N_15054);
and U15883 (N_15883,N_15048,N_14878);
and U15884 (N_15884,N_14767,N_14788);
and U15885 (N_15885,N_14677,N_14850);
xnor U15886 (N_15886,N_14812,N_14546);
or U15887 (N_15887,N_14591,N_14589);
nor U15888 (N_15888,N_15121,N_14429);
nand U15889 (N_15889,N_14990,N_15148);
and U15890 (N_15890,N_15156,N_14839);
nand U15891 (N_15891,N_15123,N_14799);
nor U15892 (N_15892,N_14619,N_14568);
xor U15893 (N_15893,N_14710,N_14609);
or U15894 (N_15894,N_15171,N_14795);
nor U15895 (N_15895,N_14980,N_15062);
nor U15896 (N_15896,N_14829,N_15052);
or U15897 (N_15897,N_14976,N_14498);
nor U15898 (N_15898,N_15133,N_15113);
and U15899 (N_15899,N_14791,N_15038);
and U15900 (N_15900,N_14641,N_14665);
and U15901 (N_15901,N_14953,N_14829);
nor U15902 (N_15902,N_14620,N_14495);
or U15903 (N_15903,N_14426,N_14858);
xnor U15904 (N_15904,N_14613,N_15199);
xnor U15905 (N_15905,N_14439,N_15143);
xnor U15906 (N_15906,N_14775,N_14738);
nor U15907 (N_15907,N_14707,N_14805);
and U15908 (N_15908,N_15081,N_14815);
xnor U15909 (N_15909,N_14828,N_14506);
xor U15910 (N_15910,N_14855,N_14596);
nand U15911 (N_15911,N_14940,N_14696);
nand U15912 (N_15912,N_14925,N_15103);
or U15913 (N_15913,N_14797,N_14600);
or U15914 (N_15914,N_15093,N_15158);
and U15915 (N_15915,N_14520,N_14624);
or U15916 (N_15916,N_14552,N_14834);
xor U15917 (N_15917,N_14469,N_15176);
nor U15918 (N_15918,N_14763,N_15020);
nor U15919 (N_15919,N_15016,N_15003);
or U15920 (N_15920,N_14921,N_14752);
nand U15921 (N_15921,N_14768,N_15042);
and U15922 (N_15922,N_14527,N_14480);
and U15923 (N_15923,N_14997,N_14467);
xnor U15924 (N_15924,N_14455,N_15064);
and U15925 (N_15925,N_14960,N_14739);
and U15926 (N_15926,N_15174,N_15064);
xor U15927 (N_15927,N_15056,N_14982);
or U15928 (N_15928,N_14745,N_14441);
nand U15929 (N_15929,N_14473,N_14959);
or U15930 (N_15930,N_14628,N_15135);
and U15931 (N_15931,N_14975,N_14731);
xor U15932 (N_15932,N_14682,N_14586);
nand U15933 (N_15933,N_14820,N_14861);
and U15934 (N_15934,N_14460,N_15067);
xnor U15935 (N_15935,N_15014,N_14709);
nand U15936 (N_15936,N_14509,N_14871);
xnor U15937 (N_15937,N_14780,N_14463);
or U15938 (N_15938,N_14653,N_15015);
nor U15939 (N_15939,N_14836,N_15185);
and U15940 (N_15940,N_14860,N_14449);
xor U15941 (N_15941,N_15139,N_14938);
and U15942 (N_15942,N_14957,N_14413);
and U15943 (N_15943,N_14852,N_14565);
nor U15944 (N_15944,N_14524,N_14818);
nor U15945 (N_15945,N_14555,N_14402);
nor U15946 (N_15946,N_14623,N_14746);
xor U15947 (N_15947,N_14871,N_14500);
or U15948 (N_15948,N_14408,N_15017);
nand U15949 (N_15949,N_15003,N_14415);
and U15950 (N_15950,N_14987,N_15077);
or U15951 (N_15951,N_15163,N_14447);
xnor U15952 (N_15952,N_14838,N_14624);
or U15953 (N_15953,N_14898,N_15026);
or U15954 (N_15954,N_14684,N_14450);
and U15955 (N_15955,N_14571,N_14656);
nor U15956 (N_15956,N_14922,N_14536);
nor U15957 (N_15957,N_14616,N_14506);
xor U15958 (N_15958,N_15075,N_14810);
and U15959 (N_15959,N_14885,N_14675);
nand U15960 (N_15960,N_14522,N_15080);
nor U15961 (N_15961,N_14453,N_14749);
nand U15962 (N_15962,N_15170,N_14608);
nor U15963 (N_15963,N_14792,N_15157);
xor U15964 (N_15964,N_14785,N_15150);
nand U15965 (N_15965,N_15172,N_14420);
and U15966 (N_15966,N_14648,N_14695);
xnor U15967 (N_15967,N_14614,N_15143);
nor U15968 (N_15968,N_15078,N_15001);
or U15969 (N_15969,N_14664,N_14448);
nor U15970 (N_15970,N_14692,N_14913);
and U15971 (N_15971,N_14941,N_14932);
nand U15972 (N_15972,N_14511,N_14622);
and U15973 (N_15973,N_15010,N_15172);
nor U15974 (N_15974,N_14443,N_14743);
or U15975 (N_15975,N_15018,N_14678);
nor U15976 (N_15976,N_14954,N_14823);
or U15977 (N_15977,N_15080,N_15021);
nor U15978 (N_15978,N_14663,N_14501);
xor U15979 (N_15979,N_14824,N_14763);
xor U15980 (N_15980,N_14510,N_14957);
nand U15981 (N_15981,N_14900,N_14723);
and U15982 (N_15982,N_14467,N_14424);
xnor U15983 (N_15983,N_14854,N_14875);
nor U15984 (N_15984,N_15159,N_15085);
nor U15985 (N_15985,N_14979,N_14653);
xor U15986 (N_15986,N_14529,N_15149);
xor U15987 (N_15987,N_15070,N_14413);
or U15988 (N_15988,N_15095,N_14875);
xor U15989 (N_15989,N_14831,N_14629);
nand U15990 (N_15990,N_15128,N_15172);
and U15991 (N_15991,N_14830,N_14805);
nor U15992 (N_15992,N_14784,N_14747);
nand U15993 (N_15993,N_14822,N_14869);
xnor U15994 (N_15994,N_15165,N_14980);
and U15995 (N_15995,N_14622,N_14899);
nor U15996 (N_15996,N_14634,N_15087);
nor U15997 (N_15997,N_15186,N_15195);
nand U15998 (N_15998,N_14515,N_15098);
xnor U15999 (N_15999,N_14727,N_14459);
xor U16000 (N_16000,N_15812,N_15737);
xor U16001 (N_16001,N_15919,N_15430);
nand U16002 (N_16002,N_15247,N_15718);
nand U16003 (N_16003,N_15921,N_15957);
xor U16004 (N_16004,N_15696,N_15372);
xor U16005 (N_16005,N_15707,N_15551);
nor U16006 (N_16006,N_15776,N_15735);
and U16007 (N_16007,N_15463,N_15782);
nand U16008 (N_16008,N_15554,N_15779);
xnor U16009 (N_16009,N_15308,N_15645);
or U16010 (N_16010,N_15964,N_15224);
nand U16011 (N_16011,N_15392,N_15997);
nand U16012 (N_16012,N_15436,N_15828);
xor U16013 (N_16013,N_15950,N_15503);
xor U16014 (N_16014,N_15780,N_15486);
or U16015 (N_16015,N_15998,N_15675);
nor U16016 (N_16016,N_15913,N_15429);
nand U16017 (N_16017,N_15709,N_15716);
and U16018 (N_16018,N_15906,N_15861);
nor U16019 (N_16019,N_15646,N_15752);
nand U16020 (N_16020,N_15984,N_15565);
or U16021 (N_16021,N_15351,N_15695);
or U16022 (N_16022,N_15830,N_15663);
nor U16023 (N_16023,N_15910,N_15664);
or U16024 (N_16024,N_15961,N_15320);
or U16025 (N_16025,N_15443,N_15728);
or U16026 (N_16026,N_15697,N_15536);
xor U16027 (N_16027,N_15840,N_15317);
xnor U16028 (N_16028,N_15264,N_15286);
or U16029 (N_16029,N_15537,N_15237);
nor U16030 (N_16030,N_15983,N_15544);
nand U16031 (N_16031,N_15454,N_15660);
nand U16032 (N_16032,N_15492,N_15472);
nand U16033 (N_16033,N_15666,N_15580);
or U16034 (N_16034,N_15754,N_15974);
xor U16035 (N_16035,N_15755,N_15494);
xor U16036 (N_16036,N_15952,N_15771);
nor U16037 (N_16037,N_15969,N_15647);
and U16038 (N_16038,N_15889,N_15618);
and U16039 (N_16039,N_15588,N_15342);
nand U16040 (N_16040,N_15956,N_15393);
or U16041 (N_16041,N_15879,N_15719);
or U16042 (N_16042,N_15382,N_15437);
xor U16043 (N_16043,N_15468,N_15909);
xor U16044 (N_16044,N_15446,N_15493);
nor U16045 (N_16045,N_15201,N_15469);
nor U16046 (N_16046,N_15642,N_15212);
and U16047 (N_16047,N_15219,N_15733);
nand U16048 (N_16048,N_15221,N_15427);
or U16049 (N_16049,N_15641,N_15778);
nor U16050 (N_16050,N_15947,N_15692);
and U16051 (N_16051,N_15586,N_15401);
xor U16052 (N_16052,N_15291,N_15757);
and U16053 (N_16053,N_15941,N_15262);
nor U16054 (N_16054,N_15614,N_15784);
nor U16055 (N_16055,N_15684,N_15220);
or U16056 (N_16056,N_15287,N_15775);
xnor U16057 (N_16057,N_15357,N_15633);
nor U16058 (N_16058,N_15585,N_15441);
nor U16059 (N_16059,N_15727,N_15943);
and U16060 (N_16060,N_15456,N_15734);
nor U16061 (N_16061,N_15878,N_15333);
nand U16062 (N_16062,N_15922,N_15994);
xor U16063 (N_16063,N_15520,N_15243);
and U16064 (N_16064,N_15606,N_15611);
nor U16065 (N_16065,N_15496,N_15751);
and U16066 (N_16066,N_15768,N_15602);
nand U16067 (N_16067,N_15990,N_15408);
xnor U16068 (N_16068,N_15944,N_15704);
or U16069 (N_16069,N_15873,N_15999);
and U16070 (N_16070,N_15439,N_15501);
nor U16071 (N_16071,N_15271,N_15434);
nor U16072 (N_16072,N_15604,N_15412);
or U16073 (N_16073,N_15265,N_15304);
xor U16074 (N_16074,N_15447,N_15289);
nor U16075 (N_16075,N_15555,N_15253);
and U16076 (N_16076,N_15531,N_15756);
and U16077 (N_16077,N_15808,N_15968);
and U16078 (N_16078,N_15859,N_15980);
or U16079 (N_16079,N_15814,N_15419);
nor U16080 (N_16080,N_15825,N_15672);
nand U16081 (N_16081,N_15698,N_15506);
xnor U16082 (N_16082,N_15683,N_15821);
nand U16083 (N_16083,N_15407,N_15440);
and U16084 (N_16084,N_15266,N_15911);
nand U16085 (N_16085,N_15785,N_15575);
xnor U16086 (N_16086,N_15661,N_15938);
xnor U16087 (N_16087,N_15970,N_15834);
nand U16088 (N_16088,N_15538,N_15526);
xnor U16089 (N_16089,N_15530,N_15324);
and U16090 (N_16090,N_15789,N_15953);
and U16091 (N_16091,N_15724,N_15206);
xor U16092 (N_16092,N_15484,N_15368);
nor U16093 (N_16093,N_15837,N_15209);
or U16094 (N_16094,N_15644,N_15676);
and U16095 (N_16095,N_15359,N_15904);
xnor U16096 (N_16096,N_15578,N_15256);
xnor U16097 (N_16097,N_15244,N_15232);
nand U16098 (N_16098,N_15270,N_15850);
nand U16099 (N_16099,N_15200,N_15745);
and U16100 (N_16100,N_15406,N_15903);
nand U16101 (N_16101,N_15819,N_15722);
nand U16102 (N_16102,N_15485,N_15205);
nand U16103 (N_16103,N_15268,N_15818);
xnor U16104 (N_16104,N_15653,N_15912);
xnor U16105 (N_16105,N_15361,N_15620);
or U16106 (N_16106,N_15582,N_15590);
or U16107 (N_16107,N_15499,N_15791);
nor U16108 (N_16108,N_15862,N_15467);
nand U16109 (N_16109,N_15344,N_15307);
and U16110 (N_16110,N_15940,N_15433);
nand U16111 (N_16111,N_15713,N_15502);
or U16112 (N_16112,N_15313,N_15881);
or U16113 (N_16113,N_15420,N_15561);
xor U16114 (N_16114,N_15240,N_15272);
xor U16115 (N_16115,N_15549,N_15885);
or U16116 (N_16116,N_15422,N_15869);
or U16117 (N_16117,N_15556,N_15758);
xor U16118 (N_16118,N_15616,N_15852);
nor U16119 (N_16119,N_15309,N_15798);
and U16120 (N_16120,N_15741,N_15431);
or U16121 (N_16121,N_15648,N_15464);
or U16122 (N_16122,N_15444,N_15915);
or U16123 (N_16123,N_15607,N_15892);
or U16124 (N_16124,N_15388,N_15877);
xor U16125 (N_16125,N_15826,N_15452);
xnor U16126 (N_16126,N_15673,N_15358);
xor U16127 (N_16127,N_15680,N_15482);
nor U16128 (N_16128,N_15227,N_15690);
and U16129 (N_16129,N_15278,N_15528);
or U16130 (N_16130,N_15742,N_15617);
nand U16131 (N_16131,N_15517,N_15928);
nor U16132 (N_16132,N_15868,N_15667);
or U16133 (N_16133,N_15935,N_15887);
or U16134 (N_16134,N_15914,N_15274);
nor U16135 (N_16135,N_15306,N_15593);
nand U16136 (N_16136,N_15527,N_15460);
nor U16137 (N_16137,N_15213,N_15383);
xor U16138 (N_16138,N_15851,N_15962);
nor U16139 (N_16139,N_15612,N_15959);
nand U16140 (N_16140,N_15466,N_15626);
or U16141 (N_16141,N_15632,N_15438);
or U16142 (N_16142,N_15366,N_15736);
nand U16143 (N_16143,N_15708,N_15966);
and U16144 (N_16144,N_15332,N_15677);
nor U16145 (N_16145,N_15609,N_15546);
nor U16146 (N_16146,N_15700,N_15410);
and U16147 (N_16147,N_15277,N_15954);
nand U16148 (N_16148,N_15965,N_15613);
nand U16149 (N_16149,N_15678,N_15988);
nand U16150 (N_16150,N_15896,N_15652);
nand U16151 (N_16151,N_15615,N_15839);
and U16152 (N_16152,N_15318,N_15490);
nor U16153 (N_16153,N_15781,N_15703);
or U16154 (N_16154,N_15263,N_15524);
and U16155 (N_16155,N_15302,N_15594);
xor U16156 (N_16156,N_15374,N_15231);
xnor U16157 (N_16157,N_15934,N_15848);
xnor U16158 (N_16158,N_15867,N_15218);
or U16159 (N_16159,N_15883,N_15638);
nor U16160 (N_16160,N_15793,N_15573);
nor U16161 (N_16161,N_15960,N_15258);
nand U16162 (N_16162,N_15557,N_15403);
and U16163 (N_16163,N_15480,N_15809);
nor U16164 (N_16164,N_15453,N_15654);
nand U16165 (N_16165,N_15399,N_15242);
nand U16166 (N_16166,N_15346,N_15764);
xor U16167 (N_16167,N_15416,N_15689);
and U16168 (N_16168,N_15587,N_15846);
xor U16169 (N_16169,N_15627,N_15509);
and U16170 (N_16170,N_15283,N_15259);
and U16171 (N_16171,N_15976,N_15827);
nand U16172 (N_16172,N_15280,N_15777);
or U16173 (N_16173,N_15624,N_15991);
or U16174 (N_16174,N_15423,N_15982);
or U16175 (N_16175,N_15856,N_15884);
or U16176 (N_16176,N_15920,N_15621);
nor U16177 (N_16177,N_15478,N_15523);
and U16178 (N_16178,N_15699,N_15569);
xnor U16179 (N_16179,N_15577,N_15933);
nor U16180 (N_16180,N_15479,N_15323);
and U16181 (N_16181,N_15335,N_15369);
nand U16182 (N_16182,N_15898,N_15766);
xnor U16183 (N_16183,N_15595,N_15842);
nand U16184 (N_16184,N_15891,N_15375);
and U16185 (N_16185,N_15749,N_15600);
and U16186 (N_16186,N_15865,N_15712);
xor U16187 (N_16187,N_15360,N_15445);
xor U16188 (N_16188,N_15636,N_15629);
or U16189 (N_16189,N_15761,N_15596);
xor U16190 (N_16190,N_15763,N_15316);
nand U16191 (N_16191,N_15269,N_15210);
nor U16192 (N_16192,N_15448,N_15251);
nor U16193 (N_16193,N_15487,N_15669);
and U16194 (N_16194,N_15236,N_15583);
or U16195 (N_16195,N_15515,N_15246);
nand U16196 (N_16196,N_15658,N_15461);
nand U16197 (N_16197,N_15414,N_15550);
xnor U16198 (N_16198,N_15514,N_15900);
nor U16199 (N_16199,N_15744,N_15477);
or U16200 (N_16200,N_15475,N_15305);
nand U16201 (N_16201,N_15923,N_15245);
xnor U16202 (N_16202,N_15671,N_15339);
and U16203 (N_16203,N_15370,N_15738);
nor U16204 (N_16204,N_15533,N_15989);
or U16205 (N_16205,N_15455,N_15384);
and U16206 (N_16206,N_15872,N_15288);
or U16207 (N_16207,N_15207,N_15936);
xor U16208 (N_16208,N_15396,N_15813);
and U16209 (N_16209,N_15760,N_15349);
nand U16210 (N_16210,N_15405,N_15917);
and U16211 (N_16211,N_15519,N_15435);
xnor U16212 (N_16212,N_15820,N_15238);
or U16213 (N_16213,N_15599,N_15378);
and U16214 (N_16214,N_15275,N_15740);
nor U16215 (N_16215,N_15888,N_15597);
and U16216 (N_16216,N_15343,N_15285);
nor U16217 (N_16217,N_15681,N_15985);
nor U16218 (N_16218,N_15327,N_15823);
and U16219 (N_16219,N_15376,N_15838);
nor U16220 (N_16220,N_15806,N_15413);
nor U16221 (N_16221,N_15832,N_15432);
and U16222 (N_16222,N_15276,N_15390);
and U16223 (N_16223,N_15576,N_15298);
nor U16224 (N_16224,N_15686,N_15824);
or U16225 (N_16225,N_15829,N_15816);
xnor U16226 (N_16226,N_15350,N_15539);
or U16227 (N_16227,N_15987,N_15901);
and U16228 (N_16228,N_15810,N_15303);
nor U16229 (N_16229,N_15337,N_15817);
nand U16230 (N_16230,N_15908,N_15552);
nor U16231 (N_16231,N_15833,N_15299);
xnor U16232 (N_16232,N_15721,N_15656);
xor U16233 (N_16233,N_15581,N_15949);
and U16234 (N_16234,N_15657,N_15292);
nor U16235 (N_16235,N_15665,N_15717);
nand U16236 (N_16236,N_15640,N_15541);
xnor U16237 (N_16237,N_15296,N_15800);
xnor U16238 (N_16238,N_15579,N_15705);
nor U16239 (N_16239,N_15971,N_15822);
nand U16240 (N_16240,N_15866,N_15326);
or U16241 (N_16241,N_15702,N_15710);
and U16242 (N_16242,N_15572,N_15267);
xor U16243 (N_16243,N_15425,N_15542);
nor U16244 (N_16244,N_15845,N_15886);
and U16245 (N_16245,N_15659,N_15458);
and U16246 (N_16246,N_15400,N_15668);
nand U16247 (N_16247,N_15202,N_15608);
nor U16248 (N_16248,N_15398,N_15226);
nand U16249 (N_16249,N_15417,N_15418);
and U16250 (N_16250,N_15863,N_15591);
and U16251 (N_16251,N_15568,N_15574);
nand U16252 (N_16252,N_15694,N_15945);
or U16253 (N_16253,N_15281,N_15409);
nand U16254 (N_16254,N_15795,N_15312);
and U16255 (N_16255,N_15516,N_15907);
nand U16256 (N_16256,N_15228,N_15282);
nand U16257 (N_16257,N_15518,N_15507);
or U16258 (N_16258,N_15729,N_15662);
nor U16259 (N_16259,N_15619,N_15635);
xnor U16260 (N_16260,N_15521,N_15948);
nand U16261 (N_16261,N_15489,N_15926);
and U16262 (N_16262,N_15462,N_15540);
nand U16263 (N_16263,N_15381,N_15630);
nor U16264 (N_16264,N_15679,N_15715);
nor U16265 (N_16265,N_15796,N_15973);
nand U16266 (N_16266,N_15746,N_15890);
or U16267 (N_16267,N_15774,N_15876);
and U16268 (N_16268,N_15849,N_15495);
and U16269 (N_16269,N_15559,N_15924);
nand U16270 (N_16270,N_15547,N_15799);
and U16271 (N_16271,N_15241,N_15753);
xor U16272 (N_16272,N_15750,N_15261);
nor U16273 (N_16273,N_15670,N_15229);
xor U16274 (N_16274,N_15655,N_15972);
xor U16275 (N_16275,N_15854,N_15598);
and U16276 (N_16276,N_15545,N_15639);
and U16277 (N_16277,N_15726,N_15603);
xor U16278 (N_16278,N_15319,N_15643);
or U16279 (N_16279,N_15631,N_15504);
or U16280 (N_16280,N_15297,N_15880);
nand U16281 (N_16281,N_15955,N_15421);
xnor U16282 (N_16282,N_15254,N_15720);
xnor U16283 (N_16283,N_15584,N_15217);
nor U16284 (N_16284,N_15293,N_15558);
and U16285 (N_16285,N_15794,N_15273);
nand U16286 (N_16286,N_15805,N_15882);
nand U16287 (N_16287,N_15442,N_15931);
nand U16288 (N_16288,N_15875,N_15605);
and U16289 (N_16289,N_15225,N_15993);
nand U16290 (N_16290,N_15279,N_15404);
and U16291 (N_16291,N_15893,N_15512);
and U16292 (N_16292,N_15844,N_15963);
xor U16293 (N_16293,N_15711,N_15772);
and U16294 (N_16294,N_15853,N_15930);
nand U16295 (N_16295,N_15802,N_15723);
nand U16296 (N_16296,N_15451,N_15394);
and U16297 (N_16297,N_15870,N_15356);
or U16298 (N_16298,N_15211,N_15767);
or U16299 (N_16299,N_15701,N_15379);
or U16300 (N_16300,N_15341,N_15770);
xnor U16301 (N_16301,N_15248,N_15411);
xnor U16302 (N_16302,N_15769,N_15927);
nor U16303 (N_16303,N_15731,N_15459);
and U16304 (N_16304,N_15601,N_15322);
nand U16305 (N_16305,N_15216,N_15743);
and U16306 (N_16306,N_15294,N_15730);
xnor U16307 (N_16307,N_15874,N_15649);
nor U16308 (N_16308,N_15801,N_15249);
xor U16309 (N_16309,N_15855,N_15996);
and U16310 (N_16310,N_15622,N_15364);
nand U16311 (N_16311,N_15363,N_15929);
nor U16312 (N_16312,N_15786,N_15858);
and U16313 (N_16313,N_15942,N_15651);
and U16314 (N_16314,N_15300,N_15811);
or U16315 (N_16315,N_15290,N_15831);
nand U16316 (N_16316,N_15566,N_15570);
and U16317 (N_16317,N_15470,N_15567);
xnor U16318 (N_16318,N_15491,N_15977);
and U16319 (N_16319,N_15932,N_15498);
xnor U16320 (N_16320,N_15804,N_15380);
nor U16321 (N_16321,N_15894,N_15706);
nor U16322 (N_16322,N_15311,N_15522);
nand U16323 (N_16323,N_15525,N_15748);
xor U16324 (N_16324,N_15321,N_15951);
and U16325 (N_16325,N_15691,N_15223);
nand U16326 (N_16326,N_15967,N_15562);
nand U16327 (N_16327,N_15807,N_15783);
nor U16328 (N_16328,N_15937,N_15239);
or U16329 (N_16329,N_15532,N_15687);
or U16330 (N_16330,N_15714,N_15402);
or U16331 (N_16331,N_15208,N_15508);
nand U16332 (N_16332,N_15843,N_15995);
xnor U16333 (N_16333,N_15510,N_15214);
nand U16334 (N_16334,N_15387,N_15428);
nand U16335 (N_16335,N_15847,N_15513);
and U16336 (N_16336,N_15314,N_15835);
or U16337 (N_16337,N_15571,N_15362);
or U16338 (N_16338,N_15230,N_15773);
nor U16339 (N_16339,N_15203,N_15331);
or U16340 (N_16340,N_15986,N_15497);
nand U16341 (N_16341,N_15978,N_15233);
or U16342 (N_16342,N_15592,N_15788);
nand U16343 (N_16343,N_15899,N_15992);
xor U16344 (N_16344,N_15365,N_15330);
nor U16345 (N_16345,N_15946,N_15347);
xnor U16346 (N_16346,N_15257,N_15348);
xor U16347 (N_16347,N_15389,N_15476);
and U16348 (N_16348,N_15553,N_15471);
or U16349 (N_16349,N_15204,N_15762);
nand U16350 (N_16350,N_15255,N_15338);
or U16351 (N_16351,N_15385,N_15415);
nand U16352 (N_16352,N_15688,N_15563);
xnor U16353 (N_16353,N_15589,N_15377);
xnor U16354 (N_16354,N_15979,N_15905);
or U16355 (N_16355,N_15395,N_15939);
nand U16356 (N_16356,N_15450,N_15260);
xnor U16357 (N_16357,N_15397,N_15925);
or U16358 (N_16358,N_15215,N_15222);
or U16359 (N_16359,N_15747,N_15765);
nand U16360 (N_16360,N_15465,N_15836);
nor U16361 (N_16361,N_15329,N_15474);
or U16362 (N_16362,N_15250,N_15871);
and U16363 (N_16363,N_15483,N_15739);
or U16364 (N_16364,N_15334,N_15386);
nor U16365 (N_16365,N_15328,N_15543);
nor U16366 (N_16366,N_15902,N_15426);
xnor U16367 (N_16367,N_15481,N_15352);
xor U16368 (N_16368,N_15916,N_15958);
nor U16369 (N_16369,N_15505,N_15535);
nor U16370 (N_16370,N_15864,N_15560);
nor U16371 (N_16371,N_15449,N_15367);
nand U16372 (N_16372,N_15860,N_15628);
xnor U16373 (N_16373,N_15548,N_15803);
or U16374 (N_16374,N_15529,N_15975);
or U16375 (N_16375,N_15564,N_15340);
nor U16376 (N_16376,N_15295,N_15792);
and U16377 (N_16377,N_15787,N_15354);
xor U16378 (N_16378,N_15895,N_15918);
nand U16379 (N_16379,N_15610,N_15345);
xnor U16380 (N_16380,N_15815,N_15897);
and U16381 (N_16381,N_15693,N_15790);
or U16382 (N_16382,N_15650,N_15682);
or U16383 (N_16383,N_15424,N_15284);
or U16384 (N_16384,N_15685,N_15797);
nand U16385 (N_16385,N_15637,N_15732);
or U16386 (N_16386,N_15981,N_15235);
and U16387 (N_16387,N_15373,N_15234);
nor U16388 (N_16388,N_15634,N_15625);
xnor U16389 (N_16389,N_15355,N_15315);
and U16390 (N_16390,N_15371,N_15857);
or U16391 (N_16391,N_15301,N_15511);
or U16392 (N_16392,N_15759,N_15674);
nand U16393 (N_16393,N_15488,N_15534);
nor U16394 (N_16394,N_15500,N_15252);
nor U16395 (N_16395,N_15457,N_15391);
nor U16396 (N_16396,N_15725,N_15841);
or U16397 (N_16397,N_15473,N_15353);
or U16398 (N_16398,N_15310,N_15336);
nor U16399 (N_16399,N_15325,N_15623);
nand U16400 (N_16400,N_15989,N_15387);
xor U16401 (N_16401,N_15566,N_15310);
or U16402 (N_16402,N_15445,N_15230);
nand U16403 (N_16403,N_15964,N_15557);
nand U16404 (N_16404,N_15855,N_15704);
or U16405 (N_16405,N_15705,N_15856);
and U16406 (N_16406,N_15380,N_15746);
xor U16407 (N_16407,N_15528,N_15252);
xor U16408 (N_16408,N_15605,N_15640);
and U16409 (N_16409,N_15396,N_15508);
and U16410 (N_16410,N_15785,N_15293);
xor U16411 (N_16411,N_15260,N_15959);
xor U16412 (N_16412,N_15982,N_15587);
nor U16413 (N_16413,N_15852,N_15518);
nor U16414 (N_16414,N_15302,N_15261);
xor U16415 (N_16415,N_15384,N_15268);
xnor U16416 (N_16416,N_15867,N_15285);
nor U16417 (N_16417,N_15726,N_15652);
and U16418 (N_16418,N_15980,N_15941);
or U16419 (N_16419,N_15280,N_15562);
nor U16420 (N_16420,N_15216,N_15720);
xor U16421 (N_16421,N_15789,N_15410);
or U16422 (N_16422,N_15323,N_15305);
and U16423 (N_16423,N_15311,N_15647);
and U16424 (N_16424,N_15519,N_15351);
xor U16425 (N_16425,N_15840,N_15906);
xnor U16426 (N_16426,N_15536,N_15701);
nand U16427 (N_16427,N_15502,N_15617);
or U16428 (N_16428,N_15811,N_15640);
nand U16429 (N_16429,N_15374,N_15423);
nor U16430 (N_16430,N_15794,N_15315);
xor U16431 (N_16431,N_15798,N_15479);
xnor U16432 (N_16432,N_15581,N_15259);
xnor U16433 (N_16433,N_15544,N_15539);
or U16434 (N_16434,N_15959,N_15261);
nor U16435 (N_16435,N_15874,N_15861);
nor U16436 (N_16436,N_15335,N_15959);
or U16437 (N_16437,N_15425,N_15806);
and U16438 (N_16438,N_15790,N_15980);
or U16439 (N_16439,N_15848,N_15581);
nor U16440 (N_16440,N_15849,N_15804);
or U16441 (N_16441,N_15589,N_15663);
xnor U16442 (N_16442,N_15714,N_15593);
or U16443 (N_16443,N_15433,N_15252);
xnor U16444 (N_16444,N_15478,N_15706);
or U16445 (N_16445,N_15912,N_15490);
nor U16446 (N_16446,N_15869,N_15867);
nand U16447 (N_16447,N_15640,N_15841);
nor U16448 (N_16448,N_15380,N_15743);
nor U16449 (N_16449,N_15570,N_15652);
and U16450 (N_16450,N_15674,N_15244);
and U16451 (N_16451,N_15252,N_15915);
nor U16452 (N_16452,N_15673,N_15992);
nand U16453 (N_16453,N_15481,N_15750);
nand U16454 (N_16454,N_15829,N_15571);
and U16455 (N_16455,N_15435,N_15516);
nand U16456 (N_16456,N_15706,N_15933);
and U16457 (N_16457,N_15738,N_15667);
nand U16458 (N_16458,N_15780,N_15280);
or U16459 (N_16459,N_15608,N_15270);
or U16460 (N_16460,N_15270,N_15898);
xnor U16461 (N_16461,N_15568,N_15304);
nand U16462 (N_16462,N_15613,N_15914);
xnor U16463 (N_16463,N_15980,N_15279);
nand U16464 (N_16464,N_15952,N_15767);
and U16465 (N_16465,N_15287,N_15352);
xor U16466 (N_16466,N_15948,N_15540);
nor U16467 (N_16467,N_15834,N_15659);
and U16468 (N_16468,N_15225,N_15387);
and U16469 (N_16469,N_15620,N_15463);
or U16470 (N_16470,N_15877,N_15369);
and U16471 (N_16471,N_15445,N_15762);
or U16472 (N_16472,N_15976,N_15457);
and U16473 (N_16473,N_15431,N_15567);
and U16474 (N_16474,N_15460,N_15452);
nor U16475 (N_16475,N_15872,N_15300);
nor U16476 (N_16476,N_15473,N_15809);
or U16477 (N_16477,N_15441,N_15761);
nand U16478 (N_16478,N_15505,N_15876);
xnor U16479 (N_16479,N_15384,N_15986);
nand U16480 (N_16480,N_15876,N_15545);
xnor U16481 (N_16481,N_15445,N_15418);
nand U16482 (N_16482,N_15605,N_15904);
and U16483 (N_16483,N_15496,N_15752);
xor U16484 (N_16484,N_15805,N_15456);
nor U16485 (N_16485,N_15459,N_15474);
nor U16486 (N_16486,N_15742,N_15714);
nor U16487 (N_16487,N_15413,N_15519);
xor U16488 (N_16488,N_15359,N_15975);
nor U16489 (N_16489,N_15525,N_15211);
and U16490 (N_16490,N_15992,N_15368);
and U16491 (N_16491,N_15552,N_15708);
nand U16492 (N_16492,N_15503,N_15705);
or U16493 (N_16493,N_15633,N_15700);
or U16494 (N_16494,N_15202,N_15217);
xor U16495 (N_16495,N_15293,N_15793);
and U16496 (N_16496,N_15562,N_15739);
nand U16497 (N_16497,N_15671,N_15346);
or U16498 (N_16498,N_15523,N_15415);
xor U16499 (N_16499,N_15634,N_15552);
xnor U16500 (N_16500,N_15463,N_15636);
or U16501 (N_16501,N_15553,N_15265);
and U16502 (N_16502,N_15586,N_15377);
nand U16503 (N_16503,N_15639,N_15539);
xor U16504 (N_16504,N_15386,N_15519);
xnor U16505 (N_16505,N_15945,N_15206);
xnor U16506 (N_16506,N_15226,N_15990);
nand U16507 (N_16507,N_15268,N_15329);
or U16508 (N_16508,N_15311,N_15815);
nor U16509 (N_16509,N_15219,N_15346);
or U16510 (N_16510,N_15616,N_15992);
nand U16511 (N_16511,N_15339,N_15290);
or U16512 (N_16512,N_15528,N_15493);
and U16513 (N_16513,N_15876,N_15675);
nand U16514 (N_16514,N_15231,N_15607);
xor U16515 (N_16515,N_15445,N_15627);
and U16516 (N_16516,N_15716,N_15648);
xnor U16517 (N_16517,N_15412,N_15674);
and U16518 (N_16518,N_15248,N_15269);
nor U16519 (N_16519,N_15323,N_15438);
or U16520 (N_16520,N_15894,N_15651);
or U16521 (N_16521,N_15713,N_15592);
nor U16522 (N_16522,N_15971,N_15779);
nand U16523 (N_16523,N_15994,N_15529);
xnor U16524 (N_16524,N_15637,N_15251);
nor U16525 (N_16525,N_15337,N_15479);
nor U16526 (N_16526,N_15454,N_15596);
or U16527 (N_16527,N_15497,N_15924);
or U16528 (N_16528,N_15470,N_15976);
and U16529 (N_16529,N_15769,N_15591);
or U16530 (N_16530,N_15415,N_15205);
nand U16531 (N_16531,N_15501,N_15390);
or U16532 (N_16532,N_15675,N_15685);
and U16533 (N_16533,N_15538,N_15916);
and U16534 (N_16534,N_15474,N_15860);
xor U16535 (N_16535,N_15434,N_15201);
xnor U16536 (N_16536,N_15254,N_15705);
nand U16537 (N_16537,N_15515,N_15343);
xnor U16538 (N_16538,N_15602,N_15937);
or U16539 (N_16539,N_15873,N_15803);
nor U16540 (N_16540,N_15493,N_15334);
nand U16541 (N_16541,N_15813,N_15561);
nand U16542 (N_16542,N_15648,N_15801);
xor U16543 (N_16543,N_15956,N_15571);
or U16544 (N_16544,N_15561,N_15971);
or U16545 (N_16545,N_15274,N_15580);
nand U16546 (N_16546,N_15979,N_15338);
xor U16547 (N_16547,N_15625,N_15374);
nor U16548 (N_16548,N_15688,N_15705);
nor U16549 (N_16549,N_15693,N_15755);
nand U16550 (N_16550,N_15833,N_15687);
nand U16551 (N_16551,N_15596,N_15694);
and U16552 (N_16552,N_15657,N_15799);
or U16553 (N_16553,N_15966,N_15560);
and U16554 (N_16554,N_15525,N_15477);
nand U16555 (N_16555,N_15537,N_15425);
and U16556 (N_16556,N_15901,N_15898);
or U16557 (N_16557,N_15721,N_15833);
nand U16558 (N_16558,N_15912,N_15717);
or U16559 (N_16559,N_15394,N_15600);
and U16560 (N_16560,N_15430,N_15279);
nand U16561 (N_16561,N_15817,N_15530);
or U16562 (N_16562,N_15962,N_15913);
xor U16563 (N_16563,N_15307,N_15629);
and U16564 (N_16564,N_15587,N_15426);
xor U16565 (N_16565,N_15694,N_15925);
or U16566 (N_16566,N_15282,N_15532);
nand U16567 (N_16567,N_15560,N_15944);
or U16568 (N_16568,N_15464,N_15761);
and U16569 (N_16569,N_15247,N_15305);
nor U16570 (N_16570,N_15908,N_15719);
nor U16571 (N_16571,N_15831,N_15661);
nand U16572 (N_16572,N_15982,N_15403);
nand U16573 (N_16573,N_15557,N_15663);
or U16574 (N_16574,N_15478,N_15293);
nor U16575 (N_16575,N_15554,N_15257);
and U16576 (N_16576,N_15417,N_15222);
nor U16577 (N_16577,N_15419,N_15834);
nand U16578 (N_16578,N_15471,N_15607);
nand U16579 (N_16579,N_15927,N_15952);
nor U16580 (N_16580,N_15424,N_15312);
and U16581 (N_16581,N_15499,N_15492);
nand U16582 (N_16582,N_15677,N_15541);
xnor U16583 (N_16583,N_15512,N_15502);
and U16584 (N_16584,N_15805,N_15965);
and U16585 (N_16585,N_15706,N_15984);
nor U16586 (N_16586,N_15533,N_15322);
and U16587 (N_16587,N_15638,N_15201);
and U16588 (N_16588,N_15792,N_15313);
or U16589 (N_16589,N_15845,N_15521);
or U16590 (N_16590,N_15870,N_15414);
nor U16591 (N_16591,N_15409,N_15836);
nand U16592 (N_16592,N_15693,N_15329);
and U16593 (N_16593,N_15522,N_15254);
or U16594 (N_16594,N_15945,N_15938);
nand U16595 (N_16595,N_15504,N_15589);
nor U16596 (N_16596,N_15968,N_15795);
nor U16597 (N_16597,N_15534,N_15992);
nor U16598 (N_16598,N_15512,N_15830);
xnor U16599 (N_16599,N_15574,N_15263);
nor U16600 (N_16600,N_15486,N_15745);
and U16601 (N_16601,N_15612,N_15597);
and U16602 (N_16602,N_15235,N_15871);
and U16603 (N_16603,N_15312,N_15831);
and U16604 (N_16604,N_15856,N_15337);
or U16605 (N_16605,N_15638,N_15353);
xor U16606 (N_16606,N_15231,N_15780);
or U16607 (N_16607,N_15770,N_15843);
xnor U16608 (N_16608,N_15529,N_15486);
and U16609 (N_16609,N_15567,N_15981);
nor U16610 (N_16610,N_15472,N_15755);
nor U16611 (N_16611,N_15719,N_15532);
or U16612 (N_16612,N_15807,N_15752);
or U16613 (N_16613,N_15499,N_15902);
nand U16614 (N_16614,N_15942,N_15582);
xnor U16615 (N_16615,N_15737,N_15877);
and U16616 (N_16616,N_15679,N_15864);
or U16617 (N_16617,N_15780,N_15666);
and U16618 (N_16618,N_15980,N_15559);
and U16619 (N_16619,N_15685,N_15554);
nand U16620 (N_16620,N_15815,N_15955);
or U16621 (N_16621,N_15856,N_15956);
and U16622 (N_16622,N_15927,N_15832);
and U16623 (N_16623,N_15248,N_15705);
and U16624 (N_16624,N_15899,N_15687);
nand U16625 (N_16625,N_15854,N_15659);
nand U16626 (N_16626,N_15540,N_15832);
nand U16627 (N_16627,N_15414,N_15377);
nor U16628 (N_16628,N_15782,N_15200);
nand U16629 (N_16629,N_15575,N_15608);
nand U16630 (N_16630,N_15938,N_15449);
and U16631 (N_16631,N_15597,N_15801);
nor U16632 (N_16632,N_15292,N_15902);
and U16633 (N_16633,N_15231,N_15406);
nor U16634 (N_16634,N_15774,N_15293);
or U16635 (N_16635,N_15592,N_15892);
nor U16636 (N_16636,N_15594,N_15938);
and U16637 (N_16637,N_15769,N_15946);
nand U16638 (N_16638,N_15608,N_15963);
xnor U16639 (N_16639,N_15712,N_15644);
and U16640 (N_16640,N_15644,N_15657);
xor U16641 (N_16641,N_15764,N_15403);
nand U16642 (N_16642,N_15339,N_15611);
xor U16643 (N_16643,N_15852,N_15298);
or U16644 (N_16644,N_15786,N_15531);
nor U16645 (N_16645,N_15347,N_15444);
xnor U16646 (N_16646,N_15749,N_15578);
xnor U16647 (N_16647,N_15379,N_15693);
or U16648 (N_16648,N_15264,N_15998);
nor U16649 (N_16649,N_15460,N_15825);
nand U16650 (N_16650,N_15231,N_15460);
nor U16651 (N_16651,N_15757,N_15449);
nand U16652 (N_16652,N_15896,N_15494);
xor U16653 (N_16653,N_15807,N_15715);
nand U16654 (N_16654,N_15242,N_15374);
nand U16655 (N_16655,N_15751,N_15523);
nand U16656 (N_16656,N_15502,N_15462);
xor U16657 (N_16657,N_15317,N_15729);
xor U16658 (N_16658,N_15449,N_15252);
or U16659 (N_16659,N_15319,N_15636);
and U16660 (N_16660,N_15694,N_15704);
or U16661 (N_16661,N_15446,N_15222);
nor U16662 (N_16662,N_15418,N_15226);
nand U16663 (N_16663,N_15283,N_15890);
xnor U16664 (N_16664,N_15970,N_15979);
xor U16665 (N_16665,N_15749,N_15617);
and U16666 (N_16666,N_15270,N_15619);
xnor U16667 (N_16667,N_15764,N_15500);
nor U16668 (N_16668,N_15934,N_15618);
nand U16669 (N_16669,N_15239,N_15711);
nor U16670 (N_16670,N_15776,N_15762);
xor U16671 (N_16671,N_15706,N_15250);
nor U16672 (N_16672,N_15770,N_15545);
or U16673 (N_16673,N_15384,N_15252);
or U16674 (N_16674,N_15729,N_15822);
nand U16675 (N_16675,N_15210,N_15620);
or U16676 (N_16676,N_15687,N_15500);
and U16677 (N_16677,N_15600,N_15785);
xnor U16678 (N_16678,N_15324,N_15283);
xor U16679 (N_16679,N_15465,N_15371);
nand U16680 (N_16680,N_15262,N_15437);
or U16681 (N_16681,N_15730,N_15985);
nand U16682 (N_16682,N_15278,N_15500);
xor U16683 (N_16683,N_15265,N_15435);
and U16684 (N_16684,N_15974,N_15619);
xnor U16685 (N_16685,N_15441,N_15640);
xor U16686 (N_16686,N_15362,N_15910);
nor U16687 (N_16687,N_15633,N_15491);
xnor U16688 (N_16688,N_15220,N_15746);
xor U16689 (N_16689,N_15666,N_15852);
or U16690 (N_16690,N_15978,N_15924);
xnor U16691 (N_16691,N_15787,N_15393);
xnor U16692 (N_16692,N_15673,N_15540);
nor U16693 (N_16693,N_15561,N_15304);
and U16694 (N_16694,N_15271,N_15950);
or U16695 (N_16695,N_15926,N_15962);
and U16696 (N_16696,N_15370,N_15629);
and U16697 (N_16697,N_15362,N_15343);
nand U16698 (N_16698,N_15642,N_15876);
and U16699 (N_16699,N_15306,N_15734);
xor U16700 (N_16700,N_15496,N_15948);
xor U16701 (N_16701,N_15557,N_15552);
and U16702 (N_16702,N_15457,N_15961);
nand U16703 (N_16703,N_15415,N_15529);
nand U16704 (N_16704,N_15577,N_15772);
nand U16705 (N_16705,N_15981,N_15874);
nor U16706 (N_16706,N_15326,N_15802);
nor U16707 (N_16707,N_15486,N_15532);
and U16708 (N_16708,N_15262,N_15734);
and U16709 (N_16709,N_15412,N_15805);
and U16710 (N_16710,N_15372,N_15834);
or U16711 (N_16711,N_15852,N_15251);
or U16712 (N_16712,N_15776,N_15937);
nor U16713 (N_16713,N_15733,N_15640);
and U16714 (N_16714,N_15605,N_15616);
and U16715 (N_16715,N_15359,N_15502);
xnor U16716 (N_16716,N_15504,N_15888);
and U16717 (N_16717,N_15907,N_15494);
xor U16718 (N_16718,N_15384,N_15769);
xor U16719 (N_16719,N_15307,N_15259);
nor U16720 (N_16720,N_15661,N_15890);
and U16721 (N_16721,N_15485,N_15542);
or U16722 (N_16722,N_15901,N_15636);
or U16723 (N_16723,N_15343,N_15677);
xor U16724 (N_16724,N_15866,N_15729);
xor U16725 (N_16725,N_15424,N_15222);
nor U16726 (N_16726,N_15854,N_15403);
and U16727 (N_16727,N_15806,N_15695);
nor U16728 (N_16728,N_15358,N_15535);
or U16729 (N_16729,N_15509,N_15603);
nand U16730 (N_16730,N_15425,N_15212);
nor U16731 (N_16731,N_15713,N_15567);
nand U16732 (N_16732,N_15327,N_15672);
or U16733 (N_16733,N_15536,N_15715);
nor U16734 (N_16734,N_15346,N_15570);
and U16735 (N_16735,N_15950,N_15933);
or U16736 (N_16736,N_15350,N_15980);
or U16737 (N_16737,N_15394,N_15931);
and U16738 (N_16738,N_15589,N_15711);
or U16739 (N_16739,N_15786,N_15392);
nor U16740 (N_16740,N_15566,N_15728);
and U16741 (N_16741,N_15842,N_15520);
nor U16742 (N_16742,N_15740,N_15954);
and U16743 (N_16743,N_15842,N_15909);
and U16744 (N_16744,N_15920,N_15362);
nor U16745 (N_16745,N_15408,N_15894);
nand U16746 (N_16746,N_15665,N_15819);
nor U16747 (N_16747,N_15247,N_15517);
and U16748 (N_16748,N_15292,N_15238);
or U16749 (N_16749,N_15369,N_15285);
nand U16750 (N_16750,N_15271,N_15496);
nand U16751 (N_16751,N_15903,N_15350);
or U16752 (N_16752,N_15585,N_15339);
nor U16753 (N_16753,N_15718,N_15928);
nor U16754 (N_16754,N_15356,N_15767);
nor U16755 (N_16755,N_15362,N_15883);
and U16756 (N_16756,N_15936,N_15448);
xor U16757 (N_16757,N_15261,N_15390);
xnor U16758 (N_16758,N_15890,N_15699);
or U16759 (N_16759,N_15973,N_15405);
nand U16760 (N_16760,N_15209,N_15916);
or U16761 (N_16761,N_15831,N_15366);
or U16762 (N_16762,N_15360,N_15278);
nand U16763 (N_16763,N_15539,N_15661);
nand U16764 (N_16764,N_15902,N_15930);
nor U16765 (N_16765,N_15410,N_15636);
nand U16766 (N_16766,N_15221,N_15444);
nand U16767 (N_16767,N_15232,N_15523);
nand U16768 (N_16768,N_15520,N_15946);
and U16769 (N_16769,N_15349,N_15837);
xor U16770 (N_16770,N_15517,N_15471);
xnor U16771 (N_16771,N_15225,N_15648);
nor U16772 (N_16772,N_15925,N_15218);
xnor U16773 (N_16773,N_15278,N_15911);
nor U16774 (N_16774,N_15387,N_15214);
or U16775 (N_16775,N_15362,N_15340);
nor U16776 (N_16776,N_15203,N_15692);
nand U16777 (N_16777,N_15276,N_15955);
nor U16778 (N_16778,N_15786,N_15854);
xor U16779 (N_16779,N_15629,N_15696);
and U16780 (N_16780,N_15353,N_15567);
nor U16781 (N_16781,N_15760,N_15917);
or U16782 (N_16782,N_15737,N_15975);
and U16783 (N_16783,N_15355,N_15740);
nor U16784 (N_16784,N_15292,N_15544);
and U16785 (N_16785,N_15647,N_15819);
nand U16786 (N_16786,N_15707,N_15784);
and U16787 (N_16787,N_15672,N_15337);
nor U16788 (N_16788,N_15995,N_15938);
nor U16789 (N_16789,N_15779,N_15858);
xnor U16790 (N_16790,N_15774,N_15782);
or U16791 (N_16791,N_15919,N_15589);
and U16792 (N_16792,N_15264,N_15844);
xor U16793 (N_16793,N_15395,N_15232);
nor U16794 (N_16794,N_15228,N_15536);
xnor U16795 (N_16795,N_15699,N_15438);
xnor U16796 (N_16796,N_15409,N_15233);
nor U16797 (N_16797,N_15611,N_15456);
xnor U16798 (N_16798,N_15551,N_15483);
xor U16799 (N_16799,N_15296,N_15408);
xnor U16800 (N_16800,N_16688,N_16136);
nand U16801 (N_16801,N_16508,N_16782);
and U16802 (N_16802,N_16784,N_16699);
nor U16803 (N_16803,N_16029,N_16668);
nor U16804 (N_16804,N_16569,N_16428);
nor U16805 (N_16805,N_16395,N_16003);
nand U16806 (N_16806,N_16289,N_16212);
and U16807 (N_16807,N_16053,N_16337);
nor U16808 (N_16808,N_16341,N_16317);
nor U16809 (N_16809,N_16272,N_16352);
nor U16810 (N_16810,N_16601,N_16764);
nand U16811 (N_16811,N_16350,N_16041);
nand U16812 (N_16812,N_16240,N_16563);
and U16813 (N_16813,N_16293,N_16179);
nand U16814 (N_16814,N_16017,N_16780);
or U16815 (N_16815,N_16708,N_16324);
or U16816 (N_16816,N_16048,N_16438);
and U16817 (N_16817,N_16538,N_16302);
xor U16818 (N_16818,N_16333,N_16363);
or U16819 (N_16819,N_16307,N_16447);
or U16820 (N_16820,N_16451,N_16799);
and U16821 (N_16821,N_16010,N_16276);
and U16822 (N_16822,N_16222,N_16541);
and U16823 (N_16823,N_16623,N_16481);
and U16824 (N_16824,N_16000,N_16594);
and U16825 (N_16825,N_16226,N_16525);
or U16826 (N_16826,N_16374,N_16087);
or U16827 (N_16827,N_16638,N_16200);
and U16828 (N_16828,N_16116,N_16076);
and U16829 (N_16829,N_16607,N_16537);
nand U16830 (N_16830,N_16731,N_16006);
xor U16831 (N_16831,N_16439,N_16037);
or U16832 (N_16832,N_16792,N_16183);
xnor U16833 (N_16833,N_16705,N_16702);
nand U16834 (N_16834,N_16507,N_16347);
xor U16835 (N_16835,N_16646,N_16194);
xnor U16836 (N_16836,N_16298,N_16167);
xor U16837 (N_16837,N_16196,N_16191);
and U16838 (N_16838,N_16744,N_16434);
xnor U16839 (N_16839,N_16489,N_16188);
nand U16840 (N_16840,N_16463,N_16288);
nand U16841 (N_16841,N_16577,N_16295);
or U16842 (N_16842,N_16444,N_16408);
xor U16843 (N_16843,N_16404,N_16138);
and U16844 (N_16844,N_16580,N_16584);
and U16845 (N_16845,N_16506,N_16736);
nand U16846 (N_16846,N_16246,N_16096);
and U16847 (N_16847,N_16484,N_16013);
nor U16848 (N_16848,N_16218,N_16264);
xnor U16849 (N_16849,N_16645,N_16223);
nor U16850 (N_16850,N_16703,N_16588);
and U16851 (N_16851,N_16763,N_16501);
nand U16852 (N_16852,N_16460,N_16380);
or U16853 (N_16853,N_16553,N_16529);
nand U16854 (N_16854,N_16252,N_16742);
and U16855 (N_16855,N_16234,N_16099);
xor U16856 (N_16856,N_16069,N_16219);
or U16857 (N_16857,N_16431,N_16312);
nand U16858 (N_16858,N_16297,N_16393);
and U16859 (N_16859,N_16065,N_16388);
or U16860 (N_16860,N_16078,N_16409);
or U16861 (N_16861,N_16661,N_16193);
xor U16862 (N_16862,N_16083,N_16278);
and U16863 (N_16863,N_16372,N_16367);
nand U16864 (N_16864,N_16560,N_16398);
and U16865 (N_16865,N_16318,N_16261);
nand U16866 (N_16866,N_16113,N_16488);
xnor U16867 (N_16867,N_16545,N_16426);
or U16868 (N_16868,N_16187,N_16299);
nor U16869 (N_16869,N_16051,N_16137);
nor U16870 (N_16870,N_16206,N_16332);
and U16871 (N_16871,N_16168,N_16734);
and U16872 (N_16872,N_16473,N_16284);
nand U16873 (N_16873,N_16464,N_16696);
or U16874 (N_16874,N_16482,N_16542);
and U16875 (N_16875,N_16241,N_16617);
and U16876 (N_16876,N_16279,N_16233);
xnor U16877 (N_16877,N_16086,N_16568);
or U16878 (N_16878,N_16391,N_16766);
or U16879 (N_16879,N_16397,N_16211);
nand U16880 (N_16880,N_16522,N_16047);
and U16881 (N_16881,N_16762,N_16059);
xor U16882 (N_16882,N_16531,N_16121);
xnor U16883 (N_16883,N_16007,N_16752);
xnor U16884 (N_16884,N_16054,N_16477);
nor U16885 (N_16885,N_16660,N_16134);
or U16886 (N_16886,N_16157,N_16609);
and U16887 (N_16887,N_16407,N_16677);
xor U16888 (N_16888,N_16469,N_16741);
xor U16889 (N_16889,N_16496,N_16758);
nor U16890 (N_16890,N_16163,N_16214);
or U16891 (N_16891,N_16729,N_16445);
nand U16892 (N_16892,N_16493,N_16512);
xor U16893 (N_16893,N_16693,N_16564);
nand U16894 (N_16894,N_16064,N_16412);
nor U16895 (N_16895,N_16282,N_16050);
nor U16896 (N_16896,N_16449,N_16127);
and U16897 (N_16897,N_16122,N_16310);
or U16898 (N_16898,N_16622,N_16381);
and U16899 (N_16899,N_16229,N_16485);
xor U16900 (N_16900,N_16558,N_16364);
or U16901 (N_16901,N_16624,N_16796);
nand U16902 (N_16902,N_16578,N_16334);
and U16903 (N_16903,N_16572,N_16361);
nor U16904 (N_16904,N_16698,N_16798);
xor U16905 (N_16905,N_16141,N_16448);
nor U16906 (N_16906,N_16110,N_16730);
xnor U16907 (N_16907,N_16290,N_16783);
nor U16908 (N_16908,N_16416,N_16062);
and U16909 (N_16909,N_16186,N_16192);
and U16910 (N_16910,N_16033,N_16467);
nor U16911 (N_16911,N_16376,N_16719);
and U16912 (N_16912,N_16678,N_16180);
xnor U16913 (N_16913,N_16402,N_16420);
nor U16914 (N_16914,N_16414,N_16230);
and U16915 (N_16915,N_16107,N_16331);
and U16916 (N_16916,N_16461,N_16596);
nor U16917 (N_16917,N_16446,N_16396);
nor U16918 (N_16918,N_16265,N_16664);
xnor U16919 (N_16919,N_16589,N_16789);
xor U16920 (N_16920,N_16123,N_16119);
nor U16921 (N_16921,N_16144,N_16253);
xor U16922 (N_16922,N_16479,N_16270);
nand U16923 (N_16923,N_16148,N_16706);
xnor U16924 (N_16924,N_16262,N_16605);
or U16925 (N_16925,N_16384,N_16385);
xor U16926 (N_16926,N_16442,N_16018);
or U16927 (N_16927,N_16345,N_16475);
xor U16928 (N_16928,N_16557,N_16478);
nand U16929 (N_16929,N_16203,N_16044);
nand U16930 (N_16930,N_16081,N_16775);
nand U16931 (N_16931,N_16399,N_16049);
or U16932 (N_16932,N_16658,N_16314);
nor U16933 (N_16933,N_16309,N_16383);
nor U16934 (N_16934,N_16684,N_16303);
or U16935 (N_16935,N_16406,N_16453);
or U16936 (N_16936,N_16714,N_16145);
and U16937 (N_16937,N_16002,N_16514);
or U16938 (N_16938,N_16527,N_16778);
nor U16939 (N_16939,N_16436,N_16057);
xnor U16940 (N_16940,N_16389,N_16235);
nor U16941 (N_16941,N_16089,N_16510);
or U16942 (N_16942,N_16008,N_16631);
nand U16943 (N_16943,N_16074,N_16548);
and U16944 (N_16944,N_16343,N_16523);
and U16945 (N_16945,N_16286,N_16737);
or U16946 (N_16946,N_16505,N_16080);
nor U16947 (N_16947,N_16131,N_16280);
xor U16948 (N_16948,N_16190,N_16169);
or U16949 (N_16949,N_16555,N_16612);
nand U16950 (N_16950,N_16067,N_16739);
nand U16951 (N_16951,N_16338,N_16178);
and U16952 (N_16952,N_16518,N_16503);
or U16953 (N_16953,N_16418,N_16632);
nand U16954 (N_16954,N_16535,N_16019);
and U16955 (N_16955,N_16432,N_16287);
nand U16956 (N_16956,N_16735,N_16056);
xnor U16957 (N_16957,N_16774,N_16329);
xor U16958 (N_16958,N_16746,N_16728);
nor U16959 (N_16959,N_16228,N_16315);
and U16960 (N_16960,N_16327,N_16452);
or U16961 (N_16961,N_16618,N_16534);
and U16962 (N_16962,N_16466,N_16648);
nand U16963 (N_16963,N_16582,N_16680);
or U16964 (N_16964,N_16595,N_16513);
xnor U16965 (N_16965,N_16429,N_16709);
or U16966 (N_16966,N_16665,N_16704);
nand U16967 (N_16967,N_16515,N_16630);
xor U16968 (N_16968,N_16585,N_16182);
nand U16969 (N_16969,N_16567,N_16304);
nand U16970 (N_16970,N_16356,N_16625);
and U16971 (N_16971,N_16401,N_16592);
nor U16972 (N_16972,N_16245,N_16369);
xnor U16973 (N_16973,N_16691,N_16026);
or U16974 (N_16974,N_16225,N_16063);
or U16975 (N_16975,N_16035,N_16351);
xnor U16976 (N_16976,N_16022,N_16546);
xnor U16977 (N_16977,N_16779,N_16635);
nand U16978 (N_16978,N_16767,N_16727);
xor U16979 (N_16979,N_16112,N_16621);
xnor U16980 (N_16980,N_16375,N_16690);
nand U16981 (N_16981,N_16034,N_16055);
and U16982 (N_16982,N_16640,N_16599);
and U16983 (N_16983,N_16435,N_16517);
xnor U16984 (N_16984,N_16770,N_16100);
nand U16985 (N_16985,N_16636,N_16330);
and U16986 (N_16986,N_16682,N_16201);
xnor U16987 (N_16987,N_16227,N_16043);
and U16988 (N_16988,N_16647,N_16058);
nand U16989 (N_16989,N_16552,N_16177);
nand U16990 (N_16990,N_16633,N_16686);
or U16991 (N_16991,N_16405,N_16591);
xor U16992 (N_16992,N_16685,N_16726);
xor U16993 (N_16993,N_16793,N_16532);
and U16994 (N_16994,N_16346,N_16732);
nor U16995 (N_16995,N_16720,N_16143);
or U16996 (N_16996,N_16118,N_16771);
xnor U16997 (N_16997,N_16785,N_16593);
nand U16998 (N_16998,N_16755,N_16095);
and U16999 (N_16999,N_16274,N_16400);
and U17000 (N_17000,N_16387,N_16259);
xnor U17001 (N_17001,N_16313,N_16511);
or U17002 (N_17002,N_16761,N_16365);
and U17003 (N_17003,N_16751,N_16207);
xor U17004 (N_17004,N_16471,N_16075);
xnor U17005 (N_17005,N_16366,N_16738);
nand U17006 (N_17006,N_16016,N_16576);
xnor U17007 (N_17007,N_16749,N_16184);
nand U17008 (N_17008,N_16249,N_16672);
or U17009 (N_17009,N_16358,N_16114);
nand U17010 (N_17010,N_16768,N_16140);
xnor U17011 (N_17011,N_16260,N_16336);
xor U17012 (N_17012,N_16483,N_16547);
or U17013 (N_17013,N_16454,N_16011);
and U17014 (N_17014,N_16519,N_16208);
xnor U17015 (N_17015,N_16486,N_16787);
nand U17016 (N_17016,N_16325,N_16300);
nand U17017 (N_17017,N_16457,N_16390);
xnor U17018 (N_17018,N_16597,N_16025);
nor U17019 (N_17019,N_16232,N_16285);
nor U17020 (N_17020,N_16371,N_16465);
or U17021 (N_17021,N_16456,N_16125);
nor U17022 (N_17022,N_16150,N_16109);
and U17023 (N_17023,N_16348,N_16419);
nand U17024 (N_17024,N_16600,N_16701);
nor U17025 (N_17025,N_16619,N_16472);
or U17026 (N_17026,N_16574,N_16681);
or U17027 (N_17027,N_16458,N_16543);
and U17028 (N_17028,N_16236,N_16733);
and U17029 (N_17029,N_16490,N_16135);
and U17030 (N_17030,N_16052,N_16643);
xnor U17031 (N_17031,N_16476,N_16256);
nor U17032 (N_17032,N_16649,N_16676);
xor U17033 (N_17033,N_16104,N_16620);
nand U17034 (N_17034,N_16210,N_16583);
nor U17035 (N_17035,N_16171,N_16772);
or U17036 (N_17036,N_16516,N_16791);
nand U17037 (N_17037,N_16711,N_16571);
or U17038 (N_17038,N_16725,N_16561);
or U17039 (N_17039,N_16674,N_16115);
or U17040 (N_17040,N_16277,N_16021);
or U17041 (N_17041,N_16267,N_16499);
or U17042 (N_17042,N_16155,N_16743);
xnor U17043 (N_17043,N_16603,N_16213);
nor U17044 (N_17044,N_16237,N_16283);
and U17045 (N_17045,N_16394,N_16129);
xor U17046 (N_17046,N_16189,N_16386);
xor U17047 (N_17047,N_16756,N_16759);
and U17048 (N_17048,N_16098,N_16321);
and U17049 (N_17049,N_16103,N_16271);
nand U17050 (N_17050,N_16250,N_16082);
nor U17051 (N_17051,N_16773,N_16653);
nand U17052 (N_17052,N_16598,N_16340);
nor U17053 (N_17053,N_16450,N_16606);
and U17054 (N_17054,N_16149,N_16224);
xnor U17055 (N_17055,N_16362,N_16637);
and U17056 (N_17056,N_16142,N_16357);
or U17057 (N_17057,N_16468,N_16269);
xor U17058 (N_17058,N_16319,N_16045);
xor U17059 (N_17059,N_16197,N_16504);
nor U17060 (N_17060,N_16164,N_16700);
and U17061 (N_17061,N_16323,N_16760);
and U17062 (N_17062,N_16328,N_16683);
nor U17063 (N_17063,N_16421,N_16378);
or U17064 (N_17064,N_16722,N_16427);
or U17065 (N_17065,N_16382,N_16377);
nor U17066 (N_17066,N_16073,N_16462);
and U17067 (N_17067,N_16117,N_16526);
xor U17068 (N_17068,N_16156,N_16258);
nor U17069 (N_17069,N_16128,N_16154);
xor U17070 (N_17070,N_16092,N_16494);
nor U17071 (N_17071,N_16255,N_16695);
or U17072 (N_17072,N_16268,N_16550);
nor U17073 (N_17073,N_16559,N_16492);
nand U17074 (N_17074,N_16368,N_16616);
and U17075 (N_17075,N_16028,N_16040);
nor U17076 (N_17076,N_16566,N_16160);
or U17077 (N_17077,N_16679,N_16248);
or U17078 (N_17078,N_16151,N_16673);
xor U17079 (N_17079,N_16320,N_16530);
and U17080 (N_17080,N_16292,N_16185);
or U17081 (N_17081,N_16536,N_16174);
xor U17082 (N_17082,N_16032,N_16788);
xnor U17083 (N_17083,N_16692,N_16379);
xnor U17084 (N_17084,N_16498,N_16296);
and U17085 (N_17085,N_16590,N_16417);
and U17086 (N_17086,N_16023,N_16216);
xnor U17087 (N_17087,N_16440,N_16721);
or U17088 (N_17088,N_16046,N_16718);
nand U17089 (N_17089,N_16159,N_16710);
nor U17090 (N_17090,N_16565,N_16088);
nand U17091 (N_17091,N_16608,N_16244);
xnor U17092 (N_17092,N_16626,N_16500);
or U17093 (N_17093,N_16757,N_16024);
xor U17094 (N_17094,N_16152,N_16639);
xnor U17095 (N_17095,N_16667,N_16797);
nand U17096 (N_17096,N_16097,N_16781);
or U17097 (N_17097,N_16671,N_16036);
xor U17098 (N_17098,N_16776,N_16102);
xor U17099 (N_17099,N_16697,N_16161);
or U17100 (N_17100,N_16602,N_16090);
nand U17101 (N_17101,N_16740,N_16166);
nor U17102 (N_17102,N_16243,N_16659);
and U17103 (N_17103,N_16392,N_16663);
nand U17104 (N_17104,N_16014,N_16004);
and U17105 (N_17105,N_16306,N_16339);
nand U17106 (N_17106,N_16215,N_16133);
xnor U17107 (N_17107,N_16355,N_16084);
or U17108 (N_17108,N_16713,N_16521);
nand U17109 (N_17109,N_16060,N_16294);
xor U17110 (N_17110,N_16422,N_16079);
and U17111 (N_17111,N_16111,N_16153);
and U17112 (N_17112,N_16424,N_16071);
xor U17113 (N_17113,N_16068,N_16611);
nand U17114 (N_17114,N_16238,N_16181);
or U17115 (N_17115,N_16675,N_16251);
nand U17116 (N_17116,N_16091,N_16644);
and U17117 (N_17117,N_16202,N_16354);
nand U17118 (N_17118,N_16132,N_16126);
nand U17119 (N_17119,N_16281,N_16433);
nor U17120 (N_17120,N_16239,N_16655);
and U17121 (N_17121,N_16410,N_16072);
and U17122 (N_17122,N_16613,N_16403);
xnor U17123 (N_17123,N_16629,N_16316);
xnor U17124 (N_17124,N_16146,N_16437);
xnor U17125 (N_17125,N_16101,N_16413);
and U17126 (N_17126,N_16165,N_16642);
xor U17127 (N_17127,N_16038,N_16652);
xor U17128 (N_17128,N_16061,N_16039);
or U17129 (N_17129,N_16195,N_16217);
and U17130 (N_17130,N_16769,N_16753);
and U17131 (N_17131,N_16441,N_16670);
xnor U17132 (N_17132,N_16031,N_16301);
or U17133 (N_17133,N_16669,N_16554);
and U17134 (N_17134,N_16015,N_16723);
or U17135 (N_17135,N_16106,N_16487);
and U17136 (N_17136,N_16308,N_16344);
or U17137 (N_17137,N_16012,N_16254);
and U17138 (N_17138,N_16231,N_16030);
nand U17139 (N_17139,N_16551,N_16750);
nor U17140 (N_17140,N_16556,N_16717);
or U17141 (N_17141,N_16273,N_16204);
nand U17142 (N_17142,N_16085,N_16747);
or U17143 (N_17143,N_16175,N_16027);
xnor U17144 (N_17144,N_16342,N_16524);
and U17145 (N_17145,N_16579,N_16587);
xnor U17146 (N_17146,N_16001,N_16497);
nor U17147 (N_17147,N_16707,N_16266);
or U17148 (N_17148,N_16474,N_16656);
xor U17149 (N_17149,N_16176,N_16139);
or U17150 (N_17150,N_16777,N_16263);
xnor U17151 (N_17151,N_16581,N_16425);
xor U17152 (N_17152,N_16533,N_16430);
nor U17153 (N_17153,N_16173,N_16687);
and U17154 (N_17154,N_16715,N_16520);
and U17155 (N_17155,N_16573,N_16205);
nand U17156 (N_17156,N_16359,N_16158);
and U17157 (N_17157,N_16005,N_16311);
nor U17158 (N_17158,N_16495,N_16480);
xor U17159 (N_17159,N_16335,N_16257);
and U17160 (N_17160,N_16562,N_16634);
nand U17161 (N_17161,N_16604,N_16162);
or U17162 (N_17162,N_16042,N_16765);
nor U17163 (N_17163,N_16650,N_16009);
or U17164 (N_17164,N_16077,N_16491);
nor U17165 (N_17165,N_16662,N_16247);
and U17166 (N_17166,N_16105,N_16370);
or U17167 (N_17167,N_16641,N_16657);
or U17168 (N_17168,N_16326,N_16198);
or U17169 (N_17169,N_16470,N_16170);
or U17170 (N_17170,N_16610,N_16627);
xor U17171 (N_17171,N_16754,N_16147);
xnor U17172 (N_17172,N_16628,N_16748);
xor U17173 (N_17173,N_16528,N_16066);
and U17174 (N_17174,N_16124,N_16614);
and U17175 (N_17175,N_16423,N_16502);
or U17176 (N_17176,N_16360,N_16570);
and U17177 (N_17177,N_16275,N_16689);
nor U17178 (N_17178,N_16120,N_16666);
and U17179 (N_17179,N_16070,N_16694);
and U17180 (N_17180,N_16549,N_16651);
nand U17181 (N_17181,N_16373,N_16586);
nor U17182 (N_17182,N_16221,N_16242);
xnor U17183 (N_17183,N_16794,N_16455);
xnor U17184 (N_17184,N_16220,N_16786);
nor U17185 (N_17185,N_16790,N_16209);
nor U17186 (N_17186,N_16130,N_16291);
nor U17187 (N_17187,N_16539,N_16415);
nor U17188 (N_17188,N_16540,N_16322);
nand U17189 (N_17189,N_16795,N_16349);
or U17190 (N_17190,N_16093,N_16575);
nor U17191 (N_17191,N_16724,N_16353);
and U17192 (N_17192,N_16615,N_16716);
xor U17193 (N_17193,N_16199,N_16509);
and U17194 (N_17194,N_16411,N_16108);
nand U17195 (N_17195,N_16745,N_16020);
nor U17196 (N_17196,N_16443,N_16712);
nand U17197 (N_17197,N_16544,N_16654);
nor U17198 (N_17198,N_16172,N_16459);
and U17199 (N_17199,N_16094,N_16305);
nor U17200 (N_17200,N_16009,N_16233);
or U17201 (N_17201,N_16746,N_16259);
and U17202 (N_17202,N_16705,N_16213);
and U17203 (N_17203,N_16192,N_16638);
or U17204 (N_17204,N_16796,N_16616);
and U17205 (N_17205,N_16338,N_16083);
nand U17206 (N_17206,N_16522,N_16605);
nand U17207 (N_17207,N_16762,N_16165);
xor U17208 (N_17208,N_16224,N_16344);
nand U17209 (N_17209,N_16630,N_16668);
xor U17210 (N_17210,N_16291,N_16732);
or U17211 (N_17211,N_16522,N_16311);
xor U17212 (N_17212,N_16348,N_16053);
and U17213 (N_17213,N_16293,N_16227);
and U17214 (N_17214,N_16522,N_16052);
and U17215 (N_17215,N_16226,N_16334);
nand U17216 (N_17216,N_16113,N_16374);
and U17217 (N_17217,N_16029,N_16390);
nand U17218 (N_17218,N_16484,N_16074);
or U17219 (N_17219,N_16082,N_16770);
nand U17220 (N_17220,N_16561,N_16255);
xor U17221 (N_17221,N_16375,N_16210);
or U17222 (N_17222,N_16762,N_16621);
xnor U17223 (N_17223,N_16493,N_16702);
and U17224 (N_17224,N_16563,N_16555);
or U17225 (N_17225,N_16609,N_16397);
xor U17226 (N_17226,N_16756,N_16321);
nand U17227 (N_17227,N_16615,N_16745);
xnor U17228 (N_17228,N_16090,N_16262);
nor U17229 (N_17229,N_16444,N_16300);
and U17230 (N_17230,N_16390,N_16234);
and U17231 (N_17231,N_16157,N_16759);
or U17232 (N_17232,N_16136,N_16419);
nand U17233 (N_17233,N_16403,N_16073);
or U17234 (N_17234,N_16180,N_16012);
or U17235 (N_17235,N_16421,N_16011);
nor U17236 (N_17236,N_16399,N_16443);
nor U17237 (N_17237,N_16187,N_16741);
and U17238 (N_17238,N_16677,N_16621);
nor U17239 (N_17239,N_16443,N_16535);
or U17240 (N_17240,N_16217,N_16062);
nand U17241 (N_17241,N_16164,N_16668);
or U17242 (N_17242,N_16169,N_16711);
or U17243 (N_17243,N_16171,N_16679);
nor U17244 (N_17244,N_16789,N_16731);
and U17245 (N_17245,N_16083,N_16201);
nor U17246 (N_17246,N_16768,N_16492);
and U17247 (N_17247,N_16544,N_16698);
or U17248 (N_17248,N_16797,N_16188);
and U17249 (N_17249,N_16598,N_16156);
xor U17250 (N_17250,N_16007,N_16310);
xor U17251 (N_17251,N_16036,N_16599);
and U17252 (N_17252,N_16767,N_16132);
and U17253 (N_17253,N_16061,N_16593);
and U17254 (N_17254,N_16682,N_16669);
nor U17255 (N_17255,N_16746,N_16270);
or U17256 (N_17256,N_16087,N_16044);
and U17257 (N_17257,N_16031,N_16371);
nor U17258 (N_17258,N_16503,N_16536);
xnor U17259 (N_17259,N_16004,N_16655);
and U17260 (N_17260,N_16090,N_16034);
xor U17261 (N_17261,N_16667,N_16768);
nand U17262 (N_17262,N_16612,N_16416);
or U17263 (N_17263,N_16301,N_16201);
or U17264 (N_17264,N_16026,N_16770);
nand U17265 (N_17265,N_16577,N_16102);
nand U17266 (N_17266,N_16131,N_16179);
xnor U17267 (N_17267,N_16034,N_16252);
or U17268 (N_17268,N_16115,N_16746);
xnor U17269 (N_17269,N_16380,N_16457);
nand U17270 (N_17270,N_16135,N_16344);
nor U17271 (N_17271,N_16310,N_16416);
or U17272 (N_17272,N_16444,N_16060);
nor U17273 (N_17273,N_16206,N_16641);
nor U17274 (N_17274,N_16431,N_16321);
nand U17275 (N_17275,N_16196,N_16684);
and U17276 (N_17276,N_16144,N_16256);
nor U17277 (N_17277,N_16443,N_16189);
nor U17278 (N_17278,N_16131,N_16649);
xnor U17279 (N_17279,N_16303,N_16384);
nor U17280 (N_17280,N_16717,N_16557);
or U17281 (N_17281,N_16630,N_16455);
nand U17282 (N_17282,N_16209,N_16734);
nor U17283 (N_17283,N_16674,N_16595);
nor U17284 (N_17284,N_16023,N_16426);
nor U17285 (N_17285,N_16625,N_16622);
xnor U17286 (N_17286,N_16095,N_16726);
nor U17287 (N_17287,N_16309,N_16191);
or U17288 (N_17288,N_16791,N_16779);
or U17289 (N_17289,N_16714,N_16125);
and U17290 (N_17290,N_16510,N_16016);
or U17291 (N_17291,N_16462,N_16442);
nand U17292 (N_17292,N_16427,N_16241);
and U17293 (N_17293,N_16071,N_16067);
xor U17294 (N_17294,N_16775,N_16589);
nor U17295 (N_17295,N_16537,N_16081);
or U17296 (N_17296,N_16545,N_16779);
or U17297 (N_17297,N_16432,N_16471);
xor U17298 (N_17298,N_16509,N_16323);
xor U17299 (N_17299,N_16069,N_16092);
nor U17300 (N_17300,N_16357,N_16565);
xnor U17301 (N_17301,N_16668,N_16118);
nor U17302 (N_17302,N_16398,N_16491);
or U17303 (N_17303,N_16200,N_16775);
nand U17304 (N_17304,N_16227,N_16609);
and U17305 (N_17305,N_16502,N_16209);
xor U17306 (N_17306,N_16475,N_16770);
and U17307 (N_17307,N_16039,N_16334);
xor U17308 (N_17308,N_16184,N_16098);
nand U17309 (N_17309,N_16678,N_16522);
xor U17310 (N_17310,N_16314,N_16641);
xor U17311 (N_17311,N_16163,N_16779);
nand U17312 (N_17312,N_16463,N_16208);
xor U17313 (N_17313,N_16401,N_16506);
nor U17314 (N_17314,N_16255,N_16368);
xnor U17315 (N_17315,N_16532,N_16760);
nand U17316 (N_17316,N_16135,N_16075);
nor U17317 (N_17317,N_16742,N_16415);
xnor U17318 (N_17318,N_16433,N_16092);
xnor U17319 (N_17319,N_16289,N_16557);
or U17320 (N_17320,N_16698,N_16263);
nor U17321 (N_17321,N_16651,N_16270);
nand U17322 (N_17322,N_16039,N_16388);
nor U17323 (N_17323,N_16620,N_16467);
and U17324 (N_17324,N_16756,N_16445);
xnor U17325 (N_17325,N_16543,N_16008);
and U17326 (N_17326,N_16602,N_16183);
and U17327 (N_17327,N_16077,N_16283);
or U17328 (N_17328,N_16420,N_16511);
nand U17329 (N_17329,N_16766,N_16154);
xnor U17330 (N_17330,N_16795,N_16087);
xor U17331 (N_17331,N_16263,N_16081);
and U17332 (N_17332,N_16228,N_16370);
and U17333 (N_17333,N_16248,N_16457);
nor U17334 (N_17334,N_16234,N_16697);
or U17335 (N_17335,N_16005,N_16799);
and U17336 (N_17336,N_16000,N_16033);
nor U17337 (N_17337,N_16205,N_16347);
nand U17338 (N_17338,N_16396,N_16060);
nor U17339 (N_17339,N_16342,N_16682);
nor U17340 (N_17340,N_16355,N_16696);
nor U17341 (N_17341,N_16706,N_16475);
nand U17342 (N_17342,N_16474,N_16559);
nand U17343 (N_17343,N_16742,N_16136);
xor U17344 (N_17344,N_16525,N_16511);
or U17345 (N_17345,N_16241,N_16665);
or U17346 (N_17346,N_16537,N_16184);
nand U17347 (N_17347,N_16523,N_16266);
nor U17348 (N_17348,N_16564,N_16243);
and U17349 (N_17349,N_16272,N_16302);
or U17350 (N_17350,N_16494,N_16146);
or U17351 (N_17351,N_16132,N_16202);
or U17352 (N_17352,N_16211,N_16199);
xnor U17353 (N_17353,N_16398,N_16395);
nand U17354 (N_17354,N_16668,N_16646);
or U17355 (N_17355,N_16747,N_16380);
nor U17356 (N_17356,N_16138,N_16393);
and U17357 (N_17357,N_16325,N_16261);
nor U17358 (N_17358,N_16637,N_16681);
xnor U17359 (N_17359,N_16146,N_16040);
and U17360 (N_17360,N_16332,N_16696);
xor U17361 (N_17361,N_16196,N_16230);
xnor U17362 (N_17362,N_16621,N_16159);
xor U17363 (N_17363,N_16598,N_16142);
nor U17364 (N_17364,N_16562,N_16063);
nand U17365 (N_17365,N_16749,N_16671);
or U17366 (N_17366,N_16192,N_16417);
nor U17367 (N_17367,N_16625,N_16357);
nand U17368 (N_17368,N_16265,N_16732);
and U17369 (N_17369,N_16089,N_16286);
and U17370 (N_17370,N_16447,N_16005);
or U17371 (N_17371,N_16330,N_16315);
xor U17372 (N_17372,N_16242,N_16407);
nand U17373 (N_17373,N_16279,N_16438);
or U17374 (N_17374,N_16365,N_16257);
nor U17375 (N_17375,N_16570,N_16490);
or U17376 (N_17376,N_16466,N_16451);
or U17377 (N_17377,N_16045,N_16625);
nand U17378 (N_17378,N_16346,N_16186);
nand U17379 (N_17379,N_16030,N_16139);
xnor U17380 (N_17380,N_16389,N_16735);
xnor U17381 (N_17381,N_16649,N_16041);
xor U17382 (N_17382,N_16755,N_16780);
or U17383 (N_17383,N_16167,N_16458);
nor U17384 (N_17384,N_16265,N_16676);
xor U17385 (N_17385,N_16599,N_16603);
or U17386 (N_17386,N_16331,N_16340);
xnor U17387 (N_17387,N_16140,N_16695);
xnor U17388 (N_17388,N_16476,N_16143);
or U17389 (N_17389,N_16360,N_16630);
or U17390 (N_17390,N_16122,N_16724);
nor U17391 (N_17391,N_16570,N_16687);
nor U17392 (N_17392,N_16585,N_16070);
and U17393 (N_17393,N_16757,N_16384);
xor U17394 (N_17394,N_16271,N_16176);
xnor U17395 (N_17395,N_16250,N_16169);
xnor U17396 (N_17396,N_16514,N_16662);
nor U17397 (N_17397,N_16527,N_16491);
xor U17398 (N_17398,N_16092,N_16588);
nand U17399 (N_17399,N_16421,N_16111);
xnor U17400 (N_17400,N_16407,N_16656);
nor U17401 (N_17401,N_16561,N_16227);
nand U17402 (N_17402,N_16729,N_16652);
xnor U17403 (N_17403,N_16244,N_16605);
and U17404 (N_17404,N_16189,N_16569);
and U17405 (N_17405,N_16783,N_16573);
or U17406 (N_17406,N_16625,N_16335);
nand U17407 (N_17407,N_16488,N_16031);
or U17408 (N_17408,N_16495,N_16246);
or U17409 (N_17409,N_16029,N_16353);
and U17410 (N_17410,N_16532,N_16233);
nand U17411 (N_17411,N_16299,N_16009);
xor U17412 (N_17412,N_16264,N_16244);
xor U17413 (N_17413,N_16472,N_16689);
nand U17414 (N_17414,N_16340,N_16547);
and U17415 (N_17415,N_16025,N_16717);
nand U17416 (N_17416,N_16167,N_16290);
and U17417 (N_17417,N_16731,N_16518);
or U17418 (N_17418,N_16438,N_16683);
xor U17419 (N_17419,N_16642,N_16450);
or U17420 (N_17420,N_16155,N_16651);
or U17421 (N_17421,N_16212,N_16014);
nand U17422 (N_17422,N_16530,N_16562);
nor U17423 (N_17423,N_16514,N_16211);
and U17424 (N_17424,N_16269,N_16558);
xnor U17425 (N_17425,N_16051,N_16459);
nor U17426 (N_17426,N_16381,N_16527);
nor U17427 (N_17427,N_16138,N_16344);
xnor U17428 (N_17428,N_16356,N_16458);
nor U17429 (N_17429,N_16075,N_16209);
and U17430 (N_17430,N_16689,N_16457);
or U17431 (N_17431,N_16487,N_16062);
nor U17432 (N_17432,N_16020,N_16606);
nand U17433 (N_17433,N_16017,N_16594);
or U17434 (N_17434,N_16125,N_16557);
xor U17435 (N_17435,N_16071,N_16707);
nor U17436 (N_17436,N_16593,N_16455);
or U17437 (N_17437,N_16599,N_16657);
or U17438 (N_17438,N_16201,N_16234);
nand U17439 (N_17439,N_16383,N_16365);
or U17440 (N_17440,N_16421,N_16504);
nor U17441 (N_17441,N_16744,N_16359);
nand U17442 (N_17442,N_16182,N_16588);
nor U17443 (N_17443,N_16743,N_16697);
xor U17444 (N_17444,N_16599,N_16790);
xnor U17445 (N_17445,N_16683,N_16023);
nand U17446 (N_17446,N_16649,N_16127);
xor U17447 (N_17447,N_16628,N_16112);
nand U17448 (N_17448,N_16650,N_16285);
nor U17449 (N_17449,N_16404,N_16683);
nor U17450 (N_17450,N_16652,N_16209);
nand U17451 (N_17451,N_16341,N_16571);
nand U17452 (N_17452,N_16264,N_16365);
and U17453 (N_17453,N_16599,N_16642);
nand U17454 (N_17454,N_16139,N_16699);
and U17455 (N_17455,N_16046,N_16396);
nor U17456 (N_17456,N_16723,N_16798);
or U17457 (N_17457,N_16220,N_16573);
xor U17458 (N_17458,N_16062,N_16452);
or U17459 (N_17459,N_16395,N_16389);
and U17460 (N_17460,N_16036,N_16605);
or U17461 (N_17461,N_16145,N_16197);
nor U17462 (N_17462,N_16345,N_16718);
nor U17463 (N_17463,N_16075,N_16689);
or U17464 (N_17464,N_16559,N_16077);
nor U17465 (N_17465,N_16768,N_16077);
nor U17466 (N_17466,N_16185,N_16797);
or U17467 (N_17467,N_16241,N_16581);
nand U17468 (N_17468,N_16675,N_16053);
nor U17469 (N_17469,N_16445,N_16319);
or U17470 (N_17470,N_16430,N_16432);
or U17471 (N_17471,N_16214,N_16747);
or U17472 (N_17472,N_16143,N_16244);
nand U17473 (N_17473,N_16538,N_16017);
xnor U17474 (N_17474,N_16071,N_16117);
or U17475 (N_17475,N_16279,N_16693);
nand U17476 (N_17476,N_16578,N_16327);
or U17477 (N_17477,N_16335,N_16203);
or U17478 (N_17478,N_16324,N_16098);
nor U17479 (N_17479,N_16258,N_16366);
or U17480 (N_17480,N_16755,N_16041);
nand U17481 (N_17481,N_16788,N_16532);
xnor U17482 (N_17482,N_16508,N_16473);
or U17483 (N_17483,N_16236,N_16793);
and U17484 (N_17484,N_16759,N_16520);
and U17485 (N_17485,N_16028,N_16507);
or U17486 (N_17486,N_16017,N_16564);
and U17487 (N_17487,N_16213,N_16541);
or U17488 (N_17488,N_16166,N_16085);
or U17489 (N_17489,N_16059,N_16500);
nor U17490 (N_17490,N_16467,N_16794);
xor U17491 (N_17491,N_16077,N_16073);
nand U17492 (N_17492,N_16017,N_16366);
and U17493 (N_17493,N_16562,N_16322);
nor U17494 (N_17494,N_16634,N_16310);
nand U17495 (N_17495,N_16544,N_16330);
and U17496 (N_17496,N_16746,N_16357);
xor U17497 (N_17497,N_16679,N_16795);
xor U17498 (N_17498,N_16665,N_16716);
nand U17499 (N_17499,N_16532,N_16369);
nand U17500 (N_17500,N_16409,N_16097);
or U17501 (N_17501,N_16445,N_16473);
and U17502 (N_17502,N_16519,N_16113);
nand U17503 (N_17503,N_16001,N_16313);
xnor U17504 (N_17504,N_16707,N_16005);
and U17505 (N_17505,N_16604,N_16113);
nand U17506 (N_17506,N_16034,N_16188);
or U17507 (N_17507,N_16551,N_16574);
nand U17508 (N_17508,N_16284,N_16484);
nor U17509 (N_17509,N_16747,N_16559);
nand U17510 (N_17510,N_16142,N_16343);
and U17511 (N_17511,N_16777,N_16160);
nor U17512 (N_17512,N_16231,N_16244);
or U17513 (N_17513,N_16726,N_16613);
and U17514 (N_17514,N_16196,N_16222);
and U17515 (N_17515,N_16270,N_16402);
xor U17516 (N_17516,N_16714,N_16430);
and U17517 (N_17517,N_16261,N_16248);
or U17518 (N_17518,N_16636,N_16301);
and U17519 (N_17519,N_16484,N_16585);
and U17520 (N_17520,N_16733,N_16214);
nor U17521 (N_17521,N_16072,N_16593);
nor U17522 (N_17522,N_16214,N_16293);
xor U17523 (N_17523,N_16418,N_16313);
nor U17524 (N_17524,N_16610,N_16137);
and U17525 (N_17525,N_16518,N_16549);
xnor U17526 (N_17526,N_16368,N_16043);
xnor U17527 (N_17527,N_16148,N_16187);
and U17528 (N_17528,N_16272,N_16050);
or U17529 (N_17529,N_16273,N_16339);
and U17530 (N_17530,N_16583,N_16294);
nor U17531 (N_17531,N_16651,N_16769);
and U17532 (N_17532,N_16009,N_16434);
and U17533 (N_17533,N_16659,N_16528);
xnor U17534 (N_17534,N_16673,N_16643);
nor U17535 (N_17535,N_16482,N_16670);
nor U17536 (N_17536,N_16620,N_16334);
or U17537 (N_17537,N_16707,N_16041);
nor U17538 (N_17538,N_16352,N_16169);
nand U17539 (N_17539,N_16015,N_16072);
xnor U17540 (N_17540,N_16243,N_16619);
or U17541 (N_17541,N_16616,N_16427);
or U17542 (N_17542,N_16262,N_16775);
and U17543 (N_17543,N_16750,N_16770);
nor U17544 (N_17544,N_16540,N_16423);
xnor U17545 (N_17545,N_16631,N_16242);
nand U17546 (N_17546,N_16648,N_16496);
and U17547 (N_17547,N_16178,N_16516);
and U17548 (N_17548,N_16491,N_16791);
nand U17549 (N_17549,N_16510,N_16741);
or U17550 (N_17550,N_16627,N_16799);
nor U17551 (N_17551,N_16263,N_16151);
and U17552 (N_17552,N_16526,N_16486);
nor U17553 (N_17553,N_16428,N_16670);
and U17554 (N_17554,N_16167,N_16179);
nor U17555 (N_17555,N_16261,N_16454);
nor U17556 (N_17556,N_16230,N_16419);
or U17557 (N_17557,N_16270,N_16653);
nand U17558 (N_17558,N_16710,N_16384);
nor U17559 (N_17559,N_16471,N_16514);
and U17560 (N_17560,N_16502,N_16462);
and U17561 (N_17561,N_16350,N_16676);
xnor U17562 (N_17562,N_16399,N_16165);
and U17563 (N_17563,N_16549,N_16018);
nand U17564 (N_17564,N_16724,N_16286);
nand U17565 (N_17565,N_16686,N_16459);
and U17566 (N_17566,N_16084,N_16711);
or U17567 (N_17567,N_16285,N_16237);
and U17568 (N_17568,N_16491,N_16764);
and U17569 (N_17569,N_16543,N_16559);
xor U17570 (N_17570,N_16159,N_16078);
xnor U17571 (N_17571,N_16416,N_16607);
nand U17572 (N_17572,N_16165,N_16207);
and U17573 (N_17573,N_16657,N_16089);
or U17574 (N_17574,N_16112,N_16048);
or U17575 (N_17575,N_16566,N_16309);
or U17576 (N_17576,N_16766,N_16299);
nor U17577 (N_17577,N_16713,N_16670);
nand U17578 (N_17578,N_16117,N_16415);
nor U17579 (N_17579,N_16350,N_16030);
and U17580 (N_17580,N_16029,N_16785);
or U17581 (N_17581,N_16147,N_16315);
and U17582 (N_17582,N_16664,N_16175);
or U17583 (N_17583,N_16570,N_16606);
and U17584 (N_17584,N_16044,N_16281);
xor U17585 (N_17585,N_16282,N_16319);
or U17586 (N_17586,N_16627,N_16274);
xor U17587 (N_17587,N_16114,N_16283);
nor U17588 (N_17588,N_16535,N_16629);
nand U17589 (N_17589,N_16402,N_16223);
nor U17590 (N_17590,N_16130,N_16461);
and U17591 (N_17591,N_16213,N_16649);
or U17592 (N_17592,N_16778,N_16158);
nand U17593 (N_17593,N_16588,N_16353);
and U17594 (N_17594,N_16575,N_16174);
or U17595 (N_17595,N_16573,N_16199);
or U17596 (N_17596,N_16728,N_16394);
or U17597 (N_17597,N_16678,N_16487);
nand U17598 (N_17598,N_16535,N_16020);
nor U17599 (N_17599,N_16439,N_16643);
nor U17600 (N_17600,N_16814,N_17518);
nand U17601 (N_17601,N_17582,N_16828);
or U17602 (N_17602,N_17234,N_17522);
or U17603 (N_17603,N_17353,N_17199);
xor U17604 (N_17604,N_17081,N_17075);
and U17605 (N_17605,N_17371,N_17528);
or U17606 (N_17606,N_16855,N_17171);
nand U17607 (N_17607,N_16801,N_17414);
or U17608 (N_17608,N_17273,N_17255);
and U17609 (N_17609,N_17423,N_17431);
xor U17610 (N_17610,N_16859,N_17027);
xnor U17611 (N_17611,N_17253,N_17091);
nor U17612 (N_17612,N_17179,N_17571);
nor U17613 (N_17613,N_17280,N_16978);
nor U17614 (N_17614,N_17326,N_16837);
nor U17615 (N_17615,N_17594,N_17087);
or U17616 (N_17616,N_17555,N_17053);
and U17617 (N_17617,N_17204,N_17543);
nand U17618 (N_17618,N_17118,N_17475);
or U17619 (N_17619,N_17206,N_17267);
or U17620 (N_17620,N_16925,N_17147);
nand U17621 (N_17621,N_17003,N_17295);
or U17622 (N_17622,N_17530,N_17078);
nand U17623 (N_17623,N_17491,N_17019);
and U17624 (N_17624,N_17464,N_17593);
nor U17625 (N_17625,N_17277,N_17224);
nand U17626 (N_17626,N_17347,N_17120);
nor U17627 (N_17627,N_16998,N_17222);
nor U17628 (N_17628,N_17346,N_17082);
xnor U17629 (N_17629,N_17237,N_17355);
xnor U17630 (N_17630,N_17070,N_16800);
and U17631 (N_17631,N_16812,N_17080);
and U17632 (N_17632,N_17203,N_16848);
xnor U17633 (N_17633,N_16880,N_16962);
nand U17634 (N_17634,N_17059,N_17592);
or U17635 (N_17635,N_16955,N_17297);
nor U17636 (N_17636,N_17545,N_17465);
and U17637 (N_17637,N_16875,N_16886);
nand U17638 (N_17638,N_17205,N_17268);
nand U17639 (N_17639,N_17497,N_17366);
nor U17640 (N_17640,N_17071,N_17260);
xnor U17641 (N_17641,N_17183,N_17215);
or U17642 (N_17642,N_17308,N_17067);
nor U17643 (N_17643,N_16988,N_17211);
nor U17644 (N_17644,N_17124,N_17453);
nand U17645 (N_17645,N_17435,N_16999);
and U17646 (N_17646,N_17228,N_17429);
xnor U17647 (N_17647,N_17021,N_17437);
xor U17648 (N_17648,N_17316,N_16900);
xor U17649 (N_17649,N_17569,N_17047);
nand U17650 (N_17650,N_17102,N_16896);
xor U17651 (N_17651,N_17046,N_17262);
nor U17652 (N_17652,N_17164,N_17135);
nor U17653 (N_17653,N_17049,N_16860);
nand U17654 (N_17654,N_17155,N_16968);
nand U17655 (N_17655,N_16845,N_17553);
or U17656 (N_17656,N_17094,N_17384);
nand U17657 (N_17657,N_17013,N_17235);
nand U17658 (N_17658,N_16909,N_16866);
and U17659 (N_17659,N_17484,N_17289);
or U17660 (N_17660,N_17542,N_17519);
nor U17661 (N_17661,N_17140,N_16937);
and U17662 (N_17662,N_17445,N_16942);
xnor U17663 (N_17663,N_17459,N_16974);
or U17664 (N_17664,N_16963,N_17559);
nand U17665 (N_17665,N_17525,N_17176);
or U17666 (N_17666,N_17424,N_17416);
nand U17667 (N_17667,N_16980,N_16873);
xor U17668 (N_17668,N_17130,N_17596);
xnor U17669 (N_17669,N_16819,N_16850);
nand U17670 (N_17670,N_17196,N_16945);
and U17671 (N_17671,N_16898,N_17101);
nand U17672 (N_17672,N_17010,N_16977);
or U17673 (N_17673,N_17270,N_17188);
nand U17674 (N_17674,N_17343,N_16882);
nand U17675 (N_17675,N_17048,N_17016);
nor U17676 (N_17676,N_17139,N_17434);
nand U17677 (N_17677,N_17396,N_17560);
xnor U17678 (N_17678,N_17551,N_16916);
nor U17679 (N_17679,N_17031,N_17402);
xnor U17680 (N_17680,N_17058,N_17441);
xnor U17681 (N_17681,N_17531,N_16894);
nor U17682 (N_17682,N_17388,N_17149);
nor U17683 (N_17683,N_17293,N_17008);
or U17684 (N_17684,N_16863,N_16893);
nand U17685 (N_17685,N_16921,N_17471);
nor U17686 (N_17686,N_16930,N_17232);
or U17687 (N_17687,N_17446,N_17291);
or U17688 (N_17688,N_16841,N_17264);
xor U17689 (N_17689,N_17061,N_17357);
or U17690 (N_17690,N_16908,N_16934);
and U17691 (N_17691,N_17391,N_17247);
or U17692 (N_17692,N_16954,N_17558);
or U17693 (N_17693,N_17045,N_17409);
nand U17694 (N_17694,N_17038,N_17202);
xor U17695 (N_17695,N_16877,N_16985);
xor U17696 (N_17696,N_17127,N_17192);
xnor U17697 (N_17697,N_17405,N_17329);
nor U17698 (N_17698,N_17482,N_17532);
nor U17699 (N_17699,N_17440,N_17461);
and U17700 (N_17700,N_16815,N_17083);
and U17701 (N_17701,N_17052,N_17447);
and U17702 (N_17702,N_17470,N_17263);
xor U17703 (N_17703,N_17397,N_17212);
and U17704 (N_17704,N_17336,N_16834);
xnor U17705 (N_17705,N_17564,N_17126);
nand U17706 (N_17706,N_17033,N_17376);
xnor U17707 (N_17707,N_17356,N_16982);
xor U17708 (N_17708,N_16917,N_16810);
nand U17709 (N_17709,N_17578,N_17546);
nand U17710 (N_17710,N_17112,N_17166);
or U17711 (N_17711,N_16804,N_17375);
xnor U17712 (N_17712,N_17244,N_16904);
nand U17713 (N_17713,N_17389,N_16947);
nor U17714 (N_17714,N_17085,N_16981);
nand U17715 (N_17715,N_17328,N_17221);
and U17716 (N_17716,N_17116,N_17442);
or U17717 (N_17717,N_16840,N_17517);
or U17718 (N_17718,N_17151,N_16933);
nand U17719 (N_17719,N_17208,N_17566);
nor U17720 (N_17720,N_17369,N_16842);
nand U17721 (N_17721,N_17495,N_17303);
nor U17722 (N_17722,N_16936,N_16984);
nand U17723 (N_17723,N_16931,N_16849);
xor U17724 (N_17724,N_17514,N_16958);
xor U17725 (N_17725,N_16990,N_17398);
or U17726 (N_17726,N_17042,N_17092);
and U17727 (N_17727,N_17349,N_17315);
and U17728 (N_17728,N_17283,N_17313);
or U17729 (N_17729,N_17536,N_17233);
xnor U17730 (N_17730,N_17039,N_16844);
nand U17731 (N_17731,N_17077,N_16961);
and U17732 (N_17732,N_17436,N_17084);
xor U17733 (N_17733,N_17143,N_17163);
nor U17734 (N_17734,N_17284,N_17055);
or U17735 (N_17735,N_17157,N_17413);
or U17736 (N_17736,N_16965,N_17590);
and U17737 (N_17737,N_17567,N_17425);
xor U17738 (N_17738,N_16976,N_16808);
xnor U17739 (N_17739,N_17090,N_17159);
xor U17740 (N_17740,N_17427,N_16878);
nor U17741 (N_17741,N_16874,N_17351);
xnor U17742 (N_17742,N_16920,N_17129);
xnor U17743 (N_17743,N_17097,N_17304);
nor U17744 (N_17744,N_17125,N_17287);
xor U17745 (N_17745,N_17462,N_17529);
and U17746 (N_17746,N_17523,N_17065);
and U17747 (N_17747,N_16870,N_16851);
and U17748 (N_17748,N_17156,N_17230);
xor U17749 (N_17749,N_16864,N_16871);
nand U17750 (N_17750,N_17219,N_17452);
or U17751 (N_17751,N_17580,N_17539);
xor U17752 (N_17752,N_16922,N_17421);
or U17753 (N_17753,N_17541,N_17223);
xor U17754 (N_17754,N_17469,N_17296);
and U17755 (N_17755,N_17152,N_17279);
or U17756 (N_17756,N_17302,N_17041);
or U17757 (N_17757,N_17526,N_17412);
or U17758 (N_17758,N_17111,N_17165);
nand U17759 (N_17759,N_16928,N_17348);
xnor U17760 (N_17760,N_17374,N_17318);
or U17761 (N_17761,N_17317,N_17261);
nand U17762 (N_17762,N_17242,N_17504);
xnor U17763 (N_17763,N_16952,N_17191);
and U17764 (N_17764,N_17554,N_17400);
and U17765 (N_17765,N_17500,N_17505);
xor U17766 (N_17766,N_17568,N_17119);
or U17767 (N_17767,N_17030,N_17521);
and U17768 (N_17768,N_16805,N_17054);
and U17769 (N_17769,N_17455,N_17494);
xor U17770 (N_17770,N_17439,N_17588);
nand U17771 (N_17771,N_17114,N_16973);
and U17772 (N_17772,N_17390,N_17319);
nand U17773 (N_17773,N_17361,N_17426);
or U17774 (N_17774,N_16979,N_17332);
or U17775 (N_17775,N_16929,N_16858);
nand U17776 (N_17776,N_17486,N_17327);
xnor U17777 (N_17777,N_17271,N_16861);
xnor U17778 (N_17778,N_17314,N_17477);
nand U17779 (N_17779,N_17066,N_16957);
xor U17780 (N_17780,N_17109,N_17385);
and U17781 (N_17781,N_17419,N_16997);
nand U17782 (N_17782,N_17586,N_17472);
nand U17783 (N_17783,N_17325,N_16983);
nand U17784 (N_17784,N_17367,N_16802);
xnor U17785 (N_17785,N_17581,N_16970);
and U17786 (N_17786,N_17018,N_17236);
nor U17787 (N_17787,N_17217,N_17024);
nor U17788 (N_17788,N_17288,N_16888);
xor U17789 (N_17789,N_16879,N_16901);
nor U17790 (N_17790,N_16852,N_17506);
xor U17791 (N_17791,N_16836,N_17474);
and U17792 (N_17792,N_17064,N_17136);
nor U17793 (N_17793,N_16902,N_16956);
nor U17794 (N_17794,N_17577,N_17345);
nand U17795 (N_17795,N_17392,N_16946);
nor U17796 (N_17796,N_17173,N_17298);
nor U17797 (N_17797,N_17103,N_16823);
nand U17798 (N_17798,N_17074,N_17487);
or U17799 (N_17799,N_17290,N_16891);
or U17800 (N_17800,N_17457,N_17073);
xor U17801 (N_17801,N_16826,N_16822);
nand U17802 (N_17802,N_17257,N_16811);
and U17803 (N_17803,N_16907,N_17556);
or U17804 (N_17804,N_17012,N_17218);
nor U17805 (N_17805,N_17323,N_17305);
xnor U17806 (N_17806,N_17256,N_17197);
nor U17807 (N_17807,N_17510,N_16996);
xor U17808 (N_17808,N_17025,N_16895);
nand U17809 (N_17809,N_17034,N_16960);
nor U17810 (N_17810,N_17020,N_17026);
or U17811 (N_17811,N_16899,N_17007);
nor U17812 (N_17812,N_17489,N_16884);
xor U17813 (N_17813,N_16969,N_16897);
xnor U17814 (N_17814,N_16918,N_17422);
and U17815 (N_17815,N_17272,N_17309);
nor U17816 (N_17816,N_17386,N_17051);
and U17817 (N_17817,N_17524,N_17002);
nand U17818 (N_17818,N_16868,N_17172);
and U17819 (N_17819,N_17372,N_17299);
and U17820 (N_17820,N_17169,N_17358);
and U17821 (N_17821,N_17117,N_16992);
nand U17822 (N_17822,N_17301,N_17285);
and U17823 (N_17823,N_17266,N_17512);
and U17824 (N_17824,N_17100,N_17170);
or U17825 (N_17825,N_17250,N_17294);
xnor U17826 (N_17826,N_17190,N_17324);
and U17827 (N_17827,N_17450,N_17340);
or U17828 (N_17828,N_17200,N_17443);
nor U17829 (N_17829,N_16943,N_17158);
and U17830 (N_17830,N_17359,N_17241);
or U17831 (N_17831,N_16989,N_16847);
nor U17832 (N_17832,N_17310,N_17570);
xnor U17833 (N_17833,N_17547,N_17338);
and U17834 (N_17834,N_17418,N_17050);
nor U17835 (N_17835,N_16915,N_17178);
or U17836 (N_17836,N_16872,N_17185);
xnor U17837 (N_17837,N_16816,N_16919);
and U17838 (N_17838,N_17036,N_16939);
nand U17839 (N_17839,N_16953,N_17468);
nand U17840 (N_17840,N_16806,N_17458);
nand U17841 (N_17841,N_17544,N_17121);
and U17842 (N_17842,N_17527,N_17311);
or U17843 (N_17843,N_16892,N_17286);
or U17844 (N_17844,N_17181,N_16830);
or U17845 (N_17845,N_17227,N_17360);
xnor U17846 (N_17846,N_16924,N_17186);
nor U17847 (N_17847,N_17395,N_17220);
xnor U17848 (N_17848,N_17043,N_17177);
nor U17849 (N_17849,N_17565,N_17509);
and U17850 (N_17850,N_17088,N_17079);
or U17851 (N_17851,N_17281,N_17122);
or U17852 (N_17852,N_17444,N_17337);
nand U17853 (N_17853,N_17193,N_17201);
nand U17854 (N_17854,N_17068,N_17467);
or U17855 (N_17855,N_17410,N_17098);
nand U17856 (N_17856,N_17584,N_17023);
nand U17857 (N_17857,N_16966,N_17005);
or U17858 (N_17858,N_17378,N_17104);
nand U17859 (N_17859,N_16987,N_17107);
nand U17860 (N_17860,N_16825,N_16890);
nand U17861 (N_17861,N_17226,N_17550);
nor U17862 (N_17862,N_17239,N_17096);
xnor U17863 (N_17863,N_16967,N_16995);
or U17864 (N_17864,N_17168,N_17520);
nor U17865 (N_17865,N_17382,N_17145);
nand U17866 (N_17866,N_17167,N_17344);
nand U17867 (N_17867,N_16994,N_17252);
or U17868 (N_17868,N_17591,N_17411);
xor U17869 (N_17869,N_17000,N_17563);
nand U17870 (N_17870,N_17404,N_17415);
xnor U17871 (N_17871,N_17175,N_16857);
or U17872 (N_17872,N_17513,N_17589);
and U17873 (N_17873,N_16843,N_17276);
nor U17874 (N_17874,N_17354,N_17274);
nor U17875 (N_17875,N_17022,N_17449);
or U17876 (N_17876,N_17093,N_17573);
nor U17877 (N_17877,N_17511,N_17456);
and U17878 (N_17878,N_17428,N_16876);
nand U17879 (N_17879,N_16862,N_17269);
and U17880 (N_17880,N_17029,N_17035);
or U17881 (N_17881,N_17032,N_17381);
and U17882 (N_17882,N_17162,N_16912);
and U17883 (N_17883,N_17306,N_17148);
and U17884 (N_17884,N_16853,N_17144);
nor U17885 (N_17885,N_17587,N_16906);
nand U17886 (N_17886,N_16832,N_17365);
nor U17887 (N_17887,N_17502,N_17417);
nor U17888 (N_17888,N_17154,N_17063);
nor U17889 (N_17889,N_17597,N_17265);
and U17890 (N_17890,N_17331,N_17072);
nand U17891 (N_17891,N_17150,N_17498);
nand U17892 (N_17892,N_17363,N_17198);
or U17893 (N_17893,N_17258,N_17420);
xnor U17894 (N_17894,N_17086,N_16865);
or U17895 (N_17895,N_17174,N_17561);
and U17896 (N_17896,N_17394,N_17161);
xnor U17897 (N_17897,N_17380,N_17599);
nand U17898 (N_17898,N_17187,N_17278);
nand U17899 (N_17899,N_17557,N_17407);
xor U17900 (N_17900,N_16951,N_16911);
and U17901 (N_17901,N_17138,N_16913);
nand U17902 (N_17902,N_17108,N_17195);
nor U17903 (N_17903,N_16941,N_17213);
and U17904 (N_17904,N_17320,N_17249);
nand U17905 (N_17905,N_17160,N_16817);
or U17906 (N_17906,N_17579,N_16940);
and U17907 (N_17907,N_17342,N_17089);
nand U17908 (N_17908,N_17399,N_17383);
nor U17909 (N_17909,N_17463,N_16867);
nand U17910 (N_17910,N_17106,N_17238);
nor U17911 (N_17911,N_17370,N_17057);
nand U17912 (N_17912,N_16910,N_16949);
nor U17913 (N_17913,N_17466,N_17387);
and U17914 (N_17914,N_17009,N_17300);
xor U17915 (N_17915,N_17460,N_17339);
or U17916 (N_17916,N_16986,N_17275);
or U17917 (N_17917,N_16883,N_17216);
and U17918 (N_17918,N_16971,N_17040);
or U17919 (N_17919,N_17379,N_17015);
and U17920 (N_17920,N_17245,N_16932);
and U17921 (N_17921,N_17056,N_17490);
or U17922 (N_17922,N_16944,N_16813);
nor U17923 (N_17923,N_17182,N_17499);
and U17924 (N_17924,N_17393,N_17246);
xnor U17925 (N_17925,N_17478,N_16824);
nor U17926 (N_17926,N_17479,N_17377);
xor U17927 (N_17927,N_17432,N_17515);
xor U17928 (N_17928,N_17480,N_17113);
nor U17929 (N_17929,N_17006,N_17503);
and U17930 (N_17930,N_17209,N_17134);
or U17931 (N_17931,N_17362,N_16948);
and U17932 (N_17932,N_17516,N_17254);
nand U17933 (N_17933,N_16927,N_17321);
or U17934 (N_17934,N_17483,N_17128);
and U17935 (N_17935,N_17194,N_17001);
nand U17936 (N_17936,N_17350,N_17534);
nand U17937 (N_17937,N_17017,N_17585);
and U17938 (N_17938,N_16838,N_17574);
nand U17939 (N_17939,N_16959,N_16885);
xnor U17940 (N_17940,N_17368,N_17481);
nand U17941 (N_17941,N_17401,N_16905);
and U17942 (N_17942,N_17501,N_17131);
xnor U17943 (N_17943,N_17110,N_17540);
and U17944 (N_17944,N_17229,N_17322);
or U17945 (N_17945,N_16846,N_17433);
nor U17946 (N_17946,N_16833,N_16975);
or U17947 (N_17947,N_17069,N_16914);
nand U17948 (N_17948,N_16972,N_17492);
xnor U17949 (N_17949,N_17341,N_17028);
or U17950 (N_17950,N_17214,N_16809);
or U17951 (N_17951,N_17248,N_17403);
nor U17952 (N_17952,N_16889,N_17307);
xnor U17953 (N_17953,N_17123,N_17240);
xnor U17954 (N_17954,N_17533,N_16923);
xor U17955 (N_17955,N_17493,N_17473);
xor U17956 (N_17956,N_17243,N_17476);
xor U17957 (N_17957,N_17312,N_17282);
xor U17958 (N_17958,N_17184,N_17583);
and U17959 (N_17959,N_17595,N_17373);
nor U17960 (N_17960,N_17364,N_17225);
and U17961 (N_17961,N_16881,N_16926);
xnor U17962 (N_17962,N_16831,N_17485);
nor U17963 (N_17963,N_16820,N_16803);
nor U17964 (N_17964,N_17231,N_17105);
nor U17965 (N_17965,N_17406,N_16827);
xor U17966 (N_17966,N_17575,N_17142);
or U17967 (N_17967,N_16821,N_17141);
and U17968 (N_17968,N_17438,N_16869);
nand U17969 (N_17969,N_16938,N_17062);
or U17970 (N_17970,N_17076,N_16950);
or U17971 (N_17971,N_17115,N_17598);
nand U17972 (N_17972,N_17095,N_17535);
xnor U17973 (N_17973,N_17549,N_17137);
nand U17974 (N_17974,N_17572,N_16964);
xnor U17975 (N_17975,N_17496,N_17552);
nor U17976 (N_17976,N_17180,N_17292);
xor U17977 (N_17977,N_17488,N_17044);
nor U17978 (N_17978,N_17451,N_16993);
or U17979 (N_17979,N_17430,N_17014);
nand U17980 (N_17980,N_17207,N_16829);
xnor U17981 (N_17981,N_17210,N_16839);
or U17982 (N_17982,N_17189,N_17334);
nor U17983 (N_17983,N_17259,N_17133);
or U17984 (N_17984,N_16903,N_17548);
or U17985 (N_17985,N_16818,N_17099);
and U17986 (N_17986,N_17448,N_17153);
nor U17987 (N_17987,N_17333,N_17330);
and U17988 (N_17988,N_17146,N_17037);
and U17989 (N_17989,N_17335,N_16807);
xnor U17990 (N_17990,N_17011,N_16835);
nand U17991 (N_17991,N_16887,N_17537);
nand U17992 (N_17992,N_16856,N_16991);
nor U17993 (N_17993,N_17538,N_17060);
or U17994 (N_17994,N_17004,N_17352);
nand U17995 (N_17995,N_17507,N_17251);
nand U17996 (N_17996,N_16935,N_17508);
nor U17997 (N_17997,N_17576,N_17562);
xnor U17998 (N_17998,N_17132,N_17454);
nor U17999 (N_17999,N_16854,N_17408);
nor U18000 (N_18000,N_16903,N_17587);
and U18001 (N_18001,N_16982,N_17312);
nor U18002 (N_18002,N_17153,N_16849);
xnor U18003 (N_18003,N_17498,N_17541);
and U18004 (N_18004,N_16856,N_17266);
and U18005 (N_18005,N_17155,N_17334);
or U18006 (N_18006,N_16950,N_16952);
nor U18007 (N_18007,N_16931,N_17356);
xnor U18008 (N_18008,N_17215,N_17197);
xnor U18009 (N_18009,N_17480,N_16884);
xor U18010 (N_18010,N_16938,N_16881);
nor U18011 (N_18011,N_17029,N_17207);
nand U18012 (N_18012,N_17515,N_16824);
nor U18013 (N_18013,N_17221,N_17246);
and U18014 (N_18014,N_17446,N_16869);
nand U18015 (N_18015,N_16875,N_17442);
nand U18016 (N_18016,N_16864,N_16817);
nor U18017 (N_18017,N_17465,N_17187);
and U18018 (N_18018,N_17298,N_17255);
xnor U18019 (N_18019,N_17334,N_17169);
or U18020 (N_18020,N_17046,N_16978);
xor U18021 (N_18021,N_16816,N_17055);
and U18022 (N_18022,N_17147,N_17066);
and U18023 (N_18023,N_17387,N_17323);
or U18024 (N_18024,N_17425,N_16900);
or U18025 (N_18025,N_17383,N_17377);
or U18026 (N_18026,N_17285,N_17161);
or U18027 (N_18027,N_17183,N_16812);
xnor U18028 (N_18028,N_16916,N_17514);
xor U18029 (N_18029,N_17158,N_17363);
nor U18030 (N_18030,N_17318,N_17164);
and U18031 (N_18031,N_17522,N_17337);
and U18032 (N_18032,N_17065,N_16943);
xor U18033 (N_18033,N_16968,N_16998);
or U18034 (N_18034,N_17593,N_17481);
xnor U18035 (N_18035,N_16809,N_17594);
xor U18036 (N_18036,N_17128,N_17270);
or U18037 (N_18037,N_17279,N_17568);
and U18038 (N_18038,N_17192,N_17348);
xnor U18039 (N_18039,N_16984,N_17308);
nand U18040 (N_18040,N_16960,N_17282);
and U18041 (N_18041,N_17382,N_17258);
and U18042 (N_18042,N_16869,N_16825);
or U18043 (N_18043,N_16865,N_16855);
nand U18044 (N_18044,N_17263,N_17521);
xnor U18045 (N_18045,N_17502,N_17052);
xnor U18046 (N_18046,N_17335,N_17136);
xnor U18047 (N_18047,N_16960,N_16806);
nand U18048 (N_18048,N_17193,N_17325);
nor U18049 (N_18049,N_17431,N_17432);
and U18050 (N_18050,N_16822,N_17285);
nor U18051 (N_18051,N_16911,N_16967);
or U18052 (N_18052,N_17555,N_17440);
or U18053 (N_18053,N_17381,N_17441);
nor U18054 (N_18054,N_16937,N_17376);
and U18055 (N_18055,N_17216,N_17376);
or U18056 (N_18056,N_16917,N_17363);
nor U18057 (N_18057,N_17574,N_17150);
and U18058 (N_18058,N_17478,N_17595);
and U18059 (N_18059,N_17403,N_17006);
nand U18060 (N_18060,N_17072,N_17541);
or U18061 (N_18061,N_17292,N_17269);
and U18062 (N_18062,N_16813,N_16977);
nor U18063 (N_18063,N_17225,N_17508);
xor U18064 (N_18064,N_17234,N_17130);
and U18065 (N_18065,N_17172,N_16972);
and U18066 (N_18066,N_17539,N_17372);
or U18067 (N_18067,N_17346,N_17278);
xnor U18068 (N_18068,N_17575,N_17106);
nor U18069 (N_18069,N_17264,N_16940);
nand U18070 (N_18070,N_16869,N_17426);
nand U18071 (N_18071,N_17233,N_16925);
nor U18072 (N_18072,N_17472,N_17391);
and U18073 (N_18073,N_16907,N_16875);
nand U18074 (N_18074,N_17389,N_17049);
nand U18075 (N_18075,N_16998,N_17025);
or U18076 (N_18076,N_16839,N_16824);
nand U18077 (N_18077,N_17278,N_16912);
nand U18078 (N_18078,N_17452,N_17123);
or U18079 (N_18079,N_17301,N_17507);
or U18080 (N_18080,N_17260,N_17225);
or U18081 (N_18081,N_17133,N_16986);
nor U18082 (N_18082,N_17383,N_16960);
nand U18083 (N_18083,N_16875,N_16839);
and U18084 (N_18084,N_16956,N_17507);
nor U18085 (N_18085,N_17541,N_16932);
nand U18086 (N_18086,N_17433,N_17229);
xor U18087 (N_18087,N_17493,N_17523);
nand U18088 (N_18088,N_16877,N_17569);
xnor U18089 (N_18089,N_17047,N_17180);
or U18090 (N_18090,N_16872,N_16943);
xor U18091 (N_18091,N_17013,N_17407);
and U18092 (N_18092,N_17379,N_17123);
or U18093 (N_18093,N_17556,N_17216);
xor U18094 (N_18094,N_17003,N_17262);
nand U18095 (N_18095,N_17313,N_16840);
and U18096 (N_18096,N_17325,N_17304);
or U18097 (N_18097,N_17279,N_17258);
and U18098 (N_18098,N_16862,N_16992);
nand U18099 (N_18099,N_16997,N_17532);
and U18100 (N_18100,N_17533,N_16884);
nand U18101 (N_18101,N_17239,N_17442);
and U18102 (N_18102,N_16827,N_17246);
xnor U18103 (N_18103,N_17261,N_17208);
or U18104 (N_18104,N_17397,N_17306);
and U18105 (N_18105,N_17319,N_17514);
and U18106 (N_18106,N_17134,N_17549);
and U18107 (N_18107,N_16968,N_17000);
and U18108 (N_18108,N_17168,N_17504);
xor U18109 (N_18109,N_17576,N_17222);
or U18110 (N_18110,N_17150,N_17589);
nand U18111 (N_18111,N_17251,N_17486);
and U18112 (N_18112,N_16858,N_17532);
and U18113 (N_18113,N_17282,N_17044);
and U18114 (N_18114,N_16895,N_16925);
and U18115 (N_18115,N_17177,N_17499);
xor U18116 (N_18116,N_17275,N_17511);
nand U18117 (N_18117,N_17554,N_16883);
nand U18118 (N_18118,N_17324,N_16861);
xor U18119 (N_18119,N_17175,N_17141);
or U18120 (N_18120,N_17476,N_16945);
nor U18121 (N_18121,N_16933,N_17484);
nor U18122 (N_18122,N_17537,N_16811);
or U18123 (N_18123,N_17414,N_17161);
or U18124 (N_18124,N_17144,N_17093);
xor U18125 (N_18125,N_17533,N_17306);
or U18126 (N_18126,N_17292,N_17095);
nand U18127 (N_18127,N_17149,N_17026);
and U18128 (N_18128,N_16827,N_17107);
and U18129 (N_18129,N_17438,N_16902);
xnor U18130 (N_18130,N_17105,N_17308);
nor U18131 (N_18131,N_17408,N_17332);
nand U18132 (N_18132,N_17479,N_17292);
nor U18133 (N_18133,N_16819,N_17220);
xor U18134 (N_18134,N_17284,N_16973);
xnor U18135 (N_18135,N_17570,N_17575);
or U18136 (N_18136,N_17569,N_17242);
or U18137 (N_18137,N_17322,N_17341);
or U18138 (N_18138,N_17145,N_17190);
xnor U18139 (N_18139,N_17150,N_17179);
or U18140 (N_18140,N_16942,N_16810);
and U18141 (N_18141,N_16975,N_17166);
nor U18142 (N_18142,N_16880,N_17094);
or U18143 (N_18143,N_17541,N_17109);
nor U18144 (N_18144,N_17562,N_16803);
or U18145 (N_18145,N_17384,N_17021);
xor U18146 (N_18146,N_17031,N_16883);
and U18147 (N_18147,N_17223,N_16908);
or U18148 (N_18148,N_17126,N_17335);
or U18149 (N_18149,N_17156,N_17002);
nand U18150 (N_18150,N_17356,N_17270);
xnor U18151 (N_18151,N_17461,N_16983);
nor U18152 (N_18152,N_17205,N_17151);
xnor U18153 (N_18153,N_16961,N_16905);
or U18154 (N_18154,N_17505,N_17413);
xnor U18155 (N_18155,N_17157,N_17421);
nand U18156 (N_18156,N_17121,N_17316);
nor U18157 (N_18157,N_16907,N_17072);
nand U18158 (N_18158,N_17272,N_17052);
xnor U18159 (N_18159,N_17027,N_16901);
or U18160 (N_18160,N_17476,N_17321);
xnor U18161 (N_18161,N_16874,N_17310);
nand U18162 (N_18162,N_17584,N_17293);
nor U18163 (N_18163,N_16922,N_17322);
xor U18164 (N_18164,N_17320,N_17415);
or U18165 (N_18165,N_16901,N_17147);
and U18166 (N_18166,N_17025,N_17010);
and U18167 (N_18167,N_17381,N_17106);
xor U18168 (N_18168,N_17293,N_17080);
and U18169 (N_18169,N_17279,N_17530);
or U18170 (N_18170,N_16895,N_17343);
nor U18171 (N_18171,N_17112,N_17060);
nand U18172 (N_18172,N_17401,N_17137);
nor U18173 (N_18173,N_17118,N_17301);
or U18174 (N_18174,N_17262,N_17424);
nor U18175 (N_18175,N_17145,N_17091);
nand U18176 (N_18176,N_17024,N_17317);
and U18177 (N_18177,N_16989,N_17324);
or U18178 (N_18178,N_16854,N_17544);
nor U18179 (N_18179,N_17364,N_16964);
nor U18180 (N_18180,N_17241,N_16838);
nand U18181 (N_18181,N_17032,N_17100);
or U18182 (N_18182,N_17155,N_17427);
nor U18183 (N_18183,N_17303,N_17177);
and U18184 (N_18184,N_17105,N_17320);
and U18185 (N_18185,N_16832,N_16898);
and U18186 (N_18186,N_17315,N_17360);
and U18187 (N_18187,N_17060,N_17040);
and U18188 (N_18188,N_17448,N_17562);
nand U18189 (N_18189,N_17361,N_17269);
nor U18190 (N_18190,N_16988,N_16826);
or U18191 (N_18191,N_17132,N_17340);
xor U18192 (N_18192,N_17083,N_17089);
or U18193 (N_18193,N_17471,N_16913);
nand U18194 (N_18194,N_17142,N_16984);
and U18195 (N_18195,N_16804,N_17397);
nor U18196 (N_18196,N_17569,N_17581);
nand U18197 (N_18197,N_17449,N_16835);
nand U18198 (N_18198,N_17181,N_17202);
nor U18199 (N_18199,N_17414,N_17502);
nand U18200 (N_18200,N_17346,N_17428);
and U18201 (N_18201,N_16838,N_17117);
xnor U18202 (N_18202,N_17265,N_17113);
and U18203 (N_18203,N_17041,N_16806);
xnor U18204 (N_18204,N_17589,N_17192);
xor U18205 (N_18205,N_17044,N_17279);
or U18206 (N_18206,N_17471,N_17308);
nand U18207 (N_18207,N_17195,N_17371);
nor U18208 (N_18208,N_16887,N_17132);
xor U18209 (N_18209,N_16960,N_17433);
and U18210 (N_18210,N_17098,N_17398);
and U18211 (N_18211,N_17287,N_17391);
xnor U18212 (N_18212,N_17509,N_17558);
or U18213 (N_18213,N_16802,N_17553);
nor U18214 (N_18214,N_17302,N_16854);
or U18215 (N_18215,N_16841,N_16844);
or U18216 (N_18216,N_17037,N_17201);
nand U18217 (N_18217,N_16980,N_17301);
or U18218 (N_18218,N_17574,N_16800);
or U18219 (N_18219,N_17334,N_17399);
or U18220 (N_18220,N_17341,N_17102);
nand U18221 (N_18221,N_17140,N_17069);
and U18222 (N_18222,N_16906,N_16824);
nor U18223 (N_18223,N_17176,N_17263);
nor U18224 (N_18224,N_17203,N_17055);
xnor U18225 (N_18225,N_17122,N_17217);
xnor U18226 (N_18226,N_16847,N_17267);
nor U18227 (N_18227,N_17234,N_16953);
nand U18228 (N_18228,N_17001,N_17142);
nand U18229 (N_18229,N_17590,N_17092);
nand U18230 (N_18230,N_17577,N_17428);
xor U18231 (N_18231,N_17076,N_17509);
nand U18232 (N_18232,N_17261,N_17492);
nor U18233 (N_18233,N_17074,N_16844);
nand U18234 (N_18234,N_17589,N_17005);
or U18235 (N_18235,N_17379,N_17083);
and U18236 (N_18236,N_16877,N_17043);
nand U18237 (N_18237,N_17202,N_16858);
nand U18238 (N_18238,N_16860,N_17348);
or U18239 (N_18239,N_17454,N_16960);
or U18240 (N_18240,N_17066,N_17508);
nor U18241 (N_18241,N_17188,N_17339);
xnor U18242 (N_18242,N_16966,N_17021);
and U18243 (N_18243,N_17122,N_17187);
xor U18244 (N_18244,N_17525,N_17545);
nor U18245 (N_18245,N_17105,N_16941);
nor U18246 (N_18246,N_17429,N_17005);
and U18247 (N_18247,N_17462,N_17551);
xor U18248 (N_18248,N_17399,N_17413);
nand U18249 (N_18249,N_17073,N_17336);
nor U18250 (N_18250,N_17293,N_17216);
nand U18251 (N_18251,N_17311,N_17127);
xnor U18252 (N_18252,N_16989,N_17245);
xnor U18253 (N_18253,N_16969,N_17141);
nand U18254 (N_18254,N_17289,N_17142);
or U18255 (N_18255,N_17368,N_17190);
or U18256 (N_18256,N_17371,N_17566);
nor U18257 (N_18257,N_17077,N_17578);
nand U18258 (N_18258,N_17327,N_17490);
nor U18259 (N_18259,N_17073,N_16906);
nor U18260 (N_18260,N_16801,N_17192);
nand U18261 (N_18261,N_17441,N_17030);
xnor U18262 (N_18262,N_17020,N_17199);
xor U18263 (N_18263,N_17527,N_16944);
and U18264 (N_18264,N_17461,N_17021);
or U18265 (N_18265,N_17463,N_16851);
xor U18266 (N_18266,N_16827,N_17276);
or U18267 (N_18267,N_17333,N_17530);
or U18268 (N_18268,N_17344,N_17535);
xor U18269 (N_18269,N_17149,N_17451);
or U18270 (N_18270,N_16930,N_17491);
nand U18271 (N_18271,N_17102,N_17354);
or U18272 (N_18272,N_17039,N_16867);
nor U18273 (N_18273,N_17326,N_17314);
xor U18274 (N_18274,N_16865,N_16990);
and U18275 (N_18275,N_17073,N_17396);
and U18276 (N_18276,N_17300,N_16964);
xnor U18277 (N_18277,N_16978,N_17300);
xnor U18278 (N_18278,N_16866,N_17271);
xnor U18279 (N_18279,N_17169,N_17314);
or U18280 (N_18280,N_17407,N_17569);
xor U18281 (N_18281,N_17341,N_17196);
nor U18282 (N_18282,N_17058,N_17394);
nand U18283 (N_18283,N_17194,N_17521);
and U18284 (N_18284,N_17188,N_17261);
or U18285 (N_18285,N_17154,N_16826);
or U18286 (N_18286,N_17170,N_17532);
nand U18287 (N_18287,N_17094,N_17005);
nand U18288 (N_18288,N_17188,N_17418);
nand U18289 (N_18289,N_17015,N_16886);
and U18290 (N_18290,N_16912,N_16864);
xnor U18291 (N_18291,N_17002,N_16907);
nand U18292 (N_18292,N_17198,N_17540);
and U18293 (N_18293,N_17208,N_17572);
and U18294 (N_18294,N_17287,N_17206);
or U18295 (N_18295,N_17164,N_17145);
and U18296 (N_18296,N_17245,N_17082);
nor U18297 (N_18297,N_16958,N_17243);
and U18298 (N_18298,N_17377,N_17546);
and U18299 (N_18299,N_16928,N_17475);
nor U18300 (N_18300,N_17194,N_17579);
nand U18301 (N_18301,N_17068,N_16850);
xor U18302 (N_18302,N_17581,N_17234);
or U18303 (N_18303,N_16818,N_17579);
xnor U18304 (N_18304,N_17564,N_17356);
and U18305 (N_18305,N_17417,N_17032);
nor U18306 (N_18306,N_17016,N_16852);
xor U18307 (N_18307,N_16993,N_16920);
xor U18308 (N_18308,N_17161,N_17167);
nor U18309 (N_18309,N_17000,N_17026);
nor U18310 (N_18310,N_16963,N_17311);
and U18311 (N_18311,N_17366,N_16912);
xor U18312 (N_18312,N_16969,N_17419);
or U18313 (N_18313,N_17420,N_17115);
and U18314 (N_18314,N_17015,N_17184);
or U18315 (N_18315,N_17255,N_17320);
xnor U18316 (N_18316,N_17073,N_17141);
or U18317 (N_18317,N_17320,N_17090);
nand U18318 (N_18318,N_16979,N_16893);
or U18319 (N_18319,N_16933,N_17399);
and U18320 (N_18320,N_17019,N_17550);
or U18321 (N_18321,N_16876,N_17385);
or U18322 (N_18322,N_17184,N_16913);
and U18323 (N_18323,N_17147,N_17369);
or U18324 (N_18324,N_16903,N_17432);
nor U18325 (N_18325,N_17205,N_17208);
and U18326 (N_18326,N_17272,N_17569);
xor U18327 (N_18327,N_17528,N_16864);
xor U18328 (N_18328,N_17406,N_17030);
and U18329 (N_18329,N_17472,N_17543);
nand U18330 (N_18330,N_16861,N_17171);
or U18331 (N_18331,N_17402,N_17533);
or U18332 (N_18332,N_16986,N_17208);
nand U18333 (N_18333,N_17484,N_17463);
and U18334 (N_18334,N_17089,N_16967);
or U18335 (N_18335,N_17038,N_16928);
and U18336 (N_18336,N_17150,N_17258);
and U18337 (N_18337,N_17076,N_17051);
and U18338 (N_18338,N_17011,N_17572);
and U18339 (N_18339,N_16898,N_16839);
nor U18340 (N_18340,N_17317,N_17396);
and U18341 (N_18341,N_16918,N_17007);
nand U18342 (N_18342,N_17124,N_17473);
or U18343 (N_18343,N_17412,N_17172);
nand U18344 (N_18344,N_16884,N_17371);
and U18345 (N_18345,N_16830,N_17172);
or U18346 (N_18346,N_17558,N_17213);
nor U18347 (N_18347,N_17104,N_17098);
xnor U18348 (N_18348,N_17591,N_17050);
nand U18349 (N_18349,N_17479,N_17552);
nor U18350 (N_18350,N_16856,N_17338);
nor U18351 (N_18351,N_16915,N_17254);
nor U18352 (N_18352,N_17483,N_17503);
and U18353 (N_18353,N_17153,N_17232);
nand U18354 (N_18354,N_17252,N_17211);
or U18355 (N_18355,N_17102,N_16809);
nor U18356 (N_18356,N_17166,N_16866);
nor U18357 (N_18357,N_17167,N_16914);
nand U18358 (N_18358,N_17071,N_17590);
xor U18359 (N_18359,N_17469,N_17555);
nand U18360 (N_18360,N_16902,N_17595);
or U18361 (N_18361,N_17321,N_17365);
and U18362 (N_18362,N_17093,N_17244);
or U18363 (N_18363,N_17014,N_17477);
xor U18364 (N_18364,N_16846,N_17058);
nand U18365 (N_18365,N_17457,N_17520);
nand U18366 (N_18366,N_16855,N_17101);
nand U18367 (N_18367,N_17542,N_16960);
nor U18368 (N_18368,N_17374,N_17105);
and U18369 (N_18369,N_16986,N_17258);
nor U18370 (N_18370,N_17030,N_16873);
or U18371 (N_18371,N_17465,N_17079);
nand U18372 (N_18372,N_17119,N_17228);
nor U18373 (N_18373,N_17254,N_17173);
nand U18374 (N_18374,N_17293,N_17096);
nand U18375 (N_18375,N_17265,N_16842);
or U18376 (N_18376,N_17219,N_17490);
nor U18377 (N_18377,N_17581,N_17295);
nand U18378 (N_18378,N_17528,N_16853);
nor U18379 (N_18379,N_17209,N_17510);
and U18380 (N_18380,N_16820,N_17585);
nand U18381 (N_18381,N_16951,N_17371);
nand U18382 (N_18382,N_17148,N_16904);
nand U18383 (N_18383,N_17590,N_17405);
or U18384 (N_18384,N_17387,N_17226);
or U18385 (N_18385,N_17308,N_16916);
and U18386 (N_18386,N_17101,N_17575);
nor U18387 (N_18387,N_16809,N_17566);
nand U18388 (N_18388,N_16916,N_16896);
or U18389 (N_18389,N_17372,N_17517);
nand U18390 (N_18390,N_17338,N_17084);
or U18391 (N_18391,N_17238,N_17340);
and U18392 (N_18392,N_17025,N_16944);
xor U18393 (N_18393,N_17115,N_17314);
nand U18394 (N_18394,N_16819,N_17212);
and U18395 (N_18395,N_17269,N_17093);
xor U18396 (N_18396,N_17257,N_17568);
and U18397 (N_18397,N_17199,N_17155);
and U18398 (N_18398,N_17483,N_17357);
nand U18399 (N_18399,N_17376,N_17036);
xor U18400 (N_18400,N_18203,N_17795);
or U18401 (N_18401,N_18068,N_18275);
nor U18402 (N_18402,N_17664,N_17810);
nor U18403 (N_18403,N_17761,N_18037);
or U18404 (N_18404,N_18289,N_18394);
nor U18405 (N_18405,N_18191,N_17684);
nor U18406 (N_18406,N_18300,N_17640);
and U18407 (N_18407,N_18237,N_17837);
and U18408 (N_18408,N_18057,N_17749);
or U18409 (N_18409,N_17843,N_17858);
nand U18410 (N_18410,N_18029,N_18109);
or U18411 (N_18411,N_17848,N_17970);
and U18412 (N_18412,N_18084,N_17708);
nor U18413 (N_18413,N_18291,N_17671);
xnor U18414 (N_18414,N_17642,N_18022);
xor U18415 (N_18415,N_18099,N_17993);
xnor U18416 (N_18416,N_18026,N_17814);
xor U18417 (N_18417,N_17672,N_17637);
nor U18418 (N_18418,N_17842,N_17887);
or U18419 (N_18419,N_17778,N_18094);
or U18420 (N_18420,N_18028,N_18149);
or U18421 (N_18421,N_17816,N_17770);
and U18422 (N_18422,N_18260,N_17994);
nand U18423 (N_18423,N_17957,N_18215);
nor U18424 (N_18424,N_17953,N_17794);
and U18425 (N_18425,N_17859,N_18176);
or U18426 (N_18426,N_18120,N_18183);
nand U18427 (N_18427,N_17905,N_17755);
nor U18428 (N_18428,N_17676,N_18238);
nor U18429 (N_18429,N_18271,N_18207);
nor U18430 (N_18430,N_18041,N_18193);
xnor U18431 (N_18431,N_17717,N_18065);
nor U18432 (N_18432,N_17720,N_17935);
and U18433 (N_18433,N_18069,N_18017);
and U18434 (N_18434,N_17906,N_18181);
and U18435 (N_18435,N_17751,N_17904);
nand U18436 (N_18436,N_18352,N_18366);
and U18437 (N_18437,N_18189,N_17765);
nor U18438 (N_18438,N_17768,N_18055);
xnor U18439 (N_18439,N_18000,N_18317);
nand U18440 (N_18440,N_17729,N_17998);
or U18441 (N_18441,N_17975,N_18110);
nor U18442 (N_18442,N_17628,N_17688);
nor U18443 (N_18443,N_17609,N_17853);
nor U18444 (N_18444,N_18249,N_18326);
nor U18445 (N_18445,N_17736,N_17883);
nor U18446 (N_18446,N_18388,N_18341);
nor U18447 (N_18447,N_18089,N_17634);
nor U18448 (N_18448,N_18395,N_18225);
and U18449 (N_18449,N_18387,N_17940);
and U18450 (N_18450,N_17682,N_18266);
xnor U18451 (N_18451,N_18383,N_17888);
nand U18452 (N_18452,N_17959,N_18036);
nand U18453 (N_18453,N_17660,N_17697);
xnor U18454 (N_18454,N_18126,N_17808);
nand U18455 (N_18455,N_18391,N_17614);
xor U18456 (N_18456,N_17833,N_18111);
and U18457 (N_18457,N_17972,N_17866);
xor U18458 (N_18458,N_18038,N_18075);
xnor U18459 (N_18459,N_18121,N_18321);
nor U18460 (N_18460,N_18081,N_18045);
xnor U18461 (N_18461,N_17695,N_17698);
nor U18462 (N_18462,N_18315,N_18286);
or U18463 (N_18463,N_17613,N_18245);
nand U18464 (N_18464,N_17659,N_17675);
nand U18465 (N_18465,N_17780,N_17629);
and U18466 (N_18466,N_18323,N_17608);
xnor U18467 (N_18467,N_18169,N_17856);
nand U18468 (N_18468,N_17707,N_18064);
nand U18469 (N_18469,N_17841,N_18370);
xnor U18470 (N_18470,N_17645,N_18309);
and U18471 (N_18471,N_18033,N_17644);
xor U18472 (N_18472,N_17889,N_18338);
and U18473 (N_18473,N_18122,N_17744);
nor U18474 (N_18474,N_18185,N_18170);
and U18475 (N_18475,N_17763,N_18293);
nand U18476 (N_18476,N_17896,N_18213);
nor U18477 (N_18477,N_17611,N_18005);
nor U18478 (N_18478,N_18374,N_18197);
xor U18479 (N_18479,N_17944,N_18124);
nor U18480 (N_18480,N_17665,N_17724);
or U18481 (N_18481,N_18337,N_18159);
nand U18482 (N_18482,N_18103,N_18048);
or U18483 (N_18483,N_17828,N_17850);
and U18484 (N_18484,N_17928,N_18231);
xor U18485 (N_18485,N_17683,N_18371);
nand U18486 (N_18486,N_17890,N_18192);
and U18487 (N_18487,N_18272,N_18161);
and U18488 (N_18488,N_17949,N_17711);
nor U18489 (N_18489,N_17908,N_18131);
xor U18490 (N_18490,N_18186,N_18102);
and U18491 (N_18491,N_18072,N_17978);
xnor U18492 (N_18492,N_18206,N_17967);
or U18493 (N_18493,N_17825,N_17867);
xor U18494 (N_18494,N_18117,N_17690);
nor U18495 (N_18495,N_17956,N_18182);
xor U18496 (N_18496,N_18001,N_18040);
or U18497 (N_18497,N_17689,N_18107);
xor U18498 (N_18498,N_17741,N_18021);
or U18499 (N_18499,N_18244,N_17855);
nand U18500 (N_18500,N_18187,N_18158);
or U18501 (N_18501,N_17982,N_17840);
nor U18502 (N_18502,N_18322,N_18018);
nor U18503 (N_18503,N_17791,N_18328);
xor U18504 (N_18504,N_17925,N_17836);
nor U18505 (N_18505,N_18228,N_18138);
xor U18506 (N_18506,N_17983,N_18344);
or U18507 (N_18507,N_17649,N_18195);
nor U18508 (N_18508,N_17678,N_18240);
nor U18509 (N_18509,N_17785,N_18091);
xnor U18510 (N_18510,N_18024,N_18135);
and U18511 (N_18511,N_17961,N_17827);
nor U18512 (N_18512,N_18320,N_17880);
nand U18513 (N_18513,N_18397,N_18178);
nand U18514 (N_18514,N_18205,N_17702);
nor U18515 (N_18515,N_18330,N_17913);
nand U18516 (N_18516,N_18252,N_18230);
nor U18517 (N_18517,N_17835,N_17705);
nand U18518 (N_18518,N_18285,N_17799);
nand U18519 (N_18519,N_17782,N_18379);
nor U18520 (N_18520,N_17803,N_18044);
nand U18521 (N_18521,N_17938,N_17726);
nand U18522 (N_18522,N_17960,N_18127);
or U18523 (N_18523,N_18118,N_18167);
or U18524 (N_18524,N_17604,N_18092);
nor U18525 (N_18525,N_18373,N_18332);
or U18526 (N_18526,N_18253,N_18292);
or U18527 (N_18527,N_18198,N_17712);
nand U18528 (N_18528,N_18232,N_17710);
nand U18529 (N_18529,N_18350,N_18058);
nor U18530 (N_18530,N_18247,N_18347);
and U18531 (N_18531,N_17945,N_17621);
and U18532 (N_18532,N_18047,N_18223);
nand U18533 (N_18533,N_17931,N_17605);
nand U18534 (N_18534,N_18273,N_18156);
nand U18535 (N_18535,N_17882,N_17876);
nand U18536 (N_18536,N_17666,N_17701);
nor U18537 (N_18537,N_17815,N_18208);
xnor U18538 (N_18538,N_18357,N_18319);
xor U18539 (N_18539,N_17654,N_17921);
and U18540 (N_18540,N_17910,N_18339);
and U18541 (N_18541,N_17631,N_18359);
nand U18542 (N_18542,N_18151,N_17679);
xor U18543 (N_18543,N_18278,N_17740);
and U18544 (N_18544,N_18296,N_17879);
and U18545 (N_18545,N_17725,N_17894);
and U18546 (N_18546,N_17977,N_17900);
or U18547 (N_18547,N_17746,N_17764);
xor U18548 (N_18548,N_17706,N_17812);
xor U18549 (N_18549,N_17811,N_18051);
and U18550 (N_18550,N_18035,N_18140);
nand U18551 (N_18551,N_18386,N_18380);
xnor U18552 (N_18552,N_17809,N_18003);
or U18553 (N_18553,N_17777,N_17694);
or U18554 (N_18554,N_17932,N_17759);
nor U18555 (N_18555,N_18087,N_17719);
xor U18556 (N_18556,N_18020,N_18025);
nand U18557 (N_18557,N_18325,N_17875);
nor U18558 (N_18558,N_18053,N_18190);
and U18559 (N_18559,N_17699,N_18175);
and U18560 (N_18560,N_18153,N_18141);
xnor U18561 (N_18561,N_17730,N_17796);
and U18562 (N_18562,N_17847,N_18262);
nor U18563 (N_18563,N_18369,N_17807);
xor U18564 (N_18564,N_18258,N_18304);
nand U18565 (N_18565,N_17832,N_17602);
or U18566 (N_18566,N_18265,N_17732);
nand U18567 (N_18567,N_17797,N_17754);
nor U18568 (N_18568,N_17926,N_18201);
nor U18569 (N_18569,N_18148,N_17692);
or U18570 (N_18570,N_18060,N_17958);
or U18571 (N_18571,N_17622,N_18168);
nor U18572 (N_18572,N_18254,N_18125);
nand U18573 (N_18573,N_17750,N_18171);
and U18574 (N_18574,N_17851,N_18200);
xor U18575 (N_18575,N_18002,N_18362);
nor U18576 (N_18576,N_18080,N_18165);
xor U18577 (N_18577,N_17618,N_18384);
nand U18578 (N_18578,N_17999,N_18105);
nand U18579 (N_18579,N_17673,N_18006);
xnor U18580 (N_18580,N_18363,N_18399);
nor U18581 (N_18581,N_18016,N_17868);
and U18582 (N_18582,N_18355,N_18222);
and U18583 (N_18583,N_18004,N_18358);
or U18584 (N_18584,N_18155,N_18160);
and U18585 (N_18585,N_18210,N_17722);
xor U18586 (N_18586,N_17947,N_18389);
nand U18587 (N_18587,N_17737,N_18385);
nand U18588 (N_18588,N_18276,N_18052);
nor U18589 (N_18589,N_17757,N_18378);
nand U18590 (N_18590,N_18137,N_17892);
xor U18591 (N_18591,N_17930,N_18219);
xor U18592 (N_18592,N_17929,N_17802);
nor U18593 (N_18593,N_17820,N_18393);
xor U18594 (N_18594,N_17728,N_17806);
and U18595 (N_18595,N_17909,N_18014);
xor U18596 (N_18596,N_17774,N_18015);
nand U18597 (N_18597,N_18318,N_18246);
xor U18598 (N_18598,N_18164,N_17919);
nor U18599 (N_18599,N_18129,N_17838);
nor U18600 (N_18600,N_18209,N_17687);
nand U18601 (N_18601,N_18039,N_17821);
nand U18602 (N_18602,N_18196,N_18177);
and U18603 (N_18603,N_17917,N_18070);
nor U18604 (N_18604,N_17893,N_17667);
and U18605 (N_18605,N_17901,N_17980);
xor U18606 (N_18606,N_17603,N_18360);
or U18607 (N_18607,N_17834,N_18263);
and U18608 (N_18608,N_18382,N_18241);
xor U18609 (N_18609,N_18180,N_17756);
nand U18610 (N_18610,N_17787,N_17996);
nand U18611 (N_18611,N_17963,N_18329);
nand U18612 (N_18612,N_18308,N_17771);
nand U18613 (N_18613,N_18216,N_18130);
xor U18614 (N_18614,N_18023,N_17647);
xnor U18615 (N_18615,N_17788,N_18335);
or U18616 (N_18616,N_18157,N_17748);
and U18617 (N_18617,N_18085,N_18088);
or U18618 (N_18618,N_18123,N_18287);
nor U18619 (N_18619,N_17624,N_18364);
and U18620 (N_18620,N_18256,N_18234);
nor U18621 (N_18621,N_17987,N_17627);
xor U18622 (N_18622,N_18143,N_17601);
and U18623 (N_18623,N_18145,N_18340);
nand U18624 (N_18624,N_18239,N_17641);
xnor U18625 (N_18625,N_18361,N_17860);
and U18626 (N_18626,N_17844,N_18007);
or U18627 (N_18627,N_17658,N_18298);
nand U18628 (N_18628,N_17669,N_18073);
xnor U18629 (N_18629,N_18257,N_17817);
or U18630 (N_18630,N_17704,N_17918);
or U18631 (N_18631,N_17826,N_17630);
nor U18632 (N_18632,N_18013,N_18199);
nor U18633 (N_18633,N_18101,N_17648);
and U18634 (N_18634,N_18316,N_17965);
or U18635 (N_18635,N_17973,N_18248);
xnor U18636 (N_18636,N_17864,N_17862);
nand U18637 (N_18637,N_17937,N_18331);
or U18638 (N_18638,N_17916,N_18349);
nand U18639 (N_18639,N_18184,N_18313);
xor U18640 (N_18640,N_17646,N_17995);
xor U18641 (N_18641,N_18348,N_18311);
nor U18642 (N_18642,N_18019,N_18056);
and U18643 (N_18643,N_18119,N_17709);
nand U18644 (N_18644,N_17985,N_17869);
or U18645 (N_18645,N_17877,N_17721);
or U18646 (N_18646,N_17952,N_18172);
or U18647 (N_18647,N_17767,N_17951);
xnor U18648 (N_18648,N_17903,N_18284);
and U18649 (N_18649,N_18297,N_17685);
nand U18650 (N_18650,N_17779,N_18303);
nor U18651 (N_18651,N_17912,N_17792);
nand U18652 (N_18652,N_18063,N_18093);
nor U18653 (N_18653,N_17992,N_17703);
xnor U18654 (N_18654,N_18220,N_17943);
xor U18655 (N_18655,N_17638,N_17619);
and U18656 (N_18656,N_17881,N_17739);
and U18657 (N_18657,N_18235,N_17784);
and U18658 (N_18658,N_17760,N_17899);
or U18659 (N_18659,N_18226,N_18031);
and U18660 (N_18660,N_18116,N_18012);
nor U18661 (N_18661,N_18142,N_17733);
and U18662 (N_18662,N_18377,N_18345);
xor U18663 (N_18663,N_17715,N_18295);
xor U18664 (N_18664,N_18146,N_17823);
nand U18665 (N_18665,N_17902,N_17924);
nor U18666 (N_18666,N_18030,N_18312);
nand U18667 (N_18667,N_18221,N_17933);
or U18668 (N_18668,N_17955,N_18283);
nor U18669 (N_18669,N_18390,N_17606);
nand U18670 (N_18670,N_17735,N_17969);
and U18671 (N_18671,N_17886,N_17773);
nor U18672 (N_18672,N_18128,N_18368);
nand U18673 (N_18673,N_18305,N_18212);
or U18674 (N_18674,N_17650,N_18067);
xnor U18675 (N_18675,N_17745,N_18071);
xnor U18676 (N_18676,N_17878,N_17623);
nand U18677 (N_18677,N_18314,N_17632);
and U18678 (N_18678,N_17873,N_17670);
and U18679 (N_18679,N_18346,N_18268);
nor U18680 (N_18680,N_18261,N_17655);
or U18681 (N_18681,N_18100,N_17661);
and U18682 (N_18682,N_18288,N_17845);
nor U18683 (N_18683,N_17793,N_18375);
nor U18684 (N_18684,N_18396,N_17968);
xor U18685 (N_18685,N_18299,N_18301);
and U18686 (N_18686,N_18162,N_17798);
nand U18687 (N_18687,N_17716,N_18367);
or U18688 (N_18688,N_17984,N_17907);
and U18689 (N_18689,N_17997,N_17936);
or U18690 (N_18690,N_17783,N_17865);
nand U18691 (N_18691,N_17942,N_18166);
nor U18692 (N_18692,N_17731,N_18062);
nand U18693 (N_18693,N_18202,N_18043);
xnor U18694 (N_18694,N_18270,N_17839);
nand U18695 (N_18695,N_17789,N_18115);
nand U18696 (N_18696,N_17686,N_18104);
or U18697 (N_18697,N_17633,N_18277);
xnor U18698 (N_18698,N_18302,N_18090);
xnor U18699 (N_18699,N_17610,N_17656);
xnor U18700 (N_18700,N_17693,N_17713);
nand U18701 (N_18701,N_18034,N_18010);
nand U18702 (N_18702,N_17822,N_18061);
and U18703 (N_18703,N_18398,N_18274);
nor U18704 (N_18704,N_17954,N_17920);
and U18705 (N_18705,N_17691,N_18133);
nand U18706 (N_18706,N_17897,N_18009);
nor U18707 (N_18707,N_17852,N_17818);
nor U18708 (N_18708,N_18174,N_18076);
nor U18709 (N_18709,N_17871,N_18327);
nand U18710 (N_18710,N_17747,N_17643);
and U18711 (N_18711,N_17800,N_18279);
or U18712 (N_18712,N_17657,N_17663);
xor U18713 (N_18713,N_18008,N_18086);
nand U18714 (N_18714,N_17941,N_18066);
xor U18715 (N_18715,N_18233,N_17762);
nor U18716 (N_18716,N_17861,N_17766);
nand U18717 (N_18717,N_17652,N_17950);
and U18718 (N_18718,N_17829,N_18097);
nor U18719 (N_18719,N_17742,N_17976);
xor U18720 (N_18720,N_17846,N_18144);
nor U18721 (N_18721,N_17769,N_17922);
or U18722 (N_18722,N_18049,N_18251);
or U18723 (N_18723,N_18334,N_18027);
xor U18724 (N_18724,N_17651,N_18333);
nand U18725 (N_18725,N_18154,N_17819);
xnor U18726 (N_18726,N_18059,N_18294);
xor U18727 (N_18727,N_18204,N_17625);
nor U18728 (N_18728,N_17989,N_18214);
or U18729 (N_18729,N_17612,N_18324);
nand U18730 (N_18730,N_18078,N_18243);
and U18731 (N_18731,N_17934,N_18163);
or U18732 (N_18732,N_18343,N_18269);
and U18733 (N_18733,N_17966,N_18113);
nor U18734 (N_18734,N_18042,N_17971);
nor U18735 (N_18735,N_18074,N_17813);
nor U18736 (N_18736,N_17991,N_17885);
nor U18737 (N_18737,N_17626,N_17636);
nor U18738 (N_18738,N_18106,N_17668);
or U18739 (N_18739,N_17915,N_17831);
nand U18740 (N_18740,N_18376,N_17653);
and U18741 (N_18741,N_17981,N_17600);
or U18742 (N_18742,N_17635,N_17734);
or U18743 (N_18743,N_18227,N_18336);
xor U18744 (N_18744,N_17979,N_17854);
xor U18745 (N_18745,N_17804,N_18306);
or U18746 (N_18746,N_18079,N_18259);
or U18747 (N_18747,N_18098,N_17617);
nor U18748 (N_18748,N_17857,N_17898);
and U18749 (N_18749,N_18342,N_18307);
xnor U18750 (N_18750,N_17988,N_18108);
or U18751 (N_18751,N_17781,N_17738);
or U18752 (N_18752,N_17946,N_17805);
or U18753 (N_18753,N_17962,N_17615);
xnor U18754 (N_18754,N_18083,N_18267);
nand U18755 (N_18755,N_17874,N_18114);
nor U18756 (N_18756,N_17700,N_17616);
xnor U18757 (N_18757,N_18372,N_17743);
nor U18758 (N_18758,N_18011,N_17986);
or U18759 (N_18759,N_18032,N_17872);
or U18760 (N_18760,N_18381,N_18281);
and U18761 (N_18761,N_18282,N_18392);
nor U18762 (N_18762,N_18136,N_18179);
or U18763 (N_18763,N_18353,N_18218);
nand U18764 (N_18764,N_18147,N_17758);
nand U18765 (N_18765,N_17753,N_17662);
nand U18766 (N_18766,N_18050,N_18236);
and U18767 (N_18767,N_18242,N_18217);
or U18768 (N_18768,N_18310,N_17775);
and U18769 (N_18769,N_17927,N_18211);
nor U18770 (N_18770,N_18264,N_17824);
xnor U18771 (N_18771,N_17891,N_18290);
nor U18772 (N_18772,N_18365,N_17849);
nor U18773 (N_18773,N_18095,N_17801);
or U18774 (N_18774,N_18112,N_17776);
or U18775 (N_18775,N_18229,N_17607);
and U18776 (N_18776,N_17727,N_17790);
xor U18777 (N_18777,N_17964,N_17639);
xnor U18778 (N_18778,N_18082,N_18152);
or U18779 (N_18779,N_18250,N_18096);
or U18780 (N_18780,N_18280,N_18139);
nand U18781 (N_18781,N_17884,N_17870);
or U18782 (N_18782,N_18150,N_17696);
or U18783 (N_18783,N_17974,N_18224);
nor U18784 (N_18784,N_17681,N_17914);
nor U18785 (N_18785,N_18354,N_18054);
nand U18786 (N_18786,N_17863,N_17752);
nand U18787 (N_18787,N_18132,N_18077);
xnor U18788 (N_18788,N_17786,N_17680);
nand U18789 (N_18789,N_17723,N_18351);
or U18790 (N_18790,N_17895,N_17911);
nand U18791 (N_18791,N_17674,N_18046);
xor U18792 (N_18792,N_18194,N_17939);
nor U18793 (N_18793,N_18356,N_17677);
xnor U18794 (N_18794,N_17923,N_18255);
nor U18795 (N_18795,N_17620,N_17714);
nand U18796 (N_18796,N_17830,N_17718);
nor U18797 (N_18797,N_18188,N_17990);
nand U18798 (N_18798,N_18134,N_17948);
and U18799 (N_18799,N_18173,N_17772);
nor U18800 (N_18800,N_18171,N_17626);
and U18801 (N_18801,N_17959,N_18147);
and U18802 (N_18802,N_17648,N_18187);
xor U18803 (N_18803,N_18189,N_18260);
xor U18804 (N_18804,N_17878,N_17792);
xnor U18805 (N_18805,N_18329,N_17872);
or U18806 (N_18806,N_18158,N_18266);
or U18807 (N_18807,N_17808,N_17947);
nor U18808 (N_18808,N_18012,N_17669);
nand U18809 (N_18809,N_17960,N_17812);
xor U18810 (N_18810,N_18323,N_17993);
xor U18811 (N_18811,N_18261,N_17870);
nor U18812 (N_18812,N_18146,N_17917);
nor U18813 (N_18813,N_17758,N_17648);
and U18814 (N_18814,N_18329,N_17628);
xnor U18815 (N_18815,N_17707,N_17845);
nor U18816 (N_18816,N_18166,N_17754);
nand U18817 (N_18817,N_18023,N_18228);
xnor U18818 (N_18818,N_17740,N_18334);
nor U18819 (N_18819,N_18284,N_18161);
or U18820 (N_18820,N_17687,N_17675);
or U18821 (N_18821,N_18083,N_17905);
xnor U18822 (N_18822,N_18055,N_18310);
nor U18823 (N_18823,N_17685,N_17953);
xnor U18824 (N_18824,N_18112,N_17976);
nand U18825 (N_18825,N_18078,N_18193);
nor U18826 (N_18826,N_18234,N_17718);
xor U18827 (N_18827,N_17661,N_17607);
nand U18828 (N_18828,N_18026,N_18130);
and U18829 (N_18829,N_17804,N_18379);
or U18830 (N_18830,N_17628,N_18144);
or U18831 (N_18831,N_17692,N_18022);
nor U18832 (N_18832,N_18058,N_18214);
and U18833 (N_18833,N_18291,N_18010);
nand U18834 (N_18834,N_17692,N_18270);
nand U18835 (N_18835,N_18228,N_18205);
or U18836 (N_18836,N_18064,N_18160);
and U18837 (N_18837,N_18367,N_18096);
or U18838 (N_18838,N_17838,N_18034);
nor U18839 (N_18839,N_18168,N_17911);
nand U18840 (N_18840,N_18331,N_17838);
nand U18841 (N_18841,N_17622,N_18395);
nor U18842 (N_18842,N_17840,N_17796);
and U18843 (N_18843,N_18288,N_17691);
nor U18844 (N_18844,N_18283,N_18323);
xor U18845 (N_18845,N_17757,N_18109);
nor U18846 (N_18846,N_18372,N_17938);
nor U18847 (N_18847,N_18019,N_18096);
and U18848 (N_18848,N_18198,N_18284);
and U18849 (N_18849,N_18182,N_17786);
or U18850 (N_18850,N_18239,N_18148);
xnor U18851 (N_18851,N_18070,N_18084);
and U18852 (N_18852,N_18141,N_17702);
nand U18853 (N_18853,N_18010,N_17688);
xnor U18854 (N_18854,N_18071,N_18235);
or U18855 (N_18855,N_18155,N_18301);
nor U18856 (N_18856,N_18392,N_18215);
xor U18857 (N_18857,N_18177,N_18230);
or U18858 (N_18858,N_17764,N_17707);
and U18859 (N_18859,N_17950,N_17853);
and U18860 (N_18860,N_17898,N_18066);
and U18861 (N_18861,N_17917,N_17797);
nand U18862 (N_18862,N_18010,N_17843);
and U18863 (N_18863,N_18205,N_17689);
and U18864 (N_18864,N_17898,N_18206);
xor U18865 (N_18865,N_17910,N_17981);
nor U18866 (N_18866,N_17732,N_17949);
and U18867 (N_18867,N_18293,N_17934);
nor U18868 (N_18868,N_17822,N_18224);
and U18869 (N_18869,N_17963,N_18312);
or U18870 (N_18870,N_18327,N_18143);
nand U18871 (N_18871,N_17676,N_17639);
and U18872 (N_18872,N_17903,N_18196);
nand U18873 (N_18873,N_17804,N_18196);
nand U18874 (N_18874,N_17602,N_18364);
xor U18875 (N_18875,N_18287,N_17613);
or U18876 (N_18876,N_17662,N_17766);
nand U18877 (N_18877,N_17759,N_18177);
xnor U18878 (N_18878,N_17771,N_17850);
nand U18879 (N_18879,N_18086,N_18285);
or U18880 (N_18880,N_17622,N_18388);
or U18881 (N_18881,N_18031,N_18186);
or U18882 (N_18882,N_18166,N_17668);
and U18883 (N_18883,N_17814,N_18149);
and U18884 (N_18884,N_17665,N_17699);
and U18885 (N_18885,N_17849,N_17652);
and U18886 (N_18886,N_18014,N_18317);
nor U18887 (N_18887,N_18160,N_18300);
xnor U18888 (N_18888,N_18235,N_18181);
xnor U18889 (N_18889,N_17663,N_17747);
nor U18890 (N_18890,N_18203,N_17658);
xnor U18891 (N_18891,N_18302,N_18185);
xor U18892 (N_18892,N_17917,N_18336);
xor U18893 (N_18893,N_17666,N_17868);
nor U18894 (N_18894,N_18057,N_17868);
xor U18895 (N_18895,N_17992,N_17711);
nor U18896 (N_18896,N_17907,N_17694);
or U18897 (N_18897,N_17943,N_17835);
nand U18898 (N_18898,N_17756,N_17638);
or U18899 (N_18899,N_17916,N_17998);
nor U18900 (N_18900,N_18072,N_17806);
xnor U18901 (N_18901,N_18209,N_17893);
and U18902 (N_18902,N_17810,N_17602);
nand U18903 (N_18903,N_18169,N_18202);
xor U18904 (N_18904,N_17793,N_17716);
nand U18905 (N_18905,N_18225,N_17756);
nand U18906 (N_18906,N_18225,N_18359);
nand U18907 (N_18907,N_18343,N_18299);
nor U18908 (N_18908,N_18341,N_18195);
or U18909 (N_18909,N_18389,N_17821);
xnor U18910 (N_18910,N_18265,N_18394);
and U18911 (N_18911,N_18133,N_18034);
xnor U18912 (N_18912,N_18077,N_17793);
and U18913 (N_18913,N_18010,N_17818);
and U18914 (N_18914,N_17763,N_18355);
nor U18915 (N_18915,N_18261,N_18106);
nand U18916 (N_18916,N_18204,N_17808);
or U18917 (N_18917,N_17667,N_18130);
or U18918 (N_18918,N_18350,N_18006);
or U18919 (N_18919,N_18142,N_18213);
xnor U18920 (N_18920,N_17688,N_18040);
xnor U18921 (N_18921,N_18103,N_17637);
nand U18922 (N_18922,N_18005,N_18041);
nor U18923 (N_18923,N_17882,N_17634);
and U18924 (N_18924,N_17645,N_17971);
nand U18925 (N_18925,N_17711,N_18250);
and U18926 (N_18926,N_17715,N_18058);
or U18927 (N_18927,N_17920,N_18259);
or U18928 (N_18928,N_17810,N_18205);
or U18929 (N_18929,N_17722,N_17774);
or U18930 (N_18930,N_18271,N_18214);
or U18931 (N_18931,N_18323,N_18377);
xor U18932 (N_18932,N_18165,N_18252);
nor U18933 (N_18933,N_18115,N_18306);
xnor U18934 (N_18934,N_17683,N_17941);
xnor U18935 (N_18935,N_17651,N_18192);
nand U18936 (N_18936,N_17873,N_17652);
nand U18937 (N_18937,N_18218,N_17774);
nor U18938 (N_18938,N_18149,N_18184);
nand U18939 (N_18939,N_18035,N_17867);
and U18940 (N_18940,N_17659,N_17782);
xor U18941 (N_18941,N_17954,N_17993);
and U18942 (N_18942,N_17627,N_17852);
and U18943 (N_18943,N_17606,N_18139);
or U18944 (N_18944,N_17762,N_18278);
nor U18945 (N_18945,N_18098,N_18254);
or U18946 (N_18946,N_17974,N_17615);
or U18947 (N_18947,N_18222,N_18179);
nor U18948 (N_18948,N_17775,N_18157);
and U18949 (N_18949,N_18394,N_17717);
xor U18950 (N_18950,N_17653,N_17795);
or U18951 (N_18951,N_18197,N_17761);
and U18952 (N_18952,N_18389,N_18032);
or U18953 (N_18953,N_17874,N_17921);
or U18954 (N_18954,N_18045,N_17990);
or U18955 (N_18955,N_17822,N_18005);
xnor U18956 (N_18956,N_18278,N_18323);
xnor U18957 (N_18957,N_17749,N_17965);
xnor U18958 (N_18958,N_17768,N_17741);
nand U18959 (N_18959,N_18341,N_17765);
nand U18960 (N_18960,N_17776,N_18171);
and U18961 (N_18961,N_18324,N_18247);
nor U18962 (N_18962,N_18085,N_18352);
xnor U18963 (N_18963,N_18190,N_18268);
or U18964 (N_18964,N_18080,N_18283);
nor U18965 (N_18965,N_18046,N_18123);
or U18966 (N_18966,N_18107,N_18385);
nand U18967 (N_18967,N_18158,N_18357);
nand U18968 (N_18968,N_18277,N_18333);
xnor U18969 (N_18969,N_17643,N_18306);
and U18970 (N_18970,N_18006,N_17649);
nand U18971 (N_18971,N_18313,N_18304);
and U18972 (N_18972,N_17801,N_17649);
nor U18973 (N_18973,N_18377,N_17880);
or U18974 (N_18974,N_17951,N_17751);
nor U18975 (N_18975,N_17896,N_17736);
or U18976 (N_18976,N_17766,N_17653);
xnor U18977 (N_18977,N_17601,N_18126);
xnor U18978 (N_18978,N_17961,N_17794);
and U18979 (N_18979,N_18343,N_17718);
and U18980 (N_18980,N_17819,N_18078);
nor U18981 (N_18981,N_18387,N_18205);
nor U18982 (N_18982,N_17674,N_18263);
nand U18983 (N_18983,N_18245,N_17905);
nor U18984 (N_18984,N_17601,N_17992);
and U18985 (N_18985,N_17743,N_17901);
or U18986 (N_18986,N_17742,N_17996);
nand U18987 (N_18987,N_17728,N_17707);
or U18988 (N_18988,N_17820,N_18227);
or U18989 (N_18989,N_17687,N_17608);
or U18990 (N_18990,N_17616,N_18253);
xnor U18991 (N_18991,N_17745,N_18298);
nor U18992 (N_18992,N_17876,N_18028);
xnor U18993 (N_18993,N_17935,N_17896);
nor U18994 (N_18994,N_18248,N_17605);
or U18995 (N_18995,N_17616,N_18032);
nor U18996 (N_18996,N_18068,N_18041);
nor U18997 (N_18997,N_17784,N_17999);
and U18998 (N_18998,N_18102,N_18193);
nand U18999 (N_18999,N_17927,N_18139);
or U19000 (N_19000,N_17910,N_18230);
or U19001 (N_19001,N_17966,N_18109);
nor U19002 (N_19002,N_17804,N_17652);
xnor U19003 (N_19003,N_18259,N_18193);
nand U19004 (N_19004,N_17710,N_17703);
nor U19005 (N_19005,N_17919,N_18241);
nand U19006 (N_19006,N_17753,N_18174);
or U19007 (N_19007,N_18251,N_17667);
and U19008 (N_19008,N_17872,N_17725);
xor U19009 (N_19009,N_18297,N_17649);
xnor U19010 (N_19010,N_17939,N_17692);
or U19011 (N_19011,N_18131,N_17807);
or U19012 (N_19012,N_17865,N_18028);
nor U19013 (N_19013,N_18082,N_17766);
nor U19014 (N_19014,N_18108,N_18055);
nand U19015 (N_19015,N_17816,N_17709);
nor U19016 (N_19016,N_18094,N_18376);
and U19017 (N_19017,N_18161,N_17925);
and U19018 (N_19018,N_17854,N_18065);
nor U19019 (N_19019,N_18268,N_17841);
or U19020 (N_19020,N_17810,N_18096);
xor U19021 (N_19021,N_17802,N_17796);
and U19022 (N_19022,N_18001,N_18200);
nor U19023 (N_19023,N_18220,N_18271);
and U19024 (N_19024,N_18007,N_18353);
or U19025 (N_19025,N_18331,N_18332);
or U19026 (N_19026,N_18220,N_17720);
nand U19027 (N_19027,N_18307,N_17876);
nor U19028 (N_19028,N_17627,N_18234);
and U19029 (N_19029,N_18228,N_18237);
and U19030 (N_19030,N_18043,N_17655);
xnor U19031 (N_19031,N_18245,N_18330);
and U19032 (N_19032,N_17662,N_17700);
nor U19033 (N_19033,N_17923,N_18349);
xnor U19034 (N_19034,N_17689,N_18022);
nand U19035 (N_19035,N_17843,N_18085);
nor U19036 (N_19036,N_18068,N_17649);
and U19037 (N_19037,N_17707,N_18334);
nand U19038 (N_19038,N_17603,N_17737);
xor U19039 (N_19039,N_17788,N_17988);
nor U19040 (N_19040,N_17812,N_17713);
xor U19041 (N_19041,N_17975,N_17924);
xor U19042 (N_19042,N_17684,N_17882);
nand U19043 (N_19043,N_17721,N_17631);
nor U19044 (N_19044,N_18202,N_17640);
or U19045 (N_19045,N_17873,N_18201);
and U19046 (N_19046,N_18109,N_18155);
xor U19047 (N_19047,N_18244,N_18323);
nand U19048 (N_19048,N_17638,N_17807);
xnor U19049 (N_19049,N_17743,N_17624);
and U19050 (N_19050,N_18270,N_18012);
nor U19051 (N_19051,N_17752,N_18223);
nor U19052 (N_19052,N_18304,N_18045);
nand U19053 (N_19053,N_18340,N_17673);
nand U19054 (N_19054,N_17966,N_17736);
or U19055 (N_19055,N_18363,N_17807);
or U19056 (N_19056,N_18288,N_18152);
nor U19057 (N_19057,N_17998,N_18031);
and U19058 (N_19058,N_17988,N_18381);
xor U19059 (N_19059,N_17860,N_17923);
nand U19060 (N_19060,N_17689,N_17634);
nor U19061 (N_19061,N_18146,N_18107);
nand U19062 (N_19062,N_17630,N_18261);
and U19063 (N_19063,N_17700,N_17901);
nand U19064 (N_19064,N_18375,N_18298);
xor U19065 (N_19065,N_18047,N_18066);
nand U19066 (N_19066,N_18336,N_17945);
nor U19067 (N_19067,N_18062,N_17850);
xnor U19068 (N_19068,N_18268,N_18367);
and U19069 (N_19069,N_18019,N_18175);
xnor U19070 (N_19070,N_18315,N_18236);
and U19071 (N_19071,N_17821,N_17729);
nor U19072 (N_19072,N_17887,N_17941);
and U19073 (N_19073,N_18277,N_18014);
nand U19074 (N_19074,N_17702,N_18151);
and U19075 (N_19075,N_18367,N_17871);
nand U19076 (N_19076,N_18345,N_17698);
nand U19077 (N_19077,N_17868,N_17733);
or U19078 (N_19078,N_17999,N_17957);
or U19079 (N_19079,N_17779,N_17919);
and U19080 (N_19080,N_17704,N_18179);
nand U19081 (N_19081,N_18098,N_17907);
xnor U19082 (N_19082,N_17744,N_18062);
xnor U19083 (N_19083,N_18078,N_18153);
nand U19084 (N_19084,N_18363,N_18108);
and U19085 (N_19085,N_17899,N_17959);
and U19086 (N_19086,N_17905,N_18032);
nor U19087 (N_19087,N_18086,N_17829);
and U19088 (N_19088,N_18096,N_18304);
or U19089 (N_19089,N_17948,N_18274);
xnor U19090 (N_19090,N_17646,N_18060);
xnor U19091 (N_19091,N_18099,N_17927);
and U19092 (N_19092,N_18115,N_17649);
xor U19093 (N_19093,N_17891,N_17711);
nor U19094 (N_19094,N_18291,N_18173);
xor U19095 (N_19095,N_18052,N_17731);
and U19096 (N_19096,N_17661,N_17695);
nand U19097 (N_19097,N_17971,N_18165);
and U19098 (N_19098,N_18207,N_18264);
or U19099 (N_19099,N_18131,N_17659);
nor U19100 (N_19100,N_17784,N_17913);
and U19101 (N_19101,N_18101,N_17818);
xor U19102 (N_19102,N_17993,N_17600);
xnor U19103 (N_19103,N_18120,N_17666);
xor U19104 (N_19104,N_18214,N_17615);
nand U19105 (N_19105,N_17969,N_17753);
or U19106 (N_19106,N_18157,N_18076);
nor U19107 (N_19107,N_17847,N_17993);
xor U19108 (N_19108,N_17699,N_18009);
nor U19109 (N_19109,N_18298,N_18110);
and U19110 (N_19110,N_18287,N_17757);
xor U19111 (N_19111,N_17982,N_18229);
nand U19112 (N_19112,N_17622,N_17913);
and U19113 (N_19113,N_18143,N_18165);
nor U19114 (N_19114,N_18372,N_18159);
or U19115 (N_19115,N_17919,N_18018);
nand U19116 (N_19116,N_18319,N_17652);
nand U19117 (N_19117,N_18323,N_18165);
nor U19118 (N_19118,N_18276,N_18341);
or U19119 (N_19119,N_18174,N_17885);
or U19120 (N_19120,N_18190,N_18373);
xor U19121 (N_19121,N_17994,N_18298);
or U19122 (N_19122,N_17637,N_18242);
xor U19123 (N_19123,N_17942,N_18138);
xor U19124 (N_19124,N_17962,N_18287);
nor U19125 (N_19125,N_18212,N_18056);
or U19126 (N_19126,N_18282,N_17737);
or U19127 (N_19127,N_17890,N_17940);
nor U19128 (N_19128,N_17632,N_18084);
nand U19129 (N_19129,N_17619,N_17839);
nor U19130 (N_19130,N_17866,N_18292);
xor U19131 (N_19131,N_18369,N_17669);
xnor U19132 (N_19132,N_17962,N_17809);
nand U19133 (N_19133,N_17665,N_18077);
nor U19134 (N_19134,N_18199,N_17962);
xnor U19135 (N_19135,N_18206,N_18245);
or U19136 (N_19136,N_18279,N_18197);
and U19137 (N_19137,N_17632,N_17810);
xnor U19138 (N_19138,N_17791,N_17922);
and U19139 (N_19139,N_18319,N_17808);
nand U19140 (N_19140,N_18062,N_18187);
or U19141 (N_19141,N_17826,N_17607);
and U19142 (N_19142,N_17677,N_18122);
nand U19143 (N_19143,N_17743,N_18064);
or U19144 (N_19144,N_17757,N_17656);
xnor U19145 (N_19145,N_18146,N_18075);
and U19146 (N_19146,N_18124,N_18396);
nand U19147 (N_19147,N_17755,N_18342);
xnor U19148 (N_19148,N_17821,N_17765);
or U19149 (N_19149,N_18139,N_18029);
nor U19150 (N_19150,N_18072,N_18390);
and U19151 (N_19151,N_18299,N_17723);
xor U19152 (N_19152,N_18281,N_17944);
xor U19153 (N_19153,N_17782,N_18165);
and U19154 (N_19154,N_17984,N_18339);
and U19155 (N_19155,N_17638,N_18377);
nor U19156 (N_19156,N_17658,N_17646);
xnor U19157 (N_19157,N_18362,N_18346);
nor U19158 (N_19158,N_18349,N_18060);
xor U19159 (N_19159,N_17974,N_17625);
nor U19160 (N_19160,N_18115,N_17718);
nor U19161 (N_19161,N_17800,N_18024);
or U19162 (N_19162,N_17832,N_17964);
xor U19163 (N_19163,N_17999,N_17858);
and U19164 (N_19164,N_17715,N_17935);
xor U19165 (N_19165,N_17954,N_18299);
xor U19166 (N_19166,N_18050,N_17813);
nor U19167 (N_19167,N_18036,N_17741);
nor U19168 (N_19168,N_18089,N_17702);
nand U19169 (N_19169,N_17914,N_17934);
nand U19170 (N_19170,N_17648,N_18366);
or U19171 (N_19171,N_17879,N_18204);
nor U19172 (N_19172,N_18125,N_17686);
nor U19173 (N_19173,N_18347,N_17918);
xnor U19174 (N_19174,N_17823,N_18262);
and U19175 (N_19175,N_17913,N_17882);
and U19176 (N_19176,N_18284,N_18075);
or U19177 (N_19177,N_17922,N_17829);
nor U19178 (N_19178,N_17839,N_18232);
and U19179 (N_19179,N_18143,N_18283);
nand U19180 (N_19180,N_17915,N_18113);
and U19181 (N_19181,N_18386,N_18006);
nand U19182 (N_19182,N_18382,N_17793);
nor U19183 (N_19183,N_17746,N_17819);
xor U19184 (N_19184,N_17882,N_18338);
nor U19185 (N_19185,N_18318,N_17930);
or U19186 (N_19186,N_18368,N_17835);
and U19187 (N_19187,N_17962,N_18349);
xnor U19188 (N_19188,N_18271,N_18317);
nand U19189 (N_19189,N_17884,N_17713);
or U19190 (N_19190,N_18366,N_18009);
and U19191 (N_19191,N_18305,N_17980);
nor U19192 (N_19192,N_17802,N_17823);
and U19193 (N_19193,N_18138,N_17835);
xnor U19194 (N_19194,N_17707,N_18388);
nor U19195 (N_19195,N_18311,N_18193);
or U19196 (N_19196,N_17873,N_17879);
nand U19197 (N_19197,N_17842,N_18335);
nor U19198 (N_19198,N_18382,N_17624);
nor U19199 (N_19199,N_18253,N_18143);
or U19200 (N_19200,N_19129,N_18876);
or U19201 (N_19201,N_19132,N_18922);
nor U19202 (N_19202,N_18677,N_18741);
and U19203 (N_19203,N_18423,N_19122);
or U19204 (N_19204,N_18436,N_19125);
nand U19205 (N_19205,N_19191,N_19195);
nor U19206 (N_19206,N_18734,N_19091);
or U19207 (N_19207,N_18755,N_18659);
nor U19208 (N_19208,N_18980,N_18526);
and U19209 (N_19209,N_18431,N_19147);
xor U19210 (N_19210,N_19134,N_18637);
or U19211 (N_19211,N_18559,N_18546);
or U19212 (N_19212,N_18548,N_18969);
xnor U19213 (N_19213,N_19040,N_18706);
xnor U19214 (N_19214,N_19184,N_18588);
nor U19215 (N_19215,N_18448,N_18433);
and U19216 (N_19216,N_19000,N_18416);
or U19217 (N_19217,N_19058,N_18949);
xnor U19218 (N_19218,N_18401,N_18855);
and U19219 (N_19219,N_18461,N_18607);
xor U19220 (N_19220,N_18952,N_18744);
nand U19221 (N_19221,N_18468,N_19112);
nor U19222 (N_19222,N_18718,N_18599);
and U19223 (N_19223,N_18560,N_18892);
or U19224 (N_19224,N_18690,N_18806);
nand U19225 (N_19225,N_19143,N_19121);
nor U19226 (N_19226,N_19066,N_18986);
xor U19227 (N_19227,N_18807,N_19187);
nand U19228 (N_19228,N_19141,N_19079);
nor U19229 (N_19229,N_19120,N_18789);
xor U19230 (N_19230,N_19092,N_19111);
nand U19231 (N_19231,N_18890,N_19131);
nor U19232 (N_19232,N_19022,N_19159);
xnor U19233 (N_19233,N_18943,N_18688);
and U19234 (N_19234,N_18711,N_18427);
nor U19235 (N_19235,N_18437,N_19196);
or U19236 (N_19236,N_19038,N_19153);
or U19237 (N_19237,N_18647,N_18603);
and U19238 (N_19238,N_18407,N_19006);
or U19239 (N_19239,N_18798,N_19019);
xnor U19240 (N_19240,N_19067,N_18780);
or U19241 (N_19241,N_18778,N_18692);
xor U19242 (N_19242,N_18749,N_18936);
or U19243 (N_19243,N_18738,N_19042);
nand U19244 (N_19244,N_18455,N_18833);
nand U19245 (N_19245,N_19062,N_19149);
or U19246 (N_19246,N_18625,N_18424);
nor U19247 (N_19247,N_18421,N_19020);
nor U19248 (N_19248,N_18730,N_19085);
xnor U19249 (N_19249,N_18618,N_18435);
xnor U19250 (N_19250,N_18914,N_18944);
nand U19251 (N_19251,N_18765,N_19048);
nand U19252 (N_19252,N_18726,N_18926);
and U19253 (N_19253,N_19059,N_18459);
nand U19254 (N_19254,N_19065,N_18545);
or U19255 (N_19255,N_18779,N_18695);
xnor U19256 (N_19256,N_18541,N_18858);
nor U19257 (N_19257,N_18739,N_18820);
nor U19258 (N_19258,N_19157,N_19004);
xor U19259 (N_19259,N_18897,N_18997);
and U19260 (N_19260,N_18796,N_18786);
and U19261 (N_19261,N_19003,N_18516);
xnor U19262 (N_19262,N_18924,N_18937);
nor U19263 (N_19263,N_18488,N_18494);
xnor U19264 (N_19264,N_18528,N_18854);
or U19265 (N_19265,N_18681,N_19130);
or U19266 (N_19266,N_18425,N_18913);
nor U19267 (N_19267,N_18624,N_18982);
nor U19268 (N_19268,N_18801,N_18841);
nand U19269 (N_19269,N_18453,N_18714);
xor U19270 (N_19270,N_19123,N_18617);
nor U19271 (N_19271,N_18863,N_19035);
and U19272 (N_19272,N_18552,N_18939);
and U19273 (N_19273,N_18990,N_18697);
xnor U19274 (N_19274,N_19156,N_18816);
and U19275 (N_19275,N_18888,N_19114);
and U19276 (N_19276,N_18877,N_18664);
nor U19277 (N_19277,N_18674,N_19009);
nor U19278 (N_19278,N_19013,N_18803);
or U19279 (N_19279,N_19174,N_19088);
xor U19280 (N_19280,N_18960,N_18585);
nor U19281 (N_19281,N_19016,N_18737);
and U19282 (N_19282,N_18752,N_18710);
xor U19283 (N_19283,N_18403,N_18645);
nor U19284 (N_19284,N_18635,N_18933);
xor U19285 (N_19285,N_18555,N_19158);
nor U19286 (N_19286,N_18483,N_18646);
xnor U19287 (N_19287,N_19098,N_18750);
and U19288 (N_19288,N_19096,N_18499);
or U19289 (N_19289,N_18747,N_18577);
and U19290 (N_19290,N_19140,N_18579);
and U19291 (N_19291,N_18497,N_18587);
or U19292 (N_19292,N_18733,N_18583);
and U19293 (N_19293,N_18686,N_18698);
xor U19294 (N_19294,N_18551,N_18853);
nand U19295 (N_19295,N_19183,N_18685);
nor U19296 (N_19296,N_18974,N_18412);
xnor U19297 (N_19297,N_19078,N_18523);
nand U19298 (N_19298,N_18650,N_18429);
and U19299 (N_19299,N_18561,N_18649);
xor U19300 (N_19300,N_18813,N_18802);
nor U19301 (N_19301,N_18929,N_19041);
or U19302 (N_19302,N_18406,N_19083);
xor U19303 (N_19303,N_18848,N_19063);
nand U19304 (N_19304,N_18763,N_18840);
nor U19305 (N_19305,N_19142,N_18604);
nor U19306 (N_19306,N_18661,N_18970);
nor U19307 (N_19307,N_18699,N_18989);
nand U19308 (N_19308,N_19181,N_18844);
xnor U19309 (N_19309,N_18812,N_18758);
xnor U19310 (N_19310,N_19115,N_19093);
or U19311 (N_19311,N_18827,N_18787);
or U19312 (N_19312,N_18931,N_19025);
nor U19313 (N_19313,N_18894,N_18794);
and U19314 (N_19314,N_19069,N_19089);
or U19315 (N_19315,N_19165,N_18482);
xnor U19316 (N_19316,N_18520,N_18769);
xnor U19317 (N_19317,N_18438,N_18622);
and U19318 (N_19318,N_18633,N_18927);
and U19319 (N_19319,N_18413,N_18768);
nand U19320 (N_19320,N_18707,N_18471);
or U19321 (N_19321,N_18977,N_18602);
xnor U19322 (N_19322,N_19194,N_18477);
or U19323 (N_19323,N_18930,N_18867);
nor U19324 (N_19324,N_18463,N_19146);
xor U19325 (N_19325,N_18484,N_18919);
nor U19326 (N_19326,N_18701,N_18613);
xnor U19327 (N_19327,N_18441,N_18689);
and U19328 (N_19328,N_18999,N_18521);
xor U19329 (N_19329,N_18605,N_19172);
and U19330 (N_19330,N_18715,N_18742);
nand U19331 (N_19331,N_18620,N_18814);
and U19332 (N_19332,N_18962,N_19007);
or U19333 (N_19333,N_18507,N_18419);
nand U19334 (N_19334,N_18479,N_18581);
xnor U19335 (N_19335,N_19014,N_18716);
xnor U19336 (N_19336,N_19077,N_18996);
and U19337 (N_19337,N_18884,N_18906);
nor U19338 (N_19338,N_18723,N_18636);
nor U19339 (N_19339,N_18793,N_18847);
nor U19340 (N_19340,N_18512,N_18683);
nor U19341 (N_19341,N_19053,N_18567);
and U19342 (N_19342,N_18800,N_19090);
or U19343 (N_19343,N_18799,N_18887);
nor U19344 (N_19344,N_18432,N_18946);
nand U19345 (N_19345,N_18729,N_18916);
xor U19346 (N_19346,N_19049,N_19164);
xor U19347 (N_19347,N_18912,N_18935);
nor U19348 (N_19348,N_19011,N_18940);
or U19349 (N_19349,N_18662,N_18880);
xnor U19350 (N_19350,N_19026,N_19010);
and U19351 (N_19351,N_18573,N_18817);
and U19352 (N_19352,N_19139,N_18684);
and U19353 (N_19353,N_19056,N_18719);
or U19354 (N_19354,N_18702,N_19137);
or U19355 (N_19355,N_18612,N_18500);
xor U19356 (N_19356,N_18776,N_19167);
and U19357 (N_19357,N_18873,N_18404);
and U19358 (N_19358,N_19099,N_18673);
and U19359 (N_19359,N_18593,N_18902);
nor U19360 (N_19360,N_18859,N_18487);
nand U19361 (N_19361,N_19168,N_18762);
and U19362 (N_19362,N_18866,N_18955);
or U19363 (N_19363,N_18964,N_18958);
xor U19364 (N_19364,N_18992,N_18703);
and U19365 (N_19365,N_18630,N_18918);
or U19366 (N_19366,N_18691,N_19145);
or U19367 (N_19367,N_19095,N_18591);
nor U19368 (N_19368,N_18449,N_18590);
nor U19369 (N_19369,N_19036,N_19073);
nor U19370 (N_19370,N_18439,N_18822);
and U19371 (N_19371,N_18910,N_18809);
nor U19372 (N_19372,N_18967,N_18558);
nor U19373 (N_19373,N_19039,N_18420);
xor U19374 (N_19374,N_18682,N_18724);
nor U19375 (N_19375,N_18988,N_18417);
xnor U19376 (N_19376,N_19150,N_18891);
xnor U19377 (N_19377,N_18889,N_19008);
nor U19378 (N_19378,N_18904,N_18643);
or U19379 (N_19379,N_18651,N_18595);
xor U19380 (N_19380,N_18712,N_19045);
nand U19381 (N_19381,N_19154,N_18469);
xor U19382 (N_19382,N_18619,N_18547);
or U19383 (N_19383,N_18510,N_18987);
xnor U19384 (N_19384,N_19185,N_18491);
and U19385 (N_19385,N_18953,N_18631);
or U19386 (N_19386,N_19199,N_19175);
or U19387 (N_19387,N_18445,N_18898);
xnor U19388 (N_19388,N_18991,N_18971);
or U19389 (N_19389,N_18524,N_19054);
nor U19390 (N_19390,N_19136,N_18456);
and U19391 (N_19391,N_19052,N_18899);
nor U19392 (N_19392,N_18648,N_18829);
nor U19393 (N_19393,N_18415,N_18443);
or U19394 (N_19394,N_18870,N_18781);
nand U19395 (N_19395,N_18422,N_18670);
or U19396 (N_19396,N_18540,N_19103);
nand U19397 (N_19397,N_18584,N_19104);
nand U19398 (N_19398,N_18920,N_18849);
nand U19399 (N_19399,N_18722,N_19117);
or U19400 (N_19400,N_18474,N_19170);
and U19401 (N_19401,N_18565,N_18735);
nand U19402 (N_19402,N_19126,N_18736);
or U19403 (N_19403,N_18728,N_19152);
nand U19404 (N_19404,N_18983,N_18917);
nor U19405 (N_19405,N_18815,N_18676);
or U19406 (N_19406,N_19138,N_18883);
or U19407 (N_19407,N_19160,N_19107);
xnor U19408 (N_19408,N_18457,N_19173);
or U19409 (N_19409,N_18489,N_18732);
xor U19410 (N_19410,N_18678,N_18608);
nand U19411 (N_19411,N_19027,N_18978);
xnor U19412 (N_19412,N_19086,N_18409);
nor U19413 (N_19413,N_18947,N_18582);
nor U19414 (N_19414,N_18490,N_18506);
nand U19415 (N_19415,N_18908,N_18578);
nor U19416 (N_19416,N_18539,N_19047);
xor U19417 (N_19417,N_18708,N_18945);
nand U19418 (N_19418,N_18868,N_18564);
xor U19419 (N_19419,N_18843,N_18550);
nor U19420 (N_19420,N_18826,N_19037);
nor U19421 (N_19421,N_18571,N_18811);
nand U19422 (N_19422,N_18570,N_18700);
nand U19423 (N_19423,N_19127,N_18616);
xor U19424 (N_19424,N_18745,N_19051);
xnor U19425 (N_19425,N_18895,N_18466);
xor U19426 (N_19426,N_18418,N_18942);
nor U19427 (N_19427,N_18666,N_18932);
and U19428 (N_19428,N_18836,N_18609);
nand U19429 (N_19429,N_18503,N_18954);
nand U19430 (N_19430,N_18549,N_19031);
nor U19431 (N_19431,N_18772,N_18472);
and U19432 (N_19432,N_18428,N_18875);
xor U19433 (N_19433,N_18632,N_18525);
xor U19434 (N_19434,N_18901,N_18852);
and U19435 (N_19435,N_18757,N_19118);
and U19436 (N_19436,N_18518,N_19068);
and U19437 (N_19437,N_19029,N_18830);
nor U19438 (N_19438,N_19023,N_18663);
and U19439 (N_19439,N_19005,N_19018);
xor U19440 (N_19440,N_18611,N_18639);
nand U19441 (N_19441,N_18675,N_18966);
nor U19442 (N_19442,N_18537,N_18821);
nand U19443 (N_19443,N_19119,N_18984);
or U19444 (N_19444,N_19148,N_18950);
xor U19445 (N_19445,N_18515,N_18601);
nand U19446 (N_19446,N_18869,N_18496);
nor U19447 (N_19447,N_19080,N_19015);
nand U19448 (N_19448,N_19071,N_19032);
nor U19449 (N_19449,N_18574,N_19179);
xor U19450 (N_19450,N_18941,N_18979);
xnor U19451 (N_19451,N_19072,N_18774);
nor U19452 (N_19452,N_18411,N_18580);
xor U19453 (N_19453,N_18782,N_18511);
nor U19454 (N_19454,N_18596,N_18717);
nand U19455 (N_19455,N_18775,N_19046);
nor U19456 (N_19456,N_18478,N_18652);
nand U19457 (N_19457,N_18544,N_18671);
or U19458 (N_19458,N_18623,N_18743);
xor U19459 (N_19459,N_18911,N_19043);
nand U19460 (N_19460,N_19024,N_18909);
and U19461 (N_19461,N_19162,N_18865);
xnor U19462 (N_19462,N_18400,N_19075);
xor U19463 (N_19463,N_18641,N_19110);
and U19464 (N_19464,N_18808,N_18956);
nor U19465 (N_19465,N_19034,N_18531);
nor U19466 (N_19466,N_18572,N_18835);
nor U19467 (N_19467,N_18556,N_19044);
and U19468 (N_19468,N_18566,N_19070);
and U19469 (N_19469,N_18740,N_18857);
and U19470 (N_19470,N_18680,N_18896);
and U19471 (N_19471,N_18864,N_18597);
xnor U19472 (N_19472,N_19012,N_19190);
or U19473 (N_19473,N_18473,N_18839);
nand U19474 (N_19474,N_18975,N_19017);
or U19475 (N_19475,N_18993,N_18961);
xor U19476 (N_19476,N_18834,N_18842);
xnor U19477 (N_19477,N_18998,N_18629);
nand U19478 (N_19478,N_18485,N_18480);
xnor U19479 (N_19479,N_18838,N_18770);
xnor U19480 (N_19480,N_18656,N_18973);
or U19481 (N_19481,N_18654,N_19188);
nand U19482 (N_19482,N_18968,N_18532);
nor U19483 (N_19483,N_18627,N_18791);
xnor U19484 (N_19484,N_19106,N_18754);
nand U19485 (N_19485,N_19176,N_18667);
nor U19486 (N_19486,N_18535,N_18938);
xnor U19487 (N_19487,N_18705,N_18783);
nor U19488 (N_19488,N_19180,N_18679);
and U19489 (N_19489,N_19057,N_19144);
nor U19490 (N_19490,N_18903,N_18492);
nor U19491 (N_19491,N_19124,N_19055);
xnor U19492 (N_19492,N_18626,N_19197);
and U19493 (N_19493,N_18907,N_18777);
or U19494 (N_19494,N_18845,N_19050);
nor U19495 (N_19495,N_19064,N_18557);
or U19496 (N_19496,N_18860,N_19100);
and U19497 (N_19497,N_18672,N_19163);
nor U19498 (N_19498,N_18576,N_18882);
and U19499 (N_19499,N_18447,N_18764);
and U19500 (N_19500,N_18562,N_18753);
and U19501 (N_19501,N_18900,N_18615);
xnor U19502 (N_19502,N_19105,N_19097);
xor U19503 (N_19503,N_18694,N_18530);
xor U19504 (N_19504,N_18759,N_19189);
or U19505 (N_19505,N_18746,N_18495);
xor U19506 (N_19506,N_19084,N_19076);
or U19507 (N_19507,N_18642,N_19192);
nor U19508 (N_19508,N_18606,N_19108);
nor U19509 (N_19509,N_18923,N_18575);
and U19510 (N_19510,N_18725,N_18767);
and U19511 (N_19511,N_18509,N_18655);
and U19512 (N_19512,N_18687,N_18948);
nand U19513 (N_19513,N_18533,N_18784);
or U19514 (N_19514,N_18959,N_18804);
xnor U19515 (N_19515,N_18788,N_18634);
nand U19516 (N_19516,N_18893,N_18886);
xnor U19517 (N_19517,N_19198,N_19128);
nand U19518 (N_19518,N_18644,N_18621);
or U19519 (N_19519,N_18825,N_18563);
or U19520 (N_19520,N_18592,N_18861);
and U19521 (N_19521,N_18467,N_18828);
and U19522 (N_19522,N_18450,N_18885);
and U19523 (N_19523,N_18536,N_18543);
and U19524 (N_19524,N_18514,N_18638);
xnor U19525 (N_19525,N_19021,N_19113);
and U19526 (N_19526,N_18810,N_18874);
xnor U19527 (N_19527,N_19001,N_18905);
xnor U19528 (N_19528,N_18410,N_18628);
and U19529 (N_19529,N_18850,N_19109);
nor U19530 (N_19530,N_18660,N_19101);
or U19531 (N_19531,N_18965,N_18505);
nand U19532 (N_19532,N_18493,N_18486);
xnor U19533 (N_19533,N_18693,N_18665);
or U19534 (N_19534,N_18542,N_18795);
nor U19535 (N_19535,N_18529,N_18957);
nor U19536 (N_19536,N_18862,N_19074);
xor U19537 (N_19537,N_18994,N_18921);
or U19538 (N_19538,N_18508,N_18451);
and U19539 (N_19539,N_18773,N_18727);
nor U19540 (N_19540,N_18879,N_18824);
and U19541 (N_19541,N_18519,N_18713);
xor U19542 (N_19542,N_18446,N_18568);
nand U19543 (N_19543,N_18668,N_18440);
nor U19544 (N_19544,N_19002,N_18709);
or U19545 (N_19545,N_18598,N_18442);
and U19546 (N_19546,N_18766,N_18653);
xnor U19547 (N_19547,N_18569,N_18831);
nor U19548 (N_19548,N_19061,N_18414);
and U19549 (N_19549,N_18513,N_18881);
and U19550 (N_19550,N_18846,N_18405);
nand U19551 (N_19551,N_18837,N_19151);
or U19552 (N_19552,N_19166,N_18925);
xor U19553 (N_19553,N_18476,N_18538);
or U19554 (N_19554,N_18498,N_18522);
and U19555 (N_19555,N_18951,N_18934);
or U19556 (N_19556,N_18851,N_18972);
xor U19557 (N_19557,N_18465,N_18452);
or U19558 (N_19558,N_18589,N_18797);
xnor U19559 (N_19559,N_18818,N_18657);
or U19560 (N_19560,N_18586,N_19102);
nand U19561 (N_19561,N_19030,N_18614);
or U19562 (N_19562,N_19182,N_19178);
or U19563 (N_19563,N_18871,N_18527);
or U19564 (N_19564,N_19161,N_18790);
or U19565 (N_19565,N_18995,N_18600);
xor U19566 (N_19566,N_18731,N_18460);
nand U19567 (N_19567,N_18430,N_18594);
and U19568 (N_19568,N_19135,N_19094);
nor U19569 (N_19569,N_18475,N_19171);
and U19570 (N_19570,N_18756,N_18760);
and U19571 (N_19571,N_18704,N_18402);
nand U19572 (N_19572,N_19087,N_18856);
xor U19573 (N_19573,N_18771,N_18470);
nand U19574 (N_19574,N_19060,N_19169);
and U19575 (N_19575,N_18434,N_18610);
xor U19576 (N_19576,N_19133,N_18792);
nand U19577 (N_19577,N_18823,N_18721);
nor U19578 (N_19578,N_18554,N_18534);
and U19579 (N_19579,N_18696,N_18669);
xor U19580 (N_19580,N_19193,N_18872);
and U19581 (N_19581,N_18761,N_18819);
nand U19582 (N_19582,N_19177,N_19033);
xor U19583 (N_19583,N_18963,N_18426);
nor U19584 (N_19584,N_18985,N_18501);
and U19585 (N_19585,N_18720,N_18462);
nor U19586 (N_19586,N_18928,N_18458);
nor U19587 (N_19587,N_18454,N_18658);
nand U19588 (N_19588,N_19155,N_18832);
and U19589 (N_19589,N_18751,N_18915);
xor U19590 (N_19590,N_18408,N_18502);
or U19591 (N_19591,N_18444,N_18481);
nand U19592 (N_19592,N_19081,N_18976);
or U19593 (N_19593,N_18878,N_18504);
nor U19594 (N_19594,N_18640,N_18517);
and U19595 (N_19595,N_18805,N_19116);
nor U19596 (N_19596,N_19082,N_18748);
and U19597 (N_19597,N_19028,N_18464);
or U19598 (N_19598,N_18553,N_18785);
or U19599 (N_19599,N_19186,N_18981);
or U19600 (N_19600,N_18632,N_18483);
or U19601 (N_19601,N_18472,N_19131);
and U19602 (N_19602,N_18471,N_18713);
and U19603 (N_19603,N_18807,N_18957);
or U19604 (N_19604,N_18993,N_18743);
xor U19605 (N_19605,N_18592,N_18920);
and U19606 (N_19606,N_18840,N_18779);
nor U19607 (N_19607,N_18895,N_18881);
or U19608 (N_19608,N_18862,N_19165);
or U19609 (N_19609,N_18403,N_18774);
nand U19610 (N_19610,N_18921,N_18782);
nor U19611 (N_19611,N_19081,N_18838);
xor U19612 (N_19612,N_19024,N_18604);
xnor U19613 (N_19613,N_19081,N_19036);
nand U19614 (N_19614,N_18616,N_18428);
xnor U19615 (N_19615,N_18513,N_18980);
xor U19616 (N_19616,N_18472,N_18565);
nand U19617 (N_19617,N_19176,N_18759);
or U19618 (N_19618,N_18479,N_18424);
nor U19619 (N_19619,N_19068,N_19154);
xnor U19620 (N_19620,N_18867,N_19173);
xnor U19621 (N_19621,N_19114,N_18901);
nor U19622 (N_19622,N_18506,N_18925);
nor U19623 (N_19623,N_18939,N_18435);
nor U19624 (N_19624,N_18707,N_18497);
xor U19625 (N_19625,N_18785,N_19093);
nor U19626 (N_19626,N_18681,N_18404);
or U19627 (N_19627,N_18761,N_18766);
nor U19628 (N_19628,N_19164,N_18927);
nor U19629 (N_19629,N_18527,N_19180);
nand U19630 (N_19630,N_18494,N_18985);
and U19631 (N_19631,N_18670,N_18769);
nand U19632 (N_19632,N_18710,N_19040);
or U19633 (N_19633,N_18442,N_19199);
and U19634 (N_19634,N_18943,N_18752);
or U19635 (N_19635,N_19102,N_18456);
xor U19636 (N_19636,N_18707,N_19164);
nand U19637 (N_19637,N_18434,N_18906);
xnor U19638 (N_19638,N_19042,N_18498);
nand U19639 (N_19639,N_18562,N_18736);
xor U19640 (N_19640,N_18519,N_18931);
xnor U19641 (N_19641,N_18428,N_18708);
nor U19642 (N_19642,N_18699,N_18649);
or U19643 (N_19643,N_18489,N_18428);
nand U19644 (N_19644,N_18965,N_19031);
nor U19645 (N_19645,N_18916,N_19012);
nand U19646 (N_19646,N_18839,N_18975);
nand U19647 (N_19647,N_19149,N_19010);
xor U19648 (N_19648,N_19153,N_18930);
xor U19649 (N_19649,N_19041,N_18558);
nand U19650 (N_19650,N_18563,N_18415);
or U19651 (N_19651,N_18402,N_19062);
and U19652 (N_19652,N_18532,N_18540);
nand U19653 (N_19653,N_18903,N_18554);
and U19654 (N_19654,N_19059,N_18860);
or U19655 (N_19655,N_19141,N_18550);
and U19656 (N_19656,N_18450,N_18675);
nor U19657 (N_19657,N_18490,N_18856);
or U19658 (N_19658,N_19002,N_18502);
nand U19659 (N_19659,N_19102,N_19063);
and U19660 (N_19660,N_18635,N_18557);
and U19661 (N_19661,N_18432,N_18437);
xor U19662 (N_19662,N_18471,N_18946);
or U19663 (N_19663,N_18500,N_18873);
nor U19664 (N_19664,N_18934,N_19088);
nand U19665 (N_19665,N_18754,N_18503);
xnor U19666 (N_19666,N_18673,N_18550);
and U19667 (N_19667,N_18613,N_18431);
nand U19668 (N_19668,N_18705,N_18965);
or U19669 (N_19669,N_18966,N_18762);
nand U19670 (N_19670,N_19122,N_19048);
nand U19671 (N_19671,N_18648,N_18931);
nor U19672 (N_19672,N_18856,N_18451);
xor U19673 (N_19673,N_19198,N_18946);
nand U19674 (N_19674,N_18507,N_18771);
and U19675 (N_19675,N_19024,N_18979);
or U19676 (N_19676,N_18986,N_18683);
nand U19677 (N_19677,N_19044,N_18988);
and U19678 (N_19678,N_19088,N_18705);
and U19679 (N_19679,N_19008,N_19183);
xor U19680 (N_19680,N_18930,N_18488);
and U19681 (N_19681,N_19099,N_18470);
and U19682 (N_19682,N_18485,N_18601);
xor U19683 (N_19683,N_18820,N_19124);
or U19684 (N_19684,N_18888,N_18497);
nor U19685 (N_19685,N_18893,N_19054);
xnor U19686 (N_19686,N_19136,N_18792);
or U19687 (N_19687,N_19044,N_18912);
or U19688 (N_19688,N_18625,N_18726);
and U19689 (N_19689,N_18452,N_18535);
or U19690 (N_19690,N_18956,N_18870);
nand U19691 (N_19691,N_19160,N_18480);
nor U19692 (N_19692,N_18556,N_18791);
and U19693 (N_19693,N_18756,N_18737);
xnor U19694 (N_19694,N_19107,N_18625);
and U19695 (N_19695,N_18557,N_18701);
and U19696 (N_19696,N_18718,N_18866);
or U19697 (N_19697,N_18628,N_18639);
xor U19698 (N_19698,N_19027,N_19059);
or U19699 (N_19699,N_18620,N_18826);
or U19700 (N_19700,N_18836,N_18892);
xor U19701 (N_19701,N_18812,N_18517);
xnor U19702 (N_19702,N_18952,N_18725);
or U19703 (N_19703,N_18690,N_19175);
nor U19704 (N_19704,N_18599,N_18443);
xor U19705 (N_19705,N_18543,N_19023);
or U19706 (N_19706,N_19060,N_18789);
nand U19707 (N_19707,N_18953,N_18978);
nand U19708 (N_19708,N_18736,N_18854);
nor U19709 (N_19709,N_18557,N_18779);
xnor U19710 (N_19710,N_18639,N_18967);
and U19711 (N_19711,N_18578,N_18646);
xnor U19712 (N_19712,N_18891,N_18566);
nand U19713 (N_19713,N_18616,N_18813);
or U19714 (N_19714,N_18687,N_18415);
nor U19715 (N_19715,N_19066,N_18461);
nand U19716 (N_19716,N_18542,N_18415);
xnor U19717 (N_19717,N_18724,N_18491);
nand U19718 (N_19718,N_19072,N_19115);
nand U19719 (N_19719,N_18560,N_18695);
nand U19720 (N_19720,N_18963,N_18563);
xor U19721 (N_19721,N_18947,N_18876);
nand U19722 (N_19722,N_18404,N_18441);
or U19723 (N_19723,N_18703,N_18450);
nor U19724 (N_19724,N_18431,N_18989);
nor U19725 (N_19725,N_18746,N_19001);
nor U19726 (N_19726,N_18565,N_19102);
and U19727 (N_19727,N_19119,N_18588);
and U19728 (N_19728,N_18926,N_18467);
xnor U19729 (N_19729,N_18473,N_19112);
nand U19730 (N_19730,N_18949,N_18871);
nand U19731 (N_19731,N_18700,N_18954);
nor U19732 (N_19732,N_18910,N_18626);
nor U19733 (N_19733,N_18605,N_18790);
nor U19734 (N_19734,N_18491,N_18461);
nor U19735 (N_19735,N_18552,N_19142);
xnor U19736 (N_19736,N_18615,N_18535);
xnor U19737 (N_19737,N_18740,N_19021);
and U19738 (N_19738,N_18420,N_19051);
or U19739 (N_19739,N_18782,N_18505);
or U19740 (N_19740,N_18968,N_18891);
or U19741 (N_19741,N_19056,N_19170);
and U19742 (N_19742,N_18804,N_19173);
nand U19743 (N_19743,N_18974,N_18574);
nor U19744 (N_19744,N_19026,N_18987);
and U19745 (N_19745,N_18690,N_18441);
nor U19746 (N_19746,N_18743,N_18862);
or U19747 (N_19747,N_19171,N_18535);
xnor U19748 (N_19748,N_18766,N_19109);
and U19749 (N_19749,N_19054,N_18556);
nand U19750 (N_19750,N_18884,N_19110);
nand U19751 (N_19751,N_18886,N_18611);
nand U19752 (N_19752,N_18629,N_18779);
xnor U19753 (N_19753,N_18535,N_19071);
nor U19754 (N_19754,N_18430,N_19177);
nand U19755 (N_19755,N_18964,N_18968);
nand U19756 (N_19756,N_18935,N_18456);
or U19757 (N_19757,N_18626,N_19088);
nor U19758 (N_19758,N_19055,N_18420);
nand U19759 (N_19759,N_19084,N_18808);
xor U19760 (N_19760,N_18856,N_18902);
nand U19761 (N_19761,N_18539,N_18705);
or U19762 (N_19762,N_18674,N_19107);
or U19763 (N_19763,N_18661,N_19188);
xor U19764 (N_19764,N_18609,N_19052);
nor U19765 (N_19765,N_18461,N_19001);
nand U19766 (N_19766,N_18568,N_18926);
nand U19767 (N_19767,N_18533,N_18788);
nand U19768 (N_19768,N_18715,N_18552);
nor U19769 (N_19769,N_19092,N_19123);
nand U19770 (N_19770,N_18948,N_19037);
xnor U19771 (N_19771,N_19090,N_19146);
nor U19772 (N_19772,N_19004,N_18894);
and U19773 (N_19773,N_18495,N_18967);
or U19774 (N_19774,N_18935,N_19052);
nand U19775 (N_19775,N_18642,N_19023);
nand U19776 (N_19776,N_18985,N_18899);
xnor U19777 (N_19777,N_18713,N_19133);
nor U19778 (N_19778,N_18759,N_18739);
or U19779 (N_19779,N_18447,N_18478);
and U19780 (N_19780,N_19026,N_19120);
nand U19781 (N_19781,N_18953,N_18845);
and U19782 (N_19782,N_19166,N_18941);
nand U19783 (N_19783,N_18653,N_19164);
nor U19784 (N_19784,N_19097,N_18986);
or U19785 (N_19785,N_18822,N_18406);
xor U19786 (N_19786,N_19110,N_18925);
nand U19787 (N_19787,N_18962,N_18487);
and U19788 (N_19788,N_18624,N_18612);
xor U19789 (N_19789,N_19073,N_18975);
nor U19790 (N_19790,N_18530,N_18735);
nor U19791 (N_19791,N_19094,N_18722);
and U19792 (N_19792,N_18535,N_19068);
nand U19793 (N_19793,N_19089,N_19098);
nor U19794 (N_19794,N_18791,N_18894);
nand U19795 (N_19795,N_18970,N_18948);
nand U19796 (N_19796,N_18756,N_19134);
or U19797 (N_19797,N_18455,N_19120);
nand U19798 (N_19798,N_18560,N_18987);
and U19799 (N_19799,N_18549,N_18630);
xnor U19800 (N_19800,N_18403,N_18914);
and U19801 (N_19801,N_18951,N_18414);
nand U19802 (N_19802,N_18583,N_18544);
and U19803 (N_19803,N_18809,N_18422);
xnor U19804 (N_19804,N_18669,N_19020);
nand U19805 (N_19805,N_19050,N_18456);
and U19806 (N_19806,N_18624,N_18765);
and U19807 (N_19807,N_18787,N_18518);
and U19808 (N_19808,N_19183,N_18570);
nor U19809 (N_19809,N_19155,N_18806);
nand U19810 (N_19810,N_19014,N_18676);
xor U19811 (N_19811,N_18735,N_18770);
nor U19812 (N_19812,N_18739,N_19127);
nor U19813 (N_19813,N_19198,N_19151);
nand U19814 (N_19814,N_19093,N_19190);
nor U19815 (N_19815,N_19132,N_19051);
nand U19816 (N_19816,N_19137,N_18924);
xnor U19817 (N_19817,N_18416,N_18467);
or U19818 (N_19818,N_18430,N_18903);
nand U19819 (N_19819,N_18623,N_18965);
or U19820 (N_19820,N_18717,N_18809);
and U19821 (N_19821,N_18991,N_19090);
and U19822 (N_19822,N_18937,N_18774);
nor U19823 (N_19823,N_19177,N_19148);
nor U19824 (N_19824,N_18883,N_18488);
or U19825 (N_19825,N_19175,N_18862);
nand U19826 (N_19826,N_18819,N_19129);
or U19827 (N_19827,N_18575,N_19142);
and U19828 (N_19828,N_18873,N_19137);
or U19829 (N_19829,N_18872,N_18582);
nand U19830 (N_19830,N_19016,N_18717);
nor U19831 (N_19831,N_18504,N_18407);
nor U19832 (N_19832,N_18762,N_19011);
or U19833 (N_19833,N_19039,N_19078);
xnor U19834 (N_19834,N_18670,N_18850);
xnor U19835 (N_19835,N_18782,N_18842);
and U19836 (N_19836,N_18992,N_18640);
nor U19837 (N_19837,N_18598,N_18731);
and U19838 (N_19838,N_18966,N_19199);
nor U19839 (N_19839,N_19093,N_19176);
nand U19840 (N_19840,N_18412,N_18629);
or U19841 (N_19841,N_18724,N_18626);
nor U19842 (N_19842,N_18497,N_18632);
or U19843 (N_19843,N_18830,N_18985);
nand U19844 (N_19844,N_18814,N_18801);
nor U19845 (N_19845,N_18859,N_18730);
nand U19846 (N_19846,N_18544,N_19116);
and U19847 (N_19847,N_18458,N_18556);
and U19848 (N_19848,N_18536,N_19023);
xnor U19849 (N_19849,N_18436,N_18632);
nor U19850 (N_19850,N_18940,N_19030);
xnor U19851 (N_19851,N_18530,N_18734);
and U19852 (N_19852,N_19178,N_18463);
or U19853 (N_19853,N_19024,N_18589);
and U19854 (N_19854,N_18641,N_18737);
xnor U19855 (N_19855,N_18845,N_18692);
nand U19856 (N_19856,N_19070,N_18486);
xnor U19857 (N_19857,N_18574,N_18891);
and U19858 (N_19858,N_18733,N_18500);
xor U19859 (N_19859,N_19025,N_18824);
xor U19860 (N_19860,N_19091,N_18907);
nand U19861 (N_19861,N_18796,N_18512);
or U19862 (N_19862,N_19041,N_18793);
nor U19863 (N_19863,N_19023,N_18924);
and U19864 (N_19864,N_19103,N_19128);
nor U19865 (N_19865,N_18526,N_18454);
nor U19866 (N_19866,N_18591,N_19183);
nor U19867 (N_19867,N_18851,N_19022);
xor U19868 (N_19868,N_18679,N_18724);
nor U19869 (N_19869,N_18789,N_18468);
nor U19870 (N_19870,N_19166,N_18608);
xnor U19871 (N_19871,N_19037,N_18941);
nand U19872 (N_19872,N_19000,N_18540);
nand U19873 (N_19873,N_18687,N_19058);
or U19874 (N_19874,N_18512,N_18632);
nand U19875 (N_19875,N_19188,N_19018);
or U19876 (N_19876,N_19181,N_19175);
nand U19877 (N_19877,N_18810,N_18663);
nand U19878 (N_19878,N_18423,N_19139);
and U19879 (N_19879,N_19153,N_18498);
and U19880 (N_19880,N_19170,N_18781);
xnor U19881 (N_19881,N_18971,N_19081);
and U19882 (N_19882,N_18683,N_18801);
or U19883 (N_19883,N_19191,N_18472);
nand U19884 (N_19884,N_18454,N_18442);
xnor U19885 (N_19885,N_19080,N_18832);
nand U19886 (N_19886,N_18953,N_18995);
and U19887 (N_19887,N_19001,N_18495);
xnor U19888 (N_19888,N_18999,N_19173);
xnor U19889 (N_19889,N_18713,N_18436);
xnor U19890 (N_19890,N_18962,N_19021);
and U19891 (N_19891,N_18730,N_18914);
nand U19892 (N_19892,N_19104,N_18411);
or U19893 (N_19893,N_18728,N_18819);
and U19894 (N_19894,N_18994,N_18512);
or U19895 (N_19895,N_18874,N_19005);
nand U19896 (N_19896,N_19100,N_18822);
nor U19897 (N_19897,N_19018,N_18578);
nor U19898 (N_19898,N_19076,N_19173);
or U19899 (N_19899,N_18928,N_18737);
nand U19900 (N_19900,N_19169,N_18584);
xnor U19901 (N_19901,N_18686,N_18975);
nand U19902 (N_19902,N_18659,N_19098);
and U19903 (N_19903,N_18401,N_18990);
xnor U19904 (N_19904,N_19016,N_18484);
nand U19905 (N_19905,N_18838,N_18414);
nor U19906 (N_19906,N_18830,N_18573);
or U19907 (N_19907,N_18644,N_18410);
and U19908 (N_19908,N_18448,N_18644);
nor U19909 (N_19909,N_19019,N_18512);
xnor U19910 (N_19910,N_18436,N_18776);
xor U19911 (N_19911,N_18453,N_19100);
or U19912 (N_19912,N_18649,N_18576);
nand U19913 (N_19913,N_18929,N_18491);
nor U19914 (N_19914,N_19025,N_18520);
nor U19915 (N_19915,N_18969,N_18630);
nor U19916 (N_19916,N_18940,N_19129);
xor U19917 (N_19917,N_18741,N_18573);
nor U19918 (N_19918,N_18857,N_18767);
and U19919 (N_19919,N_18695,N_18604);
xor U19920 (N_19920,N_18624,N_18721);
or U19921 (N_19921,N_19070,N_18997);
xnor U19922 (N_19922,N_18583,N_19023);
and U19923 (N_19923,N_18947,N_18404);
nand U19924 (N_19924,N_18772,N_18610);
or U19925 (N_19925,N_18629,N_18949);
xnor U19926 (N_19926,N_18703,N_18948);
or U19927 (N_19927,N_18676,N_18862);
xnor U19928 (N_19928,N_18629,N_19147);
or U19929 (N_19929,N_18693,N_18766);
or U19930 (N_19930,N_19118,N_19188);
xor U19931 (N_19931,N_18573,N_18439);
and U19932 (N_19932,N_18755,N_18458);
nand U19933 (N_19933,N_18587,N_18570);
nor U19934 (N_19934,N_18570,N_19099);
or U19935 (N_19935,N_18854,N_19125);
and U19936 (N_19936,N_18554,N_18843);
nand U19937 (N_19937,N_18851,N_19073);
xnor U19938 (N_19938,N_18613,N_18713);
or U19939 (N_19939,N_19107,N_18412);
nor U19940 (N_19940,N_18721,N_18596);
nand U19941 (N_19941,N_18891,N_18507);
and U19942 (N_19942,N_18740,N_18836);
xor U19943 (N_19943,N_18582,N_18850);
and U19944 (N_19944,N_18913,N_18688);
or U19945 (N_19945,N_18775,N_18673);
xnor U19946 (N_19946,N_18783,N_19043);
nor U19947 (N_19947,N_18584,N_18557);
nand U19948 (N_19948,N_19111,N_18906);
nor U19949 (N_19949,N_18918,N_18672);
nor U19950 (N_19950,N_19092,N_18421);
or U19951 (N_19951,N_19129,N_18772);
and U19952 (N_19952,N_19149,N_18965);
nor U19953 (N_19953,N_18672,N_19024);
nor U19954 (N_19954,N_18837,N_19043);
xor U19955 (N_19955,N_18748,N_18677);
and U19956 (N_19956,N_19006,N_19189);
nor U19957 (N_19957,N_18871,N_18794);
and U19958 (N_19958,N_18734,N_18867);
nand U19959 (N_19959,N_18497,N_18724);
xor U19960 (N_19960,N_18524,N_18746);
nand U19961 (N_19961,N_18549,N_18440);
and U19962 (N_19962,N_18560,N_18739);
nor U19963 (N_19963,N_19079,N_18691);
or U19964 (N_19964,N_19092,N_18400);
xor U19965 (N_19965,N_18934,N_18948);
and U19966 (N_19966,N_19060,N_19113);
and U19967 (N_19967,N_18687,N_18894);
nand U19968 (N_19968,N_19151,N_18785);
nor U19969 (N_19969,N_19158,N_18713);
nor U19970 (N_19970,N_19051,N_18841);
xnor U19971 (N_19971,N_18593,N_18691);
nand U19972 (N_19972,N_18962,N_18585);
or U19973 (N_19973,N_18603,N_18597);
nand U19974 (N_19974,N_18753,N_19044);
or U19975 (N_19975,N_18510,N_18479);
xnor U19976 (N_19976,N_18866,N_18593);
and U19977 (N_19977,N_18832,N_18638);
and U19978 (N_19978,N_18944,N_18932);
xor U19979 (N_19979,N_18602,N_19093);
xor U19980 (N_19980,N_19004,N_18663);
or U19981 (N_19981,N_18800,N_18880);
xnor U19982 (N_19982,N_18898,N_18868);
and U19983 (N_19983,N_19123,N_18706);
or U19984 (N_19984,N_18505,N_18609);
or U19985 (N_19985,N_18830,N_18507);
or U19986 (N_19986,N_18450,N_19198);
or U19987 (N_19987,N_18584,N_19140);
nor U19988 (N_19988,N_18975,N_18550);
or U19989 (N_19989,N_18883,N_18723);
nand U19990 (N_19990,N_19036,N_18984);
nand U19991 (N_19991,N_18859,N_19132);
xor U19992 (N_19992,N_18963,N_18753);
nand U19993 (N_19993,N_18442,N_19098);
and U19994 (N_19994,N_18697,N_18474);
xor U19995 (N_19995,N_18643,N_19107);
nand U19996 (N_19996,N_18599,N_18766);
and U19997 (N_19997,N_18687,N_18438);
nor U19998 (N_19998,N_18524,N_18735);
xor U19999 (N_19999,N_19037,N_19048);
and UO_0 (O_0,N_19235,N_19552);
and UO_1 (O_1,N_19938,N_19834);
and UO_2 (O_2,N_19441,N_19906);
xnor UO_3 (O_3,N_19277,N_19362);
or UO_4 (O_4,N_19639,N_19269);
or UO_5 (O_5,N_19893,N_19368);
and UO_6 (O_6,N_19206,N_19715);
or UO_7 (O_7,N_19431,N_19797);
nor UO_8 (O_8,N_19396,N_19534);
and UO_9 (O_9,N_19523,N_19201);
or UO_10 (O_10,N_19207,N_19641);
nor UO_11 (O_11,N_19788,N_19463);
nand UO_12 (O_12,N_19386,N_19587);
and UO_13 (O_13,N_19314,N_19756);
or UO_14 (O_14,N_19911,N_19495);
nor UO_15 (O_15,N_19504,N_19766);
or UO_16 (O_16,N_19230,N_19770);
and UO_17 (O_17,N_19972,N_19238);
nand UO_18 (O_18,N_19714,N_19820);
nand UO_19 (O_19,N_19814,N_19294);
nand UO_20 (O_20,N_19627,N_19633);
xor UO_21 (O_21,N_19330,N_19305);
nor UO_22 (O_22,N_19801,N_19659);
or UO_23 (O_23,N_19784,N_19620);
xnor UO_24 (O_24,N_19719,N_19537);
nor UO_25 (O_25,N_19748,N_19223);
nand UO_26 (O_26,N_19387,N_19310);
nor UO_27 (O_27,N_19607,N_19763);
nand UO_28 (O_28,N_19740,N_19264);
xor UO_29 (O_29,N_19328,N_19509);
xor UO_30 (O_30,N_19836,N_19403);
or UO_31 (O_31,N_19614,N_19650);
or UO_32 (O_32,N_19533,N_19904);
or UO_33 (O_33,N_19342,N_19329);
and UO_34 (O_34,N_19363,N_19381);
or UO_35 (O_35,N_19320,N_19578);
nor UO_36 (O_36,N_19244,N_19691);
or UO_37 (O_37,N_19525,N_19574);
nor UO_38 (O_38,N_19489,N_19675);
xnor UO_39 (O_39,N_19685,N_19648);
xor UO_40 (O_40,N_19736,N_19361);
and UO_41 (O_41,N_19324,N_19751);
or UO_42 (O_42,N_19453,N_19638);
xnor UO_43 (O_43,N_19476,N_19251);
and UO_44 (O_44,N_19432,N_19864);
xnor UO_45 (O_45,N_19390,N_19786);
nor UO_46 (O_46,N_19233,N_19592);
and UO_47 (O_47,N_19253,N_19535);
xor UO_48 (O_48,N_19848,N_19565);
nor UO_49 (O_49,N_19876,N_19618);
nor UO_50 (O_50,N_19332,N_19824);
nand UO_51 (O_51,N_19393,N_19875);
or UO_52 (O_52,N_19821,N_19566);
nor UO_53 (O_53,N_19919,N_19846);
nand UO_54 (O_54,N_19501,N_19757);
and UO_55 (O_55,N_19774,N_19389);
nor UO_56 (O_56,N_19941,N_19375);
nand UO_57 (O_57,N_19860,N_19634);
and UO_58 (O_58,N_19584,N_19494);
and UO_59 (O_59,N_19528,N_19271);
or UO_60 (O_60,N_19488,N_19512);
nor UO_61 (O_61,N_19805,N_19379);
xor UO_62 (O_62,N_19621,N_19830);
nand UO_63 (O_63,N_19210,N_19835);
and UO_64 (O_64,N_19213,N_19485);
and UO_65 (O_65,N_19540,N_19554);
nand UO_66 (O_66,N_19249,N_19200);
and UO_67 (O_67,N_19421,N_19257);
xor UO_68 (O_68,N_19203,N_19259);
and UO_69 (O_69,N_19450,N_19869);
and UO_70 (O_70,N_19349,N_19355);
nor UO_71 (O_71,N_19730,N_19908);
or UO_72 (O_72,N_19871,N_19804);
xnor UO_73 (O_73,N_19994,N_19413);
and UO_74 (O_74,N_19672,N_19872);
nand UO_75 (O_75,N_19483,N_19591);
or UO_76 (O_76,N_19988,N_19536);
xor UO_77 (O_77,N_19430,N_19302);
nand UO_78 (O_78,N_19482,N_19929);
or UO_79 (O_79,N_19724,N_19926);
xnor UO_80 (O_80,N_19378,N_19990);
nor UO_81 (O_81,N_19408,N_19885);
nor UO_82 (O_82,N_19985,N_19812);
or UO_83 (O_83,N_19412,N_19576);
nand UO_84 (O_84,N_19466,N_19597);
or UO_85 (O_85,N_19799,N_19286);
or UO_86 (O_86,N_19942,N_19753);
nor UO_87 (O_87,N_19905,N_19644);
xnor UO_88 (O_88,N_19380,N_19215);
or UO_89 (O_89,N_19603,N_19816);
nand UO_90 (O_90,N_19468,N_19833);
xor UO_91 (O_91,N_19296,N_19726);
and UO_92 (O_92,N_19910,N_19609);
and UO_93 (O_93,N_19831,N_19819);
nand UO_94 (O_94,N_19404,N_19371);
xnor UO_95 (O_95,N_19859,N_19426);
nor UO_96 (O_96,N_19987,N_19266);
nor UO_97 (O_97,N_19419,N_19612);
nand UO_98 (O_98,N_19702,N_19682);
or UO_99 (O_99,N_19745,N_19725);
and UO_100 (O_100,N_19948,N_19851);
nand UO_101 (O_101,N_19677,N_19518);
or UO_102 (O_102,N_19917,N_19918);
or UO_103 (O_103,N_19569,N_19777);
nor UO_104 (O_104,N_19307,N_19940);
or UO_105 (O_105,N_19850,N_19514);
and UO_106 (O_106,N_19478,N_19510);
nand UO_107 (O_107,N_19789,N_19274);
and UO_108 (O_108,N_19645,N_19843);
nor UO_109 (O_109,N_19626,N_19240);
nand UO_110 (O_110,N_19369,N_19418);
or UO_111 (O_111,N_19707,N_19858);
nand UO_112 (O_112,N_19300,N_19878);
nor UO_113 (O_113,N_19366,N_19664);
nand UO_114 (O_114,N_19586,N_19998);
nor UO_115 (O_115,N_19326,N_19881);
and UO_116 (O_116,N_19924,N_19734);
or UO_117 (O_117,N_19506,N_19604);
nor UO_118 (O_118,N_19713,N_19334);
and UO_119 (O_119,N_19907,N_19969);
nor UO_120 (O_120,N_19519,N_19204);
nand UO_121 (O_121,N_19628,N_19452);
and UO_122 (O_122,N_19260,N_19467);
xor UO_123 (O_123,N_19863,N_19890);
nor UO_124 (O_124,N_19856,N_19601);
nand UO_125 (O_125,N_19352,N_19477);
and UO_126 (O_126,N_19790,N_19595);
xnor UO_127 (O_127,N_19365,N_19686);
and UO_128 (O_128,N_19646,N_19538);
nand UO_129 (O_129,N_19376,N_19667);
nand UO_130 (O_130,N_19401,N_19992);
nor UO_131 (O_131,N_19471,N_19610);
xor UO_132 (O_132,N_19405,N_19921);
or UO_133 (O_133,N_19779,N_19861);
or UO_134 (O_134,N_19977,N_19311);
xor UO_135 (O_135,N_19409,N_19706);
xnor UO_136 (O_136,N_19265,N_19782);
nand UO_137 (O_137,N_19953,N_19205);
or UO_138 (O_138,N_19439,N_19986);
or UO_139 (O_139,N_19796,N_19773);
nand UO_140 (O_140,N_19950,N_19267);
xnor UO_141 (O_141,N_19752,N_19636);
nor UO_142 (O_142,N_19559,N_19807);
and UO_143 (O_143,N_19958,N_19415);
nand UO_144 (O_144,N_19712,N_19316);
nor UO_145 (O_145,N_19543,N_19547);
and UO_146 (O_146,N_19364,N_19532);
or UO_147 (O_147,N_19580,N_19935);
nor UO_148 (O_148,N_19282,N_19974);
nand UO_149 (O_149,N_19486,N_19884);
xnor UO_150 (O_150,N_19284,N_19357);
and UO_151 (O_151,N_19336,N_19960);
or UO_152 (O_152,N_19312,N_19507);
nand UO_153 (O_153,N_19397,N_19697);
nand UO_154 (O_154,N_19270,N_19778);
xnor UO_155 (O_155,N_19737,N_19594);
nor UO_156 (O_156,N_19423,N_19652);
nand UO_157 (O_157,N_19429,N_19384);
xor UO_158 (O_158,N_19695,N_19800);
or UO_159 (O_159,N_19344,N_19560);
nor UO_160 (O_160,N_19787,N_19882);
nor UO_161 (O_161,N_19643,N_19377);
xor UO_162 (O_162,N_19658,N_19629);
and UO_163 (O_163,N_19605,N_19406);
nand UO_164 (O_164,N_19451,N_19826);
and UO_165 (O_165,N_19898,N_19696);
or UO_166 (O_166,N_19530,N_19593);
and UO_167 (O_167,N_19802,N_19226);
or UO_168 (O_168,N_19337,N_19339);
or UO_169 (O_169,N_19457,N_19966);
or UO_170 (O_170,N_19600,N_19493);
and UO_171 (O_171,N_19978,N_19862);
nor UO_172 (O_172,N_19229,N_19571);
xnor UO_173 (O_173,N_19623,N_19870);
nor UO_174 (O_174,N_19964,N_19407);
nand UO_175 (O_175,N_19443,N_19520);
nor UO_176 (O_176,N_19656,N_19338);
nand UO_177 (O_177,N_19283,N_19976);
nor UO_178 (O_178,N_19359,N_19563);
or UO_179 (O_179,N_19783,N_19810);
and UO_180 (O_180,N_19733,N_19959);
nor UO_181 (O_181,N_19449,N_19982);
nor UO_182 (O_182,N_19722,N_19718);
nor UO_183 (O_183,N_19936,N_19433);
nand UO_184 (O_184,N_19553,N_19392);
nand UO_185 (O_185,N_19222,N_19301);
and UO_186 (O_186,N_19825,N_19232);
xnor UO_187 (O_187,N_19589,N_19276);
nor UO_188 (O_188,N_19687,N_19723);
or UO_189 (O_189,N_19481,N_19690);
xnor UO_190 (O_190,N_19469,N_19317);
xor UO_191 (O_191,N_19420,N_19475);
or UO_192 (O_192,N_19289,N_19221);
and UO_193 (O_193,N_19951,N_19318);
nor UO_194 (O_194,N_19746,N_19549);
or UO_195 (O_195,N_19588,N_19946);
and UO_196 (O_196,N_19996,N_19769);
and UO_197 (O_197,N_19841,N_19877);
and UO_198 (O_198,N_19304,N_19775);
nor UO_199 (O_199,N_19278,N_19382);
and UO_200 (O_200,N_19293,N_19434);
or UO_201 (O_201,N_19268,N_19704);
or UO_202 (O_202,N_19590,N_19887);
nand UO_203 (O_203,N_19930,N_19701);
xnor UO_204 (O_204,N_19981,N_19899);
and UO_205 (O_205,N_19873,N_19236);
nor UO_206 (O_206,N_19517,N_19688);
and UO_207 (O_207,N_19681,N_19557);
or UO_208 (O_208,N_19308,N_19219);
nand UO_209 (O_209,N_19732,N_19447);
xor UO_210 (O_210,N_19208,N_19497);
xnor UO_211 (O_211,N_19367,N_19546);
or UO_212 (O_212,N_19731,N_19684);
nand UO_213 (O_213,N_19303,N_19915);
xnor UO_214 (O_214,N_19671,N_19480);
xor UO_215 (O_215,N_19699,N_19741);
nor UO_216 (O_216,N_19735,N_19247);
and UO_217 (O_217,N_19853,N_19822);
nor UO_218 (O_218,N_19649,N_19490);
or UO_219 (O_219,N_19511,N_19700);
xnor UO_220 (O_220,N_19327,N_19279);
nand UO_221 (O_221,N_19716,N_19927);
nand UO_222 (O_222,N_19273,N_19388);
or UO_223 (O_223,N_19928,N_19635);
nand UO_224 (O_224,N_19579,N_19963);
nand UO_225 (O_225,N_19351,N_19250);
or UO_226 (O_226,N_19891,N_19849);
xnor UO_227 (O_227,N_19562,N_19867);
xnor UO_228 (O_228,N_19298,N_19564);
nand UO_229 (O_229,N_19903,N_19313);
nand UO_230 (O_230,N_19823,N_19622);
nand UO_231 (O_231,N_19542,N_19916);
nand UO_232 (O_232,N_19479,N_19886);
xor UO_233 (O_233,N_19484,N_19721);
nand UO_234 (O_234,N_19360,N_19943);
nand UO_235 (O_235,N_19632,N_19792);
xnor UO_236 (O_236,N_19427,N_19973);
and UO_237 (O_237,N_19492,N_19508);
nand UO_238 (O_238,N_19909,N_19570);
nor UO_239 (O_239,N_19582,N_19502);
and UO_240 (O_240,N_19496,N_19306);
nand UO_241 (O_241,N_19720,N_19583);
and UO_242 (O_242,N_19556,N_19487);
nand UO_243 (O_243,N_19262,N_19474);
nand UO_244 (O_244,N_19808,N_19442);
nand UO_245 (O_245,N_19422,N_19742);
or UO_246 (O_246,N_19347,N_19228);
and UO_247 (O_247,N_19400,N_19705);
nand UO_248 (O_248,N_19241,N_19331);
nor UO_249 (O_249,N_19984,N_19446);
or UO_250 (O_250,N_19894,N_19956);
xnor UO_251 (O_251,N_19711,N_19224);
nor UO_252 (O_252,N_19551,N_19548);
nand UO_253 (O_253,N_19568,N_19345);
xor UO_254 (O_254,N_19854,N_19617);
and UO_255 (O_255,N_19252,N_19209);
nand UO_256 (O_256,N_19738,N_19842);
and UO_257 (O_257,N_19970,N_19989);
or UO_258 (O_258,N_19353,N_19465);
or UO_259 (O_259,N_19416,N_19585);
xnor UO_260 (O_260,N_19436,N_19424);
and UO_261 (O_261,N_19611,N_19350);
nand UO_262 (O_262,N_19613,N_19945);
xor UO_263 (O_263,N_19817,N_19322);
or UO_264 (O_264,N_19955,N_19897);
nor UO_265 (O_265,N_19630,N_19944);
nand UO_266 (O_266,N_19855,N_19417);
or UO_267 (O_267,N_19428,N_19913);
nand UO_268 (O_268,N_19500,N_19678);
nor UO_269 (O_269,N_19280,N_19999);
or UO_270 (O_270,N_19608,N_19888);
nand UO_271 (O_271,N_19503,N_19470);
nor UO_272 (O_272,N_19498,N_19975);
and UO_273 (O_273,N_19794,N_19454);
nor UO_274 (O_274,N_19245,N_19642);
and UO_275 (O_275,N_19524,N_19679);
and UO_276 (O_276,N_19758,N_19811);
nand UO_277 (O_277,N_19771,N_19637);
xnor UO_278 (O_278,N_19640,N_19827);
and UO_279 (O_279,N_19768,N_19934);
xor UO_280 (O_280,N_19414,N_19728);
or UO_281 (O_281,N_19920,N_19865);
nor UO_282 (O_282,N_19914,N_19983);
nor UO_283 (O_283,N_19340,N_19654);
nor UO_284 (O_284,N_19438,N_19596);
nand UO_285 (O_285,N_19767,N_19896);
nand UO_286 (O_286,N_19791,N_19473);
nor UO_287 (O_287,N_19291,N_19965);
nand UO_288 (O_288,N_19727,N_19764);
nand UO_289 (O_289,N_19292,N_19673);
nor UO_290 (O_290,N_19995,N_19309);
or UO_291 (O_291,N_19933,N_19461);
and UO_292 (O_292,N_19818,N_19743);
nand UO_293 (O_293,N_19239,N_19615);
xnor UO_294 (O_294,N_19348,N_19866);
xor UO_295 (O_295,N_19806,N_19263);
nand UO_296 (O_296,N_19828,N_19683);
xnor UO_297 (O_297,N_19954,N_19997);
nand UO_298 (O_298,N_19925,N_19670);
and UO_299 (O_299,N_19323,N_19445);
nand UO_300 (O_300,N_19795,N_19581);
nor UO_301 (O_301,N_19435,N_19880);
and UO_302 (O_302,N_19356,N_19459);
and UO_303 (O_303,N_19341,N_19710);
nand UO_304 (O_304,N_19957,N_19460);
nand UO_305 (O_305,N_19837,N_19346);
nor UO_306 (O_306,N_19967,N_19372);
nand UO_307 (O_307,N_19922,N_19759);
xor UO_308 (O_308,N_19962,N_19980);
nor UO_309 (O_309,N_19545,N_19491);
or UO_310 (O_310,N_19321,N_19660);
nand UO_311 (O_311,N_19567,N_19709);
xnor UO_312 (O_312,N_19662,N_19674);
xor UO_313 (O_313,N_19651,N_19602);
and UO_314 (O_314,N_19772,N_19892);
nor UO_315 (O_315,N_19550,N_19395);
xnor UO_316 (O_316,N_19272,N_19932);
nand UO_317 (O_317,N_19577,N_19217);
nor UO_318 (O_318,N_19693,N_19762);
or UO_319 (O_319,N_19761,N_19968);
nand UO_320 (O_320,N_19513,N_19522);
xnor UO_321 (O_321,N_19847,N_19776);
nand UO_322 (O_322,N_19516,N_19555);
and UO_323 (O_323,N_19874,N_19243);
nor UO_324 (O_324,N_19680,N_19444);
or UO_325 (O_325,N_19971,N_19385);
xnor UO_326 (O_326,N_19297,N_19668);
nor UO_327 (O_327,N_19793,N_19211);
xor UO_328 (O_328,N_19370,N_19531);
nor UO_329 (O_329,N_19780,N_19225);
xnor UO_330 (O_330,N_19979,N_19689);
nand UO_331 (O_331,N_19676,N_19573);
and UO_332 (O_332,N_19242,N_19358);
and UO_333 (O_333,N_19394,N_19845);
xor UO_334 (O_334,N_19572,N_19868);
and UO_335 (O_335,N_19655,N_19717);
nand UO_336 (O_336,N_19299,N_19325);
xor UO_337 (O_337,N_19398,N_19526);
xnor UO_338 (O_338,N_19472,N_19993);
and UO_339 (O_339,N_19829,N_19539);
or UO_340 (O_340,N_19781,N_19335);
and UO_341 (O_341,N_19391,N_19288);
nor UO_342 (O_342,N_19561,N_19931);
xnor UO_343 (O_343,N_19505,N_19923);
nand UO_344 (O_344,N_19216,N_19529);
or UO_345 (O_345,N_19521,N_19703);
nand UO_346 (O_346,N_19661,N_19544);
nand UO_347 (O_347,N_19744,N_19458);
nor UO_348 (O_348,N_19729,N_19665);
and UO_349 (O_349,N_19437,N_19631);
or UO_350 (O_350,N_19902,N_19883);
or UO_351 (O_351,N_19220,N_19527);
nor UO_352 (O_352,N_19575,N_19947);
xnor UO_353 (O_353,N_19541,N_19889);
and UO_354 (O_354,N_19839,N_19952);
xnor UO_355 (O_355,N_19694,N_19937);
or UO_356 (O_356,N_19234,N_19750);
nor UO_357 (O_357,N_19254,N_19319);
and UO_358 (O_358,N_19809,N_19647);
xor UO_359 (O_359,N_19901,N_19803);
or UO_360 (O_360,N_19598,N_19462);
nand UO_361 (O_361,N_19895,N_19383);
and UO_362 (O_362,N_19708,N_19838);
and UO_363 (O_363,N_19456,N_19411);
xnor UO_364 (O_364,N_19798,N_19464);
nor UO_365 (O_365,N_19852,N_19515);
nand UO_366 (O_366,N_19256,N_19949);
or UO_367 (O_367,N_19832,N_19354);
and UO_368 (O_368,N_19248,N_19815);
or UO_369 (O_369,N_19912,N_19373);
nor UO_370 (O_370,N_19991,N_19961);
xnor UO_371 (O_371,N_19275,N_19448);
nor UO_372 (O_372,N_19425,N_19290);
nor UO_373 (O_373,N_19227,N_19624);
xor UO_374 (O_374,N_19315,N_19754);
and UO_375 (O_375,N_19698,N_19900);
and UO_376 (O_376,N_19558,N_19857);
nor UO_377 (O_377,N_19499,N_19844);
or UO_378 (O_378,N_19606,N_19755);
or UO_379 (O_379,N_19625,N_19255);
or UO_380 (O_380,N_19237,N_19765);
nand UO_381 (O_381,N_19785,N_19258);
xnor UO_382 (O_382,N_19939,N_19261);
and UO_383 (O_383,N_19739,N_19214);
nor UO_384 (O_384,N_19879,N_19231);
xor UO_385 (O_385,N_19747,N_19287);
or UO_386 (O_386,N_19281,N_19599);
xor UO_387 (O_387,N_19285,N_19669);
and UO_388 (O_388,N_19616,N_19749);
nor UO_389 (O_389,N_19212,N_19399);
xor UO_390 (O_390,N_19333,N_19666);
or UO_391 (O_391,N_19840,N_19218);
or UO_392 (O_392,N_19440,N_19410);
xnor UO_393 (O_393,N_19619,N_19663);
nor UO_394 (O_394,N_19295,N_19657);
nand UO_395 (O_395,N_19653,N_19246);
xnor UO_396 (O_396,N_19343,N_19692);
nor UO_397 (O_397,N_19402,N_19455);
xnor UO_398 (O_398,N_19813,N_19374);
xnor UO_399 (O_399,N_19760,N_19202);
or UO_400 (O_400,N_19316,N_19756);
or UO_401 (O_401,N_19985,N_19933);
and UO_402 (O_402,N_19788,N_19326);
xnor UO_403 (O_403,N_19807,N_19992);
nor UO_404 (O_404,N_19296,N_19299);
nand UO_405 (O_405,N_19532,N_19294);
and UO_406 (O_406,N_19862,N_19607);
nor UO_407 (O_407,N_19380,N_19598);
nand UO_408 (O_408,N_19973,N_19864);
nand UO_409 (O_409,N_19461,N_19347);
nand UO_410 (O_410,N_19689,N_19429);
nor UO_411 (O_411,N_19380,N_19935);
and UO_412 (O_412,N_19729,N_19580);
nor UO_413 (O_413,N_19875,N_19441);
nand UO_414 (O_414,N_19493,N_19526);
nor UO_415 (O_415,N_19227,N_19270);
xnor UO_416 (O_416,N_19961,N_19974);
xnor UO_417 (O_417,N_19863,N_19962);
xnor UO_418 (O_418,N_19421,N_19546);
xnor UO_419 (O_419,N_19753,N_19968);
or UO_420 (O_420,N_19952,N_19932);
or UO_421 (O_421,N_19796,N_19853);
nand UO_422 (O_422,N_19958,N_19344);
nand UO_423 (O_423,N_19398,N_19542);
nor UO_424 (O_424,N_19299,N_19268);
nand UO_425 (O_425,N_19922,N_19561);
nor UO_426 (O_426,N_19760,N_19270);
and UO_427 (O_427,N_19373,N_19926);
nand UO_428 (O_428,N_19522,N_19630);
nand UO_429 (O_429,N_19689,N_19499);
or UO_430 (O_430,N_19380,N_19834);
or UO_431 (O_431,N_19456,N_19395);
and UO_432 (O_432,N_19752,N_19477);
nand UO_433 (O_433,N_19978,N_19959);
and UO_434 (O_434,N_19436,N_19842);
and UO_435 (O_435,N_19698,N_19530);
and UO_436 (O_436,N_19544,N_19464);
or UO_437 (O_437,N_19997,N_19558);
and UO_438 (O_438,N_19668,N_19866);
or UO_439 (O_439,N_19572,N_19601);
nor UO_440 (O_440,N_19438,N_19541);
or UO_441 (O_441,N_19927,N_19595);
or UO_442 (O_442,N_19794,N_19484);
xor UO_443 (O_443,N_19696,N_19777);
xor UO_444 (O_444,N_19292,N_19404);
nand UO_445 (O_445,N_19583,N_19496);
xnor UO_446 (O_446,N_19780,N_19272);
nand UO_447 (O_447,N_19699,N_19915);
xnor UO_448 (O_448,N_19689,N_19326);
nor UO_449 (O_449,N_19687,N_19276);
and UO_450 (O_450,N_19504,N_19873);
and UO_451 (O_451,N_19476,N_19346);
and UO_452 (O_452,N_19620,N_19901);
nor UO_453 (O_453,N_19876,N_19573);
nor UO_454 (O_454,N_19827,N_19680);
or UO_455 (O_455,N_19819,N_19528);
nand UO_456 (O_456,N_19506,N_19998);
xnor UO_457 (O_457,N_19442,N_19451);
nor UO_458 (O_458,N_19671,N_19553);
nor UO_459 (O_459,N_19357,N_19453);
and UO_460 (O_460,N_19238,N_19588);
or UO_461 (O_461,N_19621,N_19694);
nor UO_462 (O_462,N_19536,N_19457);
xnor UO_463 (O_463,N_19977,N_19751);
and UO_464 (O_464,N_19302,N_19907);
or UO_465 (O_465,N_19341,N_19650);
xnor UO_466 (O_466,N_19303,N_19654);
or UO_467 (O_467,N_19429,N_19839);
or UO_468 (O_468,N_19473,N_19461);
nor UO_469 (O_469,N_19404,N_19735);
nand UO_470 (O_470,N_19863,N_19301);
nor UO_471 (O_471,N_19281,N_19863);
and UO_472 (O_472,N_19904,N_19843);
and UO_473 (O_473,N_19692,N_19334);
nor UO_474 (O_474,N_19648,N_19926);
nor UO_475 (O_475,N_19881,N_19407);
nand UO_476 (O_476,N_19202,N_19559);
nor UO_477 (O_477,N_19281,N_19234);
and UO_478 (O_478,N_19278,N_19616);
nand UO_479 (O_479,N_19634,N_19798);
and UO_480 (O_480,N_19736,N_19639);
nand UO_481 (O_481,N_19716,N_19206);
or UO_482 (O_482,N_19679,N_19256);
nand UO_483 (O_483,N_19720,N_19765);
and UO_484 (O_484,N_19615,N_19202);
or UO_485 (O_485,N_19574,N_19876);
and UO_486 (O_486,N_19888,N_19953);
nor UO_487 (O_487,N_19928,N_19531);
nand UO_488 (O_488,N_19281,N_19237);
nand UO_489 (O_489,N_19205,N_19689);
and UO_490 (O_490,N_19698,N_19972);
and UO_491 (O_491,N_19888,N_19973);
xnor UO_492 (O_492,N_19557,N_19272);
nand UO_493 (O_493,N_19721,N_19863);
and UO_494 (O_494,N_19740,N_19286);
nand UO_495 (O_495,N_19441,N_19760);
and UO_496 (O_496,N_19716,N_19999);
or UO_497 (O_497,N_19978,N_19951);
and UO_498 (O_498,N_19417,N_19510);
and UO_499 (O_499,N_19355,N_19779);
nand UO_500 (O_500,N_19712,N_19721);
and UO_501 (O_501,N_19267,N_19922);
xnor UO_502 (O_502,N_19782,N_19387);
xor UO_503 (O_503,N_19432,N_19938);
nor UO_504 (O_504,N_19965,N_19520);
xnor UO_505 (O_505,N_19679,N_19699);
and UO_506 (O_506,N_19280,N_19927);
nand UO_507 (O_507,N_19876,N_19901);
and UO_508 (O_508,N_19662,N_19403);
or UO_509 (O_509,N_19604,N_19536);
nor UO_510 (O_510,N_19368,N_19581);
nand UO_511 (O_511,N_19403,N_19331);
xnor UO_512 (O_512,N_19718,N_19853);
nor UO_513 (O_513,N_19422,N_19230);
and UO_514 (O_514,N_19717,N_19492);
and UO_515 (O_515,N_19302,N_19961);
nor UO_516 (O_516,N_19554,N_19813);
and UO_517 (O_517,N_19467,N_19428);
nand UO_518 (O_518,N_19310,N_19639);
nand UO_519 (O_519,N_19278,N_19977);
nor UO_520 (O_520,N_19477,N_19859);
or UO_521 (O_521,N_19637,N_19423);
or UO_522 (O_522,N_19378,N_19517);
nand UO_523 (O_523,N_19894,N_19760);
xor UO_524 (O_524,N_19378,N_19391);
nand UO_525 (O_525,N_19611,N_19898);
nand UO_526 (O_526,N_19766,N_19608);
and UO_527 (O_527,N_19208,N_19939);
nor UO_528 (O_528,N_19572,N_19660);
or UO_529 (O_529,N_19853,N_19481);
nand UO_530 (O_530,N_19882,N_19600);
xnor UO_531 (O_531,N_19379,N_19779);
and UO_532 (O_532,N_19328,N_19272);
nor UO_533 (O_533,N_19539,N_19802);
nor UO_534 (O_534,N_19758,N_19402);
nand UO_535 (O_535,N_19675,N_19635);
or UO_536 (O_536,N_19985,N_19336);
xnor UO_537 (O_537,N_19993,N_19315);
nor UO_538 (O_538,N_19849,N_19922);
nand UO_539 (O_539,N_19518,N_19220);
and UO_540 (O_540,N_19587,N_19846);
and UO_541 (O_541,N_19736,N_19892);
xor UO_542 (O_542,N_19604,N_19299);
or UO_543 (O_543,N_19941,N_19659);
nand UO_544 (O_544,N_19625,N_19983);
xor UO_545 (O_545,N_19635,N_19956);
or UO_546 (O_546,N_19308,N_19731);
xnor UO_547 (O_547,N_19699,N_19301);
nor UO_548 (O_548,N_19958,N_19680);
nand UO_549 (O_549,N_19228,N_19346);
nand UO_550 (O_550,N_19215,N_19315);
and UO_551 (O_551,N_19408,N_19840);
xor UO_552 (O_552,N_19297,N_19712);
or UO_553 (O_553,N_19924,N_19327);
xor UO_554 (O_554,N_19222,N_19980);
nand UO_555 (O_555,N_19817,N_19765);
or UO_556 (O_556,N_19813,N_19819);
nand UO_557 (O_557,N_19378,N_19379);
nand UO_558 (O_558,N_19606,N_19795);
xnor UO_559 (O_559,N_19530,N_19426);
or UO_560 (O_560,N_19799,N_19228);
xnor UO_561 (O_561,N_19557,N_19487);
nand UO_562 (O_562,N_19227,N_19833);
or UO_563 (O_563,N_19969,N_19927);
xnor UO_564 (O_564,N_19810,N_19605);
and UO_565 (O_565,N_19726,N_19232);
or UO_566 (O_566,N_19263,N_19484);
and UO_567 (O_567,N_19327,N_19546);
nor UO_568 (O_568,N_19491,N_19554);
and UO_569 (O_569,N_19866,N_19443);
xor UO_570 (O_570,N_19285,N_19566);
nor UO_571 (O_571,N_19699,N_19396);
or UO_572 (O_572,N_19211,N_19573);
nand UO_573 (O_573,N_19690,N_19634);
nor UO_574 (O_574,N_19724,N_19656);
nand UO_575 (O_575,N_19242,N_19464);
nor UO_576 (O_576,N_19616,N_19912);
nand UO_577 (O_577,N_19547,N_19258);
nand UO_578 (O_578,N_19596,N_19495);
nor UO_579 (O_579,N_19732,N_19224);
xor UO_580 (O_580,N_19494,N_19539);
or UO_581 (O_581,N_19919,N_19397);
or UO_582 (O_582,N_19470,N_19448);
or UO_583 (O_583,N_19702,N_19237);
or UO_584 (O_584,N_19726,N_19719);
xnor UO_585 (O_585,N_19730,N_19525);
nor UO_586 (O_586,N_19437,N_19275);
or UO_587 (O_587,N_19988,N_19455);
nand UO_588 (O_588,N_19372,N_19259);
nand UO_589 (O_589,N_19915,N_19550);
xor UO_590 (O_590,N_19768,N_19394);
and UO_591 (O_591,N_19361,N_19689);
xnor UO_592 (O_592,N_19948,N_19937);
nand UO_593 (O_593,N_19444,N_19257);
nand UO_594 (O_594,N_19539,N_19524);
or UO_595 (O_595,N_19838,N_19874);
or UO_596 (O_596,N_19633,N_19873);
nand UO_597 (O_597,N_19465,N_19593);
or UO_598 (O_598,N_19871,N_19980);
xor UO_599 (O_599,N_19555,N_19275);
or UO_600 (O_600,N_19693,N_19899);
xnor UO_601 (O_601,N_19972,N_19591);
or UO_602 (O_602,N_19575,N_19267);
nand UO_603 (O_603,N_19812,N_19286);
nand UO_604 (O_604,N_19727,N_19302);
and UO_605 (O_605,N_19220,N_19422);
xor UO_606 (O_606,N_19958,N_19261);
and UO_607 (O_607,N_19605,N_19294);
and UO_608 (O_608,N_19433,N_19259);
nor UO_609 (O_609,N_19205,N_19344);
xor UO_610 (O_610,N_19244,N_19649);
or UO_611 (O_611,N_19237,N_19256);
and UO_612 (O_612,N_19852,N_19356);
and UO_613 (O_613,N_19428,N_19545);
and UO_614 (O_614,N_19511,N_19631);
xnor UO_615 (O_615,N_19308,N_19978);
xor UO_616 (O_616,N_19864,N_19488);
xnor UO_617 (O_617,N_19449,N_19902);
nor UO_618 (O_618,N_19220,N_19302);
nand UO_619 (O_619,N_19961,N_19864);
nor UO_620 (O_620,N_19947,N_19527);
xor UO_621 (O_621,N_19955,N_19484);
xor UO_622 (O_622,N_19378,N_19535);
and UO_623 (O_623,N_19777,N_19500);
nand UO_624 (O_624,N_19271,N_19455);
xor UO_625 (O_625,N_19997,N_19596);
or UO_626 (O_626,N_19562,N_19632);
nand UO_627 (O_627,N_19520,N_19675);
xnor UO_628 (O_628,N_19877,N_19749);
and UO_629 (O_629,N_19307,N_19571);
or UO_630 (O_630,N_19705,N_19264);
nor UO_631 (O_631,N_19447,N_19854);
and UO_632 (O_632,N_19452,N_19757);
nor UO_633 (O_633,N_19716,N_19478);
nand UO_634 (O_634,N_19626,N_19327);
xnor UO_635 (O_635,N_19867,N_19555);
nand UO_636 (O_636,N_19270,N_19789);
or UO_637 (O_637,N_19755,N_19824);
nand UO_638 (O_638,N_19936,N_19638);
nor UO_639 (O_639,N_19771,N_19826);
and UO_640 (O_640,N_19476,N_19954);
xnor UO_641 (O_641,N_19312,N_19332);
xor UO_642 (O_642,N_19905,N_19529);
nor UO_643 (O_643,N_19249,N_19240);
or UO_644 (O_644,N_19882,N_19611);
or UO_645 (O_645,N_19347,N_19979);
and UO_646 (O_646,N_19689,N_19768);
nand UO_647 (O_647,N_19472,N_19632);
xnor UO_648 (O_648,N_19297,N_19996);
nand UO_649 (O_649,N_19250,N_19563);
or UO_650 (O_650,N_19724,N_19481);
nand UO_651 (O_651,N_19554,N_19228);
nor UO_652 (O_652,N_19538,N_19512);
nor UO_653 (O_653,N_19274,N_19803);
nand UO_654 (O_654,N_19807,N_19880);
or UO_655 (O_655,N_19589,N_19957);
nor UO_656 (O_656,N_19507,N_19672);
xnor UO_657 (O_657,N_19349,N_19409);
xor UO_658 (O_658,N_19950,N_19838);
nor UO_659 (O_659,N_19876,N_19675);
nor UO_660 (O_660,N_19800,N_19558);
nor UO_661 (O_661,N_19395,N_19720);
xnor UO_662 (O_662,N_19723,N_19757);
nand UO_663 (O_663,N_19857,N_19797);
nor UO_664 (O_664,N_19332,N_19502);
or UO_665 (O_665,N_19964,N_19719);
xnor UO_666 (O_666,N_19669,N_19431);
xnor UO_667 (O_667,N_19460,N_19503);
xnor UO_668 (O_668,N_19559,N_19490);
and UO_669 (O_669,N_19757,N_19529);
xor UO_670 (O_670,N_19721,N_19465);
and UO_671 (O_671,N_19219,N_19565);
and UO_672 (O_672,N_19921,N_19991);
xnor UO_673 (O_673,N_19766,N_19209);
nor UO_674 (O_674,N_19823,N_19742);
nor UO_675 (O_675,N_19425,N_19417);
and UO_676 (O_676,N_19296,N_19435);
or UO_677 (O_677,N_19314,N_19612);
nand UO_678 (O_678,N_19391,N_19270);
xnor UO_679 (O_679,N_19792,N_19849);
nand UO_680 (O_680,N_19993,N_19649);
nand UO_681 (O_681,N_19760,N_19998);
nand UO_682 (O_682,N_19301,N_19546);
and UO_683 (O_683,N_19395,N_19713);
and UO_684 (O_684,N_19464,N_19624);
nand UO_685 (O_685,N_19222,N_19544);
nor UO_686 (O_686,N_19928,N_19468);
or UO_687 (O_687,N_19471,N_19906);
nor UO_688 (O_688,N_19365,N_19965);
or UO_689 (O_689,N_19393,N_19835);
nor UO_690 (O_690,N_19477,N_19380);
nand UO_691 (O_691,N_19694,N_19853);
xnor UO_692 (O_692,N_19966,N_19608);
nor UO_693 (O_693,N_19201,N_19208);
xor UO_694 (O_694,N_19885,N_19403);
nand UO_695 (O_695,N_19852,N_19231);
xnor UO_696 (O_696,N_19597,N_19251);
or UO_697 (O_697,N_19400,N_19880);
nand UO_698 (O_698,N_19691,N_19815);
or UO_699 (O_699,N_19683,N_19803);
nand UO_700 (O_700,N_19933,N_19968);
and UO_701 (O_701,N_19823,N_19364);
nand UO_702 (O_702,N_19743,N_19451);
nor UO_703 (O_703,N_19530,N_19933);
xor UO_704 (O_704,N_19341,N_19400);
or UO_705 (O_705,N_19277,N_19697);
or UO_706 (O_706,N_19865,N_19436);
or UO_707 (O_707,N_19801,N_19293);
or UO_708 (O_708,N_19580,N_19381);
xor UO_709 (O_709,N_19314,N_19350);
xnor UO_710 (O_710,N_19219,N_19669);
nor UO_711 (O_711,N_19466,N_19416);
nor UO_712 (O_712,N_19449,N_19255);
nor UO_713 (O_713,N_19409,N_19243);
nand UO_714 (O_714,N_19870,N_19313);
xnor UO_715 (O_715,N_19542,N_19908);
nand UO_716 (O_716,N_19784,N_19320);
or UO_717 (O_717,N_19372,N_19709);
xnor UO_718 (O_718,N_19498,N_19471);
nor UO_719 (O_719,N_19466,N_19854);
xnor UO_720 (O_720,N_19897,N_19836);
xnor UO_721 (O_721,N_19485,N_19336);
nand UO_722 (O_722,N_19679,N_19950);
or UO_723 (O_723,N_19425,N_19406);
or UO_724 (O_724,N_19386,N_19942);
nor UO_725 (O_725,N_19476,N_19784);
and UO_726 (O_726,N_19829,N_19869);
or UO_727 (O_727,N_19690,N_19473);
nand UO_728 (O_728,N_19411,N_19755);
nor UO_729 (O_729,N_19667,N_19982);
or UO_730 (O_730,N_19334,N_19745);
nor UO_731 (O_731,N_19992,N_19436);
and UO_732 (O_732,N_19506,N_19302);
nand UO_733 (O_733,N_19667,N_19372);
nor UO_734 (O_734,N_19338,N_19347);
nor UO_735 (O_735,N_19752,N_19221);
xor UO_736 (O_736,N_19274,N_19548);
or UO_737 (O_737,N_19225,N_19421);
nor UO_738 (O_738,N_19219,N_19384);
or UO_739 (O_739,N_19362,N_19484);
and UO_740 (O_740,N_19273,N_19955);
nor UO_741 (O_741,N_19609,N_19513);
nand UO_742 (O_742,N_19757,N_19579);
nor UO_743 (O_743,N_19445,N_19691);
and UO_744 (O_744,N_19319,N_19519);
and UO_745 (O_745,N_19252,N_19315);
and UO_746 (O_746,N_19806,N_19365);
nand UO_747 (O_747,N_19393,N_19986);
nor UO_748 (O_748,N_19811,N_19440);
xor UO_749 (O_749,N_19999,N_19678);
and UO_750 (O_750,N_19896,N_19846);
or UO_751 (O_751,N_19391,N_19756);
nand UO_752 (O_752,N_19305,N_19761);
or UO_753 (O_753,N_19753,N_19772);
xor UO_754 (O_754,N_19499,N_19486);
xor UO_755 (O_755,N_19856,N_19423);
xor UO_756 (O_756,N_19376,N_19924);
nor UO_757 (O_757,N_19526,N_19375);
and UO_758 (O_758,N_19908,N_19740);
and UO_759 (O_759,N_19724,N_19299);
xor UO_760 (O_760,N_19996,N_19941);
nor UO_761 (O_761,N_19450,N_19957);
xor UO_762 (O_762,N_19576,N_19229);
xnor UO_763 (O_763,N_19246,N_19720);
xor UO_764 (O_764,N_19974,N_19944);
nor UO_765 (O_765,N_19430,N_19380);
xnor UO_766 (O_766,N_19843,N_19203);
nor UO_767 (O_767,N_19690,N_19608);
nor UO_768 (O_768,N_19274,N_19592);
or UO_769 (O_769,N_19970,N_19256);
and UO_770 (O_770,N_19847,N_19975);
nor UO_771 (O_771,N_19645,N_19428);
nor UO_772 (O_772,N_19867,N_19773);
nand UO_773 (O_773,N_19582,N_19466);
and UO_774 (O_774,N_19632,N_19254);
and UO_775 (O_775,N_19553,N_19509);
xnor UO_776 (O_776,N_19241,N_19838);
and UO_777 (O_777,N_19359,N_19320);
and UO_778 (O_778,N_19610,N_19978);
nor UO_779 (O_779,N_19947,N_19454);
xnor UO_780 (O_780,N_19222,N_19944);
and UO_781 (O_781,N_19972,N_19302);
xor UO_782 (O_782,N_19777,N_19400);
xnor UO_783 (O_783,N_19243,N_19649);
nand UO_784 (O_784,N_19915,N_19482);
xor UO_785 (O_785,N_19330,N_19575);
xnor UO_786 (O_786,N_19714,N_19291);
and UO_787 (O_787,N_19444,N_19902);
nand UO_788 (O_788,N_19620,N_19656);
and UO_789 (O_789,N_19652,N_19874);
and UO_790 (O_790,N_19863,N_19865);
xor UO_791 (O_791,N_19886,N_19281);
xnor UO_792 (O_792,N_19509,N_19711);
nand UO_793 (O_793,N_19587,N_19532);
or UO_794 (O_794,N_19368,N_19699);
xor UO_795 (O_795,N_19379,N_19376);
nor UO_796 (O_796,N_19632,N_19339);
xor UO_797 (O_797,N_19257,N_19316);
nand UO_798 (O_798,N_19353,N_19218);
xor UO_799 (O_799,N_19914,N_19778);
nor UO_800 (O_800,N_19782,N_19914);
or UO_801 (O_801,N_19215,N_19424);
or UO_802 (O_802,N_19942,N_19610);
or UO_803 (O_803,N_19204,N_19747);
nor UO_804 (O_804,N_19957,N_19855);
and UO_805 (O_805,N_19852,N_19512);
nand UO_806 (O_806,N_19971,N_19244);
nor UO_807 (O_807,N_19587,N_19739);
or UO_808 (O_808,N_19406,N_19635);
xnor UO_809 (O_809,N_19883,N_19632);
or UO_810 (O_810,N_19954,N_19985);
and UO_811 (O_811,N_19877,N_19643);
and UO_812 (O_812,N_19852,N_19855);
nor UO_813 (O_813,N_19640,N_19262);
nor UO_814 (O_814,N_19883,N_19228);
nand UO_815 (O_815,N_19663,N_19869);
nor UO_816 (O_816,N_19339,N_19284);
nand UO_817 (O_817,N_19831,N_19820);
or UO_818 (O_818,N_19517,N_19474);
nand UO_819 (O_819,N_19357,N_19396);
nor UO_820 (O_820,N_19393,N_19303);
xnor UO_821 (O_821,N_19272,N_19790);
and UO_822 (O_822,N_19584,N_19353);
nand UO_823 (O_823,N_19254,N_19531);
nand UO_824 (O_824,N_19907,N_19755);
xnor UO_825 (O_825,N_19392,N_19544);
xor UO_826 (O_826,N_19730,N_19255);
or UO_827 (O_827,N_19227,N_19599);
or UO_828 (O_828,N_19639,N_19803);
or UO_829 (O_829,N_19642,N_19414);
xnor UO_830 (O_830,N_19777,N_19973);
nand UO_831 (O_831,N_19912,N_19645);
nand UO_832 (O_832,N_19548,N_19246);
nor UO_833 (O_833,N_19730,N_19644);
and UO_834 (O_834,N_19247,N_19978);
and UO_835 (O_835,N_19763,N_19506);
nand UO_836 (O_836,N_19513,N_19610);
nand UO_837 (O_837,N_19322,N_19263);
or UO_838 (O_838,N_19349,N_19777);
or UO_839 (O_839,N_19395,N_19406);
or UO_840 (O_840,N_19343,N_19442);
and UO_841 (O_841,N_19641,N_19236);
nand UO_842 (O_842,N_19522,N_19687);
and UO_843 (O_843,N_19623,N_19478);
xor UO_844 (O_844,N_19336,N_19791);
nand UO_845 (O_845,N_19300,N_19768);
xor UO_846 (O_846,N_19917,N_19466);
and UO_847 (O_847,N_19389,N_19668);
nor UO_848 (O_848,N_19253,N_19994);
nand UO_849 (O_849,N_19883,N_19928);
and UO_850 (O_850,N_19308,N_19456);
nor UO_851 (O_851,N_19325,N_19603);
xnor UO_852 (O_852,N_19880,N_19263);
xor UO_853 (O_853,N_19951,N_19700);
nand UO_854 (O_854,N_19489,N_19249);
or UO_855 (O_855,N_19979,N_19340);
and UO_856 (O_856,N_19353,N_19342);
xor UO_857 (O_857,N_19889,N_19617);
nand UO_858 (O_858,N_19345,N_19717);
and UO_859 (O_859,N_19272,N_19871);
nand UO_860 (O_860,N_19702,N_19373);
nand UO_861 (O_861,N_19851,N_19840);
and UO_862 (O_862,N_19433,N_19469);
or UO_863 (O_863,N_19467,N_19964);
xnor UO_864 (O_864,N_19297,N_19755);
nor UO_865 (O_865,N_19618,N_19696);
and UO_866 (O_866,N_19934,N_19505);
xnor UO_867 (O_867,N_19695,N_19502);
nor UO_868 (O_868,N_19913,N_19772);
nand UO_869 (O_869,N_19679,N_19424);
nand UO_870 (O_870,N_19352,N_19698);
or UO_871 (O_871,N_19747,N_19347);
nand UO_872 (O_872,N_19847,N_19281);
nand UO_873 (O_873,N_19396,N_19413);
nand UO_874 (O_874,N_19973,N_19720);
nand UO_875 (O_875,N_19705,N_19805);
xnor UO_876 (O_876,N_19533,N_19815);
xor UO_877 (O_877,N_19378,N_19436);
and UO_878 (O_878,N_19532,N_19777);
xnor UO_879 (O_879,N_19935,N_19786);
nor UO_880 (O_880,N_19651,N_19641);
xnor UO_881 (O_881,N_19619,N_19544);
or UO_882 (O_882,N_19839,N_19633);
or UO_883 (O_883,N_19204,N_19705);
nor UO_884 (O_884,N_19968,N_19263);
xor UO_885 (O_885,N_19513,N_19306);
nand UO_886 (O_886,N_19210,N_19947);
nand UO_887 (O_887,N_19824,N_19205);
or UO_888 (O_888,N_19256,N_19280);
nor UO_889 (O_889,N_19813,N_19281);
nor UO_890 (O_890,N_19244,N_19797);
or UO_891 (O_891,N_19735,N_19691);
xor UO_892 (O_892,N_19708,N_19795);
nor UO_893 (O_893,N_19763,N_19649);
or UO_894 (O_894,N_19535,N_19254);
xor UO_895 (O_895,N_19953,N_19428);
and UO_896 (O_896,N_19425,N_19459);
xnor UO_897 (O_897,N_19355,N_19605);
or UO_898 (O_898,N_19349,N_19981);
xor UO_899 (O_899,N_19847,N_19308);
nor UO_900 (O_900,N_19419,N_19616);
xnor UO_901 (O_901,N_19929,N_19853);
and UO_902 (O_902,N_19676,N_19411);
and UO_903 (O_903,N_19813,N_19730);
and UO_904 (O_904,N_19351,N_19972);
and UO_905 (O_905,N_19430,N_19765);
or UO_906 (O_906,N_19735,N_19405);
or UO_907 (O_907,N_19855,N_19734);
nand UO_908 (O_908,N_19845,N_19277);
and UO_909 (O_909,N_19258,N_19504);
nand UO_910 (O_910,N_19628,N_19508);
and UO_911 (O_911,N_19858,N_19650);
nor UO_912 (O_912,N_19908,N_19944);
nand UO_913 (O_913,N_19610,N_19537);
and UO_914 (O_914,N_19227,N_19243);
xnor UO_915 (O_915,N_19899,N_19243);
nor UO_916 (O_916,N_19397,N_19805);
nand UO_917 (O_917,N_19789,N_19658);
or UO_918 (O_918,N_19825,N_19491);
or UO_919 (O_919,N_19554,N_19314);
and UO_920 (O_920,N_19895,N_19856);
or UO_921 (O_921,N_19247,N_19768);
xor UO_922 (O_922,N_19771,N_19781);
or UO_923 (O_923,N_19298,N_19221);
or UO_924 (O_924,N_19408,N_19434);
or UO_925 (O_925,N_19264,N_19532);
or UO_926 (O_926,N_19781,N_19471);
or UO_927 (O_927,N_19922,N_19205);
xnor UO_928 (O_928,N_19456,N_19859);
nand UO_929 (O_929,N_19588,N_19573);
xnor UO_930 (O_930,N_19254,N_19468);
xor UO_931 (O_931,N_19695,N_19838);
nand UO_932 (O_932,N_19642,N_19231);
or UO_933 (O_933,N_19222,N_19380);
and UO_934 (O_934,N_19454,N_19240);
xor UO_935 (O_935,N_19848,N_19704);
and UO_936 (O_936,N_19647,N_19822);
or UO_937 (O_937,N_19776,N_19916);
xnor UO_938 (O_938,N_19739,N_19349);
nor UO_939 (O_939,N_19827,N_19495);
nor UO_940 (O_940,N_19292,N_19826);
nand UO_941 (O_941,N_19419,N_19858);
xor UO_942 (O_942,N_19652,N_19953);
and UO_943 (O_943,N_19945,N_19765);
nor UO_944 (O_944,N_19456,N_19686);
xnor UO_945 (O_945,N_19761,N_19491);
and UO_946 (O_946,N_19698,N_19580);
nand UO_947 (O_947,N_19247,N_19854);
nand UO_948 (O_948,N_19987,N_19356);
xor UO_949 (O_949,N_19242,N_19688);
nand UO_950 (O_950,N_19755,N_19786);
nand UO_951 (O_951,N_19328,N_19494);
nor UO_952 (O_952,N_19559,N_19798);
and UO_953 (O_953,N_19870,N_19299);
nand UO_954 (O_954,N_19483,N_19779);
or UO_955 (O_955,N_19453,N_19919);
and UO_956 (O_956,N_19773,N_19872);
nand UO_957 (O_957,N_19201,N_19519);
nor UO_958 (O_958,N_19694,N_19398);
xor UO_959 (O_959,N_19859,N_19421);
xnor UO_960 (O_960,N_19539,N_19879);
xor UO_961 (O_961,N_19299,N_19435);
or UO_962 (O_962,N_19389,N_19219);
xnor UO_963 (O_963,N_19440,N_19647);
xor UO_964 (O_964,N_19442,N_19970);
xor UO_965 (O_965,N_19551,N_19831);
nor UO_966 (O_966,N_19274,N_19514);
nor UO_967 (O_967,N_19905,N_19421);
nor UO_968 (O_968,N_19392,N_19313);
and UO_969 (O_969,N_19774,N_19706);
nand UO_970 (O_970,N_19378,N_19615);
and UO_971 (O_971,N_19874,N_19293);
and UO_972 (O_972,N_19984,N_19467);
or UO_973 (O_973,N_19796,N_19626);
nand UO_974 (O_974,N_19401,N_19802);
nor UO_975 (O_975,N_19837,N_19573);
or UO_976 (O_976,N_19484,N_19594);
xor UO_977 (O_977,N_19753,N_19383);
and UO_978 (O_978,N_19371,N_19376);
and UO_979 (O_979,N_19930,N_19516);
xor UO_980 (O_980,N_19465,N_19976);
xnor UO_981 (O_981,N_19767,N_19798);
xor UO_982 (O_982,N_19464,N_19917);
nor UO_983 (O_983,N_19457,N_19916);
or UO_984 (O_984,N_19519,N_19464);
nor UO_985 (O_985,N_19982,N_19950);
nand UO_986 (O_986,N_19501,N_19235);
nor UO_987 (O_987,N_19728,N_19270);
xor UO_988 (O_988,N_19617,N_19942);
nor UO_989 (O_989,N_19658,N_19902);
nand UO_990 (O_990,N_19568,N_19808);
and UO_991 (O_991,N_19329,N_19671);
xnor UO_992 (O_992,N_19412,N_19371);
nand UO_993 (O_993,N_19411,N_19417);
nand UO_994 (O_994,N_19621,N_19841);
nand UO_995 (O_995,N_19732,N_19857);
xor UO_996 (O_996,N_19435,N_19850);
and UO_997 (O_997,N_19500,N_19536);
nand UO_998 (O_998,N_19926,N_19737);
xnor UO_999 (O_999,N_19749,N_19839);
xnor UO_1000 (O_1000,N_19601,N_19567);
xor UO_1001 (O_1001,N_19745,N_19324);
or UO_1002 (O_1002,N_19327,N_19933);
and UO_1003 (O_1003,N_19961,N_19984);
or UO_1004 (O_1004,N_19232,N_19247);
and UO_1005 (O_1005,N_19537,N_19699);
and UO_1006 (O_1006,N_19941,N_19466);
and UO_1007 (O_1007,N_19586,N_19867);
xnor UO_1008 (O_1008,N_19715,N_19585);
nor UO_1009 (O_1009,N_19541,N_19393);
nand UO_1010 (O_1010,N_19711,N_19229);
nor UO_1011 (O_1011,N_19863,N_19774);
and UO_1012 (O_1012,N_19857,N_19605);
nor UO_1013 (O_1013,N_19976,N_19288);
and UO_1014 (O_1014,N_19227,N_19697);
nand UO_1015 (O_1015,N_19391,N_19639);
or UO_1016 (O_1016,N_19602,N_19834);
xnor UO_1017 (O_1017,N_19957,N_19285);
or UO_1018 (O_1018,N_19492,N_19751);
nor UO_1019 (O_1019,N_19855,N_19823);
xor UO_1020 (O_1020,N_19840,N_19420);
and UO_1021 (O_1021,N_19380,N_19328);
nand UO_1022 (O_1022,N_19976,N_19363);
nor UO_1023 (O_1023,N_19317,N_19840);
and UO_1024 (O_1024,N_19570,N_19583);
nor UO_1025 (O_1025,N_19615,N_19872);
or UO_1026 (O_1026,N_19718,N_19568);
xor UO_1027 (O_1027,N_19756,N_19996);
xor UO_1028 (O_1028,N_19294,N_19318);
nand UO_1029 (O_1029,N_19475,N_19684);
xor UO_1030 (O_1030,N_19397,N_19996);
or UO_1031 (O_1031,N_19309,N_19819);
nor UO_1032 (O_1032,N_19355,N_19747);
nand UO_1033 (O_1033,N_19560,N_19462);
or UO_1034 (O_1034,N_19399,N_19380);
xor UO_1035 (O_1035,N_19510,N_19846);
nand UO_1036 (O_1036,N_19692,N_19520);
or UO_1037 (O_1037,N_19764,N_19716);
nor UO_1038 (O_1038,N_19517,N_19406);
nand UO_1039 (O_1039,N_19786,N_19804);
xor UO_1040 (O_1040,N_19807,N_19740);
or UO_1041 (O_1041,N_19331,N_19906);
xnor UO_1042 (O_1042,N_19733,N_19410);
nor UO_1043 (O_1043,N_19349,N_19293);
nand UO_1044 (O_1044,N_19248,N_19599);
xor UO_1045 (O_1045,N_19586,N_19736);
or UO_1046 (O_1046,N_19465,N_19626);
and UO_1047 (O_1047,N_19803,N_19727);
nand UO_1048 (O_1048,N_19931,N_19995);
xor UO_1049 (O_1049,N_19657,N_19519);
nor UO_1050 (O_1050,N_19821,N_19852);
nor UO_1051 (O_1051,N_19241,N_19515);
and UO_1052 (O_1052,N_19755,N_19805);
nand UO_1053 (O_1053,N_19407,N_19301);
xnor UO_1054 (O_1054,N_19643,N_19806);
xnor UO_1055 (O_1055,N_19858,N_19503);
or UO_1056 (O_1056,N_19695,N_19868);
and UO_1057 (O_1057,N_19351,N_19550);
nand UO_1058 (O_1058,N_19615,N_19265);
and UO_1059 (O_1059,N_19900,N_19849);
xnor UO_1060 (O_1060,N_19235,N_19982);
xor UO_1061 (O_1061,N_19737,N_19205);
or UO_1062 (O_1062,N_19256,N_19569);
xnor UO_1063 (O_1063,N_19358,N_19213);
nand UO_1064 (O_1064,N_19802,N_19805);
or UO_1065 (O_1065,N_19553,N_19798);
xnor UO_1066 (O_1066,N_19756,N_19915);
and UO_1067 (O_1067,N_19485,N_19529);
and UO_1068 (O_1068,N_19440,N_19769);
nand UO_1069 (O_1069,N_19923,N_19693);
or UO_1070 (O_1070,N_19605,N_19892);
and UO_1071 (O_1071,N_19323,N_19359);
nand UO_1072 (O_1072,N_19714,N_19861);
nand UO_1073 (O_1073,N_19359,N_19395);
nor UO_1074 (O_1074,N_19838,N_19221);
nand UO_1075 (O_1075,N_19803,N_19706);
or UO_1076 (O_1076,N_19292,N_19206);
and UO_1077 (O_1077,N_19256,N_19975);
or UO_1078 (O_1078,N_19422,N_19513);
xnor UO_1079 (O_1079,N_19419,N_19274);
and UO_1080 (O_1080,N_19710,N_19555);
xnor UO_1081 (O_1081,N_19739,N_19521);
nand UO_1082 (O_1082,N_19576,N_19232);
or UO_1083 (O_1083,N_19257,N_19605);
and UO_1084 (O_1084,N_19209,N_19910);
xor UO_1085 (O_1085,N_19892,N_19806);
and UO_1086 (O_1086,N_19667,N_19637);
xnor UO_1087 (O_1087,N_19330,N_19304);
xnor UO_1088 (O_1088,N_19971,N_19540);
xor UO_1089 (O_1089,N_19287,N_19704);
nand UO_1090 (O_1090,N_19845,N_19782);
and UO_1091 (O_1091,N_19694,N_19670);
and UO_1092 (O_1092,N_19528,N_19596);
xnor UO_1093 (O_1093,N_19448,N_19900);
and UO_1094 (O_1094,N_19878,N_19269);
xor UO_1095 (O_1095,N_19768,N_19502);
or UO_1096 (O_1096,N_19507,N_19828);
xnor UO_1097 (O_1097,N_19932,N_19745);
and UO_1098 (O_1098,N_19673,N_19714);
nor UO_1099 (O_1099,N_19247,N_19544);
nor UO_1100 (O_1100,N_19881,N_19413);
nand UO_1101 (O_1101,N_19363,N_19941);
and UO_1102 (O_1102,N_19723,N_19396);
nor UO_1103 (O_1103,N_19427,N_19974);
nor UO_1104 (O_1104,N_19763,N_19522);
and UO_1105 (O_1105,N_19273,N_19553);
nor UO_1106 (O_1106,N_19878,N_19787);
or UO_1107 (O_1107,N_19823,N_19332);
nor UO_1108 (O_1108,N_19819,N_19341);
or UO_1109 (O_1109,N_19576,N_19678);
nor UO_1110 (O_1110,N_19350,N_19934);
xnor UO_1111 (O_1111,N_19785,N_19568);
nand UO_1112 (O_1112,N_19909,N_19828);
xor UO_1113 (O_1113,N_19786,N_19257);
and UO_1114 (O_1114,N_19908,N_19692);
xor UO_1115 (O_1115,N_19344,N_19345);
nor UO_1116 (O_1116,N_19791,N_19777);
xnor UO_1117 (O_1117,N_19737,N_19252);
nor UO_1118 (O_1118,N_19791,N_19566);
or UO_1119 (O_1119,N_19289,N_19483);
or UO_1120 (O_1120,N_19701,N_19984);
nand UO_1121 (O_1121,N_19465,N_19440);
nor UO_1122 (O_1122,N_19856,N_19583);
nor UO_1123 (O_1123,N_19699,N_19732);
or UO_1124 (O_1124,N_19720,N_19484);
xor UO_1125 (O_1125,N_19880,N_19852);
and UO_1126 (O_1126,N_19684,N_19687);
xnor UO_1127 (O_1127,N_19947,N_19987);
and UO_1128 (O_1128,N_19711,N_19855);
and UO_1129 (O_1129,N_19388,N_19896);
nor UO_1130 (O_1130,N_19365,N_19284);
nor UO_1131 (O_1131,N_19815,N_19895);
nand UO_1132 (O_1132,N_19453,N_19499);
nor UO_1133 (O_1133,N_19709,N_19405);
nand UO_1134 (O_1134,N_19914,N_19422);
nor UO_1135 (O_1135,N_19726,N_19763);
nand UO_1136 (O_1136,N_19465,N_19300);
and UO_1137 (O_1137,N_19749,N_19848);
nor UO_1138 (O_1138,N_19393,N_19976);
or UO_1139 (O_1139,N_19742,N_19894);
or UO_1140 (O_1140,N_19860,N_19840);
nand UO_1141 (O_1141,N_19599,N_19508);
or UO_1142 (O_1142,N_19890,N_19969);
or UO_1143 (O_1143,N_19321,N_19543);
and UO_1144 (O_1144,N_19200,N_19424);
nand UO_1145 (O_1145,N_19670,N_19754);
or UO_1146 (O_1146,N_19960,N_19890);
and UO_1147 (O_1147,N_19989,N_19926);
and UO_1148 (O_1148,N_19585,N_19429);
nor UO_1149 (O_1149,N_19253,N_19266);
nand UO_1150 (O_1150,N_19294,N_19820);
xnor UO_1151 (O_1151,N_19367,N_19765);
and UO_1152 (O_1152,N_19712,N_19815);
and UO_1153 (O_1153,N_19720,N_19616);
nor UO_1154 (O_1154,N_19912,N_19788);
and UO_1155 (O_1155,N_19824,N_19735);
nand UO_1156 (O_1156,N_19893,N_19320);
nand UO_1157 (O_1157,N_19912,N_19354);
nand UO_1158 (O_1158,N_19548,N_19410);
and UO_1159 (O_1159,N_19411,N_19938);
and UO_1160 (O_1160,N_19986,N_19420);
or UO_1161 (O_1161,N_19206,N_19812);
xor UO_1162 (O_1162,N_19686,N_19594);
and UO_1163 (O_1163,N_19907,N_19642);
nor UO_1164 (O_1164,N_19385,N_19980);
nor UO_1165 (O_1165,N_19553,N_19861);
xnor UO_1166 (O_1166,N_19393,N_19363);
xnor UO_1167 (O_1167,N_19633,N_19754);
or UO_1168 (O_1168,N_19862,N_19578);
nand UO_1169 (O_1169,N_19998,N_19466);
and UO_1170 (O_1170,N_19335,N_19419);
nand UO_1171 (O_1171,N_19336,N_19853);
nand UO_1172 (O_1172,N_19415,N_19864);
xor UO_1173 (O_1173,N_19953,N_19214);
xor UO_1174 (O_1174,N_19856,N_19514);
xnor UO_1175 (O_1175,N_19405,N_19224);
and UO_1176 (O_1176,N_19965,N_19382);
nor UO_1177 (O_1177,N_19290,N_19582);
nand UO_1178 (O_1178,N_19821,N_19206);
nor UO_1179 (O_1179,N_19616,N_19855);
nor UO_1180 (O_1180,N_19274,N_19387);
nor UO_1181 (O_1181,N_19674,N_19971);
xnor UO_1182 (O_1182,N_19396,N_19336);
xor UO_1183 (O_1183,N_19746,N_19612);
nor UO_1184 (O_1184,N_19579,N_19411);
xor UO_1185 (O_1185,N_19201,N_19997);
nor UO_1186 (O_1186,N_19463,N_19483);
nand UO_1187 (O_1187,N_19710,N_19890);
and UO_1188 (O_1188,N_19548,N_19711);
nand UO_1189 (O_1189,N_19508,N_19683);
and UO_1190 (O_1190,N_19411,N_19935);
or UO_1191 (O_1191,N_19308,N_19807);
xnor UO_1192 (O_1192,N_19251,N_19818);
nand UO_1193 (O_1193,N_19229,N_19549);
nand UO_1194 (O_1194,N_19962,N_19796);
nand UO_1195 (O_1195,N_19982,N_19995);
or UO_1196 (O_1196,N_19585,N_19327);
xor UO_1197 (O_1197,N_19526,N_19249);
nand UO_1198 (O_1198,N_19774,N_19810);
nor UO_1199 (O_1199,N_19691,N_19876);
nor UO_1200 (O_1200,N_19970,N_19938);
xor UO_1201 (O_1201,N_19805,N_19523);
and UO_1202 (O_1202,N_19902,N_19275);
nand UO_1203 (O_1203,N_19648,N_19489);
nand UO_1204 (O_1204,N_19328,N_19650);
xnor UO_1205 (O_1205,N_19573,N_19741);
nand UO_1206 (O_1206,N_19813,N_19419);
and UO_1207 (O_1207,N_19567,N_19360);
nand UO_1208 (O_1208,N_19333,N_19692);
or UO_1209 (O_1209,N_19568,N_19499);
nor UO_1210 (O_1210,N_19859,N_19957);
and UO_1211 (O_1211,N_19539,N_19774);
or UO_1212 (O_1212,N_19761,N_19234);
or UO_1213 (O_1213,N_19954,N_19444);
nor UO_1214 (O_1214,N_19910,N_19530);
nand UO_1215 (O_1215,N_19517,N_19520);
or UO_1216 (O_1216,N_19619,N_19607);
nand UO_1217 (O_1217,N_19761,N_19910);
xnor UO_1218 (O_1218,N_19674,N_19979);
or UO_1219 (O_1219,N_19526,N_19977);
xnor UO_1220 (O_1220,N_19964,N_19595);
xnor UO_1221 (O_1221,N_19307,N_19630);
nor UO_1222 (O_1222,N_19926,N_19819);
xnor UO_1223 (O_1223,N_19226,N_19243);
nor UO_1224 (O_1224,N_19504,N_19491);
and UO_1225 (O_1225,N_19769,N_19765);
or UO_1226 (O_1226,N_19317,N_19812);
nor UO_1227 (O_1227,N_19295,N_19212);
nor UO_1228 (O_1228,N_19483,N_19447);
nand UO_1229 (O_1229,N_19736,N_19452);
nand UO_1230 (O_1230,N_19372,N_19577);
or UO_1231 (O_1231,N_19924,N_19639);
or UO_1232 (O_1232,N_19402,N_19893);
nor UO_1233 (O_1233,N_19784,N_19762);
and UO_1234 (O_1234,N_19888,N_19983);
xor UO_1235 (O_1235,N_19440,N_19969);
or UO_1236 (O_1236,N_19911,N_19753);
nor UO_1237 (O_1237,N_19252,N_19261);
or UO_1238 (O_1238,N_19918,N_19409);
and UO_1239 (O_1239,N_19855,N_19342);
nor UO_1240 (O_1240,N_19453,N_19205);
and UO_1241 (O_1241,N_19605,N_19290);
nand UO_1242 (O_1242,N_19728,N_19230);
nand UO_1243 (O_1243,N_19472,N_19908);
and UO_1244 (O_1244,N_19289,N_19512);
and UO_1245 (O_1245,N_19928,N_19899);
and UO_1246 (O_1246,N_19893,N_19287);
nor UO_1247 (O_1247,N_19974,N_19858);
and UO_1248 (O_1248,N_19374,N_19243);
or UO_1249 (O_1249,N_19663,N_19940);
or UO_1250 (O_1250,N_19379,N_19510);
nor UO_1251 (O_1251,N_19697,N_19878);
xnor UO_1252 (O_1252,N_19509,N_19421);
nor UO_1253 (O_1253,N_19469,N_19815);
nor UO_1254 (O_1254,N_19789,N_19998);
nor UO_1255 (O_1255,N_19386,N_19564);
and UO_1256 (O_1256,N_19578,N_19896);
nor UO_1257 (O_1257,N_19225,N_19306);
nand UO_1258 (O_1258,N_19523,N_19560);
nand UO_1259 (O_1259,N_19798,N_19597);
xor UO_1260 (O_1260,N_19604,N_19683);
nor UO_1261 (O_1261,N_19333,N_19563);
and UO_1262 (O_1262,N_19966,N_19680);
nand UO_1263 (O_1263,N_19269,N_19418);
and UO_1264 (O_1264,N_19700,N_19739);
xnor UO_1265 (O_1265,N_19373,N_19611);
or UO_1266 (O_1266,N_19364,N_19785);
or UO_1267 (O_1267,N_19712,N_19520);
xnor UO_1268 (O_1268,N_19772,N_19613);
nor UO_1269 (O_1269,N_19333,N_19961);
or UO_1270 (O_1270,N_19380,N_19928);
xnor UO_1271 (O_1271,N_19433,N_19895);
or UO_1272 (O_1272,N_19729,N_19344);
nand UO_1273 (O_1273,N_19398,N_19493);
nand UO_1274 (O_1274,N_19749,N_19844);
nor UO_1275 (O_1275,N_19668,N_19827);
nor UO_1276 (O_1276,N_19442,N_19880);
or UO_1277 (O_1277,N_19842,N_19826);
nand UO_1278 (O_1278,N_19512,N_19547);
nor UO_1279 (O_1279,N_19613,N_19741);
and UO_1280 (O_1280,N_19328,N_19737);
or UO_1281 (O_1281,N_19414,N_19689);
and UO_1282 (O_1282,N_19434,N_19468);
nand UO_1283 (O_1283,N_19730,N_19243);
xnor UO_1284 (O_1284,N_19874,N_19735);
nand UO_1285 (O_1285,N_19633,N_19855);
nand UO_1286 (O_1286,N_19395,N_19202);
xor UO_1287 (O_1287,N_19842,N_19388);
and UO_1288 (O_1288,N_19935,N_19641);
xnor UO_1289 (O_1289,N_19672,N_19337);
or UO_1290 (O_1290,N_19341,N_19619);
and UO_1291 (O_1291,N_19605,N_19521);
or UO_1292 (O_1292,N_19719,N_19645);
and UO_1293 (O_1293,N_19704,N_19476);
and UO_1294 (O_1294,N_19291,N_19225);
nor UO_1295 (O_1295,N_19787,N_19757);
nand UO_1296 (O_1296,N_19699,N_19581);
or UO_1297 (O_1297,N_19449,N_19677);
xnor UO_1298 (O_1298,N_19782,N_19365);
nand UO_1299 (O_1299,N_19394,N_19778);
nand UO_1300 (O_1300,N_19586,N_19768);
xor UO_1301 (O_1301,N_19706,N_19248);
and UO_1302 (O_1302,N_19411,N_19401);
xor UO_1303 (O_1303,N_19575,N_19790);
or UO_1304 (O_1304,N_19370,N_19256);
or UO_1305 (O_1305,N_19267,N_19785);
xor UO_1306 (O_1306,N_19869,N_19530);
or UO_1307 (O_1307,N_19599,N_19428);
or UO_1308 (O_1308,N_19367,N_19539);
and UO_1309 (O_1309,N_19874,N_19562);
nand UO_1310 (O_1310,N_19694,N_19768);
xor UO_1311 (O_1311,N_19510,N_19781);
nand UO_1312 (O_1312,N_19910,N_19234);
nor UO_1313 (O_1313,N_19984,N_19371);
nand UO_1314 (O_1314,N_19479,N_19513);
and UO_1315 (O_1315,N_19762,N_19907);
or UO_1316 (O_1316,N_19331,N_19255);
xnor UO_1317 (O_1317,N_19543,N_19419);
and UO_1318 (O_1318,N_19358,N_19831);
nor UO_1319 (O_1319,N_19705,N_19345);
or UO_1320 (O_1320,N_19536,N_19795);
xor UO_1321 (O_1321,N_19624,N_19999);
and UO_1322 (O_1322,N_19237,N_19391);
xor UO_1323 (O_1323,N_19844,N_19416);
xnor UO_1324 (O_1324,N_19553,N_19305);
xnor UO_1325 (O_1325,N_19487,N_19426);
nand UO_1326 (O_1326,N_19676,N_19703);
nand UO_1327 (O_1327,N_19630,N_19557);
or UO_1328 (O_1328,N_19461,N_19950);
nand UO_1329 (O_1329,N_19998,N_19898);
xnor UO_1330 (O_1330,N_19670,N_19611);
xor UO_1331 (O_1331,N_19827,N_19296);
or UO_1332 (O_1332,N_19545,N_19993);
nand UO_1333 (O_1333,N_19932,N_19665);
nor UO_1334 (O_1334,N_19263,N_19876);
and UO_1335 (O_1335,N_19702,N_19522);
nor UO_1336 (O_1336,N_19587,N_19697);
nand UO_1337 (O_1337,N_19289,N_19494);
xor UO_1338 (O_1338,N_19633,N_19430);
xnor UO_1339 (O_1339,N_19454,N_19261);
and UO_1340 (O_1340,N_19300,N_19593);
nand UO_1341 (O_1341,N_19961,N_19846);
xnor UO_1342 (O_1342,N_19934,N_19787);
nor UO_1343 (O_1343,N_19305,N_19961);
and UO_1344 (O_1344,N_19587,N_19753);
nand UO_1345 (O_1345,N_19641,N_19447);
and UO_1346 (O_1346,N_19767,N_19326);
and UO_1347 (O_1347,N_19685,N_19288);
and UO_1348 (O_1348,N_19552,N_19273);
nand UO_1349 (O_1349,N_19739,N_19863);
nor UO_1350 (O_1350,N_19335,N_19350);
xnor UO_1351 (O_1351,N_19722,N_19285);
nand UO_1352 (O_1352,N_19693,N_19643);
or UO_1353 (O_1353,N_19819,N_19883);
and UO_1354 (O_1354,N_19728,N_19397);
and UO_1355 (O_1355,N_19316,N_19612);
nand UO_1356 (O_1356,N_19298,N_19529);
or UO_1357 (O_1357,N_19548,N_19896);
nand UO_1358 (O_1358,N_19733,N_19485);
xor UO_1359 (O_1359,N_19803,N_19769);
or UO_1360 (O_1360,N_19715,N_19755);
nand UO_1361 (O_1361,N_19698,N_19286);
nand UO_1362 (O_1362,N_19994,N_19928);
nor UO_1363 (O_1363,N_19665,N_19712);
nor UO_1364 (O_1364,N_19847,N_19468);
or UO_1365 (O_1365,N_19954,N_19638);
nor UO_1366 (O_1366,N_19648,N_19832);
nand UO_1367 (O_1367,N_19974,N_19895);
and UO_1368 (O_1368,N_19482,N_19216);
nand UO_1369 (O_1369,N_19966,N_19482);
and UO_1370 (O_1370,N_19796,N_19821);
or UO_1371 (O_1371,N_19222,N_19356);
or UO_1372 (O_1372,N_19574,N_19561);
nand UO_1373 (O_1373,N_19845,N_19593);
nor UO_1374 (O_1374,N_19558,N_19724);
and UO_1375 (O_1375,N_19785,N_19866);
or UO_1376 (O_1376,N_19749,N_19798);
nand UO_1377 (O_1377,N_19633,N_19529);
nor UO_1378 (O_1378,N_19330,N_19854);
nor UO_1379 (O_1379,N_19569,N_19799);
nand UO_1380 (O_1380,N_19986,N_19841);
nor UO_1381 (O_1381,N_19897,N_19499);
nand UO_1382 (O_1382,N_19869,N_19222);
and UO_1383 (O_1383,N_19729,N_19246);
nor UO_1384 (O_1384,N_19905,N_19963);
and UO_1385 (O_1385,N_19874,N_19414);
and UO_1386 (O_1386,N_19702,N_19291);
xnor UO_1387 (O_1387,N_19407,N_19787);
or UO_1388 (O_1388,N_19980,N_19420);
nand UO_1389 (O_1389,N_19348,N_19484);
nor UO_1390 (O_1390,N_19293,N_19810);
nor UO_1391 (O_1391,N_19798,N_19534);
xnor UO_1392 (O_1392,N_19248,N_19401);
xnor UO_1393 (O_1393,N_19419,N_19828);
nand UO_1394 (O_1394,N_19653,N_19967);
or UO_1395 (O_1395,N_19786,N_19922);
nor UO_1396 (O_1396,N_19557,N_19697);
xnor UO_1397 (O_1397,N_19808,N_19500);
and UO_1398 (O_1398,N_19741,N_19620);
nor UO_1399 (O_1399,N_19262,N_19389);
nand UO_1400 (O_1400,N_19421,N_19929);
nand UO_1401 (O_1401,N_19524,N_19748);
or UO_1402 (O_1402,N_19716,N_19625);
nor UO_1403 (O_1403,N_19456,N_19319);
nand UO_1404 (O_1404,N_19516,N_19819);
xor UO_1405 (O_1405,N_19616,N_19200);
or UO_1406 (O_1406,N_19327,N_19859);
nor UO_1407 (O_1407,N_19779,N_19374);
nand UO_1408 (O_1408,N_19532,N_19717);
or UO_1409 (O_1409,N_19323,N_19823);
or UO_1410 (O_1410,N_19592,N_19606);
xor UO_1411 (O_1411,N_19978,N_19580);
and UO_1412 (O_1412,N_19936,N_19471);
and UO_1413 (O_1413,N_19556,N_19538);
nor UO_1414 (O_1414,N_19704,N_19883);
or UO_1415 (O_1415,N_19790,N_19471);
and UO_1416 (O_1416,N_19300,N_19212);
nand UO_1417 (O_1417,N_19524,N_19243);
or UO_1418 (O_1418,N_19732,N_19958);
and UO_1419 (O_1419,N_19275,N_19919);
nand UO_1420 (O_1420,N_19730,N_19670);
nand UO_1421 (O_1421,N_19545,N_19421);
nor UO_1422 (O_1422,N_19908,N_19900);
xnor UO_1423 (O_1423,N_19310,N_19467);
or UO_1424 (O_1424,N_19973,N_19748);
or UO_1425 (O_1425,N_19578,N_19979);
and UO_1426 (O_1426,N_19587,N_19717);
or UO_1427 (O_1427,N_19606,N_19499);
or UO_1428 (O_1428,N_19589,N_19575);
nor UO_1429 (O_1429,N_19338,N_19595);
nand UO_1430 (O_1430,N_19880,N_19428);
nor UO_1431 (O_1431,N_19950,N_19870);
nand UO_1432 (O_1432,N_19601,N_19383);
xnor UO_1433 (O_1433,N_19706,N_19730);
nor UO_1434 (O_1434,N_19454,N_19746);
xor UO_1435 (O_1435,N_19394,N_19288);
or UO_1436 (O_1436,N_19448,N_19285);
or UO_1437 (O_1437,N_19243,N_19571);
or UO_1438 (O_1438,N_19877,N_19506);
nand UO_1439 (O_1439,N_19953,N_19207);
nor UO_1440 (O_1440,N_19978,N_19483);
nand UO_1441 (O_1441,N_19391,N_19951);
nand UO_1442 (O_1442,N_19623,N_19695);
and UO_1443 (O_1443,N_19500,N_19389);
or UO_1444 (O_1444,N_19811,N_19792);
nor UO_1445 (O_1445,N_19448,N_19915);
xor UO_1446 (O_1446,N_19319,N_19555);
and UO_1447 (O_1447,N_19320,N_19415);
or UO_1448 (O_1448,N_19548,N_19310);
nand UO_1449 (O_1449,N_19512,N_19670);
nand UO_1450 (O_1450,N_19868,N_19663);
or UO_1451 (O_1451,N_19433,N_19889);
xnor UO_1452 (O_1452,N_19641,N_19764);
or UO_1453 (O_1453,N_19298,N_19522);
nand UO_1454 (O_1454,N_19696,N_19805);
and UO_1455 (O_1455,N_19547,N_19624);
and UO_1456 (O_1456,N_19297,N_19966);
xnor UO_1457 (O_1457,N_19813,N_19549);
and UO_1458 (O_1458,N_19580,N_19578);
or UO_1459 (O_1459,N_19967,N_19629);
nand UO_1460 (O_1460,N_19236,N_19337);
and UO_1461 (O_1461,N_19345,N_19522);
and UO_1462 (O_1462,N_19261,N_19637);
and UO_1463 (O_1463,N_19399,N_19930);
or UO_1464 (O_1464,N_19600,N_19989);
nor UO_1465 (O_1465,N_19980,N_19933);
nor UO_1466 (O_1466,N_19471,N_19415);
or UO_1467 (O_1467,N_19359,N_19215);
and UO_1468 (O_1468,N_19342,N_19478);
xnor UO_1469 (O_1469,N_19419,N_19969);
and UO_1470 (O_1470,N_19795,N_19521);
or UO_1471 (O_1471,N_19664,N_19416);
xor UO_1472 (O_1472,N_19289,N_19507);
nor UO_1473 (O_1473,N_19832,N_19815);
xor UO_1474 (O_1474,N_19463,N_19536);
nand UO_1475 (O_1475,N_19305,N_19464);
or UO_1476 (O_1476,N_19394,N_19795);
xnor UO_1477 (O_1477,N_19556,N_19944);
nand UO_1478 (O_1478,N_19733,N_19728);
xnor UO_1479 (O_1479,N_19907,N_19882);
nor UO_1480 (O_1480,N_19344,N_19630);
nand UO_1481 (O_1481,N_19383,N_19734);
or UO_1482 (O_1482,N_19561,N_19696);
and UO_1483 (O_1483,N_19787,N_19370);
and UO_1484 (O_1484,N_19878,N_19756);
xnor UO_1485 (O_1485,N_19741,N_19736);
and UO_1486 (O_1486,N_19391,N_19620);
or UO_1487 (O_1487,N_19891,N_19777);
xnor UO_1488 (O_1488,N_19950,N_19539);
nor UO_1489 (O_1489,N_19494,N_19389);
xnor UO_1490 (O_1490,N_19715,N_19440);
and UO_1491 (O_1491,N_19941,N_19311);
nor UO_1492 (O_1492,N_19242,N_19850);
and UO_1493 (O_1493,N_19888,N_19400);
nor UO_1494 (O_1494,N_19413,N_19522);
and UO_1495 (O_1495,N_19900,N_19817);
xor UO_1496 (O_1496,N_19406,N_19831);
xor UO_1497 (O_1497,N_19687,N_19863);
nand UO_1498 (O_1498,N_19954,N_19975);
and UO_1499 (O_1499,N_19970,N_19754);
or UO_1500 (O_1500,N_19623,N_19966);
nand UO_1501 (O_1501,N_19238,N_19908);
nor UO_1502 (O_1502,N_19534,N_19718);
nor UO_1503 (O_1503,N_19971,N_19944);
nor UO_1504 (O_1504,N_19685,N_19388);
and UO_1505 (O_1505,N_19842,N_19378);
xor UO_1506 (O_1506,N_19384,N_19354);
xor UO_1507 (O_1507,N_19494,N_19956);
nor UO_1508 (O_1508,N_19952,N_19471);
xnor UO_1509 (O_1509,N_19666,N_19782);
nor UO_1510 (O_1510,N_19858,N_19989);
xor UO_1511 (O_1511,N_19597,N_19793);
nand UO_1512 (O_1512,N_19503,N_19555);
nor UO_1513 (O_1513,N_19905,N_19600);
xor UO_1514 (O_1514,N_19660,N_19807);
xor UO_1515 (O_1515,N_19438,N_19602);
nand UO_1516 (O_1516,N_19745,N_19234);
nand UO_1517 (O_1517,N_19429,N_19457);
or UO_1518 (O_1518,N_19552,N_19829);
and UO_1519 (O_1519,N_19933,N_19423);
nor UO_1520 (O_1520,N_19906,N_19645);
or UO_1521 (O_1521,N_19902,N_19283);
xor UO_1522 (O_1522,N_19297,N_19373);
xnor UO_1523 (O_1523,N_19253,N_19335);
nor UO_1524 (O_1524,N_19930,N_19519);
or UO_1525 (O_1525,N_19898,N_19999);
xnor UO_1526 (O_1526,N_19411,N_19399);
nand UO_1527 (O_1527,N_19959,N_19383);
xnor UO_1528 (O_1528,N_19351,N_19580);
nor UO_1529 (O_1529,N_19797,N_19796);
nand UO_1530 (O_1530,N_19606,N_19825);
nand UO_1531 (O_1531,N_19921,N_19754);
xnor UO_1532 (O_1532,N_19399,N_19341);
xor UO_1533 (O_1533,N_19718,N_19844);
or UO_1534 (O_1534,N_19684,N_19455);
and UO_1535 (O_1535,N_19977,N_19736);
nor UO_1536 (O_1536,N_19250,N_19378);
xor UO_1537 (O_1537,N_19871,N_19213);
and UO_1538 (O_1538,N_19960,N_19887);
and UO_1539 (O_1539,N_19311,N_19863);
or UO_1540 (O_1540,N_19687,N_19214);
or UO_1541 (O_1541,N_19650,N_19304);
and UO_1542 (O_1542,N_19739,N_19933);
or UO_1543 (O_1543,N_19340,N_19787);
nand UO_1544 (O_1544,N_19415,N_19547);
and UO_1545 (O_1545,N_19636,N_19915);
or UO_1546 (O_1546,N_19521,N_19533);
nor UO_1547 (O_1547,N_19764,N_19843);
and UO_1548 (O_1548,N_19554,N_19703);
nand UO_1549 (O_1549,N_19668,N_19730);
or UO_1550 (O_1550,N_19238,N_19321);
xnor UO_1551 (O_1551,N_19309,N_19844);
or UO_1552 (O_1552,N_19522,N_19332);
and UO_1553 (O_1553,N_19687,N_19751);
nand UO_1554 (O_1554,N_19668,N_19838);
nor UO_1555 (O_1555,N_19674,N_19360);
xor UO_1556 (O_1556,N_19537,N_19876);
xnor UO_1557 (O_1557,N_19292,N_19704);
and UO_1558 (O_1558,N_19386,N_19264);
nand UO_1559 (O_1559,N_19345,N_19239);
nand UO_1560 (O_1560,N_19770,N_19594);
nand UO_1561 (O_1561,N_19529,N_19589);
or UO_1562 (O_1562,N_19279,N_19681);
xnor UO_1563 (O_1563,N_19668,N_19989);
and UO_1564 (O_1564,N_19766,N_19973);
nor UO_1565 (O_1565,N_19946,N_19253);
or UO_1566 (O_1566,N_19843,N_19316);
or UO_1567 (O_1567,N_19775,N_19675);
nor UO_1568 (O_1568,N_19658,N_19533);
xnor UO_1569 (O_1569,N_19247,N_19895);
nand UO_1570 (O_1570,N_19526,N_19528);
nor UO_1571 (O_1571,N_19379,N_19213);
xnor UO_1572 (O_1572,N_19531,N_19759);
nand UO_1573 (O_1573,N_19971,N_19862);
or UO_1574 (O_1574,N_19513,N_19879);
nor UO_1575 (O_1575,N_19726,N_19383);
nor UO_1576 (O_1576,N_19852,N_19228);
nor UO_1577 (O_1577,N_19892,N_19915);
and UO_1578 (O_1578,N_19207,N_19404);
nand UO_1579 (O_1579,N_19816,N_19249);
xor UO_1580 (O_1580,N_19458,N_19424);
or UO_1581 (O_1581,N_19753,N_19616);
nand UO_1582 (O_1582,N_19453,N_19756);
nor UO_1583 (O_1583,N_19627,N_19654);
nand UO_1584 (O_1584,N_19978,N_19773);
and UO_1585 (O_1585,N_19826,N_19639);
and UO_1586 (O_1586,N_19648,N_19898);
nand UO_1587 (O_1587,N_19774,N_19895);
nor UO_1588 (O_1588,N_19591,N_19678);
nand UO_1589 (O_1589,N_19852,N_19758);
nor UO_1590 (O_1590,N_19262,N_19346);
nand UO_1591 (O_1591,N_19447,N_19833);
and UO_1592 (O_1592,N_19237,N_19879);
xnor UO_1593 (O_1593,N_19904,N_19866);
nand UO_1594 (O_1594,N_19887,N_19435);
nor UO_1595 (O_1595,N_19529,N_19482);
and UO_1596 (O_1596,N_19260,N_19539);
or UO_1597 (O_1597,N_19860,N_19935);
and UO_1598 (O_1598,N_19821,N_19648);
xor UO_1599 (O_1599,N_19605,N_19482);
nor UO_1600 (O_1600,N_19965,N_19235);
and UO_1601 (O_1601,N_19869,N_19391);
nand UO_1602 (O_1602,N_19961,N_19779);
or UO_1603 (O_1603,N_19704,N_19763);
xnor UO_1604 (O_1604,N_19890,N_19314);
xnor UO_1605 (O_1605,N_19886,N_19389);
xor UO_1606 (O_1606,N_19759,N_19861);
or UO_1607 (O_1607,N_19578,N_19847);
xnor UO_1608 (O_1608,N_19942,N_19246);
nand UO_1609 (O_1609,N_19338,N_19377);
and UO_1610 (O_1610,N_19867,N_19365);
nand UO_1611 (O_1611,N_19485,N_19470);
and UO_1612 (O_1612,N_19555,N_19799);
xor UO_1613 (O_1613,N_19252,N_19336);
and UO_1614 (O_1614,N_19347,N_19733);
xnor UO_1615 (O_1615,N_19677,N_19477);
and UO_1616 (O_1616,N_19269,N_19249);
nand UO_1617 (O_1617,N_19713,N_19815);
or UO_1618 (O_1618,N_19269,N_19737);
nand UO_1619 (O_1619,N_19510,N_19572);
or UO_1620 (O_1620,N_19468,N_19401);
or UO_1621 (O_1621,N_19502,N_19744);
xor UO_1622 (O_1622,N_19778,N_19388);
nand UO_1623 (O_1623,N_19741,N_19981);
or UO_1624 (O_1624,N_19936,N_19507);
nor UO_1625 (O_1625,N_19421,N_19837);
or UO_1626 (O_1626,N_19889,N_19459);
xor UO_1627 (O_1627,N_19442,N_19547);
xor UO_1628 (O_1628,N_19646,N_19797);
xor UO_1629 (O_1629,N_19585,N_19912);
nand UO_1630 (O_1630,N_19487,N_19933);
nor UO_1631 (O_1631,N_19408,N_19788);
and UO_1632 (O_1632,N_19542,N_19834);
or UO_1633 (O_1633,N_19936,N_19337);
xor UO_1634 (O_1634,N_19352,N_19476);
or UO_1635 (O_1635,N_19593,N_19291);
xor UO_1636 (O_1636,N_19543,N_19514);
nand UO_1637 (O_1637,N_19300,N_19794);
nor UO_1638 (O_1638,N_19487,N_19755);
or UO_1639 (O_1639,N_19975,N_19717);
nor UO_1640 (O_1640,N_19543,N_19515);
or UO_1641 (O_1641,N_19358,N_19628);
and UO_1642 (O_1642,N_19400,N_19589);
or UO_1643 (O_1643,N_19612,N_19838);
xor UO_1644 (O_1644,N_19264,N_19929);
and UO_1645 (O_1645,N_19962,N_19525);
nor UO_1646 (O_1646,N_19898,N_19370);
and UO_1647 (O_1647,N_19355,N_19395);
or UO_1648 (O_1648,N_19913,N_19766);
nand UO_1649 (O_1649,N_19690,N_19965);
or UO_1650 (O_1650,N_19833,N_19653);
nor UO_1651 (O_1651,N_19872,N_19576);
or UO_1652 (O_1652,N_19662,N_19956);
nand UO_1653 (O_1653,N_19635,N_19295);
and UO_1654 (O_1654,N_19741,N_19447);
nor UO_1655 (O_1655,N_19666,N_19263);
nand UO_1656 (O_1656,N_19405,N_19872);
nor UO_1657 (O_1657,N_19326,N_19821);
xor UO_1658 (O_1658,N_19794,N_19498);
or UO_1659 (O_1659,N_19934,N_19936);
or UO_1660 (O_1660,N_19930,N_19748);
and UO_1661 (O_1661,N_19476,N_19436);
nor UO_1662 (O_1662,N_19285,N_19821);
nor UO_1663 (O_1663,N_19655,N_19930);
nor UO_1664 (O_1664,N_19211,N_19415);
or UO_1665 (O_1665,N_19206,N_19815);
and UO_1666 (O_1666,N_19521,N_19648);
xnor UO_1667 (O_1667,N_19755,N_19348);
or UO_1668 (O_1668,N_19743,N_19536);
xnor UO_1669 (O_1669,N_19500,N_19344);
nand UO_1670 (O_1670,N_19434,N_19400);
and UO_1671 (O_1671,N_19715,N_19801);
or UO_1672 (O_1672,N_19429,N_19571);
xnor UO_1673 (O_1673,N_19730,N_19874);
nand UO_1674 (O_1674,N_19649,N_19879);
xor UO_1675 (O_1675,N_19410,N_19942);
nor UO_1676 (O_1676,N_19244,N_19741);
and UO_1677 (O_1677,N_19674,N_19993);
xnor UO_1678 (O_1678,N_19988,N_19210);
or UO_1679 (O_1679,N_19393,N_19983);
nor UO_1680 (O_1680,N_19536,N_19930);
nand UO_1681 (O_1681,N_19437,N_19863);
nand UO_1682 (O_1682,N_19340,N_19662);
and UO_1683 (O_1683,N_19404,N_19214);
nand UO_1684 (O_1684,N_19959,N_19807);
or UO_1685 (O_1685,N_19256,N_19620);
or UO_1686 (O_1686,N_19433,N_19697);
and UO_1687 (O_1687,N_19913,N_19874);
nand UO_1688 (O_1688,N_19972,N_19822);
nor UO_1689 (O_1689,N_19422,N_19535);
xnor UO_1690 (O_1690,N_19917,N_19330);
nand UO_1691 (O_1691,N_19761,N_19767);
or UO_1692 (O_1692,N_19270,N_19403);
nor UO_1693 (O_1693,N_19809,N_19543);
nand UO_1694 (O_1694,N_19963,N_19634);
nor UO_1695 (O_1695,N_19235,N_19679);
xnor UO_1696 (O_1696,N_19335,N_19997);
nand UO_1697 (O_1697,N_19503,N_19549);
nand UO_1698 (O_1698,N_19222,N_19231);
and UO_1699 (O_1699,N_19942,N_19270);
xnor UO_1700 (O_1700,N_19386,N_19735);
xnor UO_1701 (O_1701,N_19888,N_19267);
and UO_1702 (O_1702,N_19584,N_19983);
nor UO_1703 (O_1703,N_19866,N_19310);
and UO_1704 (O_1704,N_19751,N_19425);
nor UO_1705 (O_1705,N_19395,N_19465);
nand UO_1706 (O_1706,N_19948,N_19943);
and UO_1707 (O_1707,N_19404,N_19205);
and UO_1708 (O_1708,N_19217,N_19872);
or UO_1709 (O_1709,N_19683,N_19634);
or UO_1710 (O_1710,N_19684,N_19948);
nor UO_1711 (O_1711,N_19849,N_19681);
nand UO_1712 (O_1712,N_19511,N_19472);
nand UO_1713 (O_1713,N_19892,N_19288);
and UO_1714 (O_1714,N_19889,N_19835);
xnor UO_1715 (O_1715,N_19993,N_19729);
nand UO_1716 (O_1716,N_19267,N_19208);
or UO_1717 (O_1717,N_19588,N_19255);
xor UO_1718 (O_1718,N_19258,N_19271);
xnor UO_1719 (O_1719,N_19697,N_19876);
nand UO_1720 (O_1720,N_19532,N_19995);
xnor UO_1721 (O_1721,N_19617,N_19671);
or UO_1722 (O_1722,N_19861,N_19213);
or UO_1723 (O_1723,N_19468,N_19761);
nand UO_1724 (O_1724,N_19397,N_19667);
and UO_1725 (O_1725,N_19389,N_19546);
nor UO_1726 (O_1726,N_19513,N_19496);
xor UO_1727 (O_1727,N_19920,N_19568);
xnor UO_1728 (O_1728,N_19956,N_19941);
or UO_1729 (O_1729,N_19381,N_19611);
xor UO_1730 (O_1730,N_19375,N_19396);
xnor UO_1731 (O_1731,N_19957,N_19766);
nor UO_1732 (O_1732,N_19893,N_19764);
nand UO_1733 (O_1733,N_19296,N_19734);
or UO_1734 (O_1734,N_19971,N_19558);
nand UO_1735 (O_1735,N_19426,N_19816);
and UO_1736 (O_1736,N_19760,N_19777);
and UO_1737 (O_1737,N_19504,N_19712);
nand UO_1738 (O_1738,N_19260,N_19487);
or UO_1739 (O_1739,N_19722,N_19865);
nor UO_1740 (O_1740,N_19218,N_19876);
nand UO_1741 (O_1741,N_19576,N_19453);
xnor UO_1742 (O_1742,N_19456,N_19303);
nand UO_1743 (O_1743,N_19265,N_19944);
nor UO_1744 (O_1744,N_19648,N_19641);
or UO_1745 (O_1745,N_19427,N_19677);
xnor UO_1746 (O_1746,N_19865,N_19785);
or UO_1747 (O_1747,N_19757,N_19378);
xor UO_1748 (O_1748,N_19446,N_19221);
xor UO_1749 (O_1749,N_19269,N_19316);
or UO_1750 (O_1750,N_19378,N_19891);
nand UO_1751 (O_1751,N_19553,N_19534);
or UO_1752 (O_1752,N_19346,N_19893);
nor UO_1753 (O_1753,N_19249,N_19783);
or UO_1754 (O_1754,N_19534,N_19387);
xnor UO_1755 (O_1755,N_19752,N_19744);
nor UO_1756 (O_1756,N_19646,N_19714);
nor UO_1757 (O_1757,N_19987,N_19455);
or UO_1758 (O_1758,N_19825,N_19999);
and UO_1759 (O_1759,N_19955,N_19322);
nor UO_1760 (O_1760,N_19661,N_19946);
nand UO_1761 (O_1761,N_19833,N_19370);
and UO_1762 (O_1762,N_19981,N_19474);
nand UO_1763 (O_1763,N_19441,N_19255);
and UO_1764 (O_1764,N_19769,N_19735);
and UO_1765 (O_1765,N_19559,N_19989);
nand UO_1766 (O_1766,N_19788,N_19980);
or UO_1767 (O_1767,N_19930,N_19401);
and UO_1768 (O_1768,N_19741,N_19515);
xor UO_1769 (O_1769,N_19921,N_19768);
nand UO_1770 (O_1770,N_19496,N_19311);
nor UO_1771 (O_1771,N_19506,N_19514);
or UO_1772 (O_1772,N_19671,N_19702);
and UO_1773 (O_1773,N_19370,N_19885);
nand UO_1774 (O_1774,N_19378,N_19538);
xor UO_1775 (O_1775,N_19599,N_19506);
and UO_1776 (O_1776,N_19904,N_19789);
nand UO_1777 (O_1777,N_19895,N_19752);
and UO_1778 (O_1778,N_19476,N_19406);
nor UO_1779 (O_1779,N_19574,N_19623);
or UO_1780 (O_1780,N_19462,N_19361);
nor UO_1781 (O_1781,N_19822,N_19627);
and UO_1782 (O_1782,N_19436,N_19612);
xor UO_1783 (O_1783,N_19298,N_19767);
nor UO_1784 (O_1784,N_19665,N_19385);
nand UO_1785 (O_1785,N_19369,N_19506);
nor UO_1786 (O_1786,N_19908,N_19757);
nand UO_1787 (O_1787,N_19235,N_19705);
and UO_1788 (O_1788,N_19625,N_19567);
or UO_1789 (O_1789,N_19601,N_19579);
xor UO_1790 (O_1790,N_19567,N_19451);
or UO_1791 (O_1791,N_19461,N_19690);
or UO_1792 (O_1792,N_19374,N_19546);
or UO_1793 (O_1793,N_19433,N_19553);
or UO_1794 (O_1794,N_19202,N_19508);
nand UO_1795 (O_1795,N_19560,N_19522);
nor UO_1796 (O_1796,N_19904,N_19936);
xor UO_1797 (O_1797,N_19746,N_19820);
and UO_1798 (O_1798,N_19709,N_19378);
and UO_1799 (O_1799,N_19633,N_19488);
nand UO_1800 (O_1800,N_19421,N_19565);
nor UO_1801 (O_1801,N_19326,N_19820);
nor UO_1802 (O_1802,N_19641,N_19232);
nor UO_1803 (O_1803,N_19645,N_19384);
and UO_1804 (O_1804,N_19327,N_19896);
nor UO_1805 (O_1805,N_19445,N_19605);
or UO_1806 (O_1806,N_19814,N_19210);
nand UO_1807 (O_1807,N_19314,N_19437);
or UO_1808 (O_1808,N_19955,N_19689);
nor UO_1809 (O_1809,N_19816,N_19834);
xor UO_1810 (O_1810,N_19200,N_19740);
xor UO_1811 (O_1811,N_19200,N_19956);
xnor UO_1812 (O_1812,N_19652,N_19897);
nor UO_1813 (O_1813,N_19723,N_19763);
xor UO_1814 (O_1814,N_19936,N_19517);
nor UO_1815 (O_1815,N_19591,N_19485);
or UO_1816 (O_1816,N_19835,N_19891);
nand UO_1817 (O_1817,N_19454,N_19547);
or UO_1818 (O_1818,N_19686,N_19573);
or UO_1819 (O_1819,N_19581,N_19855);
nor UO_1820 (O_1820,N_19942,N_19735);
or UO_1821 (O_1821,N_19758,N_19738);
and UO_1822 (O_1822,N_19902,N_19218);
nor UO_1823 (O_1823,N_19736,N_19737);
or UO_1824 (O_1824,N_19879,N_19969);
xnor UO_1825 (O_1825,N_19869,N_19503);
nand UO_1826 (O_1826,N_19982,N_19874);
nand UO_1827 (O_1827,N_19422,N_19678);
xnor UO_1828 (O_1828,N_19658,N_19914);
or UO_1829 (O_1829,N_19927,N_19636);
and UO_1830 (O_1830,N_19204,N_19959);
nand UO_1831 (O_1831,N_19794,N_19348);
and UO_1832 (O_1832,N_19470,N_19781);
nand UO_1833 (O_1833,N_19341,N_19440);
or UO_1834 (O_1834,N_19309,N_19567);
nor UO_1835 (O_1835,N_19525,N_19726);
and UO_1836 (O_1836,N_19234,N_19456);
xnor UO_1837 (O_1837,N_19645,N_19618);
or UO_1838 (O_1838,N_19679,N_19642);
or UO_1839 (O_1839,N_19303,N_19309);
and UO_1840 (O_1840,N_19516,N_19909);
nor UO_1841 (O_1841,N_19353,N_19743);
xnor UO_1842 (O_1842,N_19552,N_19824);
and UO_1843 (O_1843,N_19815,N_19616);
or UO_1844 (O_1844,N_19648,N_19324);
xor UO_1845 (O_1845,N_19360,N_19253);
xor UO_1846 (O_1846,N_19925,N_19951);
or UO_1847 (O_1847,N_19461,N_19666);
and UO_1848 (O_1848,N_19503,N_19266);
nor UO_1849 (O_1849,N_19646,N_19975);
nor UO_1850 (O_1850,N_19334,N_19913);
and UO_1851 (O_1851,N_19754,N_19700);
xnor UO_1852 (O_1852,N_19713,N_19492);
nand UO_1853 (O_1853,N_19715,N_19467);
xor UO_1854 (O_1854,N_19978,N_19301);
and UO_1855 (O_1855,N_19680,N_19644);
nand UO_1856 (O_1856,N_19259,N_19470);
or UO_1857 (O_1857,N_19346,N_19221);
nand UO_1858 (O_1858,N_19734,N_19601);
xnor UO_1859 (O_1859,N_19886,N_19600);
or UO_1860 (O_1860,N_19664,N_19445);
xor UO_1861 (O_1861,N_19589,N_19462);
and UO_1862 (O_1862,N_19975,N_19977);
nand UO_1863 (O_1863,N_19224,N_19539);
or UO_1864 (O_1864,N_19642,N_19960);
xnor UO_1865 (O_1865,N_19626,N_19598);
xor UO_1866 (O_1866,N_19494,N_19490);
nor UO_1867 (O_1867,N_19407,N_19329);
nand UO_1868 (O_1868,N_19566,N_19839);
nand UO_1869 (O_1869,N_19803,N_19233);
xnor UO_1870 (O_1870,N_19599,N_19226);
xnor UO_1871 (O_1871,N_19205,N_19270);
nor UO_1872 (O_1872,N_19700,N_19853);
nor UO_1873 (O_1873,N_19797,N_19251);
nor UO_1874 (O_1874,N_19976,N_19892);
and UO_1875 (O_1875,N_19706,N_19258);
and UO_1876 (O_1876,N_19736,N_19345);
xnor UO_1877 (O_1877,N_19426,N_19971);
and UO_1878 (O_1878,N_19262,N_19726);
or UO_1879 (O_1879,N_19786,N_19576);
or UO_1880 (O_1880,N_19486,N_19835);
nor UO_1881 (O_1881,N_19634,N_19749);
or UO_1882 (O_1882,N_19484,N_19365);
nor UO_1883 (O_1883,N_19547,N_19653);
nor UO_1884 (O_1884,N_19847,N_19821);
xnor UO_1885 (O_1885,N_19701,N_19753);
nand UO_1886 (O_1886,N_19426,N_19336);
nand UO_1887 (O_1887,N_19874,N_19280);
nand UO_1888 (O_1888,N_19958,N_19695);
nor UO_1889 (O_1889,N_19984,N_19820);
and UO_1890 (O_1890,N_19875,N_19406);
xor UO_1891 (O_1891,N_19449,N_19656);
nand UO_1892 (O_1892,N_19932,N_19373);
nand UO_1893 (O_1893,N_19675,N_19644);
nand UO_1894 (O_1894,N_19977,N_19342);
nor UO_1895 (O_1895,N_19391,N_19838);
nand UO_1896 (O_1896,N_19926,N_19338);
xor UO_1897 (O_1897,N_19997,N_19530);
xnor UO_1898 (O_1898,N_19310,N_19691);
xor UO_1899 (O_1899,N_19610,N_19430);
nor UO_1900 (O_1900,N_19607,N_19775);
nand UO_1901 (O_1901,N_19510,N_19626);
or UO_1902 (O_1902,N_19612,N_19392);
nand UO_1903 (O_1903,N_19200,N_19477);
or UO_1904 (O_1904,N_19389,N_19709);
nand UO_1905 (O_1905,N_19949,N_19830);
or UO_1906 (O_1906,N_19672,N_19664);
xor UO_1907 (O_1907,N_19814,N_19670);
or UO_1908 (O_1908,N_19374,N_19967);
or UO_1909 (O_1909,N_19403,N_19895);
nand UO_1910 (O_1910,N_19724,N_19767);
nand UO_1911 (O_1911,N_19997,N_19885);
nor UO_1912 (O_1912,N_19766,N_19495);
nor UO_1913 (O_1913,N_19515,N_19324);
and UO_1914 (O_1914,N_19230,N_19758);
and UO_1915 (O_1915,N_19614,N_19909);
nand UO_1916 (O_1916,N_19463,N_19529);
and UO_1917 (O_1917,N_19273,N_19351);
and UO_1918 (O_1918,N_19646,N_19920);
and UO_1919 (O_1919,N_19899,N_19450);
or UO_1920 (O_1920,N_19230,N_19257);
nor UO_1921 (O_1921,N_19538,N_19845);
nand UO_1922 (O_1922,N_19690,N_19431);
xor UO_1923 (O_1923,N_19999,N_19808);
nor UO_1924 (O_1924,N_19773,N_19476);
xnor UO_1925 (O_1925,N_19951,N_19712);
nand UO_1926 (O_1926,N_19807,N_19220);
nor UO_1927 (O_1927,N_19648,N_19210);
xor UO_1928 (O_1928,N_19351,N_19516);
xnor UO_1929 (O_1929,N_19413,N_19530);
xor UO_1930 (O_1930,N_19715,N_19358);
nor UO_1931 (O_1931,N_19644,N_19467);
nand UO_1932 (O_1932,N_19836,N_19586);
or UO_1933 (O_1933,N_19614,N_19225);
xnor UO_1934 (O_1934,N_19701,N_19582);
xnor UO_1935 (O_1935,N_19857,N_19899);
or UO_1936 (O_1936,N_19749,N_19593);
nand UO_1937 (O_1937,N_19424,N_19688);
or UO_1938 (O_1938,N_19739,N_19284);
xnor UO_1939 (O_1939,N_19630,N_19801);
and UO_1940 (O_1940,N_19814,N_19449);
xnor UO_1941 (O_1941,N_19270,N_19409);
and UO_1942 (O_1942,N_19450,N_19317);
nor UO_1943 (O_1943,N_19215,N_19831);
nand UO_1944 (O_1944,N_19501,N_19499);
nor UO_1945 (O_1945,N_19961,N_19300);
or UO_1946 (O_1946,N_19428,N_19654);
nand UO_1947 (O_1947,N_19689,N_19832);
nor UO_1948 (O_1948,N_19978,N_19725);
nand UO_1949 (O_1949,N_19825,N_19353);
and UO_1950 (O_1950,N_19816,N_19896);
or UO_1951 (O_1951,N_19687,N_19382);
nor UO_1952 (O_1952,N_19281,N_19207);
or UO_1953 (O_1953,N_19648,N_19655);
xor UO_1954 (O_1954,N_19328,N_19589);
nor UO_1955 (O_1955,N_19646,N_19309);
xnor UO_1956 (O_1956,N_19496,N_19738);
xor UO_1957 (O_1957,N_19947,N_19372);
nor UO_1958 (O_1958,N_19923,N_19597);
nand UO_1959 (O_1959,N_19395,N_19446);
xor UO_1960 (O_1960,N_19742,N_19292);
or UO_1961 (O_1961,N_19958,N_19956);
nor UO_1962 (O_1962,N_19987,N_19908);
nor UO_1963 (O_1963,N_19707,N_19883);
nor UO_1964 (O_1964,N_19389,N_19440);
and UO_1965 (O_1965,N_19913,N_19603);
nand UO_1966 (O_1966,N_19884,N_19300);
or UO_1967 (O_1967,N_19302,N_19486);
xnor UO_1968 (O_1968,N_19728,N_19560);
xor UO_1969 (O_1969,N_19618,N_19659);
or UO_1970 (O_1970,N_19793,N_19380);
xnor UO_1971 (O_1971,N_19957,N_19504);
nor UO_1972 (O_1972,N_19375,N_19470);
and UO_1973 (O_1973,N_19220,N_19496);
nand UO_1974 (O_1974,N_19954,N_19326);
or UO_1975 (O_1975,N_19986,N_19369);
nand UO_1976 (O_1976,N_19712,N_19663);
nor UO_1977 (O_1977,N_19558,N_19575);
or UO_1978 (O_1978,N_19461,N_19476);
nand UO_1979 (O_1979,N_19459,N_19256);
and UO_1980 (O_1980,N_19225,N_19761);
or UO_1981 (O_1981,N_19239,N_19629);
xnor UO_1982 (O_1982,N_19326,N_19359);
xnor UO_1983 (O_1983,N_19450,N_19337);
nor UO_1984 (O_1984,N_19574,N_19559);
and UO_1985 (O_1985,N_19459,N_19388);
xor UO_1986 (O_1986,N_19554,N_19968);
nand UO_1987 (O_1987,N_19776,N_19855);
nor UO_1988 (O_1988,N_19326,N_19253);
or UO_1989 (O_1989,N_19671,N_19368);
or UO_1990 (O_1990,N_19546,N_19319);
xnor UO_1991 (O_1991,N_19618,N_19903);
and UO_1992 (O_1992,N_19984,N_19737);
xor UO_1993 (O_1993,N_19527,N_19875);
or UO_1994 (O_1994,N_19341,N_19749);
nand UO_1995 (O_1995,N_19946,N_19592);
nand UO_1996 (O_1996,N_19534,N_19371);
and UO_1997 (O_1997,N_19322,N_19846);
nor UO_1998 (O_1998,N_19654,N_19338);
xnor UO_1999 (O_1999,N_19905,N_19346);
nor UO_2000 (O_2000,N_19218,N_19577);
and UO_2001 (O_2001,N_19932,N_19208);
and UO_2002 (O_2002,N_19222,N_19982);
and UO_2003 (O_2003,N_19753,N_19366);
xor UO_2004 (O_2004,N_19592,N_19658);
xnor UO_2005 (O_2005,N_19967,N_19837);
xnor UO_2006 (O_2006,N_19782,N_19846);
or UO_2007 (O_2007,N_19814,N_19232);
and UO_2008 (O_2008,N_19671,N_19681);
and UO_2009 (O_2009,N_19657,N_19402);
or UO_2010 (O_2010,N_19623,N_19280);
or UO_2011 (O_2011,N_19222,N_19253);
nor UO_2012 (O_2012,N_19240,N_19321);
nand UO_2013 (O_2013,N_19620,N_19430);
nand UO_2014 (O_2014,N_19912,N_19935);
xor UO_2015 (O_2015,N_19869,N_19938);
or UO_2016 (O_2016,N_19899,N_19337);
xor UO_2017 (O_2017,N_19345,N_19860);
xor UO_2018 (O_2018,N_19235,N_19553);
nor UO_2019 (O_2019,N_19482,N_19679);
nand UO_2020 (O_2020,N_19714,N_19549);
nand UO_2021 (O_2021,N_19864,N_19543);
or UO_2022 (O_2022,N_19446,N_19378);
nor UO_2023 (O_2023,N_19540,N_19546);
xnor UO_2024 (O_2024,N_19979,N_19781);
xnor UO_2025 (O_2025,N_19907,N_19414);
xnor UO_2026 (O_2026,N_19797,N_19428);
or UO_2027 (O_2027,N_19206,N_19796);
xnor UO_2028 (O_2028,N_19704,N_19558);
nand UO_2029 (O_2029,N_19993,N_19795);
and UO_2030 (O_2030,N_19411,N_19908);
nor UO_2031 (O_2031,N_19895,N_19445);
xnor UO_2032 (O_2032,N_19701,N_19915);
nor UO_2033 (O_2033,N_19981,N_19921);
xor UO_2034 (O_2034,N_19822,N_19690);
nand UO_2035 (O_2035,N_19368,N_19248);
and UO_2036 (O_2036,N_19210,N_19781);
xor UO_2037 (O_2037,N_19656,N_19874);
nand UO_2038 (O_2038,N_19411,N_19358);
xnor UO_2039 (O_2039,N_19202,N_19664);
and UO_2040 (O_2040,N_19544,N_19611);
nor UO_2041 (O_2041,N_19467,N_19314);
xnor UO_2042 (O_2042,N_19294,N_19724);
nand UO_2043 (O_2043,N_19322,N_19463);
nand UO_2044 (O_2044,N_19734,N_19985);
xor UO_2045 (O_2045,N_19437,N_19418);
xor UO_2046 (O_2046,N_19684,N_19740);
nand UO_2047 (O_2047,N_19338,N_19614);
or UO_2048 (O_2048,N_19569,N_19240);
or UO_2049 (O_2049,N_19263,N_19801);
nor UO_2050 (O_2050,N_19415,N_19544);
nand UO_2051 (O_2051,N_19833,N_19538);
or UO_2052 (O_2052,N_19497,N_19343);
nor UO_2053 (O_2053,N_19938,N_19990);
or UO_2054 (O_2054,N_19764,N_19602);
nor UO_2055 (O_2055,N_19225,N_19514);
xor UO_2056 (O_2056,N_19446,N_19501);
xnor UO_2057 (O_2057,N_19548,N_19555);
nand UO_2058 (O_2058,N_19773,N_19578);
nor UO_2059 (O_2059,N_19513,N_19401);
nand UO_2060 (O_2060,N_19441,N_19823);
and UO_2061 (O_2061,N_19755,N_19695);
nand UO_2062 (O_2062,N_19210,N_19540);
xor UO_2063 (O_2063,N_19535,N_19467);
or UO_2064 (O_2064,N_19753,N_19660);
xnor UO_2065 (O_2065,N_19311,N_19209);
xor UO_2066 (O_2066,N_19669,N_19947);
nor UO_2067 (O_2067,N_19913,N_19409);
nand UO_2068 (O_2068,N_19341,N_19386);
nor UO_2069 (O_2069,N_19213,N_19973);
or UO_2070 (O_2070,N_19805,N_19442);
and UO_2071 (O_2071,N_19788,N_19291);
nor UO_2072 (O_2072,N_19425,N_19996);
xor UO_2073 (O_2073,N_19689,N_19927);
nor UO_2074 (O_2074,N_19389,N_19821);
or UO_2075 (O_2075,N_19602,N_19207);
nand UO_2076 (O_2076,N_19600,N_19804);
and UO_2077 (O_2077,N_19269,N_19385);
or UO_2078 (O_2078,N_19658,N_19214);
nor UO_2079 (O_2079,N_19875,N_19599);
nor UO_2080 (O_2080,N_19719,N_19386);
nand UO_2081 (O_2081,N_19888,N_19975);
nand UO_2082 (O_2082,N_19448,N_19248);
nand UO_2083 (O_2083,N_19885,N_19976);
nand UO_2084 (O_2084,N_19937,N_19727);
xnor UO_2085 (O_2085,N_19519,N_19639);
or UO_2086 (O_2086,N_19645,N_19346);
and UO_2087 (O_2087,N_19950,N_19617);
or UO_2088 (O_2088,N_19529,N_19719);
xor UO_2089 (O_2089,N_19844,N_19272);
nor UO_2090 (O_2090,N_19916,N_19236);
and UO_2091 (O_2091,N_19451,N_19499);
xor UO_2092 (O_2092,N_19681,N_19521);
nor UO_2093 (O_2093,N_19733,N_19926);
or UO_2094 (O_2094,N_19706,N_19681);
xor UO_2095 (O_2095,N_19981,N_19789);
and UO_2096 (O_2096,N_19722,N_19595);
nand UO_2097 (O_2097,N_19315,N_19543);
xor UO_2098 (O_2098,N_19515,N_19722);
or UO_2099 (O_2099,N_19839,N_19328);
or UO_2100 (O_2100,N_19369,N_19665);
nor UO_2101 (O_2101,N_19421,N_19857);
nor UO_2102 (O_2102,N_19258,N_19434);
nand UO_2103 (O_2103,N_19640,N_19554);
nand UO_2104 (O_2104,N_19966,N_19509);
xor UO_2105 (O_2105,N_19949,N_19969);
nor UO_2106 (O_2106,N_19256,N_19671);
or UO_2107 (O_2107,N_19465,N_19840);
and UO_2108 (O_2108,N_19238,N_19486);
and UO_2109 (O_2109,N_19574,N_19916);
nor UO_2110 (O_2110,N_19234,N_19290);
nand UO_2111 (O_2111,N_19340,N_19982);
nand UO_2112 (O_2112,N_19408,N_19374);
xnor UO_2113 (O_2113,N_19239,N_19908);
or UO_2114 (O_2114,N_19339,N_19800);
or UO_2115 (O_2115,N_19591,N_19542);
nand UO_2116 (O_2116,N_19712,N_19731);
nand UO_2117 (O_2117,N_19310,N_19213);
nor UO_2118 (O_2118,N_19778,N_19485);
nand UO_2119 (O_2119,N_19568,N_19543);
and UO_2120 (O_2120,N_19831,N_19465);
and UO_2121 (O_2121,N_19401,N_19494);
or UO_2122 (O_2122,N_19773,N_19382);
and UO_2123 (O_2123,N_19662,N_19687);
xnor UO_2124 (O_2124,N_19638,N_19608);
nor UO_2125 (O_2125,N_19417,N_19695);
nor UO_2126 (O_2126,N_19881,N_19306);
nor UO_2127 (O_2127,N_19469,N_19242);
nor UO_2128 (O_2128,N_19278,N_19918);
and UO_2129 (O_2129,N_19713,N_19364);
xor UO_2130 (O_2130,N_19265,N_19537);
nor UO_2131 (O_2131,N_19223,N_19717);
or UO_2132 (O_2132,N_19767,N_19283);
xnor UO_2133 (O_2133,N_19300,N_19425);
nand UO_2134 (O_2134,N_19755,N_19526);
and UO_2135 (O_2135,N_19899,N_19335);
or UO_2136 (O_2136,N_19865,N_19475);
xor UO_2137 (O_2137,N_19244,N_19693);
nand UO_2138 (O_2138,N_19655,N_19582);
nor UO_2139 (O_2139,N_19822,N_19916);
or UO_2140 (O_2140,N_19508,N_19337);
nor UO_2141 (O_2141,N_19414,N_19570);
xor UO_2142 (O_2142,N_19647,N_19922);
xor UO_2143 (O_2143,N_19446,N_19835);
or UO_2144 (O_2144,N_19490,N_19221);
nor UO_2145 (O_2145,N_19897,N_19425);
and UO_2146 (O_2146,N_19269,N_19610);
nor UO_2147 (O_2147,N_19553,N_19908);
xnor UO_2148 (O_2148,N_19991,N_19541);
xor UO_2149 (O_2149,N_19968,N_19800);
or UO_2150 (O_2150,N_19670,N_19995);
or UO_2151 (O_2151,N_19594,N_19235);
nor UO_2152 (O_2152,N_19615,N_19504);
nor UO_2153 (O_2153,N_19305,N_19767);
and UO_2154 (O_2154,N_19450,N_19505);
or UO_2155 (O_2155,N_19226,N_19957);
nor UO_2156 (O_2156,N_19263,N_19338);
xnor UO_2157 (O_2157,N_19572,N_19414);
nand UO_2158 (O_2158,N_19968,N_19542);
nand UO_2159 (O_2159,N_19323,N_19877);
and UO_2160 (O_2160,N_19586,N_19641);
or UO_2161 (O_2161,N_19312,N_19811);
nor UO_2162 (O_2162,N_19475,N_19914);
and UO_2163 (O_2163,N_19904,N_19998);
or UO_2164 (O_2164,N_19643,N_19922);
or UO_2165 (O_2165,N_19857,N_19777);
and UO_2166 (O_2166,N_19658,N_19470);
nand UO_2167 (O_2167,N_19680,N_19447);
xor UO_2168 (O_2168,N_19369,N_19985);
xnor UO_2169 (O_2169,N_19323,N_19913);
nand UO_2170 (O_2170,N_19959,N_19498);
nor UO_2171 (O_2171,N_19583,N_19470);
xnor UO_2172 (O_2172,N_19913,N_19985);
nor UO_2173 (O_2173,N_19458,N_19522);
and UO_2174 (O_2174,N_19947,N_19362);
or UO_2175 (O_2175,N_19766,N_19496);
or UO_2176 (O_2176,N_19632,N_19654);
xnor UO_2177 (O_2177,N_19832,N_19538);
nor UO_2178 (O_2178,N_19344,N_19730);
xnor UO_2179 (O_2179,N_19452,N_19726);
nand UO_2180 (O_2180,N_19678,N_19854);
nor UO_2181 (O_2181,N_19357,N_19603);
and UO_2182 (O_2182,N_19457,N_19575);
nor UO_2183 (O_2183,N_19511,N_19584);
xnor UO_2184 (O_2184,N_19571,N_19491);
nand UO_2185 (O_2185,N_19524,N_19673);
xor UO_2186 (O_2186,N_19705,N_19455);
nor UO_2187 (O_2187,N_19924,N_19314);
or UO_2188 (O_2188,N_19606,N_19381);
nand UO_2189 (O_2189,N_19492,N_19332);
and UO_2190 (O_2190,N_19519,N_19978);
xor UO_2191 (O_2191,N_19472,N_19502);
nand UO_2192 (O_2192,N_19691,N_19698);
and UO_2193 (O_2193,N_19288,N_19966);
nor UO_2194 (O_2194,N_19893,N_19770);
or UO_2195 (O_2195,N_19862,N_19884);
nand UO_2196 (O_2196,N_19243,N_19514);
and UO_2197 (O_2197,N_19929,N_19258);
or UO_2198 (O_2198,N_19676,N_19578);
nand UO_2199 (O_2199,N_19979,N_19453);
nand UO_2200 (O_2200,N_19348,N_19724);
xor UO_2201 (O_2201,N_19859,N_19812);
xor UO_2202 (O_2202,N_19802,N_19780);
nor UO_2203 (O_2203,N_19438,N_19958);
and UO_2204 (O_2204,N_19685,N_19922);
nand UO_2205 (O_2205,N_19926,N_19760);
and UO_2206 (O_2206,N_19267,N_19288);
or UO_2207 (O_2207,N_19610,N_19350);
xor UO_2208 (O_2208,N_19339,N_19887);
nand UO_2209 (O_2209,N_19397,N_19302);
and UO_2210 (O_2210,N_19438,N_19467);
nor UO_2211 (O_2211,N_19260,N_19521);
and UO_2212 (O_2212,N_19274,N_19215);
nand UO_2213 (O_2213,N_19938,N_19804);
or UO_2214 (O_2214,N_19226,N_19613);
and UO_2215 (O_2215,N_19239,N_19886);
xnor UO_2216 (O_2216,N_19961,N_19514);
nand UO_2217 (O_2217,N_19683,N_19614);
and UO_2218 (O_2218,N_19505,N_19322);
nand UO_2219 (O_2219,N_19566,N_19705);
nand UO_2220 (O_2220,N_19897,N_19273);
or UO_2221 (O_2221,N_19890,N_19984);
xnor UO_2222 (O_2222,N_19414,N_19827);
or UO_2223 (O_2223,N_19314,N_19841);
and UO_2224 (O_2224,N_19679,N_19227);
xor UO_2225 (O_2225,N_19239,N_19413);
xor UO_2226 (O_2226,N_19884,N_19282);
xnor UO_2227 (O_2227,N_19219,N_19781);
xnor UO_2228 (O_2228,N_19652,N_19313);
and UO_2229 (O_2229,N_19755,N_19336);
nand UO_2230 (O_2230,N_19933,N_19224);
nand UO_2231 (O_2231,N_19215,N_19802);
and UO_2232 (O_2232,N_19217,N_19383);
nand UO_2233 (O_2233,N_19423,N_19302);
or UO_2234 (O_2234,N_19742,N_19938);
nand UO_2235 (O_2235,N_19528,N_19247);
nor UO_2236 (O_2236,N_19484,N_19565);
and UO_2237 (O_2237,N_19657,N_19443);
nand UO_2238 (O_2238,N_19237,N_19904);
and UO_2239 (O_2239,N_19479,N_19407);
and UO_2240 (O_2240,N_19687,N_19737);
or UO_2241 (O_2241,N_19583,N_19790);
or UO_2242 (O_2242,N_19507,N_19695);
nand UO_2243 (O_2243,N_19342,N_19948);
and UO_2244 (O_2244,N_19953,N_19735);
nand UO_2245 (O_2245,N_19380,N_19779);
nor UO_2246 (O_2246,N_19324,N_19551);
xnor UO_2247 (O_2247,N_19235,N_19777);
nand UO_2248 (O_2248,N_19508,N_19949);
and UO_2249 (O_2249,N_19810,N_19905);
xor UO_2250 (O_2250,N_19651,N_19832);
nand UO_2251 (O_2251,N_19882,N_19968);
or UO_2252 (O_2252,N_19566,N_19642);
or UO_2253 (O_2253,N_19827,N_19402);
and UO_2254 (O_2254,N_19344,N_19333);
and UO_2255 (O_2255,N_19209,N_19367);
nand UO_2256 (O_2256,N_19835,N_19716);
xnor UO_2257 (O_2257,N_19493,N_19222);
nand UO_2258 (O_2258,N_19911,N_19392);
nor UO_2259 (O_2259,N_19688,N_19765);
or UO_2260 (O_2260,N_19675,N_19962);
xnor UO_2261 (O_2261,N_19249,N_19382);
xnor UO_2262 (O_2262,N_19886,N_19858);
or UO_2263 (O_2263,N_19381,N_19436);
xnor UO_2264 (O_2264,N_19626,N_19687);
and UO_2265 (O_2265,N_19243,N_19248);
and UO_2266 (O_2266,N_19762,N_19312);
nor UO_2267 (O_2267,N_19612,N_19855);
or UO_2268 (O_2268,N_19730,N_19411);
nand UO_2269 (O_2269,N_19585,N_19400);
and UO_2270 (O_2270,N_19344,N_19314);
xnor UO_2271 (O_2271,N_19772,N_19207);
nand UO_2272 (O_2272,N_19426,N_19618);
nand UO_2273 (O_2273,N_19956,N_19253);
nand UO_2274 (O_2274,N_19315,N_19928);
and UO_2275 (O_2275,N_19521,N_19289);
xor UO_2276 (O_2276,N_19513,N_19732);
xor UO_2277 (O_2277,N_19953,N_19763);
nor UO_2278 (O_2278,N_19559,N_19516);
or UO_2279 (O_2279,N_19420,N_19722);
nor UO_2280 (O_2280,N_19502,N_19314);
or UO_2281 (O_2281,N_19810,N_19719);
xnor UO_2282 (O_2282,N_19212,N_19828);
and UO_2283 (O_2283,N_19806,N_19617);
nor UO_2284 (O_2284,N_19361,N_19914);
xor UO_2285 (O_2285,N_19851,N_19849);
or UO_2286 (O_2286,N_19654,N_19897);
nand UO_2287 (O_2287,N_19245,N_19526);
xor UO_2288 (O_2288,N_19200,N_19240);
or UO_2289 (O_2289,N_19778,N_19834);
and UO_2290 (O_2290,N_19395,N_19520);
and UO_2291 (O_2291,N_19727,N_19864);
nand UO_2292 (O_2292,N_19960,N_19854);
or UO_2293 (O_2293,N_19721,N_19729);
and UO_2294 (O_2294,N_19773,N_19351);
xor UO_2295 (O_2295,N_19645,N_19350);
nor UO_2296 (O_2296,N_19401,N_19534);
and UO_2297 (O_2297,N_19846,N_19583);
and UO_2298 (O_2298,N_19531,N_19436);
or UO_2299 (O_2299,N_19828,N_19762);
or UO_2300 (O_2300,N_19992,N_19369);
nand UO_2301 (O_2301,N_19629,N_19246);
and UO_2302 (O_2302,N_19834,N_19456);
and UO_2303 (O_2303,N_19921,N_19481);
xnor UO_2304 (O_2304,N_19419,N_19628);
nand UO_2305 (O_2305,N_19832,N_19731);
nor UO_2306 (O_2306,N_19476,N_19687);
or UO_2307 (O_2307,N_19895,N_19661);
or UO_2308 (O_2308,N_19762,N_19510);
and UO_2309 (O_2309,N_19522,N_19403);
nor UO_2310 (O_2310,N_19616,N_19211);
or UO_2311 (O_2311,N_19494,N_19898);
and UO_2312 (O_2312,N_19208,N_19906);
nand UO_2313 (O_2313,N_19581,N_19418);
nand UO_2314 (O_2314,N_19204,N_19847);
nand UO_2315 (O_2315,N_19740,N_19448);
and UO_2316 (O_2316,N_19963,N_19387);
xor UO_2317 (O_2317,N_19629,N_19655);
xnor UO_2318 (O_2318,N_19694,N_19944);
nand UO_2319 (O_2319,N_19854,N_19272);
or UO_2320 (O_2320,N_19717,N_19853);
and UO_2321 (O_2321,N_19645,N_19482);
or UO_2322 (O_2322,N_19861,N_19570);
nor UO_2323 (O_2323,N_19756,N_19773);
or UO_2324 (O_2324,N_19691,N_19296);
xor UO_2325 (O_2325,N_19770,N_19919);
nor UO_2326 (O_2326,N_19687,N_19225);
nor UO_2327 (O_2327,N_19279,N_19563);
xor UO_2328 (O_2328,N_19618,N_19466);
xnor UO_2329 (O_2329,N_19695,N_19619);
and UO_2330 (O_2330,N_19600,N_19329);
nand UO_2331 (O_2331,N_19620,N_19512);
xor UO_2332 (O_2332,N_19411,N_19976);
or UO_2333 (O_2333,N_19357,N_19820);
xnor UO_2334 (O_2334,N_19621,N_19434);
and UO_2335 (O_2335,N_19427,N_19497);
nand UO_2336 (O_2336,N_19403,N_19906);
or UO_2337 (O_2337,N_19278,N_19429);
nand UO_2338 (O_2338,N_19465,N_19599);
nand UO_2339 (O_2339,N_19712,N_19257);
nor UO_2340 (O_2340,N_19315,N_19259);
and UO_2341 (O_2341,N_19666,N_19845);
nor UO_2342 (O_2342,N_19600,N_19840);
or UO_2343 (O_2343,N_19651,N_19756);
nand UO_2344 (O_2344,N_19738,N_19455);
and UO_2345 (O_2345,N_19688,N_19261);
and UO_2346 (O_2346,N_19529,N_19864);
and UO_2347 (O_2347,N_19243,N_19842);
nand UO_2348 (O_2348,N_19746,N_19423);
xor UO_2349 (O_2349,N_19983,N_19242);
or UO_2350 (O_2350,N_19685,N_19352);
and UO_2351 (O_2351,N_19857,N_19320);
xnor UO_2352 (O_2352,N_19756,N_19907);
nand UO_2353 (O_2353,N_19622,N_19931);
and UO_2354 (O_2354,N_19793,N_19654);
nor UO_2355 (O_2355,N_19998,N_19383);
and UO_2356 (O_2356,N_19285,N_19454);
or UO_2357 (O_2357,N_19420,N_19376);
xor UO_2358 (O_2358,N_19416,N_19371);
xnor UO_2359 (O_2359,N_19523,N_19334);
nand UO_2360 (O_2360,N_19870,N_19983);
or UO_2361 (O_2361,N_19262,N_19823);
xnor UO_2362 (O_2362,N_19214,N_19467);
nand UO_2363 (O_2363,N_19587,N_19715);
or UO_2364 (O_2364,N_19511,N_19906);
nand UO_2365 (O_2365,N_19473,N_19315);
or UO_2366 (O_2366,N_19853,N_19763);
xnor UO_2367 (O_2367,N_19479,N_19731);
and UO_2368 (O_2368,N_19491,N_19791);
nand UO_2369 (O_2369,N_19656,N_19595);
or UO_2370 (O_2370,N_19768,N_19706);
nor UO_2371 (O_2371,N_19910,N_19890);
or UO_2372 (O_2372,N_19331,N_19809);
xor UO_2373 (O_2373,N_19813,N_19220);
nand UO_2374 (O_2374,N_19877,N_19836);
and UO_2375 (O_2375,N_19520,N_19289);
nand UO_2376 (O_2376,N_19210,N_19412);
nor UO_2377 (O_2377,N_19955,N_19681);
nand UO_2378 (O_2378,N_19939,N_19847);
xnor UO_2379 (O_2379,N_19215,N_19861);
and UO_2380 (O_2380,N_19324,N_19667);
xor UO_2381 (O_2381,N_19574,N_19513);
xnor UO_2382 (O_2382,N_19281,N_19317);
and UO_2383 (O_2383,N_19521,N_19550);
and UO_2384 (O_2384,N_19867,N_19483);
or UO_2385 (O_2385,N_19352,N_19959);
or UO_2386 (O_2386,N_19265,N_19417);
and UO_2387 (O_2387,N_19914,N_19454);
or UO_2388 (O_2388,N_19631,N_19626);
and UO_2389 (O_2389,N_19239,N_19694);
or UO_2390 (O_2390,N_19980,N_19691);
and UO_2391 (O_2391,N_19708,N_19780);
nor UO_2392 (O_2392,N_19896,N_19577);
nor UO_2393 (O_2393,N_19986,N_19435);
and UO_2394 (O_2394,N_19976,N_19449);
xor UO_2395 (O_2395,N_19243,N_19811);
nand UO_2396 (O_2396,N_19256,N_19548);
and UO_2397 (O_2397,N_19720,N_19972);
xnor UO_2398 (O_2398,N_19732,N_19952);
and UO_2399 (O_2399,N_19906,N_19553);
nor UO_2400 (O_2400,N_19477,N_19301);
nor UO_2401 (O_2401,N_19772,N_19635);
nand UO_2402 (O_2402,N_19603,N_19492);
nor UO_2403 (O_2403,N_19391,N_19987);
and UO_2404 (O_2404,N_19450,N_19693);
nand UO_2405 (O_2405,N_19389,N_19338);
nor UO_2406 (O_2406,N_19980,N_19283);
or UO_2407 (O_2407,N_19859,N_19822);
xnor UO_2408 (O_2408,N_19719,N_19687);
nor UO_2409 (O_2409,N_19469,N_19608);
and UO_2410 (O_2410,N_19242,N_19593);
nand UO_2411 (O_2411,N_19258,N_19311);
and UO_2412 (O_2412,N_19752,N_19718);
or UO_2413 (O_2413,N_19322,N_19465);
nand UO_2414 (O_2414,N_19584,N_19300);
xor UO_2415 (O_2415,N_19993,N_19286);
or UO_2416 (O_2416,N_19982,N_19621);
and UO_2417 (O_2417,N_19548,N_19851);
xnor UO_2418 (O_2418,N_19656,N_19280);
or UO_2419 (O_2419,N_19817,N_19630);
nand UO_2420 (O_2420,N_19907,N_19679);
and UO_2421 (O_2421,N_19368,N_19293);
nor UO_2422 (O_2422,N_19729,N_19463);
nor UO_2423 (O_2423,N_19560,N_19602);
and UO_2424 (O_2424,N_19894,N_19270);
nor UO_2425 (O_2425,N_19655,N_19859);
xor UO_2426 (O_2426,N_19710,N_19846);
nor UO_2427 (O_2427,N_19995,N_19529);
nor UO_2428 (O_2428,N_19646,N_19554);
xor UO_2429 (O_2429,N_19567,N_19802);
or UO_2430 (O_2430,N_19683,N_19509);
xnor UO_2431 (O_2431,N_19205,N_19798);
and UO_2432 (O_2432,N_19775,N_19468);
and UO_2433 (O_2433,N_19935,N_19514);
xor UO_2434 (O_2434,N_19935,N_19588);
nand UO_2435 (O_2435,N_19775,N_19679);
and UO_2436 (O_2436,N_19642,N_19276);
and UO_2437 (O_2437,N_19986,N_19479);
and UO_2438 (O_2438,N_19558,N_19346);
and UO_2439 (O_2439,N_19798,N_19248);
xor UO_2440 (O_2440,N_19382,N_19988);
nor UO_2441 (O_2441,N_19924,N_19221);
and UO_2442 (O_2442,N_19328,N_19498);
nand UO_2443 (O_2443,N_19339,N_19245);
or UO_2444 (O_2444,N_19627,N_19363);
xnor UO_2445 (O_2445,N_19845,N_19780);
nand UO_2446 (O_2446,N_19403,N_19379);
nand UO_2447 (O_2447,N_19848,N_19693);
nor UO_2448 (O_2448,N_19732,N_19466);
and UO_2449 (O_2449,N_19271,N_19812);
nor UO_2450 (O_2450,N_19447,N_19296);
or UO_2451 (O_2451,N_19496,N_19358);
or UO_2452 (O_2452,N_19468,N_19334);
xnor UO_2453 (O_2453,N_19576,N_19246);
and UO_2454 (O_2454,N_19615,N_19953);
nand UO_2455 (O_2455,N_19243,N_19865);
or UO_2456 (O_2456,N_19494,N_19653);
and UO_2457 (O_2457,N_19543,N_19755);
xnor UO_2458 (O_2458,N_19314,N_19499);
nor UO_2459 (O_2459,N_19220,N_19596);
xnor UO_2460 (O_2460,N_19308,N_19793);
xnor UO_2461 (O_2461,N_19735,N_19555);
xor UO_2462 (O_2462,N_19718,N_19644);
xor UO_2463 (O_2463,N_19803,N_19728);
xor UO_2464 (O_2464,N_19241,N_19786);
and UO_2465 (O_2465,N_19557,N_19700);
or UO_2466 (O_2466,N_19866,N_19827);
nand UO_2467 (O_2467,N_19512,N_19234);
or UO_2468 (O_2468,N_19795,N_19725);
or UO_2469 (O_2469,N_19540,N_19218);
or UO_2470 (O_2470,N_19873,N_19562);
xor UO_2471 (O_2471,N_19250,N_19664);
nand UO_2472 (O_2472,N_19767,N_19647);
xnor UO_2473 (O_2473,N_19956,N_19316);
or UO_2474 (O_2474,N_19287,N_19973);
nand UO_2475 (O_2475,N_19560,N_19654);
and UO_2476 (O_2476,N_19968,N_19393);
and UO_2477 (O_2477,N_19808,N_19236);
or UO_2478 (O_2478,N_19986,N_19352);
or UO_2479 (O_2479,N_19760,N_19635);
or UO_2480 (O_2480,N_19314,N_19886);
nand UO_2481 (O_2481,N_19274,N_19444);
nand UO_2482 (O_2482,N_19512,N_19714);
or UO_2483 (O_2483,N_19256,N_19447);
or UO_2484 (O_2484,N_19854,N_19987);
or UO_2485 (O_2485,N_19394,N_19436);
xor UO_2486 (O_2486,N_19339,N_19745);
or UO_2487 (O_2487,N_19567,N_19556);
nand UO_2488 (O_2488,N_19223,N_19273);
or UO_2489 (O_2489,N_19993,N_19405);
nor UO_2490 (O_2490,N_19236,N_19832);
nor UO_2491 (O_2491,N_19988,N_19365);
or UO_2492 (O_2492,N_19594,N_19756);
or UO_2493 (O_2493,N_19773,N_19483);
and UO_2494 (O_2494,N_19241,N_19614);
or UO_2495 (O_2495,N_19704,N_19481);
nor UO_2496 (O_2496,N_19400,N_19692);
nand UO_2497 (O_2497,N_19456,N_19874);
and UO_2498 (O_2498,N_19574,N_19691);
and UO_2499 (O_2499,N_19466,N_19592);
endmodule