module basic_2500_25000_3000_125_levels_10xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999;
xnor U0 (N_0,In_1579,In_734);
or U1 (N_1,In_613,In_2067);
xnor U2 (N_2,In_1212,In_549);
nand U3 (N_3,In_179,In_1498);
nand U4 (N_4,In_1986,In_544);
nand U5 (N_5,In_1588,In_1358);
nor U6 (N_6,In_2112,In_1297);
nor U7 (N_7,In_1442,In_2047);
nand U8 (N_8,In_2341,In_1476);
nand U9 (N_9,In_500,In_2488);
or U10 (N_10,In_749,In_581);
and U11 (N_11,In_986,In_635);
nand U12 (N_12,In_1062,In_1437);
and U13 (N_13,In_125,In_2147);
xor U14 (N_14,In_2043,In_389);
or U15 (N_15,In_2242,In_675);
or U16 (N_16,In_1159,In_1727);
or U17 (N_17,In_1886,In_1866);
xor U18 (N_18,In_601,In_1049);
nor U19 (N_19,In_484,In_832);
and U20 (N_20,In_1783,In_1618);
nor U21 (N_21,In_2044,In_2444);
or U22 (N_22,In_470,In_386);
nand U23 (N_23,In_2118,In_1336);
xor U24 (N_24,In_474,In_283);
and U25 (N_25,In_1822,In_933);
or U26 (N_26,In_981,In_2421);
xor U27 (N_27,In_918,In_1814);
or U28 (N_28,In_1142,In_1348);
xnor U29 (N_29,In_54,In_2066);
nor U30 (N_30,In_1120,In_604);
nor U31 (N_31,In_392,In_203);
xnor U32 (N_32,In_1842,In_62);
xnor U33 (N_33,In_1636,In_2373);
or U34 (N_34,In_547,In_1298);
or U35 (N_35,In_709,In_415);
nor U36 (N_36,In_209,In_2259);
xnor U37 (N_37,In_148,In_871);
and U38 (N_38,In_1207,In_1211);
and U39 (N_39,In_946,In_1792);
nor U40 (N_40,In_2498,In_1058);
nand U41 (N_41,In_331,In_1321);
nand U42 (N_42,In_1518,In_1675);
nand U43 (N_43,In_1703,In_2185);
xor U44 (N_44,In_2055,In_1768);
nor U45 (N_45,In_2134,In_1455);
nor U46 (N_46,In_2022,In_991);
nand U47 (N_47,In_2039,In_2056);
xor U48 (N_48,In_605,In_2273);
nand U49 (N_49,In_575,In_901);
xnor U50 (N_50,In_523,In_497);
and U51 (N_51,In_2361,In_1411);
and U52 (N_52,In_88,In_517);
nand U53 (N_53,In_760,In_2386);
or U54 (N_54,In_446,In_1691);
nor U55 (N_55,In_2179,In_457);
nor U56 (N_56,In_1405,In_2340);
or U57 (N_57,In_896,In_1373);
or U58 (N_58,In_2367,In_1807);
xor U59 (N_59,In_2369,In_127);
nand U60 (N_60,In_2431,In_1831);
or U61 (N_61,In_813,In_132);
xor U62 (N_62,In_65,In_2450);
or U63 (N_63,In_2192,In_1909);
xor U64 (N_64,In_910,In_514);
xnor U65 (N_65,In_182,In_1755);
nor U66 (N_66,In_2019,In_248);
or U67 (N_67,In_2283,In_1135);
or U68 (N_68,In_1491,In_2114);
nand U69 (N_69,In_984,In_5);
nor U70 (N_70,In_473,In_453);
xor U71 (N_71,In_365,In_2336);
or U72 (N_72,In_465,In_1493);
nand U73 (N_73,In_2175,In_258);
xnor U74 (N_74,In_1994,In_1045);
and U75 (N_75,In_1610,In_1585);
and U76 (N_76,In_2327,In_1464);
and U77 (N_77,In_414,In_2364);
nor U78 (N_78,In_1533,In_2424);
and U79 (N_79,In_1996,In_1984);
and U80 (N_80,In_451,In_1262);
or U81 (N_81,In_724,In_2487);
and U82 (N_82,In_752,In_1126);
xor U83 (N_83,In_1527,In_2042);
xor U84 (N_84,In_1429,In_2462);
xnor U85 (N_85,In_1393,In_486);
and U86 (N_86,In_2158,In_1540);
and U87 (N_87,In_740,In_2209);
nand U88 (N_88,In_1470,In_1739);
xor U89 (N_89,In_876,In_922);
or U90 (N_90,In_704,In_1421);
nor U91 (N_91,In_1927,In_1754);
and U92 (N_92,In_2142,In_1323);
xnor U93 (N_93,In_134,In_1704);
xor U94 (N_94,In_1760,In_1102);
nor U95 (N_95,In_1095,In_46);
nor U96 (N_96,In_1530,In_2272);
nand U97 (N_97,In_1804,In_758);
nor U98 (N_98,In_512,In_313);
nor U99 (N_99,In_2306,In_2086);
nor U100 (N_100,In_771,In_788);
nor U101 (N_101,In_767,In_585);
nor U102 (N_102,In_2267,In_250);
nand U103 (N_103,In_1271,In_2049);
nand U104 (N_104,In_1177,In_1320);
xnor U105 (N_105,In_1114,In_492);
or U106 (N_106,In_1017,In_1073);
nand U107 (N_107,In_176,In_1427);
or U108 (N_108,In_1634,In_228);
nor U109 (N_109,In_1712,In_94);
or U110 (N_110,In_1976,In_1823);
nand U111 (N_111,In_1125,In_235);
and U112 (N_112,In_1274,In_2024);
or U113 (N_113,In_2346,In_2411);
or U114 (N_114,In_137,In_1454);
xor U115 (N_115,In_2208,In_1709);
xnor U116 (N_116,In_270,In_1035);
nor U117 (N_117,In_2429,In_1410);
nor U118 (N_118,In_1957,In_421);
xnor U119 (N_119,In_2268,In_1884);
or U120 (N_120,In_582,In_2366);
or U121 (N_121,In_269,In_849);
xnor U122 (N_122,In_1631,In_2157);
nor U123 (N_123,In_1197,In_669);
xnor U124 (N_124,In_1632,In_2223);
nand U125 (N_125,In_2081,In_2345);
xor U126 (N_126,In_2352,In_1622);
nand U127 (N_127,In_1677,In_1985);
nor U128 (N_128,In_703,In_1332);
or U129 (N_129,In_2439,In_271);
or U130 (N_130,In_2491,In_698);
nand U131 (N_131,In_1728,In_1507);
nor U132 (N_132,In_1742,In_1970);
and U133 (N_133,In_1901,In_923);
xnor U134 (N_134,In_959,In_1551);
and U135 (N_135,In_1749,In_2377);
nor U136 (N_136,In_485,In_455);
nand U137 (N_137,In_681,In_2417);
nand U138 (N_138,In_1987,In_561);
and U139 (N_139,In_318,In_304);
xnor U140 (N_140,In_1419,In_2382);
or U141 (N_141,In_815,In_2383);
or U142 (N_142,In_1591,In_354);
nor U143 (N_143,In_744,In_244);
and U144 (N_144,In_2122,In_1828);
xnor U145 (N_145,In_1565,In_95);
or U146 (N_146,In_563,In_2412);
nor U147 (N_147,In_1714,In_2213);
xor U148 (N_148,In_216,In_1925);
and U149 (N_149,In_567,In_74);
nand U150 (N_150,In_2057,In_818);
or U151 (N_151,In_1771,In_489);
xnor U152 (N_152,In_35,In_1553);
or U153 (N_153,In_1524,In_1911);
xnor U154 (N_154,In_1782,In_2160);
and U155 (N_155,In_2410,In_2245);
or U156 (N_156,In_1293,In_1449);
nor U157 (N_157,In_2129,In_2082);
xor U158 (N_158,In_381,In_1645);
nand U159 (N_159,In_2091,In_1010);
nand U160 (N_160,In_1791,In_1388);
xnor U161 (N_161,In_1450,In_1821);
or U162 (N_162,In_1357,In_1397);
xnor U163 (N_163,In_1295,In_1174);
or U164 (N_164,In_2230,In_1029);
or U165 (N_165,In_762,In_12);
xor U166 (N_166,In_2198,In_1600);
and U167 (N_167,In_1510,In_653);
xor U168 (N_168,In_1309,In_210);
or U169 (N_169,In_2416,In_1700);
nand U170 (N_170,In_506,In_2319);
xor U171 (N_171,In_401,In_663);
nand U172 (N_172,In_129,In_593);
or U173 (N_173,In_784,In_2479);
and U174 (N_174,In_1906,In_1558);
nor U175 (N_175,In_305,In_469);
or U176 (N_176,In_797,In_89);
nand U177 (N_177,In_1269,In_776);
xnor U178 (N_178,In_2187,In_962);
nand U179 (N_179,In_443,In_2497);
nor U180 (N_180,In_260,In_1952);
or U181 (N_181,In_861,In_1576);
nor U182 (N_182,In_1939,In_2362);
xor U183 (N_183,In_1857,In_2282);
nor U184 (N_184,In_388,In_495);
or U185 (N_185,In_33,In_1148);
nand U186 (N_186,In_1578,In_2275);
nor U187 (N_187,In_1686,In_2342);
nor U188 (N_188,In_532,In_149);
and U189 (N_189,In_2100,In_1627);
xnor U190 (N_190,In_1960,In_292);
xnor U191 (N_191,In_2298,In_348);
or U192 (N_192,In_2217,In_1151);
nand U193 (N_193,In_434,In_2418);
and U194 (N_194,In_294,In_513);
or U195 (N_195,In_1398,In_2257);
or U196 (N_196,In_1376,In_422);
nand U197 (N_197,In_2481,In_721);
and U198 (N_198,In_2222,In_1228);
and U199 (N_199,In_580,In_2096);
and U200 (N_200,In_1333,N_13);
xor U201 (N_201,In_1587,In_1878);
xor U202 (N_202,In_814,In_2372);
nor U203 (N_203,In_1995,In_1733);
or U204 (N_204,In_183,In_1575);
or U205 (N_205,In_1453,In_1961);
nand U206 (N_206,In_130,In_10);
nand U207 (N_207,In_369,N_193);
or U208 (N_208,In_878,In_915);
or U209 (N_209,In_1949,In_1637);
nor U210 (N_210,In_741,In_2263);
nor U211 (N_211,In_620,In_2476);
or U212 (N_212,N_88,In_1719);
and U213 (N_213,In_2265,N_131);
xnor U214 (N_214,In_1290,In_2406);
and U215 (N_215,In_649,In_1758);
and U216 (N_216,In_1299,In_448);
nor U217 (N_217,In_110,N_55);
and U218 (N_218,In_1690,In_131);
and U219 (N_219,N_126,In_2105);
or U220 (N_220,In_1832,In_1799);
nand U221 (N_221,In_1276,In_403);
and U222 (N_222,In_2464,In_521);
nand U223 (N_223,In_1077,In_1094);
or U224 (N_224,In_1140,In_1966);
nand U225 (N_225,In_2323,In_1115);
xnor U226 (N_226,In_116,In_1698);
or U227 (N_227,In_53,In_1054);
and U228 (N_228,In_2428,In_763);
and U229 (N_229,In_1283,In_548);
xnor U230 (N_230,In_646,In_808);
nand U231 (N_231,In_945,In_79);
or U232 (N_232,In_976,In_126);
xnor U233 (N_233,In_967,In_1999);
nand U234 (N_234,In_219,In_2374);
and U235 (N_235,In_201,In_1541);
xor U236 (N_236,In_2127,In_1221);
nand U237 (N_237,In_2068,In_1347);
and U238 (N_238,In_1097,In_124);
and U239 (N_239,In_2101,In_2280);
or U240 (N_240,In_2204,In_2457);
nor U241 (N_241,In_786,In_217);
and U242 (N_242,In_2161,In_1013);
and U243 (N_243,In_1412,In_987);
xnor U244 (N_244,N_48,In_112);
xor U245 (N_245,In_1201,In_977);
or U246 (N_246,In_1294,In_2008);
xnor U247 (N_247,N_97,In_425);
or U248 (N_248,In_1292,In_667);
nor U249 (N_249,In_1403,In_2201);
nor U250 (N_250,In_1552,In_2284);
and U251 (N_251,In_1803,In_1231);
nand U252 (N_252,In_2391,N_127);
and U253 (N_253,In_2207,In_2305);
nand U254 (N_254,In_1764,In_1688);
and U255 (N_255,In_822,In_1511);
nand U256 (N_256,N_194,In_845);
or U257 (N_257,In_769,In_1667);
xor U258 (N_258,In_2063,In_2474);
or U259 (N_259,In_690,In_2069);
nor U260 (N_260,In_2005,In_2136);
and U261 (N_261,In_895,In_693);
or U262 (N_262,In_2485,In_2388);
and U263 (N_263,In_545,In_1338);
nand U264 (N_264,In_1781,In_412);
nor U265 (N_265,In_983,In_1351);
nor U266 (N_266,In_1545,In_2451);
xor U267 (N_267,In_207,In_793);
and U268 (N_268,In_276,In_1001);
and U269 (N_269,In_1875,In_1430);
and U270 (N_270,In_1273,In_799);
or U271 (N_271,In_155,N_24);
nand U272 (N_272,In_834,In_995);
nor U273 (N_273,N_70,N_154);
or U274 (N_274,In_2227,In_1215);
xnor U275 (N_275,In_1773,N_68);
nand U276 (N_276,In_2343,N_51);
nand U277 (N_277,In_2041,N_77);
nor U278 (N_278,In_138,In_2235);
nor U279 (N_279,In_522,In_1989);
nand U280 (N_280,In_829,In_1128);
nor U281 (N_281,In_1752,In_1117);
and U282 (N_282,In_1008,In_2107);
nand U283 (N_283,In_1007,In_2455);
xnor U284 (N_284,In_2050,N_91);
or U285 (N_285,In_483,In_1586);
xor U286 (N_286,In_1404,In_1639);
nor U287 (N_287,In_2435,In_2409);
nor U288 (N_288,In_1457,In_1055);
or U289 (N_289,In_1383,In_597);
xor U290 (N_290,In_2301,In_1152);
nand U291 (N_291,In_782,In_877);
and U292 (N_292,In_2300,In_1103);
nand U293 (N_293,In_2381,In_1892);
nand U294 (N_294,In_889,In_2116);
and U295 (N_295,In_916,In_1560);
and U296 (N_296,N_22,N_112);
nor U297 (N_297,In_2243,N_195);
nand U298 (N_298,In_2133,In_2335);
or U299 (N_299,In_687,In_1078);
xor U300 (N_300,N_17,In_2200);
xor U301 (N_301,In_2103,In_9);
nor U302 (N_302,In_11,N_102);
nor U303 (N_303,In_1057,N_164);
or U304 (N_304,In_1063,In_2333);
or U305 (N_305,In_1475,In_1890);
nand U306 (N_306,In_1034,In_333);
nor U307 (N_307,In_925,N_168);
nand U308 (N_308,In_2074,In_1669);
and U309 (N_309,In_316,In_196);
xnor U310 (N_310,In_2325,In_1721);
nor U311 (N_311,In_533,In_156);
and U312 (N_312,In_1039,In_2309);
or U313 (N_313,In_2385,In_1267);
nor U314 (N_314,In_2430,N_34);
nand U315 (N_315,In_1959,In_1325);
nor U316 (N_316,In_1248,In_1047);
and U317 (N_317,In_1829,In_800);
and U318 (N_318,In_163,In_97);
nor U319 (N_319,In_1439,N_74);
or U320 (N_320,In_2033,In_325);
nand U321 (N_321,N_121,In_1656);
or U322 (N_322,In_1362,In_2226);
nand U323 (N_323,In_1431,In_1443);
or U324 (N_324,In_1064,In_1529);
and U325 (N_325,In_57,In_2031);
xnor U326 (N_326,In_1873,In_1238);
nor U327 (N_327,In_1834,In_1793);
nand U328 (N_328,In_764,In_1731);
and U329 (N_329,In_2083,N_109);
nand U330 (N_330,In_144,In_1253);
and U331 (N_331,In_2270,In_543);
xor U332 (N_332,In_1982,N_113);
nor U333 (N_333,In_1659,In_1184);
and U334 (N_334,In_1127,In_2210);
nor U335 (N_335,In_24,In_98);
xnor U336 (N_336,In_1106,In_718);
xnor U337 (N_337,In_321,N_31);
nor U338 (N_338,In_1573,In_900);
nand U339 (N_339,In_1921,In_1256);
xnor U340 (N_340,In_2166,In_2153);
or U341 (N_341,In_402,In_2130);
and U342 (N_342,In_43,In_1196);
nand U343 (N_343,In_1820,In_802);
nand U344 (N_344,In_1434,In_323);
xnor U345 (N_345,In_1655,In_790);
or U346 (N_346,In_2131,In_266);
or U347 (N_347,In_873,N_186);
and U348 (N_348,In_2493,In_1706);
xnor U349 (N_349,N_110,In_45);
xnor U350 (N_350,In_1124,In_1282);
nor U351 (N_351,In_2348,In_1798);
nor U352 (N_352,In_754,In_1022);
nor U353 (N_353,In_1914,In_328);
nor U354 (N_354,In_1843,In_751);
and U355 (N_355,N_160,In_314);
and U356 (N_356,N_108,In_2018);
and U357 (N_357,In_570,In_1896);
nand U358 (N_358,In_851,In_1156);
and U359 (N_359,In_1048,In_838);
or U360 (N_360,In_76,In_101);
xor U361 (N_361,In_122,In_1602);
or U362 (N_362,In_32,N_123);
or U363 (N_363,In_937,In_939);
xor U364 (N_364,In_2357,In_1665);
nor U365 (N_365,In_344,In_1327);
xnor U366 (N_366,In_816,N_72);
and U367 (N_367,In_2135,In_2326);
nand U368 (N_368,In_75,In_1436);
nor U369 (N_369,In_966,In_633);
xnor U370 (N_370,In_1004,In_730);
or U371 (N_371,In_1683,N_189);
nor U372 (N_372,In_1301,In_376);
xnor U373 (N_373,In_2013,In_1318);
and U374 (N_374,In_1460,In_1104);
nor U375 (N_375,In_963,In_332);
or U376 (N_376,In_796,In_441);
nand U377 (N_377,In_39,In_831);
nand U378 (N_378,In_774,In_2237);
nor U379 (N_379,In_2191,In_2070);
xnor U380 (N_380,In_424,In_993);
or U381 (N_381,In_285,In_622);
xor U382 (N_382,In_657,In_2007);
nand U383 (N_383,In_380,In_2218);
nand U384 (N_384,In_1974,In_1465);
and U385 (N_385,In_1462,In_843);
or U386 (N_386,In_2304,In_1413);
xnor U387 (N_387,In_1233,In_2111);
nand U388 (N_388,In_1990,In_980);
xor U389 (N_389,In_145,In_639);
or U390 (N_390,In_1471,In_1812);
nor U391 (N_391,In_827,In_650);
nand U392 (N_392,In_172,In_1879);
nand U393 (N_393,In_594,In_1713);
and U394 (N_394,In_1644,In_801);
or U395 (N_395,In_1037,In_2020);
xnor U396 (N_396,In_1509,In_2197);
nand U397 (N_397,In_919,In_1801);
nor U398 (N_398,In_1963,In_290);
xor U399 (N_399,In_969,In_1474);
or U400 (N_400,In_1192,In_595);
and U401 (N_401,N_165,In_111);
nand U402 (N_402,In_1105,In_118);
or U403 (N_403,In_1784,N_285);
nor U404 (N_404,In_282,In_275);
xnor U405 (N_405,In_2490,In_1361);
nor U406 (N_406,In_884,In_1147);
nand U407 (N_407,In_1111,N_261);
and U408 (N_408,N_101,In_1222);
xor U409 (N_409,In_159,N_84);
and U410 (N_410,In_2169,In_944);
and U411 (N_411,In_1936,In_903);
nand U412 (N_412,N_33,N_47);
or U413 (N_413,In_2225,In_1672);
or U414 (N_414,In_972,In_1891);
and U415 (N_415,In_2466,In_638);
or U416 (N_416,In_281,In_340);
nor U417 (N_417,In_197,In_885);
nor U418 (N_418,In_1854,In_1825);
xor U419 (N_419,In_2151,In_1694);
xnor U420 (N_420,In_1658,In_181);
or U421 (N_421,In_2496,N_140);
or U422 (N_422,In_865,N_49);
and U423 (N_423,N_294,In_565);
xnor U424 (N_424,In_229,In_631);
nor U425 (N_425,In_554,In_1945);
or U426 (N_426,N_50,In_572);
xnor U427 (N_427,N_202,In_586);
or U428 (N_428,In_1108,In_353);
xnor U429 (N_429,In_1236,In_278);
xor U430 (N_430,In_1550,N_387);
nand U431 (N_431,In_1086,N_252);
nor U432 (N_432,In_1015,In_326);
or U433 (N_433,In_2094,In_187);
and U434 (N_434,In_34,In_558);
or U435 (N_435,In_2017,In_2137);
or U436 (N_436,In_614,In_864);
and U437 (N_437,In_1613,In_1905);
xnor U438 (N_438,In_1840,In_1993);
nor U439 (N_439,In_2150,In_102);
or U440 (N_440,In_1753,N_146);
or U441 (N_441,In_367,In_1286);
nand U442 (N_442,In_2363,In_1630);
or U443 (N_443,In_2486,In_224);
xnor U444 (N_444,In_2454,In_1467);
nand U445 (N_445,In_1387,N_214);
nor U446 (N_446,N_159,In_783);
nand U447 (N_447,In_2475,In_1679);
and U448 (N_448,In_1696,N_283);
and U449 (N_449,In_1305,In_1423);
xor U450 (N_450,In_91,In_920);
and U451 (N_451,N_0,In_1701);
or U452 (N_452,In_2311,In_1946);
nor U453 (N_453,In_1191,In_2171);
nor U454 (N_454,In_1466,N_342);
xnor U455 (N_455,N_95,In_629);
nor U456 (N_456,In_175,In_1265);
and U457 (N_457,In_58,In_1445);
or U458 (N_458,In_329,In_259);
nor U459 (N_459,In_1975,In_1572);
xnor U460 (N_460,In_1024,In_1189);
and U461 (N_461,In_180,In_2419);
xor U462 (N_462,In_230,In_68);
xnor U463 (N_463,In_2184,In_2467);
xor U464 (N_464,In_311,In_538);
or U465 (N_465,In_1209,In_2249);
nand U466 (N_466,N_248,In_898);
and U467 (N_467,In_694,In_378);
or U468 (N_468,In_1900,In_550);
xor U469 (N_469,N_215,In_2437);
xor U470 (N_470,In_630,In_1153);
xor U471 (N_471,N_208,N_171);
nand U472 (N_472,In_1935,In_1075);
and U473 (N_473,In_2426,In_1514);
and U474 (N_474,In_539,In_3);
and U475 (N_475,In_2089,In_569);
nor U476 (N_476,In_1761,In_296);
nor U477 (N_477,In_1000,In_1146);
and U478 (N_478,In_277,In_1623);
or U479 (N_479,N_312,N_311);
nand U480 (N_480,In_1870,In_645);
or U481 (N_481,N_309,In_234);
nand U482 (N_482,In_1796,In_1848);
nand U483 (N_483,In_1885,In_2167);
or U484 (N_484,In_706,In_936);
and U485 (N_485,In_1463,In_2165);
nand U486 (N_486,In_2046,In_464);
nor U487 (N_487,In_860,In_850);
nand U488 (N_488,In_1894,In_2220);
nor U489 (N_489,N_398,In_1160);
xnor U490 (N_490,In_1469,In_307);
nor U491 (N_491,In_371,In_1328);
and U492 (N_492,In_472,In_1523);
nand U493 (N_493,In_1635,In_578);
xnor U494 (N_494,N_185,In_1847);
or U495 (N_495,N_346,N_19);
nand U496 (N_496,In_1084,In_239);
or U497 (N_497,In_2211,In_1036);
nand U498 (N_498,N_217,N_173);
nand U499 (N_499,In_295,In_1252);
or U500 (N_500,In_454,N_330);
nand U501 (N_501,N_369,In_1458);
nor U502 (N_502,In_1609,In_691);
nor U503 (N_503,In_1889,In_1554);
nor U504 (N_504,In_2,In_2312);
nand U505 (N_505,In_14,N_59);
and U506 (N_506,In_1426,N_397);
nor U507 (N_507,In_2287,N_359);
and U508 (N_508,In_2189,In_1289);
or U509 (N_509,In_1389,In_2308);
and U510 (N_510,In_1194,In_2278);
nor U511 (N_511,In_1777,In_1304);
xor U512 (N_512,N_44,In_1206);
nand U513 (N_513,In_1931,In_1416);
or U514 (N_514,In_358,In_1488);
xnor U515 (N_515,N_75,In_71);
nor U516 (N_516,In_988,In_1947);
nand U517 (N_517,In_950,In_1313);
or U518 (N_518,In_510,In_1943);
nand U519 (N_519,In_1499,In_682);
nor U520 (N_520,In_1090,N_343);
nor U521 (N_521,In_1649,In_1296);
nand U522 (N_522,In_1089,In_1490);
and U523 (N_523,N_341,In_1446);
or U524 (N_524,N_273,In_2307);
nand U525 (N_525,In_1391,In_1992);
nand U526 (N_526,In_2036,In_1687);
and U527 (N_527,In_1249,In_1693);
xor U528 (N_528,In_2229,N_203);
nand U529 (N_529,In_2396,In_1537);
and U530 (N_530,In_642,In_735);
and U531 (N_531,In_249,In_1131);
xnor U532 (N_532,In_2252,In_1281);
nand U533 (N_533,In_73,In_6);
nand U534 (N_534,In_2138,N_268);
and U535 (N_535,In_2459,In_1213);
nand U536 (N_536,In_165,In_2276);
or U537 (N_537,In_1202,In_1258);
xnor U538 (N_538,In_1853,In_1406);
and U539 (N_539,In_842,In_610);
nand U540 (N_540,In_753,N_30);
nand U541 (N_541,In_1882,In_1264);
and U542 (N_542,N_265,In_36);
xnor U543 (N_543,In_1079,N_223);
or U544 (N_544,N_132,N_289);
xor U545 (N_545,In_427,In_2052);
nor U546 (N_546,In_2215,In_1860);
or U547 (N_547,In_688,In_406);
xnor U548 (N_548,In_2318,In_770);
nor U549 (N_549,In_356,In_70);
and U550 (N_550,In_493,In_847);
or U551 (N_551,In_509,In_1122);
xnor U552 (N_552,N_111,In_372);
xnor U553 (N_553,In_1042,N_32);
xor U554 (N_554,In_504,In_1478);
and U555 (N_555,In_1651,In_785);
or U556 (N_556,In_1392,In_2291);
nand U557 (N_557,N_46,In_1762);
xor U558 (N_558,In_2427,In_634);
nand U559 (N_559,N_155,In_1692);
nand U560 (N_560,In_820,In_869);
nor U561 (N_561,In_37,N_38);
nor U562 (N_562,In_902,In_1018);
xor U563 (N_563,In_2080,In_1893);
nor U564 (N_564,In_2277,N_178);
xor U565 (N_565,In_80,In_1951);
or U566 (N_566,In_1582,N_384);
or U567 (N_567,In_826,In_1592);
or U568 (N_568,In_1897,In_1339);
nor U569 (N_569,In_719,N_170);
and U570 (N_570,N_209,In_2402);
and U571 (N_571,In_2389,In_1536);
xor U572 (N_572,In_2104,N_82);
nor U573 (N_573,In_750,In_2285);
nand U574 (N_574,N_180,In_828);
xor U575 (N_575,In_198,In_1756);
or U576 (N_576,In_1208,In_1750);
xnor U577 (N_577,N_96,In_1616);
nor U578 (N_578,In_20,N_291);
xor U579 (N_579,In_623,In_576);
nand U580 (N_580,In_2026,In_7);
nor U581 (N_581,In_1051,In_83);
or U582 (N_582,N_381,In_1808);
and U583 (N_583,In_245,In_1978);
nand U584 (N_584,In_1626,In_16);
or U585 (N_585,In_2356,N_11);
xor U586 (N_586,In_1779,In_1020);
nand U587 (N_587,In_930,In_480);
and U588 (N_588,In_1528,In_564);
nor U589 (N_589,In_1797,In_1118);
nor U590 (N_590,In_481,In_674);
and U591 (N_591,N_63,In_117);
or U592 (N_592,In_1353,In_913);
xor U593 (N_593,In_893,In_120);
xnor U594 (N_594,In_2120,N_364);
or U595 (N_595,In_1259,N_357);
or U596 (N_596,N_259,In_947);
xnor U597 (N_597,N_191,In_1707);
nor U598 (N_598,N_175,N_237);
or U599 (N_599,In_2401,In_1019);
xnor U600 (N_600,In_419,In_1827);
or U601 (N_601,In_717,In_475);
xnor U602 (N_602,In_1210,In_1928);
xnor U603 (N_603,In_738,In_1083);
or U604 (N_604,In_1272,In_2269);
nor U605 (N_605,In_2274,In_72);
nor U606 (N_606,N_505,In_1377);
nor U607 (N_607,N_457,In_1132);
or U608 (N_608,In_1830,In_1076);
and U609 (N_609,In_1942,In_2365);
nand U610 (N_610,N_362,N_372);
and U611 (N_611,In_315,In_1517);
nor U612 (N_612,In_343,In_1386);
and U613 (N_613,N_409,In_1604);
nor U614 (N_614,N_527,In_1926);
xor U615 (N_615,N_349,In_1907);
or U616 (N_616,In_420,In_743);
or U617 (N_617,In_833,In_2338);
and U618 (N_618,In_1133,In_1137);
nor U619 (N_619,N_272,In_1718);
or U620 (N_620,In_789,In_1861);
nand U621 (N_621,In_2489,In_795);
xnor U622 (N_622,N_424,In_1326);
xnor U623 (N_623,In_713,N_469);
or U624 (N_624,In_2214,In_1883);
xnor U625 (N_625,In_218,In_152);
and U626 (N_626,In_2290,In_695);
and U627 (N_627,N_141,In_2358);
nand U628 (N_628,In_810,In_773);
and U629 (N_629,N_506,N_495);
and U630 (N_630,In_1171,N_533);
or U631 (N_631,In_1819,In_1717);
or U632 (N_632,In_1395,In_445);
nor U633 (N_633,In_195,In_1324);
nand U634 (N_634,In_1868,In_609);
nand U635 (N_635,In_113,In_1408);
nand U636 (N_636,N_43,In_212);
xnor U637 (N_637,N_485,In_899);
xnor U638 (N_638,N_324,N_264);
nand U639 (N_639,In_1331,In_943);
nand U640 (N_640,In_625,In_659);
and U641 (N_641,In_685,In_2027);
nand U642 (N_642,In_2021,In_2087);
and U643 (N_643,N_543,In_607);
and U644 (N_644,N_148,N_348);
nand U645 (N_645,In_2288,N_496);
and U646 (N_646,In_1620,N_56);
xnor U647 (N_647,In_2075,N_256);
nand U648 (N_648,In_732,In_647);
or U649 (N_649,In_2144,In_303);
or U650 (N_650,N_318,In_1031);
and U651 (N_651,In_2143,N_340);
xor U652 (N_652,In_1790,N_487);
or U653 (N_653,In_1337,In_542);
or U654 (N_654,In_632,N_572);
xnor U655 (N_655,N_100,In_496);
nand U656 (N_656,In_100,In_1016);
or U657 (N_657,In_2076,In_1765);
and U658 (N_658,In_2244,In_1163);
xnor U659 (N_659,In_222,In_596);
nor U660 (N_660,In_1162,In_2231);
or U661 (N_661,In_55,In_1730);
xor U662 (N_662,N_515,In_192);
nor U663 (N_663,In_2190,In_1082);
xor U664 (N_664,In_1695,In_541);
or U665 (N_665,N_516,In_2403);
nand U666 (N_666,N_422,N_29);
nor U667 (N_667,In_1307,In_1065);
xnor U668 (N_668,In_2010,N_275);
nor U669 (N_669,In_505,N_197);
or U670 (N_670,N_1,In_2332);
and U671 (N_671,In_2359,N_458);
xnor U672 (N_672,In_904,In_206);
nand U673 (N_673,N_7,N_408);
nor U674 (N_674,N_472,In_256);
nand U675 (N_675,In_433,In_1811);
and U676 (N_676,In_608,N_228);
and U677 (N_677,In_2492,N_588);
nand U678 (N_678,N_128,In_317);
or U679 (N_679,N_89,In_2177);
xor U680 (N_680,In_52,In_1134);
and U681 (N_681,N_69,In_194);
nand U682 (N_682,N_388,In_2482);
nor U683 (N_683,N_517,In_44);
nand U684 (N_684,In_664,N_481);
xor U685 (N_685,In_2194,In_1504);
nand U686 (N_686,In_2392,In_77);
nor U687 (N_687,In_723,N_243);
nand U688 (N_688,In_29,In_87);
nand U689 (N_689,In_1367,In_1415);
and U690 (N_690,In_1539,In_2212);
xor U691 (N_691,In_440,In_787);
and U692 (N_692,In_267,In_1030);
or U693 (N_693,In_779,In_996);
nor U694 (N_694,N_162,N_445);
nor U695 (N_695,In_2347,In_1597);
nor U696 (N_696,In_2289,In_142);
and U697 (N_697,In_400,In_1237);
xnor U698 (N_698,In_2499,In_1543);
xor U699 (N_699,N_419,In_1555);
or U700 (N_700,In_819,In_186);
or U701 (N_701,N_2,In_1227);
and U702 (N_702,In_686,N_332);
and U703 (N_703,In_1846,In_1345);
or U704 (N_704,In_755,In_51);
and U705 (N_705,In_574,In_956);
or U706 (N_706,In_839,In_310);
and U707 (N_707,N_448,In_374);
or U708 (N_708,In_1066,In_2293);
xnor U709 (N_709,In_2296,In_49);
or U710 (N_710,In_164,In_530);
xor U711 (N_711,In_677,In_1741);
nand U712 (N_712,N_60,In_1220);
nand U713 (N_713,In_2115,In_1858);
and U714 (N_714,In_2380,In_2084);
nor U715 (N_715,In_161,N_306);
nor U716 (N_716,In_853,In_1599);
and U717 (N_717,N_172,In_1245);
and U718 (N_718,In_1188,N_580);
nand U719 (N_719,In_359,In_2099);
or U720 (N_720,In_1816,In_894);
and U721 (N_721,In_1569,In_2423);
nand U722 (N_722,In_2195,In_1723);
nand U723 (N_723,In_520,N_236);
and U724 (N_724,In_1815,In_1287);
or U725 (N_725,In_2000,In_952);
and U726 (N_726,In_1110,In_949);
nor U727 (N_727,In_611,N_329);
and U728 (N_728,N_486,In_1372);
nor U729 (N_729,In_399,In_1736);
xor U730 (N_730,N_42,N_383);
and U731 (N_731,In_598,In_1369);
and U732 (N_732,In_96,In_2483);
or U733 (N_733,In_1967,In_26);
and U734 (N_734,In_2090,In_2219);
or U735 (N_735,In_990,In_1751);
xnor U736 (N_736,N_577,In_886);
nand U737 (N_737,In_858,In_1944);
and U738 (N_738,N_81,In_1648);
nand U739 (N_739,N_339,In_1335);
and U740 (N_740,In_602,In_350);
xor U741 (N_741,In_1662,In_1869);
xor U742 (N_742,In_748,In_1226);
xor U743 (N_743,In_1595,N_354);
nor U744 (N_744,N_376,In_1080);
or U745 (N_745,N_454,In_426);
or U746 (N_746,In_1862,In_1375);
xnor U747 (N_747,In_589,N_455);
nor U748 (N_748,In_2251,In_1044);
or U749 (N_749,In_92,N_122);
or U750 (N_750,N_322,In_2453);
nand U751 (N_751,In_351,In_324);
xnor U752 (N_752,In_1670,In_2404);
xor U753 (N_753,N_73,N_64);
nor U754 (N_754,In_836,In_1681);
xor U755 (N_755,In_255,In_263);
nor U756 (N_756,N_594,In_456);
and U757 (N_757,In_370,In_1178);
and U758 (N_758,In_438,N_276);
or U759 (N_759,In_1214,N_246);
and U760 (N_760,N_503,In_516);
nor U761 (N_761,In_213,In_1689);
xor U762 (N_762,N_468,In_1414);
xnor U763 (N_763,In_1917,In_1577);
nand U764 (N_764,In_1568,N_67);
nand U765 (N_765,In_2478,In_18);
nor U766 (N_766,In_1187,In_240);
nand U767 (N_767,N_134,N_447);
nor U768 (N_768,N_254,N_62);
nor U769 (N_769,In_2266,In_951);
xor U770 (N_770,N_94,In_379);
xnor U771 (N_771,N_476,N_35);
nand U772 (N_772,In_1433,N_80);
and U773 (N_773,In_2098,In_2495);
and U774 (N_774,In_1109,In_531);
and U775 (N_775,N_597,In_626);
nand U776 (N_776,In_2286,In_169);
nand U777 (N_777,In_1364,In_1316);
or U778 (N_778,In_1574,In_1881);
and U779 (N_779,In_107,In_1583);
and U780 (N_780,In_1279,In_364);
nand U781 (N_781,In_395,In_2407);
and U782 (N_782,In_1341,N_292);
and U783 (N_783,N_494,In_1515);
nor U784 (N_784,N_181,In_803);
and U785 (N_785,In_1012,In_2032);
and U786 (N_786,In_167,In_60);
and U787 (N_787,In_119,In_221);
and U788 (N_788,In_927,N_104);
xnor U789 (N_789,In_1519,In_19);
or U790 (N_790,In_1107,In_246);
nor U791 (N_791,In_90,In_1284);
nand U792 (N_792,In_2458,In_823);
and U793 (N_793,N_437,N_53);
xnor U794 (N_794,In_1181,In_1472);
nand U795 (N_795,In_349,In_1876);
nor U796 (N_796,In_160,In_1230);
nand U797 (N_797,In_511,In_1350);
nor U798 (N_798,N_57,In_1009);
xnor U799 (N_799,In_284,In_1871);
and U800 (N_800,N_117,N_737);
nor U801 (N_801,In_2170,In_1580);
nor U802 (N_802,In_2316,In_1481);
and U803 (N_803,In_556,In_189);
nand U804 (N_804,In_1021,In_30);
nor U805 (N_805,In_701,In_1778);
and U806 (N_806,In_2148,In_619);
or U807 (N_807,N_799,N_41);
and U808 (N_808,In_1563,N_575);
or U809 (N_809,N_28,In_862);
nor U810 (N_810,In_1129,In_1547);
nand U811 (N_811,N_656,In_2465);
and U812 (N_812,In_897,N_789);
and U813 (N_813,In_908,In_2048);
nor U814 (N_814,In_2422,N_589);
and U815 (N_815,N_463,In_1855);
xnor U816 (N_816,In_498,N_305);
xor U817 (N_817,In_1158,In_1950);
nor U818 (N_818,N_708,In_1938);
or U819 (N_819,In_1607,N_761);
nor U820 (N_820,In_2059,N_714);
nand U821 (N_821,N_619,N_415);
or U822 (N_822,In_1958,In_238);
and U823 (N_823,N_617,In_2233);
nor U824 (N_824,In_1138,In_710);
nor U825 (N_825,In_1139,In_1141);
or U826 (N_826,In_1661,N_459);
and U827 (N_827,N_207,In_887);
xnor U828 (N_828,In_1205,In_587);
or U829 (N_829,N_395,N_724);
xnor U830 (N_830,In_413,N_764);
or U831 (N_831,In_1571,N_512);
nor U832 (N_832,In_2093,In_93);
nor U833 (N_833,N_747,In_243);
nand U834 (N_834,In_147,N_765);
nor U835 (N_835,In_766,N_336);
xor U836 (N_836,In_2037,In_525);
nand U837 (N_837,In_728,In_975);
or U838 (N_838,N_271,N_436);
nor U839 (N_839,In_804,N_556);
or U840 (N_840,In_1769,In_726);
xnor U841 (N_841,N_599,N_61);
nand U842 (N_842,In_56,In_528);
xor U843 (N_843,In_1255,In_2329);
and U844 (N_844,In_432,In_288);
xor U845 (N_845,In_612,N_338);
nand U846 (N_846,N_382,N_370);
or U847 (N_847,In_1087,In_1813);
and U848 (N_848,N_514,N_466);
nor U849 (N_849,In_720,In_1904);
or U850 (N_850,In_1308,N_713);
and U851 (N_851,N_478,In_1566);
nand U852 (N_852,In_2140,N_532);
nor U853 (N_853,In_2248,In_1027);
and U854 (N_854,N_610,In_184);
nand U855 (N_855,N_728,N_757);
nor U856 (N_856,In_2351,In_637);
and U857 (N_857,In_2324,In_105);
and U858 (N_858,In_1052,In_1251);
nand U859 (N_859,N_755,N_366);
and U860 (N_860,In_463,N_337);
nor U861 (N_861,In_1480,N_634);
or U862 (N_862,In_2480,N_93);
xnor U863 (N_863,In_2078,N_333);
and U864 (N_864,In_2262,In_1006);
and U865 (N_865,In_368,In_711);
nor U866 (N_866,In_1997,N_721);
xnor U867 (N_867,N_151,N_702);
nor U868 (N_868,In_1402,N_769);
or U869 (N_869,N_547,In_2178);
xor U870 (N_870,In_535,N_351);
or U871 (N_871,In_591,N_603);
nand U872 (N_872,N_578,In_59);
nor U873 (N_873,In_1346,In_109);
nor U874 (N_874,In_1606,N_161);
or U875 (N_875,In_2109,N_736);
or U876 (N_876,N_20,In_428);
nand U877 (N_877,N_86,In_1934);
xor U878 (N_878,In_99,N_54);
xnor U879 (N_879,N_184,In_2350);
or U880 (N_880,In_941,In_1849);
and U881 (N_881,N_566,N_199);
or U882 (N_882,In_792,In_1520);
or U883 (N_883,In_86,N_742);
xor U884 (N_884,In_2317,In_436);
xnor U885 (N_885,N_483,In_1888);
nand U886 (N_886,In_487,N_71);
or U887 (N_887,N_731,In_2119);
or U888 (N_888,In_868,In_375);
or U889 (N_889,In_583,In_1732);
and U890 (N_890,In_846,In_1785);
or U891 (N_891,In_817,N_373);
xnor U892 (N_892,In_2468,In_1239);
nand U893 (N_893,In_2484,In_729);
and U894 (N_894,N_591,In_362);
and U895 (N_895,In_665,In_2353);
or U896 (N_896,N_792,N_327);
nor U897 (N_897,In_1535,In_361);
or U898 (N_898,In_2172,N_555);
and U899 (N_899,N_260,In_1746);
nand U900 (N_900,N_326,In_765);
xor U901 (N_901,N_200,In_337);
nor U902 (N_902,In_1266,In_888);
xor U903 (N_903,N_360,N_106);
nand U904 (N_904,In_8,N_353);
or U905 (N_905,In_1772,N_773);
nand U906 (N_906,In_606,N_645);
and U907 (N_907,In_628,In_377);
and U908 (N_908,In_158,N_686);
nand U909 (N_909,N_606,In_1584);
xnor U910 (N_910,N_438,N_600);
and U911 (N_911,In_1014,In_1069);
nand U912 (N_912,N_609,In_1810);
xnor U913 (N_913,N_701,In_133);
nand U914 (N_914,N_423,In_241);
nand U915 (N_915,In_1302,In_863);
or U916 (N_916,In_2446,N_411);
xnor U917 (N_917,In_970,In_1865);
nand U918 (N_918,In_1863,N_546);
xnor U919 (N_919,N_551,In_226);
nor U920 (N_920,N_676,In_121);
or U921 (N_921,In_791,In_1447);
or U922 (N_922,In_23,In_78);
nor U923 (N_923,N_559,In_1638);
xnor U924 (N_924,In_1023,In_652);
or U925 (N_925,In_1242,In_2294);
xnor U926 (N_926,In_616,In_1734);
xor U927 (N_927,In_1382,N_695);
and U928 (N_928,In_1641,In_640);
and U929 (N_929,N_432,N_491);
and U930 (N_930,In_725,N_697);
or U931 (N_931,In_2181,In_387);
xor U932 (N_932,N_783,In_1241);
and U933 (N_933,In_1850,N_157);
nand U934 (N_934,In_1092,N_797);
or U935 (N_935,In_1185,N_255);
and U936 (N_936,In_1219,In_2344);
nand U937 (N_937,N_150,In_1038);
or U938 (N_938,In_1601,N_287);
and U939 (N_939,In_188,N_632);
xor U940 (N_940,N_277,In_1317);
nor U941 (N_941,In_2394,In_2240);
and U942 (N_942,N_174,In_2149);
xnor U943 (N_943,N_14,In_1399);
or U944 (N_944,N_776,In_1170);
xnor U945 (N_945,In_1244,N_601);
nand U946 (N_946,In_1441,In_171);
xor U947 (N_947,In_2443,In_103);
xor U948 (N_948,In_1041,In_1154);
nand U949 (N_949,In_2420,In_482);
and U950 (N_950,N_745,In_1176);
xnor U951 (N_951,In_1101,In_293);
nor U952 (N_952,N_270,N_355);
and U953 (N_953,In_1093,In_2077);
nand U954 (N_954,N_760,In_929);
or U955 (N_955,In_2064,N_386);
and U956 (N_956,In_28,In_1941);
nor U957 (N_957,In_1175,N_446);
nor U958 (N_958,N_213,In_1724);
nor U959 (N_959,In_1729,In_0);
and U960 (N_960,N_136,N_471);
nand U961 (N_961,In_2088,In_857);
and U962 (N_962,N_220,In_1310);
xnor U963 (N_963,In_1311,N_4);
xnor U964 (N_964,N_153,In_2255);
or U965 (N_965,In_1224,N_499);
or U966 (N_966,In_2206,In_1005);
nor U967 (N_967,In_824,In_660);
and U968 (N_968,In_579,In_17);
nand U969 (N_969,N_229,In_924);
xor U970 (N_970,In_1,In_1371);
nor U971 (N_971,N_687,N_752);
nand U972 (N_972,N_119,N_490);
and U973 (N_973,N_477,In_1826);
nand U974 (N_974,In_2015,In_2051);
nand U975 (N_975,N_560,In_859);
xnor U976 (N_976,In_627,N_290);
or U977 (N_977,In_935,N_641);
and U978 (N_978,N_753,N_210);
xnor U979 (N_979,N_206,In_592);
nor U980 (N_980,N_689,In_1912);
nor U981 (N_981,In_555,In_1123);
nand U982 (N_982,In_1699,In_2040);
nand U983 (N_983,In_911,N_103);
nand U984 (N_984,In_2472,In_672);
xor U985 (N_985,N_421,In_1306);
or U986 (N_986,In_2106,N_429);
nand U987 (N_987,In_1501,N_76);
xor U988 (N_988,In_716,N_639);
and U989 (N_989,N_612,In_335);
or U990 (N_990,In_410,In_346);
xor U991 (N_991,In_1223,N_673);
and U992 (N_992,N_710,In_1198);
and U993 (N_993,In_1570,N_664);
xnor U994 (N_994,In_1715,In_696);
nor U995 (N_995,N_754,N_201);
nor U996 (N_996,N_460,In_1818);
xnor U997 (N_997,In_236,N_586);
and U998 (N_998,N_412,N_314);
or U999 (N_999,In_821,In_1562);
or U1000 (N_1000,In_1098,N_977);
nor U1001 (N_1001,In_1763,N_320);
or U1002 (N_1002,N_280,In_1081);
xnor U1003 (N_1003,N_667,In_775);
nor U1004 (N_1004,N_894,In_2292);
or U1005 (N_1005,In_2473,In_553);
nor U1006 (N_1006,N_258,In_1567);
xor U1007 (N_1007,N_520,In_460);
or U1008 (N_1008,In_466,In_985);
or U1009 (N_1009,In_524,In_2413);
xor U1010 (N_1010,N_808,N_830);
and U1011 (N_1011,N_800,N_39);
xor U1012 (N_1012,N_216,In_1182);
nor U1013 (N_1013,N_786,N_492);
or U1014 (N_1014,N_809,In_232);
nand U1015 (N_1015,In_746,In_1040);
and U1016 (N_1016,N_970,In_64);
and U1017 (N_1017,N_680,N_870);
and U1018 (N_1018,In_2355,In_2011);
xnor U1019 (N_1019,N_827,In_867);
xor U1020 (N_1020,N_288,N_425);
and U1021 (N_1021,In_2060,In_643);
nand U1022 (N_1022,In_562,In_1363);
nand U1023 (N_1023,In_416,In_1708);
or U1024 (N_1024,In_508,In_501);
xnor U1025 (N_1025,In_1461,N_250);
nor U1026 (N_1026,N_565,N_462);
and U1027 (N_1027,In_737,In_742);
xnor U1028 (N_1028,N_456,N_130);
or U1029 (N_1029,In_2141,In_805);
or U1030 (N_1030,In_673,N_875);
xnor U1031 (N_1031,In_588,N_537);
and U1032 (N_1032,In_2110,N_616);
nand U1033 (N_1033,In_1954,In_708);
xnor U1034 (N_1034,N_759,N_748);
xnor U1035 (N_1035,N_8,In_1342);
nor U1036 (N_1036,In_931,N_115);
and U1037 (N_1037,N_867,N_756);
and U1038 (N_1038,In_2264,In_1505);
nor U1039 (N_1039,In_1650,In_1956);
and U1040 (N_1040,In_1061,N_367);
or U1041 (N_1041,N_981,In_84);
and U1042 (N_1042,In_1268,In_1642);
or U1043 (N_1043,In_2432,In_727);
or U1044 (N_1044,N_553,N_984);
and U1045 (N_1045,In_1444,In_2146);
nand U1046 (N_1046,N_823,In_2387);
and U1047 (N_1047,In_1841,N_444);
nor U1048 (N_1048,In_2065,In_1564);
nor U1049 (N_1049,In_69,In_417);
nor U1050 (N_1050,In_1173,In_247);
nand U1051 (N_1051,N_895,In_992);
xnor U1052 (N_1052,N_819,In_1671);
xor U1053 (N_1053,In_1593,In_1216);
and U1054 (N_1054,N_877,In_1060);
or U1055 (N_1055,In_731,In_345);
nor U1056 (N_1056,In_928,In_253);
nor U1057 (N_1057,In_2322,In_2095);
or U1058 (N_1058,N_484,In_114);
nor U1059 (N_1059,N_832,N_441);
xor U1060 (N_1060,N_707,In_2314);
nor U1061 (N_1061,In_2174,N_147);
xnor U1062 (N_1062,In_398,N_717);
xnor U1063 (N_1063,In_1254,N_855);
xor U1064 (N_1064,In_2399,N_10);
nor U1065 (N_1065,In_2378,N_933);
or U1066 (N_1066,N_638,N_574);
and U1067 (N_1067,In_141,In_678);
and U1068 (N_1068,N_25,N_674);
or U1069 (N_1069,In_958,In_1845);
nand U1070 (N_1070,In_423,In_745);
or U1071 (N_1071,In_942,In_1418);
nand U1072 (N_1072,In_840,In_1150);
and U1073 (N_1073,In_2445,N_344);
xor U1074 (N_1074,N_521,In_1484);
nand U1075 (N_1075,N_733,In_2456);
xnor U1076 (N_1076,N_940,In_736);
and U1077 (N_1077,N_805,N_205);
nor U1078 (N_1078,N_451,In_1136);
xor U1079 (N_1079,N_677,In_1612);
or U1080 (N_1080,N_107,N_893);
or U1081 (N_1081,In_1340,In_1933);
xnor U1082 (N_1082,In_811,In_1180);
and U1083 (N_1083,N_987,In_1071);
nand U1084 (N_1084,In_13,In_954);
nand U1085 (N_1085,In_1225,In_1534);
nor U1086 (N_1086,N_951,In_1330);
nor U1087 (N_1087,In_462,In_1247);
xnor U1088 (N_1088,In_2028,In_599);
or U1089 (N_1089,N_5,N_544);
nor U1090 (N_1090,N_953,In_527);
nor U1091 (N_1091,In_1962,In_444);
and U1092 (N_1092,In_390,In_932);
and U1093 (N_1093,In_1379,N_740);
and U1094 (N_1094,In_1542,N_935);
xnor U1095 (N_1095,In_1531,N_605);
nand U1096 (N_1096,N_406,N_906);
nor U1097 (N_1097,N_297,In_1285);
xor U1098 (N_1098,In_733,N_973);
xor U1099 (N_1099,In_812,In_2471);
or U1100 (N_1100,In_479,In_2328);
or U1101 (N_1101,In_1874,In_2162);
nand U1102 (N_1102,N_440,In_768);
xnor U1103 (N_1103,N_834,In_1099);
xor U1104 (N_1104,In_537,N_803);
nor U1105 (N_1105,In_1195,In_41);
or U1106 (N_1106,In_2012,In_274);
or U1107 (N_1107,In_2034,In_306);
nand U1108 (N_1108,In_2002,In_2180);
xor U1109 (N_1109,N_964,In_1344);
xor U1110 (N_1110,In_1143,In_1400);
nor U1111 (N_1111,N_278,N_622);
nor U1112 (N_1112,N_835,In_1968);
nor U1113 (N_1113,In_2368,N_644);
or U1114 (N_1114,N_439,N_831);
xnor U1115 (N_1115,In_467,In_1972);
nand U1116 (N_1116,N_716,In_856);
nor U1117 (N_1117,N_642,N_671);
or U1118 (N_1118,In_2176,N_853);
nor U1119 (N_1119,N_584,N_941);
xnor U1120 (N_1120,N_804,In_1011);
nand U1121 (N_1121,In_641,In_1685);
nor U1122 (N_1122,In_1998,In_2236);
xnor U1123 (N_1123,N_418,In_27);
xor U1124 (N_1124,In_2139,In_1839);
xnor U1125 (N_1125,N_420,In_756);
xor U1126 (N_1126,In_1380,In_507);
and U1127 (N_1127,N_582,In_529);
and U1128 (N_1128,N_182,N_696);
and U1129 (N_1129,N_907,N_399);
and U1130 (N_1130,In_590,N_240);
nor U1131 (N_1131,N_851,In_692);
nand U1132 (N_1132,N_298,In_204);
or U1133 (N_1133,N_822,In_477);
nor U1134 (N_1134,In_352,In_494);
and U1135 (N_1135,N_852,In_2117);
and U1136 (N_1136,N_528,N_909);
or U1137 (N_1137,In_1795,N_238);
and U1138 (N_1138,In_700,N_635);
and U1139 (N_1139,In_1740,N_807);
xnor U1140 (N_1140,N_188,N_375);
xnor U1141 (N_1141,In_2113,In_2221);
or U1142 (N_1142,In_1521,N_400);
and U1143 (N_1143,In_2281,In_1887);
nand U1144 (N_1144,In_989,In_411);
nor U1145 (N_1145,N_230,In_1908);
or U1146 (N_1146,In_170,N_380);
nor U1147 (N_1147,In_566,N_510);
or U1148 (N_1148,N_675,N_901);
xor U1149 (N_1149,N_347,N_682);
or U1150 (N_1150,In_759,N_166);
xor U1151 (N_1151,N_461,N_307);
nand U1152 (N_1152,In_220,N_666);
and U1153 (N_1153,N_531,In_31);
and U1154 (N_1154,N_262,In_357);
nor U1155 (N_1155,N_613,In_968);
and U1156 (N_1156,N_836,N_669);
or U1157 (N_1157,N_365,N_524);
nand U1158 (N_1158,N_433,In_2145);
nor U1159 (N_1159,In_1260,N_286);
and U1160 (N_1160,In_1451,In_1824);
nand U1161 (N_1161,In_1835,In_2448);
xor U1162 (N_1162,In_1113,In_1496);
or U1163 (N_1163,In_405,In_957);
nand U1164 (N_1164,N_467,In_298);
nor U1165 (N_1165,In_355,N_665);
or U1166 (N_1166,In_104,N_684);
nand U1167 (N_1167,In_336,In_2062);
or U1168 (N_1168,In_670,In_25);
or U1169 (N_1169,N_653,In_1922);
nand U1170 (N_1170,N_464,In_1438);
and U1171 (N_1171,In_191,In_655);
and U1172 (N_1172,In_342,N_390);
and U1173 (N_1173,In_2016,In_1805);
or U1174 (N_1174,In_978,In_1770);
nand U1175 (N_1175,In_202,N_889);
nand U1176 (N_1176,In_1428,N_976);
nand U1177 (N_1177,In_568,N_92);
nand U1178 (N_1178,N_845,N_848);
nand U1179 (N_1179,In_973,N_898);
or U1180 (N_1180,In_225,In_1263);
or U1181 (N_1181,In_1468,In_689);
nor U1182 (N_1182,In_2126,N_317);
or U1183 (N_1183,N_690,In_739);
and U1184 (N_1184,In_2313,In_1155);
nand U1185 (N_1185,N_892,N_497);
nor U1186 (N_1186,In_1983,N_52);
nand U1187 (N_1187,N_120,N_529);
xor U1188 (N_1188,In_953,N_871);
or U1189 (N_1189,In_777,In_2469);
or U1190 (N_1190,In_658,In_1663);
and U1191 (N_1191,N_267,N_65);
nor U1192 (N_1192,In_168,In_2085);
xnor U1193 (N_1193,In_1844,N_604);
and U1194 (N_1194,In_1640,In_651);
or U1195 (N_1195,N_114,In_515);
xnor U1196 (N_1196,N_959,In_257);
nor U1197 (N_1197,In_1349,In_1277);
nor U1198 (N_1198,In_394,N_954);
nand U1199 (N_1199,N_762,N_573);
nand U1200 (N_1200,In_1722,In_781);
or U1201 (N_1201,In_193,In_2260);
nor U1202 (N_1202,N_1096,In_1100);
and U1203 (N_1203,In_1485,N_1129);
xor U1204 (N_1204,In_844,N_303);
nand U1205 (N_1205,N_741,In_1343);
and U1206 (N_1206,In_883,N_498);
or U1207 (N_1207,N_699,N_921);
xnor U1208 (N_1208,N_1027,In_366);
nor U1209 (N_1209,In_2295,In_1598);
or U1210 (N_1210,In_1425,N_231);
xnor U1211 (N_1211,In_1119,N_825);
and U1212 (N_1212,N_1181,N_1002);
nor U1213 (N_1213,N_405,In_1261);
and U1214 (N_1214,N_980,In_2250);
or U1215 (N_1215,In_1930,In_1743);
xnor U1216 (N_1216,In_264,In_435);
xor U1217 (N_1217,In_1396,In_1969);
or U1218 (N_1218,N_1109,In_2433);
nand U1219 (N_1219,N_474,N_135);
and U1220 (N_1220,N_221,N_919);
xnor U1221 (N_1221,In_407,In_1697);
nand U1222 (N_1222,N_1038,In_273);
xor U1223 (N_1223,N_715,N_923);
nand U1224 (N_1224,In_948,In_617);
nor U1225 (N_1225,In_1851,In_2186);
xnor U1226 (N_1226,In_546,N_1166);
or U1227 (N_1227,N_1118,N_513);
xor U1228 (N_1228,In_662,N_1052);
and U1229 (N_1229,In_291,N_903);
nand U1230 (N_1230,In_1621,In_1788);
and U1231 (N_1231,In_430,In_251);
xor U1232 (N_1232,In_383,N_624);
or U1233 (N_1233,N_1095,N_672);
nand U1234 (N_1234,In_2375,N_518);
and U1235 (N_1235,In_1144,In_1168);
and U1236 (N_1236,N_993,N_900);
nor U1237 (N_1237,In_1747,In_2182);
or U1238 (N_1238,N_361,In_747);
xor U1239 (N_1239,In_429,N_887);
nand U1240 (N_1240,In_404,In_1766);
or U1241 (N_1241,N_846,N_567);
nand U1242 (N_1242,In_1711,N_718);
nand U1243 (N_1243,In_806,N_861);
xor U1244 (N_1244,In_1964,N_997);
and U1245 (N_1245,In_299,In_1116);
nor U1246 (N_1246,In_1594,In_2238);
and U1247 (N_1247,N_149,N_269);
or U1248 (N_1248,N_15,N_394);
nand U1249 (N_1249,N_1090,N_723);
nor U1250 (N_1250,In_2321,N_1099);
and U1251 (N_1251,N_963,N_1034);
nor U1252 (N_1252,In_2470,N_1145);
nand U1253 (N_1253,N_969,N_585);
xnor U1254 (N_1254,In_2302,In_2425);
nor U1255 (N_1255,In_85,N_847);
xnor U1256 (N_1256,N_842,In_1940);
nand U1257 (N_1257,In_48,N_854);
nand U1258 (N_1258,In_1003,In_1217);
nand U1259 (N_1259,N_1169,In_2337);
xor U1260 (N_1260,In_1660,N_1110);
and U1261 (N_1261,In_1902,N_1150);
nor U1262 (N_1262,In_115,N_955);
nor U1263 (N_1263,In_280,N_1089);
xnor U1264 (N_1264,N_1175,N_948);
xnor U1265 (N_1265,N_1199,N_1008);
and U1266 (N_1266,In_2261,N_711);
nor U1267 (N_1267,N_1033,In_1059);
nand U1268 (N_1268,In_2360,In_1270);
and U1269 (N_1269,N_781,In_1300);
nand U1270 (N_1270,In_965,In_2025);
xnor U1271 (N_1271,In_1744,N_192);
xnor U1272 (N_1272,N_608,N_253);
nor U1273 (N_1273,In_1028,In_308);
or U1274 (N_1274,N_234,In_852);
nor U1275 (N_1275,In_1121,In_2299);
nor U1276 (N_1276,N_501,In_1833);
nor U1277 (N_1277,N_1079,In_146);
and U1278 (N_1278,N_620,N_417);
and U1279 (N_1279,N_1160,N_1015);
and U1280 (N_1280,N_1108,In_926);
and U1281 (N_1281,N_21,In_2132);
and U1282 (N_1282,N_924,N_974);
xnor U1283 (N_1283,N_124,N_137);
nor U1284 (N_1284,N_1063,In_2128);
nor U1285 (N_1285,N_782,N_1147);
xnor U1286 (N_1286,N_975,In_1497);
or U1287 (N_1287,In_2152,N_899);
nand U1288 (N_1288,In_1502,In_2205);
xor U1289 (N_1289,N_204,N_659);
or U1290 (N_1290,In_892,N_334);
xor U1291 (N_1291,N_1026,In_1053);
or U1292 (N_1292,In_661,N_960);
nor U1293 (N_1293,N_1050,N_576);
and U1294 (N_1294,N_650,In_2379);
xnor U1295 (N_1295,In_644,In_2079);
nand U1296 (N_1296,In_906,N_627);
nand U1297 (N_1297,N_118,In_600);
or U1298 (N_1298,In_1422,N_1000);
or U1299 (N_1299,In_526,N_758);
xor U1300 (N_1300,N_631,In_178);
and U1301 (N_1301,In_302,In_1374);
nand U1302 (N_1302,N_139,In_1955);
xnor U1303 (N_1303,In_1166,In_312);
nand U1304 (N_1304,In_205,N_295);
nor U1305 (N_1305,In_1165,In_1647);
nor U1306 (N_1306,N_435,N_1020);
or U1307 (N_1307,N_660,N_79);
xor U1308 (N_1308,In_1145,N_377);
nand U1309 (N_1309,In_1033,In_208);
nor U1310 (N_1310,In_2125,N_569);
and U1311 (N_1311,In_1817,N_850);
nand U1312 (N_1312,N_636,In_809);
and U1313 (N_1313,In_136,N_145);
xnor U1314 (N_1314,In_2183,In_21);
and U1315 (N_1315,In_2023,In_2038);
xor U1316 (N_1316,N_946,N_1152);
or U1317 (N_1317,In_2159,N_570);
or U1318 (N_1318,In_396,In_714);
nand U1319 (N_1319,N_525,In_2408);
and U1320 (N_1320,N_939,N_607);
and U1321 (N_1321,In_2228,N_862);
nor U1322 (N_1322,In_982,N_1177);
nor U1323 (N_1323,In_680,N_908);
and U1324 (N_1324,In_1780,N_350);
nand U1325 (N_1325,In_40,In_2001);
nand U1326 (N_1326,In_2370,N_1135);
nor U1327 (N_1327,In_1355,In_1250);
or U1328 (N_1328,In_2405,N_1045);
nor U1329 (N_1329,N_679,N_772);
nand U1330 (N_1330,N_725,In_2072);
nor U1331 (N_1331,N_957,In_997);
and U1332 (N_1332,N_167,In_2320);
or U1333 (N_1333,In_382,In_1193);
nor U1334 (N_1334,N_581,In_1971);
xor U1335 (N_1335,In_1257,In_1522);
and U1336 (N_1336,In_1608,In_684);
nand U1337 (N_1337,N_226,In_2246);
or U1338 (N_1338,N_1087,N_1161);
and U1339 (N_1339,N_885,In_2058);
xor U1340 (N_1340,In_143,In_778);
and U1341 (N_1341,N_1056,In_478);
xor U1342 (N_1342,N_233,N_1071);
nor U1343 (N_1343,In_1169,In_1315);
or U1344 (N_1344,N_225,N_179);
nor U1345 (N_1345,N_625,N_9);
or U1346 (N_1346,N_863,N_661);
and U1347 (N_1347,In_1988,In_418);
nor U1348 (N_1348,In_654,N_662);
and U1349 (N_1349,N_828,In_2253);
nand U1350 (N_1350,In_1657,In_1204);
and U1351 (N_1351,In_1167,N_785);
and U1352 (N_1352,In_409,N_985);
nor U1353 (N_1353,N_1068,In_265);
nor U1354 (N_1354,N_595,N_404);
nor U1355 (N_1355,In_22,In_552);
or U1356 (N_1356,N_507,In_2102);
nand U1357 (N_1357,In_1384,In_1486);
or U1358 (N_1358,N_693,In_1513);
nand U1359 (N_1359,In_1643,N_232);
xnor U1360 (N_1360,N_105,In_2234);
or U1361 (N_1361,N_368,N_379);
or U1362 (N_1362,N_1055,In_2438);
nand U1363 (N_1363,N_814,In_135);
nand U1364 (N_1364,In_452,N_995);
nor U1365 (N_1365,N_352,N_775);
and U1366 (N_1366,In_2452,N_224);
and U1367 (N_1367,N_583,N_1005);
nand U1368 (N_1368,N_947,N_1070);
xor U1369 (N_1369,In_1859,In_1615);
xor U1370 (N_1370,N_66,N_750);
and U1371 (N_1371,N_602,In_2156);
xnor U1372 (N_1372,In_679,N_550);
nor U1373 (N_1373,In_1161,In_1668);
or U1374 (N_1374,In_1278,N_1174);
and U1375 (N_1375,N_1168,In_1991);
or U1376 (N_1376,N_143,In_154);
xnor U1377 (N_1377,N_967,N_389);
nand U1378 (N_1378,In_1559,N_450);
nor U1379 (N_1379,In_2447,N_502);
or U1380 (N_1380,In_1280,N_952);
nand U1381 (N_1381,N_1073,N_144);
nor U1382 (N_1382,N_864,N_878);
xor U1383 (N_1383,N_1084,N_668);
or U1384 (N_1384,In_1025,N_1031);
nand U1385 (N_1385,In_798,In_2398);
or U1386 (N_1386,N_1192,In_1183);
xnor U1387 (N_1387,N_416,In_979);
and U1388 (N_1388,In_540,N_242);
xnor U1389 (N_1389,N_488,In_1920);
nor U1390 (N_1390,N_843,In_391);
nor U1391 (N_1391,In_2442,N_880);
or U1392 (N_1392,In_964,N_628);
nand U1393 (N_1393,N_651,N_1018);
or U1394 (N_1394,In_1617,N_1148);
or U1395 (N_1395,In_173,In_1370);
and U1396 (N_1396,In_50,N_1014);
and U1397 (N_1397,N_593,In_286);
nand U1398 (N_1398,N_826,N_489);
nor U1399 (N_1399,In_761,N_18);
xnor U1400 (N_1400,N_691,In_1043);
nor U1401 (N_1401,N_1296,N_548);
nor U1402 (N_1402,N_780,N_308);
xor U1403 (N_1403,In_2124,In_1899);
nand U1404 (N_1404,N_385,N_1378);
or U1405 (N_1405,N_1158,In_1726);
or U1406 (N_1406,In_2073,In_1366);
xnor U1407 (N_1407,N_1080,In_1448);
nor U1408 (N_1408,In_2384,N_1338);
or U1409 (N_1409,N_1316,In_488);
or U1410 (N_1410,N_1128,N_1365);
or U1411 (N_1411,In_2203,N_378);
nand U1412 (N_1412,N_744,N_1083);
and U1413 (N_1413,N_1315,N_1359);
and U1414 (N_1414,N_1346,In_1032);
nand U1415 (N_1415,N_1167,In_559);
or U1416 (N_1416,N_227,In_1508);
xor U1417 (N_1417,N_358,In_1495);
xor U1418 (N_1418,N_1142,N_879);
and U1419 (N_1419,In_1633,In_2202);
and U1420 (N_1420,In_1684,N_1250);
nand U1421 (N_1421,In_1417,N_1368);
and U1422 (N_1422,In_2154,N_1042);
nand U1423 (N_1423,In_1526,N_244);
and U1424 (N_1424,N_1356,N_1279);
nor U1425 (N_1425,N_363,N_1206);
and U1426 (N_1426,N_540,In_1680);
or U1427 (N_1427,N_839,N_562);
nor U1428 (N_1428,In_439,N_860);
nand U1429 (N_1429,N_1114,In_1666);
xnor U1430 (N_1430,N_1007,N_1342);
nor U1431 (N_1431,In_1619,N_568);
nand U1432 (N_1432,In_2397,N_1054);
nand U1433 (N_1433,N_1057,N_905);
nor U1434 (N_1434,In_272,N_1143);
nor U1435 (N_1435,In_1046,In_1759);
nor U1436 (N_1436,In_2163,N_685);
and U1437 (N_1437,In_1489,N_1335);
nand U1438 (N_1438,In_1424,In_1673);
nand U1439 (N_1439,N_1322,N_1264);
xnor U1440 (N_1440,In_1164,In_1243);
nor U1441 (N_1441,N_1301,N_1249);
nor U1442 (N_1442,In_1319,N_6);
nor U1443 (N_1443,N_475,N_1106);
or U1444 (N_1444,N_1124,In_917);
and U1445 (N_1445,N_927,N_986);
nand U1446 (N_1446,N_1139,N_1115);
or U1447 (N_1447,N_991,N_956);
nor U1448 (N_1448,In_712,N_300);
xor U1449 (N_1449,In_1895,In_874);
xor U1450 (N_1450,N_473,In_1748);
or U1451 (N_1451,N_934,N_1091);
nor U1452 (N_1452,In_1378,In_1716);
nor U1453 (N_1453,In_707,In_994);
nand U1454 (N_1454,N_1260,In_1735);
or U1455 (N_1455,N_1350,N_729);
nand U1456 (N_1456,In_393,N_1207);
xor U1457 (N_1457,N_1218,N_1019);
xor U1458 (N_1458,N_470,N_1004);
nand U1459 (N_1459,N_838,N_868);
xor U1460 (N_1460,N_658,In_666);
xnor U1461 (N_1461,In_676,N_396);
or U1462 (N_1462,N_962,In_322);
nor U1463 (N_1463,N_1154,In_1149);
xor U1464 (N_1464,In_848,In_1538);
nand U1465 (N_1465,In_2390,N_99);
xor U1466 (N_1466,N_1049,N_1387);
xnor U1467 (N_1467,N_796,N_1277);
or U1468 (N_1468,N_1347,N_1329);
nand U1469 (N_1469,N_1337,N_798);
xnor U1470 (N_1470,In_1877,N_1006);
and U1471 (N_1471,N_1185,N_614);
or U1472 (N_1472,N_883,N_996);
nor U1473 (N_1473,N_703,In_1420);
and U1474 (N_1474,N_428,In_1085);
nor U1475 (N_1475,In_279,N_1372);
nand U1476 (N_1476,N_743,N_1251);
nor U1477 (N_1477,N_881,N_771);
xnor U1478 (N_1478,N_1190,N_1183);
or U1479 (N_1479,N_1395,N_169);
or U1480 (N_1480,N_897,In_1856);
nor U1481 (N_1481,In_1199,N_40);
and U1482 (N_1482,N_1292,In_4);
nand U1483 (N_1483,N_1321,N_1320);
and U1484 (N_1484,N_1088,N_500);
or U1485 (N_1485,In_2258,N_534);
nor U1486 (N_1486,In_1838,In_905);
nor U1487 (N_1487,N_1360,N_211);
xor U1488 (N_1488,In_153,N_1029);
nand U1489 (N_1489,In_1056,In_837);
nand U1490 (N_1490,N_282,In_1915);
or U1491 (N_1491,N_1352,In_1487);
nand U1492 (N_1492,N_535,In_603);
xor U1493 (N_1493,N_1241,N_27);
xor U1494 (N_1494,N_681,N_787);
and U1495 (N_1495,In_1664,In_1401);
and U1496 (N_1496,N_426,N_936);
xnor U1497 (N_1497,N_239,In_1789);
and U1498 (N_1498,N_630,In_1172);
or U1499 (N_1499,In_1802,In_2339);
nand U1500 (N_1500,In_447,In_1203);
and U1501 (N_1501,N_945,In_1596);
nand U1502 (N_1502,In_880,N_1238);
xor U1503 (N_1503,N_1276,N_647);
xor U1504 (N_1504,In_1898,N_403);
nor U1505 (N_1505,N_874,N_1119);
xnor U1506 (N_1506,N_328,N_813);
nand U1507 (N_1507,In_1557,In_854);
nor U1508 (N_1508,N_1032,N_1333);
nand U1509 (N_1509,N_833,N_1282);
nand U1510 (N_1510,N_1155,N_1170);
or U1511 (N_1511,In_2393,N_431);
nand U1512 (N_1512,In_1200,In_1549);
xnor U1513 (N_1513,N_1269,N_1266);
or U1514 (N_1514,In_2247,N_904);
nand U1515 (N_1515,In_780,In_2224);
nor U1516 (N_1516,N_442,N_801);
nor U1517 (N_1517,N_402,N_1103);
nor U1518 (N_1518,N_869,In_128);
and U1519 (N_1519,N_794,N_1343);
xnor U1520 (N_1520,In_1973,In_319);
and U1521 (N_1521,N_1116,In_2477);
nor U1522 (N_1522,In_1919,N_1384);
nor U1523 (N_1523,N_1284,N_1328);
xnor U1524 (N_1524,N_1178,N_1246);
and U1525 (N_1525,In_1190,N_316);
nand U1526 (N_1526,N_1105,N_430);
nor U1527 (N_1527,In_2239,N_777);
nor U1528 (N_1528,N_590,In_190);
and U1529 (N_1529,In_2334,N_263);
nand U1530 (N_1530,In_1924,N_929);
and U1531 (N_1531,In_1234,N_1123);
xor U1532 (N_1532,N_856,In_214);
or U1533 (N_1533,N_1332,N_116);
or U1534 (N_1534,In_1581,N_1289);
nand U1535 (N_1535,N_746,In_1852);
nand U1536 (N_1536,N_493,In_2030);
nand U1537 (N_1537,N_1125,N_183);
nor U1538 (N_1538,In_1561,In_875);
nor U1539 (N_1539,N_784,In_1738);
or U1540 (N_1540,N_1393,N_774);
and U1541 (N_1541,N_479,N_1326);
nand U1542 (N_1542,In_618,In_301);
nor U1543 (N_1543,In_397,In_108);
and U1544 (N_1544,N_1309,N_722);
and U1545 (N_1545,In_2168,N_1157);
nand U1546 (N_1546,In_1654,In_2232);
xnor U1547 (N_1547,N_414,N_1120);
nor U1548 (N_1548,N_1137,N_1285);
xor U1549 (N_1549,N_712,In_668);
or U1550 (N_1550,N_1180,N_218);
and U1551 (N_1551,In_2045,In_458);
xor U1552 (N_1552,In_1091,N_1041);
nand U1553 (N_1553,N_504,In_624);
and U1554 (N_1554,N_1272,N_434);
or U1555 (N_1555,In_1218,N_633);
xor U1556 (N_1556,N_482,N_1369);
nand U1557 (N_1557,N_1225,In_471);
xnor U1558 (N_1558,N_598,N_1194);
xnor U1559 (N_1559,N_1317,N_706);
xnor U1560 (N_1560,N_1366,N_1304);
nor U1561 (N_1561,In_1720,In_347);
nand U1562 (N_1562,N_1274,N_942);
xor U1563 (N_1563,N_1062,In_1757);
and U1564 (N_1564,N_1243,In_999);
and U1565 (N_1565,N_371,N_931);
nand U1566 (N_1566,In_1786,N_1028);
xor U1567 (N_1567,N_1001,N_511);
xor U1568 (N_1568,In_1948,N_1340);
and U1569 (N_1569,N_890,In_1409);
nand U1570 (N_1570,In_1246,N_971);
and U1571 (N_1571,In_334,In_1916);
and U1572 (N_1572,N_58,N_1361);
or U1573 (N_1573,N_932,In_955);
or U1574 (N_1574,N_818,N_592);
and U1575 (N_1575,N_872,In_2061);
xnor U1576 (N_1576,In_921,In_1329);
or U1577 (N_1577,N_1209,N_545);
or U1578 (N_1578,N_1270,N_1235);
xnor U1579 (N_1579,In_807,N_817);
xnor U1580 (N_1580,In_287,N_734);
nand U1581 (N_1581,N_1156,N_1003);
or U1582 (N_1582,N_196,N_1345);
and U1583 (N_1583,N_1363,In_2354);
or U1584 (N_1584,N_413,N_508);
nand U1585 (N_1585,N_911,In_15);
or U1586 (N_1586,N_1037,In_1745);
nor U1587 (N_1587,N_1287,In_1556);
or U1588 (N_1588,In_242,In_450);
xnor U1589 (N_1589,N_1201,N_407);
nor U1590 (N_1590,N_1247,N_1308);
nor U1591 (N_1591,N_749,N_561);
or U1592 (N_1592,N_1275,In_2303);
nor U1593 (N_1593,N_1021,In_66);
nor U1594 (N_1594,N_1104,N_1223);
xor U1595 (N_1595,N_1377,N_1046);
nor U1596 (N_1596,In_1435,N_961);
nand U1597 (N_1597,N_465,N_1127);
or U1598 (N_1598,In_1652,N_886);
nor U1599 (N_1599,N_1390,N_873);
or U1600 (N_1600,In_571,N_1010);
xor U1601 (N_1601,N_1531,In_2297);
xor U1602 (N_1602,N_1134,N_663);
and U1603 (N_1603,N_1402,In_1590);
or U1604 (N_1604,N_579,In_2092);
nand U1605 (N_1605,N_944,In_1394);
nor U1606 (N_1606,In_2097,N_1205);
xnor U1607 (N_1607,N_1558,N_1196);
and U1608 (N_1608,In_757,In_1322);
nand U1609 (N_1609,In_442,N_1440);
nor U1610 (N_1610,N_1509,In_2123);
nand U1611 (N_1611,N_1173,N_698);
nand U1612 (N_1612,N_1483,N_1072);
or U1613 (N_1613,N_1252,N_1576);
or U1614 (N_1614,N_1462,In_360);
and U1615 (N_1615,N_1484,N_1051);
or U1616 (N_1616,N_1519,N_1460);
nor U1617 (N_1617,N_790,N_1258);
or U1618 (N_1618,In_1186,N_1546);
or U1619 (N_1619,N_1300,N_806);
nand U1620 (N_1620,In_1492,In_384);
xor U1621 (N_1621,N_1478,N_1396);
and U1622 (N_1622,N_821,N_1231);
nand U1623 (N_1623,N_621,N_1438);
and U1624 (N_1624,N_1461,In_320);
nor U1625 (N_1625,N_1319,N_1086);
nand U1626 (N_1626,N_965,N_979);
xnor U1627 (N_1627,In_1312,N_1064);
and U1628 (N_1628,N_1397,N_1581);
xnor U1629 (N_1629,In_934,In_1923);
and U1630 (N_1630,N_1291,N_1392);
xnor U1631 (N_1631,N_704,N_1548);
xnor U1632 (N_1632,N_1597,In_940);
xor U1633 (N_1633,N_509,N_1524);
nand U1634 (N_1634,N_1591,In_2173);
xnor U1635 (N_1635,In_1980,N_1455);
nor U1636 (N_1636,N_1491,In_1074);
xnor U1637 (N_1637,N_235,N_1324);
xor U1638 (N_1638,In_879,In_914);
xnor U1639 (N_1639,In_262,In_2279);
xnor U1640 (N_1640,N_1217,N_1144);
and U1641 (N_1641,In_1506,N_1570);
xnor U1642 (N_1642,In_1628,In_1112);
xor U1643 (N_1643,N_1434,N_1248);
or U1644 (N_1644,In_835,N_549);
and U1645 (N_1645,N_1358,N_1433);
xnor U1646 (N_1646,In_1787,In_162);
nand U1647 (N_1647,In_449,N_1327);
nand U1648 (N_1648,N_643,N_1528);
and U1649 (N_1649,N_990,N_1526);
nand U1650 (N_1650,N_87,N_1439);
or U1651 (N_1651,In_1977,N_700);
and U1652 (N_1652,N_1458,N_374);
nor U1653 (N_1653,N_876,In_2188);
nand U1654 (N_1654,In_1473,N_1405);
nor U1655 (N_1655,N_1030,In_1674);
and U1656 (N_1656,N_829,N_1288);
nor U1657 (N_1657,In_42,N_1573);
nand U1658 (N_1658,N_1515,In_1157);
nand U1659 (N_1659,N_1593,In_1179);
or U1660 (N_1660,N_1543,N_678);
nor U1661 (N_1661,In_503,N_649);
and U1662 (N_1662,N_1236,N_1025);
xor U1663 (N_1663,N_1513,N_1100);
xnor U1664 (N_1664,In_1880,N_1182);
xnor U1665 (N_1665,N_648,N_1575);
xor U1666 (N_1666,N_811,In_2415);
nand U1667 (N_1667,N_284,N_1432);
or U1668 (N_1668,N_1081,N_1061);
and U1669 (N_1669,In_166,N_1424);
nand U1670 (N_1670,N_1482,N_1349);
nor U1671 (N_1671,N_296,N_1149);
nand U1672 (N_1672,N_626,N_1481);
nor U1673 (N_1673,N_1471,N_1496);
xor U1674 (N_1674,In_2108,N_1508);
nand U1675 (N_1675,In_1354,In_177);
nor U1676 (N_1676,N_1228,In_2014);
or U1677 (N_1677,N_1133,N_1564);
and U1678 (N_1678,In_577,N_335);
or U1679 (N_1679,In_1352,N_90);
or U1680 (N_1680,N_1268,N_480);
or U1681 (N_1681,In_2054,In_1456);
and U1682 (N_1682,N_925,N_1075);
nor U1683 (N_1683,N_3,N_1584);
nand U1684 (N_1684,In_2196,In_1682);
and U1685 (N_1685,In_2494,N_1210);
and U1686 (N_1686,N_1443,N_926);
and U1687 (N_1687,In_683,In_2256);
nor U1688 (N_1688,N_1556,N_1039);
and U1689 (N_1689,In_1050,N_1043);
nor U1690 (N_1690,N_1585,N_1547);
and U1691 (N_1691,N_1549,In_199);
and U1692 (N_1692,N_1354,N_1588);
nand U1693 (N_1693,N_1280,N_1409);
nor U1694 (N_1694,N_302,N_1213);
nor U1695 (N_1695,In_2315,N_1572);
and U1696 (N_1696,N_1518,N_1497);
or U1697 (N_1697,N_1331,In_174);
xor U1698 (N_1698,N_356,In_81);
nor U1699 (N_1699,N_937,N_950);
xnor U1700 (N_1700,N_1431,N_1348);
and U1701 (N_1701,N_1085,N_778);
nor U1702 (N_1702,In_1605,In_1235);
xor U1703 (N_1703,N_989,N_16);
and U1704 (N_1704,N_1253,In_385);
or U1705 (N_1705,N_1536,In_621);
nor U1706 (N_1706,N_727,In_573);
and U1707 (N_1707,N_1164,N_1244);
xor U1708 (N_1708,N_219,In_459);
and U1709 (N_1709,In_1953,N_1569);
or U1710 (N_1710,N_319,N_1487);
nand U1711 (N_1711,N_910,N_1388);
or U1712 (N_1712,N_596,N_523);
xor U1713 (N_1713,N_176,N_1381);
nor U1714 (N_1714,N_1485,In_1589);
and U1715 (N_1715,N_1353,In_536);
xnor U1716 (N_1716,N_958,In_2371);
or U1717 (N_1717,N_1215,N_249);
nor U1718 (N_1718,N_266,N_655);
and U1719 (N_1719,N_1323,N_1211);
or U1720 (N_1720,N_1227,N_1430);
and U1721 (N_1721,N_552,In_1872);
nand U1722 (N_1722,N_1362,N_1097);
nor U1723 (N_1723,N_1131,N_1102);
nand U1724 (N_1724,In_1929,N_1093);
or U1725 (N_1725,N_1382,N_623);
xor U1726 (N_1726,N_1560,N_1441);
nand U1727 (N_1727,N_241,In_1864);
nor U1728 (N_1728,N_918,In_309);
or U1729 (N_1729,N_293,In_1452);
nor U1730 (N_1730,N_1112,N_1262);
and U1731 (N_1731,N_453,In_705);
or U1732 (N_1732,In_1314,N_1013);
xor U1733 (N_1733,In_461,N_251);
xor U1734 (N_1734,In_2440,N_902);
xnor U1735 (N_1735,In_699,In_534);
or U1736 (N_1736,N_26,N_1498);
nor U1737 (N_1737,N_1172,In_468);
nor U1738 (N_1738,In_1482,N_1414);
or U1739 (N_1739,In_437,In_1910);
and U1740 (N_1740,N_1449,N_720);
nor U1741 (N_1741,In_1913,N_1259);
and U1742 (N_1742,N_331,In_254);
xnor U1743 (N_1743,N_1574,N_1141);
and U1744 (N_1744,In_2460,N_1219);
or U1745 (N_1745,In_297,N_1488);
and U1746 (N_1746,N_849,In_140);
or U1747 (N_1747,In_551,In_1067);
or U1748 (N_1748,N_1297,N_1416);
nand U1749 (N_1749,N_1489,N_1078);
nand U1750 (N_1750,N_1425,N_1436);
and U1751 (N_1751,In_1624,N_1077);
and U1752 (N_1752,In_2400,N_1076);
xor U1753 (N_1753,In_2121,N_1394);
or U1754 (N_1754,N_1525,N_891);
nor U1755 (N_1755,N_1239,N_1512);
and U1756 (N_1756,In_1229,N_1121);
and U1757 (N_1757,N_1163,In_1360);
xnor U1758 (N_1758,N_1179,In_237);
nand U1759 (N_1759,In_722,N_994);
nor U1760 (N_1760,N_1463,N_1391);
and U1761 (N_1761,N_912,N_896);
nand U1762 (N_1762,N_1464,N_1290);
xnor U1763 (N_1763,N_1281,N_1263);
and U1764 (N_1764,In_1365,N_1579);
xnor U1765 (N_1765,N_770,N_726);
or U1766 (N_1766,In_1088,N_1171);
xor U1767 (N_1767,N_187,In_1096);
nor U1768 (N_1768,N_999,N_558);
nor U1769 (N_1769,N_1023,In_185);
xnor U1770 (N_1770,N_198,N_1273);
or U1771 (N_1771,N_779,N_1364);
xor U1772 (N_1772,In_2006,N_1522);
and U1773 (N_1773,In_1653,In_1385);
xnor U1774 (N_1774,N_972,In_123);
nor U1775 (N_1775,In_1288,N_1011);
nor U1776 (N_1776,N_587,N_1493);
nor U1777 (N_1777,N_705,In_1512);
nor U1778 (N_1778,N_646,In_502);
and U1779 (N_1779,N_1470,N_865);
nor U1780 (N_1780,In_1629,N_1310);
nor U1781 (N_1781,N_1479,N_917);
and U1782 (N_1782,In_2434,N_1370);
or U1783 (N_1783,In_1232,N_1186);
and U1784 (N_1784,N_1468,N_683);
and U1785 (N_1785,N_1530,N_888);
nor U1786 (N_1786,In_518,In_1546);
nand U1787 (N_1787,N_1501,In_63);
xnor U1788 (N_1788,N_1307,N_1562);
and U1789 (N_1789,N_767,In_1483);
nor U1790 (N_1790,In_67,N_1429);
and U1791 (N_1791,N_1299,N_1400);
nor U1792 (N_1792,N_1197,In_1459);
and U1793 (N_1793,In_872,In_289);
nand U1794 (N_1794,N_1107,N_1082);
and U1795 (N_1795,In_338,N_1159);
nor U1796 (N_1796,N_998,N_522);
nor U1797 (N_1797,N_247,In_339);
nor U1798 (N_1798,N_1473,N_992);
or U1799 (N_1799,N_1339,In_2271);
xnor U1800 (N_1800,In_1303,N_1606);
or U1801 (N_1801,N_1036,N_1417);
nor U1802 (N_1802,In_2071,N_1035);
xor U1803 (N_1803,In_1836,N_1374);
nor U1804 (N_1804,N_563,N_1603);
nand U1805 (N_1805,In_476,N_1040);
and U1806 (N_1806,N_1667,N_1571);
nand U1807 (N_1807,N_812,N_1216);
or U1808 (N_1808,N_1589,N_1306);
and U1809 (N_1809,N_142,N_1647);
nand U1810 (N_1810,N_611,N_1696);
or U1811 (N_1811,N_1587,N_1779);
xnor U1812 (N_1812,N_859,N_1744);
nor U1813 (N_1813,N_1198,In_2199);
and U1814 (N_1814,N_1255,In_1603);
or U1815 (N_1815,In_648,N_709);
or U1816 (N_1816,N_1615,N_1786);
xnor U1817 (N_1817,N_1480,N_37);
nand U1818 (N_1818,N_1474,N_1446);
nor U1819 (N_1819,N_1221,N_966);
xnor U1820 (N_1820,N_125,N_1665);
nand U1821 (N_1821,N_1661,N_222);
or U1822 (N_1822,N_928,N_1798);
nor U1823 (N_1823,N_1234,In_1774);
xor U1824 (N_1824,N_837,N_788);
nand U1825 (N_1825,In_1725,N_1720);
and U1826 (N_1826,N_1413,N_1772);
and U1827 (N_1827,N_1286,N_1444);
and U1828 (N_1828,N_1751,N_1502);
nand U1829 (N_1829,N_1151,N_530);
or U1830 (N_1830,In_519,N_1465);
or U1831 (N_1831,N_1233,N_190);
nand U1832 (N_1832,N_1723,N_1653);
nand U1833 (N_1833,N_538,N_1017);
or U1834 (N_1834,N_1686,N_1592);
xor U1835 (N_1835,N_1202,In_2155);
nor U1836 (N_1836,N_536,N_1224);
xnor U1837 (N_1837,N_98,N_1642);
xor U1838 (N_1838,In_373,N_1762);
and U1839 (N_1839,N_1419,In_300);
xor U1840 (N_1840,N_1466,N_12);
and U1841 (N_1841,In_636,N_1699);
nand U1842 (N_1842,In_491,N_1614);
or U1843 (N_1843,N_526,N_1640);
or U1844 (N_1844,N_1795,N_1666);
nand U1845 (N_1845,N_1537,N_1355);
nor U1846 (N_1846,In_408,N_735);
or U1847 (N_1847,N_1684,N_840);
xnor U1848 (N_1848,N_279,N_694);
nand U1849 (N_1849,N_652,N_1203);
and U1850 (N_1850,N_23,N_1427);
and U1851 (N_1851,In_223,N_281);
and U1852 (N_1852,N_1645,N_1351);
nand U1853 (N_1853,N_1494,N_1208);
xnor U1854 (N_1854,N_1453,In_938);
nor U1855 (N_1855,N_1490,In_1494);
nand U1856 (N_1856,N_1283,N_85);
or U1857 (N_1857,N_1680,N_1520);
nor U1858 (N_1858,N_1278,N_1657);
and U1859 (N_1859,In_1611,N_1691);
xor U1860 (N_1860,N_1176,N_1655);
or U1861 (N_1861,In_671,N_1499);
nor U1862 (N_1862,N_156,In_1981);
xor U1863 (N_1863,N_1697,In_1837);
xnor U1864 (N_1864,N_1672,N_1752);
xor U1865 (N_1865,N_1618,In_1705);
and U1866 (N_1866,N_1710,In_891);
nor U1867 (N_1867,In_1646,In_1702);
xor U1868 (N_1868,N_1608,N_1718);
nor U1869 (N_1869,N_1616,N_1230);
and U1870 (N_1870,N_1624,In_1368);
xnor U1871 (N_1871,N_1566,N_1379);
and U1872 (N_1872,In_1500,In_200);
nand U1873 (N_1873,In_252,N_1643);
nor U1874 (N_1874,N_1738,N_1641);
or U1875 (N_1875,N_1707,N_1044);
nor U1876 (N_1876,N_1637,N_1226);
or U1877 (N_1877,N_1122,N_1009);
xor U1878 (N_1878,In_1334,N_1717);
nor U1879 (N_1879,N_1713,N_1782);
and U1880 (N_1880,N_1242,N_1621);
nor U1881 (N_1881,N_1475,N_1698);
and U1882 (N_1882,N_1787,N_163);
nor U1883 (N_1883,N_1767,N_1764);
and U1884 (N_1884,In_1903,N_1312);
nor U1885 (N_1885,In_909,In_341);
nand U1886 (N_1886,N_968,N_1634);
or U1887 (N_1887,N_763,N_1701);
xnor U1888 (N_1888,N_1220,N_922);
nand U1889 (N_1889,N_1638,N_1758);
nand U1890 (N_1890,N_1741,N_1617);
or U1891 (N_1891,N_1797,N_1542);
xor U1892 (N_1892,N_1704,N_1687);
or U1893 (N_1893,In_2436,N_1646);
xor U1894 (N_1894,N_1442,N_1314);
or U1895 (N_1895,In_881,N_1399);
or U1896 (N_1896,N_1648,N_1763);
nor U1897 (N_1897,N_564,N_1714);
nand U1898 (N_1898,In_1676,N_1734);
xor U1899 (N_1899,N_1627,N_1724);
or U1900 (N_1900,In_2009,In_431);
nand U1901 (N_1901,In_2241,N_1222);
xnor U1902 (N_1902,N_1635,N_670);
nand U1903 (N_1903,In_1918,N_1675);
xnor U1904 (N_1904,N_1469,N_1334);
and U1905 (N_1905,N_1745,In_106);
nand U1906 (N_1906,N_914,N_815);
nand U1907 (N_1907,N_810,N_1789);
xnor U1908 (N_1908,N_1298,N_1165);
or U1909 (N_1909,In_912,N_1193);
xnor U1910 (N_1910,N_1674,In_1516);
nor U1911 (N_1911,N_539,N_1098);
and U1912 (N_1912,N_1357,N_1067);
xor U1913 (N_1913,N_1625,In_2331);
and U1914 (N_1914,In_327,In_697);
and U1915 (N_1915,N_884,N_1578);
and U1916 (N_1916,N_1412,N_1735);
and U1917 (N_1917,N_1658,N_730);
xor U1918 (N_1918,In_2310,N_1683);
nor U1919 (N_1919,N_795,N_1557);
xor U1920 (N_1920,In_2441,N_916);
nand U1921 (N_1921,N_766,N_692);
nand U1922 (N_1922,N_1768,In_2254);
xor U1923 (N_1923,N_1459,N_1728);
nor U1924 (N_1924,N_1792,N_1725);
nand U1925 (N_1925,N_1521,N_1418);
nand U1926 (N_1926,N_882,N_1731);
nand U1927 (N_1927,N_1507,In_2053);
and U1928 (N_1928,N_1318,In_841);
xnor U1929 (N_1929,N_1229,N_1660);
or U1930 (N_1930,In_231,In_1432);
and U1931 (N_1931,In_211,In_2035);
or U1932 (N_1932,N_1670,N_1212);
nor U1933 (N_1933,In_1240,N_913);
nor U1934 (N_1934,N_816,In_615);
nand U1935 (N_1935,N_345,N_1730);
xnor U1936 (N_1936,N_1561,In_830);
or U1937 (N_1937,N_1240,N_1060);
nor U1938 (N_1938,N_1599,N_1799);
and U1939 (N_1939,N_1305,In_1979);
nand U1940 (N_1940,In_233,N_391);
xor U1941 (N_1941,N_1777,N_1457);
nand U1942 (N_1942,N_1437,In_1130);
nand U1943 (N_1943,In_1002,N_615);
xor U1944 (N_1944,N_1788,N_1721);
nand U1945 (N_1945,N_1746,N_1662);
and U1946 (N_1946,N_1583,N_1668);
or U1947 (N_1947,N_1631,N_1341);
and U1948 (N_1948,In_560,In_971);
xnor U1949 (N_1949,N_1059,In_330);
nor U1950 (N_1950,N_1620,N_820);
nor U1951 (N_1951,N_1411,N_1184);
and U1952 (N_1952,N_1517,In_855);
or U1953 (N_1953,N_1628,N_315);
and U1954 (N_1954,N_1380,N_1545);
nor U1955 (N_1955,N_1705,N_1232);
nand U1956 (N_1956,N_1595,N_1604);
nand U1957 (N_1957,N_640,N_1047);
nand U1958 (N_1958,N_1373,N_299);
and U1959 (N_1959,N_1626,N_301);
nand U1960 (N_1960,In_907,In_1867);
xnor U1961 (N_1961,N_138,N_1293);
xor U1962 (N_1962,N_1739,N_1692);
and U1963 (N_1963,N_657,In_1806);
or U1964 (N_1964,N_1775,N_1630);
nand U1965 (N_1965,In_1937,N_1477);
nor U1966 (N_1966,N_1563,N_1689);
and U1967 (N_1967,N_1773,In_1532);
nor U1968 (N_1968,N_1765,In_2463);
nor U1969 (N_1969,N_1770,In_702);
or U1970 (N_1970,N_1729,N_443);
nand U1971 (N_1971,N_1650,N_988);
and U1972 (N_1972,In_2193,In_998);
xnor U1973 (N_1973,N_1551,N_1423);
nor U1974 (N_1974,N_637,N_732);
nand U1975 (N_1975,N_1527,N_1693);
and U1976 (N_1976,N_1407,In_227);
xor U1977 (N_1977,In_1776,N_1553);
or U1978 (N_1978,N_1633,N_1245);
and U1979 (N_1979,In_151,N_1656);
nand U1980 (N_1980,In_215,N_1510);
or U1981 (N_1981,N_1565,In_890);
nor U1982 (N_1982,N_1644,N_1622);
nand U1983 (N_1983,N_1607,N_1376);
xor U1984 (N_1984,In_870,In_150);
nor U1985 (N_1985,N_1456,N_1130);
nor U1986 (N_1986,N_1639,N_1448);
and U1987 (N_1987,N_824,N_212);
xnor U1988 (N_1988,In_1767,N_1092);
or U1989 (N_1989,N_1708,N_325);
nand U1990 (N_1990,N_1612,N_1733);
xor U1991 (N_1991,N_571,N_791);
nor U1992 (N_1992,In_825,N_1580);
xnor U1993 (N_1993,N_554,N_1554);
xnor U1994 (N_1994,N_1700,In_157);
nand U1995 (N_1995,N_1594,In_2029);
or U1996 (N_1996,N_1586,N_768);
or U1997 (N_1997,In_656,N_1420);
xnor U1998 (N_1998,N_618,N_1535);
and U1999 (N_1999,N_1451,N_393);
and U2000 (N_2000,N_452,N_1146);
nor U2001 (N_2001,In_1068,In_1678);
xor U2002 (N_2002,N_1544,N_1938);
nand U2003 (N_2003,N_1866,N_1671);
or U2004 (N_2004,N_1204,N_1859);
nor U2005 (N_2005,N_1596,N_1888);
nor U2006 (N_2006,In_1544,In_1407);
nand U2007 (N_2007,N_1847,N_1401);
and U2008 (N_2008,N_1022,In_715);
nor U2009 (N_2009,N_1939,N_1933);
nor U2010 (N_2010,N_1934,N_1891);
and U2011 (N_2011,N_1254,In_794);
nor U2012 (N_2012,N_449,N_1936);
xnor U2013 (N_2013,N_1965,N_1856);
nor U2014 (N_2014,N_1908,N_1890);
or U2015 (N_2015,In_2216,N_1766);
or U2016 (N_2016,N_1539,N_1840);
or U2017 (N_2017,N_1822,N_1998);
or U2018 (N_2018,N_1831,In_1479);
nand U2019 (N_2019,N_1966,In_490);
xnor U2020 (N_2020,In_2164,N_1445);
nand U2021 (N_2021,N_1947,N_1652);
or U2022 (N_2022,In_1932,N_1138);
or U2023 (N_2023,N_1711,N_1949);
nor U2024 (N_2024,In_1381,N_1855);
or U2025 (N_2025,N_1790,N_1793);
or U2026 (N_2026,N_1611,N_274);
xor U2027 (N_2027,N_719,In_866);
and U2028 (N_2028,N_1886,N_1367);
nand U2029 (N_2029,N_1761,In_584);
and U2030 (N_2030,N_158,N_1960);
and U2031 (N_2031,N_949,N_1774);
or U2032 (N_2032,N_1832,N_1778);
xor U2033 (N_2033,N_1781,N_1726);
nand U2034 (N_2034,N_1132,N_1256);
nor U2035 (N_2035,In_1503,N_1807);
nand U2036 (N_2036,N_1523,In_974);
nor U2037 (N_2037,N_1977,N_1944);
and U2038 (N_2038,N_1975,In_261);
or U2039 (N_2039,N_1932,N_1937);
xnor U2040 (N_2040,N_177,N_1065);
nand U2041 (N_2041,N_1796,N_1845);
xor U2042 (N_2042,N_1828,In_1026);
and U2043 (N_2043,N_245,N_1383);
or U2044 (N_2044,N_1552,In_139);
and U2045 (N_2045,N_1024,N_1999);
and U2046 (N_2046,In_961,N_1162);
nand U2047 (N_2047,In_1965,N_1988);
and U2048 (N_2048,N_257,N_1435);
and U2049 (N_2049,N_1804,N_1897);
and U2050 (N_2050,N_1830,N_983);
nand U2051 (N_2051,N_1712,N_1946);
and U2052 (N_2052,N_1740,N_1706);
or U2053 (N_2053,N_1870,N_1113);
or U2054 (N_2054,N_1732,N_45);
nor U2055 (N_2055,N_1540,N_1913);
and U2056 (N_2056,N_1421,N_1875);
or U2057 (N_2057,N_1743,N_1943);
xnor U2058 (N_2058,N_1716,N_1538);
nand U2059 (N_2059,N_1702,N_1901);
xor U2060 (N_2060,N_1970,In_2376);
or U2061 (N_2061,N_1906,N_1504);
nor U2062 (N_2062,N_1905,N_1899);
and U2063 (N_2063,N_1907,N_978);
xor U2064 (N_2064,N_1747,N_1818);
xor U2065 (N_2065,N_1837,N_1824);
or U2066 (N_2066,N_920,In_82);
nor U2067 (N_2067,N_1887,N_1500);
nor U2068 (N_2068,N_392,N_1214);
xor U2069 (N_2069,N_688,N_1058);
or U2070 (N_2070,N_1568,N_1750);
nand U2071 (N_2071,N_1894,In_363);
nor U2072 (N_2072,N_1651,In_499);
nor U2073 (N_2073,N_1016,N_1911);
and U2074 (N_2074,N_1609,In_882);
xnor U2075 (N_2075,N_1598,N_1995);
nand U2076 (N_2076,N_1195,N_1514);
and U2077 (N_2077,N_1902,N_1935);
or U2078 (N_2078,N_1467,In_38);
and U2079 (N_2079,In_1291,N_1841);
nor U2080 (N_2080,N_1450,N_1991);
xnor U2081 (N_2081,N_1629,N_1816);
or U2082 (N_2082,N_313,In_2449);
nor U2083 (N_2083,In_1775,N_1685);
nor U2084 (N_2084,N_1989,N_1885);
xor U2085 (N_2085,N_1930,N_1835);
nor U2086 (N_2086,N_1813,N_1590);
xnor U2087 (N_2087,N_857,N_1957);
nand U2088 (N_2088,N_1408,N_1812);
xor U2089 (N_2089,N_1839,N_1868);
nand U2090 (N_2090,N_1187,N_1981);
nand U2091 (N_2091,N_1690,In_268);
nor U2092 (N_2092,N_1344,In_1710);
nand U2093 (N_2093,N_1111,N_1664);
xnor U2094 (N_2094,N_557,N_1426);
nor U2095 (N_2095,In_1390,N_36);
nor U2096 (N_2096,N_1889,N_1844);
nor U2097 (N_2097,N_1914,N_1783);
xnor U2098 (N_2098,N_1094,N_938);
nand U2099 (N_2099,N_304,N_1958);
nand U2100 (N_2100,N_1994,N_1964);
nor U2101 (N_2101,In_2349,N_1878);
nand U2102 (N_2102,N_1967,N_1827);
nor U2103 (N_2103,N_1271,N_1452);
xor U2104 (N_2104,N_1857,N_1703);
xor U2105 (N_2105,N_1505,N_1916);
and U2106 (N_2106,N_1140,N_1753);
xnor U2107 (N_2107,N_1742,In_2003);
nand U2108 (N_2108,N_1834,N_1189);
or U2109 (N_2109,N_1759,N_519);
and U2110 (N_2110,N_1926,N_1313);
nor U2111 (N_2111,N_1582,N_1694);
or U2112 (N_2112,N_1810,In_47);
nor U2113 (N_2113,In_1070,N_1973);
nor U2114 (N_2114,N_858,N_1748);
or U2115 (N_2115,In_1359,N_1969);
nand U2116 (N_2116,In_960,N_1982);
nor U2117 (N_2117,N_1678,N_1404);
nor U2118 (N_2118,N_1987,N_542);
or U2119 (N_2119,N_1867,N_866);
or U2120 (N_2120,N_1601,N_1854);
nor U2121 (N_2121,N_943,N_1385);
nand U2122 (N_2122,N_1996,N_1923);
or U2123 (N_2123,N_1941,N_401);
nand U2124 (N_2124,N_1821,N_133);
and U2125 (N_2125,N_1267,N_1838);
nand U2126 (N_2126,N_1600,N_1925);
or U2127 (N_2127,N_1863,N_1952);
and U2128 (N_2128,N_1492,N_1336);
nand U2129 (N_2129,N_1993,N_1909);
xor U2130 (N_2130,N_1066,N_1757);
and U2131 (N_2131,N_1188,N_1410);
and U2132 (N_2132,N_1532,N_1237);
nor U2133 (N_2133,N_915,N_1303);
and U2134 (N_2134,N_1727,N_1971);
and U2135 (N_2135,N_1928,N_1917);
and U2136 (N_2136,N_1858,N_1846);
nor U2137 (N_2137,N_321,N_1681);
or U2138 (N_2138,N_1968,N_1892);
nor U2139 (N_2139,N_1850,N_1673);
nand U2140 (N_2140,In_1477,N_1861);
nand U2141 (N_2141,N_1688,N_1048);
and U2142 (N_2142,N_1801,N_1200);
nand U2143 (N_2143,N_1415,N_1910);
nor U2144 (N_2144,N_844,N_1871);
nor U2145 (N_2145,N_1983,N_1980);
and U2146 (N_2146,N_1806,N_1819);
nor U2147 (N_2147,N_1929,In_772);
and U2148 (N_2148,N_1884,In_1548);
xor U2149 (N_2149,N_1371,N_1942);
nor U2150 (N_2150,N_1869,N_930);
and U2151 (N_2151,N_1719,N_1862);
xnor U2152 (N_2152,N_1803,N_1940);
nand U2153 (N_2153,N_1541,N_1755);
nand U2154 (N_2154,N_1881,N_1715);
nor U2155 (N_2155,N_1842,N_1191);
nor U2156 (N_2156,N_1814,N_1985);
or U2157 (N_2157,N_1922,N_1476);
nor U2158 (N_2158,N_1074,N_1992);
and U2159 (N_2159,N_1826,N_1516);
and U2160 (N_2160,N_1882,N_1919);
xnor U2161 (N_2161,N_1809,N_1860);
and U2162 (N_2162,N_1760,N_1695);
xnor U2163 (N_2163,N_1776,N_1529);
nand U2164 (N_2164,In_557,N_1403);
xor U2165 (N_2165,N_1924,N_1900);
xnor U2166 (N_2166,N_1447,N_1811);
and U2167 (N_2167,N_310,N_1780);
and U2168 (N_2168,N_1873,N_1984);
nand U2169 (N_2169,N_1679,N_1997);
nor U2170 (N_2170,N_1559,N_1785);
nor U2171 (N_2171,N_1823,N_1808);
nor U2172 (N_2172,N_1883,N_1663);
nand U2173 (N_2173,N_1976,N_152);
nor U2174 (N_2174,N_1153,N_1613);
or U2175 (N_2175,N_1879,N_1577);
xor U2176 (N_2176,N_410,N_1495);
nor U2177 (N_2177,N_1053,N_841);
nor U2178 (N_2178,N_1986,N_1676);
or U2179 (N_2179,N_1659,N_1853);
or U2180 (N_2180,N_1948,N_83);
xor U2181 (N_2181,In_1356,N_1945);
nand U2182 (N_2182,N_751,N_1864);
and U2183 (N_2183,N_738,N_1117);
and U2184 (N_2184,N_1486,N_1619);
or U2185 (N_2185,N_1843,N_1794);
nor U2186 (N_2186,In_2004,N_1722);
xnor U2187 (N_2187,N_1954,N_1896);
nand U2188 (N_2188,N_129,N_1428);
and U2189 (N_2189,In_2461,N_1012);
nor U2190 (N_2190,N_1800,N_1865);
nand U2191 (N_2191,In_61,N_1820);
and U2192 (N_2192,N_982,N_1511);
xnor U2193 (N_2193,N_1567,N_1669);
xor U2194 (N_2194,N_1972,N_1955);
nor U2195 (N_2195,N_541,N_1877);
and U2196 (N_2196,N_1805,N_1294);
and U2197 (N_2197,N_1956,N_1769);
and U2198 (N_2198,N_1295,N_1974);
or U2199 (N_2199,N_1962,N_1895);
xnor U2200 (N_2200,N_2115,N_1311);
or U2201 (N_2201,N_2063,N_1330);
nand U2202 (N_2202,N_1872,N_2000);
xnor U2203 (N_2203,N_1265,N_2023);
xor U2204 (N_2204,N_2021,N_2102);
nand U2205 (N_2205,N_2038,N_2147);
nor U2206 (N_2206,N_2031,N_1749);
nor U2207 (N_2207,N_2174,N_2129);
and U2208 (N_2208,N_2032,N_2026);
nor U2209 (N_2209,N_2166,N_2035);
nand U2210 (N_2210,N_1990,N_2022);
or U2211 (N_2211,N_2168,N_1623);
nor U2212 (N_2212,N_2088,N_2016);
nand U2213 (N_2213,N_2110,N_2153);
nor U2214 (N_2214,N_2086,N_2082);
or U2215 (N_2215,N_2085,N_2101);
or U2216 (N_2216,N_1848,N_2078);
and U2217 (N_2217,N_2111,N_2064);
nor U2218 (N_2218,N_2199,N_1784);
xnor U2219 (N_2219,N_2036,N_427);
nand U2220 (N_2220,N_2161,N_1677);
or U2221 (N_2221,N_2155,N_1791);
or U2222 (N_2222,N_2178,N_323);
xnor U2223 (N_2223,N_2140,N_1101);
nor U2224 (N_2224,N_1325,N_1709);
xor U2225 (N_2225,N_2165,N_2027);
xor U2226 (N_2226,N_2141,N_1454);
or U2227 (N_2227,N_2044,N_2100);
or U2228 (N_2228,N_2003,N_2041);
nor U2229 (N_2229,N_2122,N_2107);
xor U2230 (N_2230,N_1963,N_2198);
or U2231 (N_2231,In_1525,N_2179);
or U2232 (N_2232,N_1534,N_2182);
nor U2233 (N_2233,In_2414,N_78);
xor U2234 (N_2234,N_2172,N_2113);
xor U2235 (N_2235,N_1506,N_1903);
nand U2236 (N_2236,N_1550,N_1756);
xor U2237 (N_2237,In_2330,N_2095);
or U2238 (N_2238,N_2049,N_1874);
or U2239 (N_2239,N_1953,N_1771);
nor U2240 (N_2240,N_2066,N_2145);
or U2241 (N_2241,N_1927,N_1126);
nor U2242 (N_2242,N_2152,N_2005);
and U2243 (N_2243,N_2008,N_2159);
nor U2244 (N_2244,N_1136,N_2099);
nor U2245 (N_2245,N_1961,N_2014);
or U2246 (N_2246,N_2120,N_1978);
or U2247 (N_2247,N_1829,N_2181);
and U2248 (N_2248,N_2057,N_2185);
or U2249 (N_2249,N_2090,N_2163);
xnor U2250 (N_2250,N_2097,N_2013);
nand U2251 (N_2251,N_2071,N_2029);
and U2252 (N_2252,N_2131,N_2191);
nor U2253 (N_2253,N_1632,N_1386);
and U2254 (N_2254,N_1959,N_2067);
xnor U2255 (N_2255,N_2127,N_2195);
nor U2256 (N_2256,N_1375,N_2083);
nand U2257 (N_2257,N_1533,N_2070);
or U2258 (N_2258,N_2184,N_2076);
or U2259 (N_2259,N_1555,N_2092);
or U2260 (N_2260,N_1920,N_2148);
nor U2261 (N_2261,N_2108,In_1800);
nor U2262 (N_2262,N_2059,N_2117);
nand U2263 (N_2263,N_2137,N_2146);
nor U2264 (N_2264,N_2080,N_2012);
and U2265 (N_2265,N_2024,N_1817);
or U2266 (N_2266,N_2010,In_1275);
nor U2267 (N_2267,N_1904,N_1503);
xor U2268 (N_2268,N_2170,N_2156);
nand U2269 (N_2269,N_2134,N_2048);
nand U2270 (N_2270,N_1654,N_2173);
and U2271 (N_2271,N_2002,N_2125);
nand U2272 (N_2272,N_1921,N_1849);
xor U2273 (N_2273,N_1422,N_1852);
nor U2274 (N_2274,N_2052,N_793);
and U2275 (N_2275,N_2054,N_2194);
xor U2276 (N_2276,In_1440,N_1893);
and U2277 (N_2277,N_2196,N_2087);
and U2278 (N_2278,In_1737,N_1836);
nor U2279 (N_2279,N_2158,N_2039);
xor U2280 (N_2280,N_2160,N_2142);
xnor U2281 (N_2281,N_1605,N_2190);
nand U2282 (N_2282,N_1912,N_2116);
nand U2283 (N_2283,N_1754,N_1610);
or U2284 (N_2284,N_1880,N_2043);
nor U2285 (N_2285,N_2004,N_2069);
nor U2286 (N_2286,N_1815,N_2033);
nand U2287 (N_2287,N_1915,N_654);
or U2288 (N_2288,N_2094,N_2068);
nand U2289 (N_2289,N_2167,N_2074);
or U2290 (N_2290,N_2180,N_2042);
and U2291 (N_2291,N_1257,N_2109);
xor U2292 (N_2292,N_1069,N_2055);
nor U2293 (N_2293,N_2188,N_2053);
nand U2294 (N_2294,N_2025,N_1261);
nand U2295 (N_2295,N_2130,N_2015);
and U2296 (N_2296,N_1302,N_2034);
nor U2297 (N_2297,N_1682,N_1398);
nand U2298 (N_2298,N_2135,N_2132);
nand U2299 (N_2299,N_2192,N_2175);
nor U2300 (N_2300,In_1072,N_2126);
xnor U2301 (N_2301,N_2123,N_629);
nand U2302 (N_2302,N_2164,N_2128);
or U2303 (N_2303,N_1602,N_2058);
xnor U2304 (N_2304,In_1614,N_2112);
nand U2305 (N_2305,N_2103,N_2119);
or U2306 (N_2306,N_2060,N_2183);
or U2307 (N_2307,N_2037,N_2124);
nor U2308 (N_2308,N_2084,N_1876);
nand U2309 (N_2309,N_1389,N_2187);
or U2310 (N_2310,N_2193,N_2093);
xor U2311 (N_2311,N_2091,N_2075);
nand U2312 (N_2312,N_1851,N_2020);
and U2313 (N_2313,N_2089,N_2143);
xnor U2314 (N_2314,N_2157,N_1472);
nor U2315 (N_2315,N_739,N_2162);
nand U2316 (N_2316,N_2050,N_2062);
xor U2317 (N_2317,N_1950,N_2006);
nor U2318 (N_2318,N_2045,N_2073);
xor U2319 (N_2319,N_2104,N_2098);
nand U2320 (N_2320,N_2149,In_1625);
or U2321 (N_2321,N_802,N_2154);
or U2322 (N_2322,N_2011,N_2065);
xnor U2323 (N_2323,N_2176,N_2056);
nand U2324 (N_2324,N_2138,N_2030);
xor U2325 (N_2325,N_2114,N_2061);
xnor U2326 (N_2326,N_2105,N_2072);
or U2327 (N_2327,N_2139,N_1918);
and U2328 (N_2328,N_1979,N_2136);
or U2329 (N_2329,N_2144,N_2189);
or U2330 (N_2330,N_2019,N_2009);
nand U2331 (N_2331,N_1636,N_1833);
or U2332 (N_2332,N_2051,N_2040);
nand U2333 (N_2333,N_2169,N_1931);
and U2334 (N_2334,N_2007,N_1406);
and U2335 (N_2335,N_2106,N_2079);
xnor U2336 (N_2336,N_2047,N_1649);
nor U2337 (N_2337,N_2077,N_1737);
xnor U2338 (N_2338,N_1898,N_2096);
or U2339 (N_2339,N_2118,N_2028);
nor U2340 (N_2340,N_2197,N_2017);
and U2341 (N_2341,N_2081,N_2133);
or U2342 (N_2342,N_2018,N_2186);
xnor U2343 (N_2343,N_1825,N_1736);
nor U2344 (N_2344,N_1951,N_2001);
nand U2345 (N_2345,In_1809,N_2151);
nor U2346 (N_2346,N_2121,In_1794);
xnor U2347 (N_2347,N_2171,In_2395);
nor U2348 (N_2348,N_2150,N_2177);
nor U2349 (N_2349,N_1802,N_2046);
nor U2350 (N_2350,N_2076,In_1614);
and U2351 (N_2351,N_2059,N_2102);
nand U2352 (N_2352,N_1898,N_2130);
nand U2353 (N_2353,N_1829,N_2117);
or U2354 (N_2354,N_2124,N_2170);
nor U2355 (N_2355,N_2115,N_2125);
or U2356 (N_2356,N_2021,N_2023);
xor U2357 (N_2357,N_2030,N_2097);
and U2358 (N_2358,N_2030,N_2096);
or U2359 (N_2359,N_2121,N_2037);
nor U2360 (N_2360,N_2056,N_1872);
xor U2361 (N_2361,N_1602,N_1904);
xor U2362 (N_2362,N_2160,N_2096);
xor U2363 (N_2363,N_2109,N_2010);
nor U2364 (N_2364,N_2197,N_2077);
nand U2365 (N_2365,N_2172,N_1506);
nor U2366 (N_2366,N_2045,N_2054);
nor U2367 (N_2367,N_2001,N_2107);
and U2368 (N_2368,N_2094,N_1636);
nand U2369 (N_2369,N_2099,N_427);
nor U2370 (N_2370,N_2078,N_2004);
nor U2371 (N_2371,N_2014,N_1848);
xor U2372 (N_2372,N_2032,N_1915);
or U2373 (N_2373,N_2005,N_739);
nor U2374 (N_2374,N_1961,N_1610);
nand U2375 (N_2375,N_1330,N_2139);
nor U2376 (N_2376,N_2133,N_2030);
nand U2377 (N_2377,N_2169,N_2039);
nand U2378 (N_2378,N_2021,N_2072);
and U2379 (N_2379,N_1649,N_1636);
nand U2380 (N_2380,N_1880,N_2113);
nor U2381 (N_2381,N_1963,N_2150);
and U2382 (N_2382,N_1654,N_1951);
nor U2383 (N_2383,N_2085,N_2075);
xor U2384 (N_2384,N_1709,N_2048);
nor U2385 (N_2385,N_2180,N_2000);
nand U2386 (N_2386,N_2073,N_1912);
xnor U2387 (N_2387,N_2164,N_2013);
or U2388 (N_2388,N_2109,N_2058);
or U2389 (N_2389,N_739,N_2107);
or U2390 (N_2390,N_2173,N_1605);
nor U2391 (N_2391,N_2081,In_1440);
nand U2392 (N_2392,N_2050,N_2160);
and U2393 (N_2393,N_1682,N_2085);
nand U2394 (N_2394,In_1625,N_2043);
and U2395 (N_2395,N_2165,N_2049);
or U2396 (N_2396,N_2029,N_2074);
xnor U2397 (N_2397,N_2174,N_2167);
xnor U2398 (N_2398,N_2029,N_2105);
or U2399 (N_2399,N_1302,N_2194);
nor U2400 (N_2400,N_2396,N_2296);
nand U2401 (N_2401,N_2287,N_2248);
nor U2402 (N_2402,N_2315,N_2355);
nor U2403 (N_2403,N_2346,N_2395);
xor U2404 (N_2404,N_2292,N_2399);
xor U2405 (N_2405,N_2358,N_2232);
nor U2406 (N_2406,N_2290,N_2328);
nand U2407 (N_2407,N_2392,N_2370);
nor U2408 (N_2408,N_2271,N_2238);
xnor U2409 (N_2409,N_2249,N_2230);
xor U2410 (N_2410,N_2326,N_2267);
nor U2411 (N_2411,N_2211,N_2217);
or U2412 (N_2412,N_2372,N_2240);
or U2413 (N_2413,N_2378,N_2377);
nor U2414 (N_2414,N_2288,N_2386);
nor U2415 (N_2415,N_2255,N_2317);
nand U2416 (N_2416,N_2283,N_2269);
nor U2417 (N_2417,N_2209,N_2339);
or U2418 (N_2418,N_2345,N_2273);
xnor U2419 (N_2419,N_2384,N_2254);
nand U2420 (N_2420,N_2264,N_2281);
nor U2421 (N_2421,N_2237,N_2272);
xnor U2422 (N_2422,N_2352,N_2329);
and U2423 (N_2423,N_2213,N_2261);
xnor U2424 (N_2424,N_2312,N_2349);
and U2425 (N_2425,N_2212,N_2245);
and U2426 (N_2426,N_2357,N_2375);
xor U2427 (N_2427,N_2222,N_2298);
nand U2428 (N_2428,N_2311,N_2233);
and U2429 (N_2429,N_2360,N_2201);
or U2430 (N_2430,N_2369,N_2314);
nor U2431 (N_2431,N_2323,N_2258);
nand U2432 (N_2432,N_2389,N_2259);
and U2433 (N_2433,N_2330,N_2205);
nor U2434 (N_2434,N_2341,N_2268);
xnor U2435 (N_2435,N_2342,N_2282);
nand U2436 (N_2436,N_2313,N_2367);
and U2437 (N_2437,N_2320,N_2302);
nand U2438 (N_2438,N_2241,N_2231);
nand U2439 (N_2439,N_2291,N_2277);
xnor U2440 (N_2440,N_2351,N_2293);
xnor U2441 (N_2441,N_2280,N_2247);
nand U2442 (N_2442,N_2274,N_2356);
xor U2443 (N_2443,N_2295,N_2206);
nand U2444 (N_2444,N_2361,N_2340);
or U2445 (N_2445,N_2275,N_2307);
xor U2446 (N_2446,N_2327,N_2348);
or U2447 (N_2447,N_2236,N_2229);
nor U2448 (N_2448,N_2368,N_2344);
nand U2449 (N_2449,N_2226,N_2353);
nand U2450 (N_2450,N_2242,N_2391);
or U2451 (N_2451,N_2303,N_2397);
nor U2452 (N_2452,N_2207,N_2208);
xor U2453 (N_2453,N_2221,N_2239);
nor U2454 (N_2454,N_2252,N_2336);
xor U2455 (N_2455,N_2214,N_2362);
nor U2456 (N_2456,N_2376,N_2289);
and U2457 (N_2457,N_2380,N_2322);
nor U2458 (N_2458,N_2219,N_2347);
xor U2459 (N_2459,N_2210,N_2363);
xor U2460 (N_2460,N_2260,N_2334);
nor U2461 (N_2461,N_2308,N_2265);
nand U2462 (N_2462,N_2388,N_2337);
xnor U2463 (N_2463,N_2333,N_2263);
or U2464 (N_2464,N_2338,N_2227);
and U2465 (N_2465,N_2278,N_2216);
xnor U2466 (N_2466,N_2223,N_2343);
nand U2467 (N_2467,N_2256,N_2228);
xor U2468 (N_2468,N_2364,N_2203);
xnor U2469 (N_2469,N_2225,N_2262);
nand U2470 (N_2470,N_2306,N_2285);
xor U2471 (N_2471,N_2279,N_2276);
xor U2472 (N_2472,N_2266,N_2382);
nand U2473 (N_2473,N_2284,N_2332);
xnor U2474 (N_2474,N_2385,N_2359);
nand U2475 (N_2475,N_2253,N_2354);
or U2476 (N_2476,N_2390,N_2286);
nor U2477 (N_2477,N_2374,N_2250);
and U2478 (N_2478,N_2310,N_2202);
xor U2479 (N_2479,N_2299,N_2224);
and U2480 (N_2480,N_2251,N_2220);
nor U2481 (N_2481,N_2379,N_2204);
and U2482 (N_2482,N_2325,N_2383);
or U2483 (N_2483,N_2301,N_2319);
xnor U2484 (N_2484,N_2270,N_2294);
nand U2485 (N_2485,N_2331,N_2381);
nor U2486 (N_2486,N_2297,N_2387);
xor U2487 (N_2487,N_2304,N_2373);
or U2488 (N_2488,N_2324,N_2371);
nand U2489 (N_2489,N_2366,N_2394);
or U2490 (N_2490,N_2393,N_2235);
nand U2491 (N_2491,N_2316,N_2305);
nor U2492 (N_2492,N_2234,N_2200);
nand U2493 (N_2493,N_2215,N_2398);
or U2494 (N_2494,N_2243,N_2318);
nor U2495 (N_2495,N_2244,N_2350);
nand U2496 (N_2496,N_2321,N_2218);
and U2497 (N_2497,N_2300,N_2365);
nand U2498 (N_2498,N_2257,N_2335);
nor U2499 (N_2499,N_2246,N_2309);
and U2500 (N_2500,N_2282,N_2292);
nand U2501 (N_2501,N_2359,N_2322);
and U2502 (N_2502,N_2216,N_2281);
and U2503 (N_2503,N_2399,N_2283);
nor U2504 (N_2504,N_2361,N_2241);
or U2505 (N_2505,N_2226,N_2297);
nand U2506 (N_2506,N_2286,N_2253);
xor U2507 (N_2507,N_2269,N_2321);
and U2508 (N_2508,N_2378,N_2342);
and U2509 (N_2509,N_2261,N_2360);
or U2510 (N_2510,N_2244,N_2222);
xor U2511 (N_2511,N_2389,N_2368);
and U2512 (N_2512,N_2278,N_2315);
xnor U2513 (N_2513,N_2206,N_2331);
nor U2514 (N_2514,N_2389,N_2327);
or U2515 (N_2515,N_2398,N_2364);
or U2516 (N_2516,N_2347,N_2342);
nor U2517 (N_2517,N_2312,N_2251);
and U2518 (N_2518,N_2261,N_2254);
and U2519 (N_2519,N_2291,N_2397);
and U2520 (N_2520,N_2335,N_2266);
or U2521 (N_2521,N_2300,N_2302);
nor U2522 (N_2522,N_2315,N_2399);
or U2523 (N_2523,N_2387,N_2352);
and U2524 (N_2524,N_2390,N_2296);
and U2525 (N_2525,N_2251,N_2205);
xor U2526 (N_2526,N_2274,N_2201);
xor U2527 (N_2527,N_2363,N_2389);
nand U2528 (N_2528,N_2386,N_2295);
or U2529 (N_2529,N_2316,N_2360);
xnor U2530 (N_2530,N_2252,N_2306);
and U2531 (N_2531,N_2248,N_2358);
xor U2532 (N_2532,N_2331,N_2244);
nand U2533 (N_2533,N_2241,N_2330);
and U2534 (N_2534,N_2237,N_2275);
xor U2535 (N_2535,N_2267,N_2257);
nand U2536 (N_2536,N_2339,N_2207);
nand U2537 (N_2537,N_2230,N_2340);
nand U2538 (N_2538,N_2399,N_2243);
nor U2539 (N_2539,N_2256,N_2206);
and U2540 (N_2540,N_2388,N_2287);
nor U2541 (N_2541,N_2266,N_2237);
xnor U2542 (N_2542,N_2377,N_2362);
and U2543 (N_2543,N_2226,N_2323);
xor U2544 (N_2544,N_2328,N_2315);
nor U2545 (N_2545,N_2259,N_2213);
nor U2546 (N_2546,N_2303,N_2302);
xnor U2547 (N_2547,N_2210,N_2293);
or U2548 (N_2548,N_2297,N_2262);
and U2549 (N_2549,N_2228,N_2274);
xor U2550 (N_2550,N_2342,N_2224);
or U2551 (N_2551,N_2293,N_2284);
nand U2552 (N_2552,N_2237,N_2239);
or U2553 (N_2553,N_2273,N_2282);
or U2554 (N_2554,N_2329,N_2345);
and U2555 (N_2555,N_2371,N_2206);
nor U2556 (N_2556,N_2269,N_2383);
xor U2557 (N_2557,N_2257,N_2352);
and U2558 (N_2558,N_2361,N_2369);
and U2559 (N_2559,N_2288,N_2392);
xnor U2560 (N_2560,N_2301,N_2254);
or U2561 (N_2561,N_2392,N_2218);
and U2562 (N_2562,N_2240,N_2262);
or U2563 (N_2563,N_2369,N_2306);
xor U2564 (N_2564,N_2298,N_2308);
nand U2565 (N_2565,N_2331,N_2376);
nand U2566 (N_2566,N_2359,N_2241);
and U2567 (N_2567,N_2272,N_2212);
nand U2568 (N_2568,N_2206,N_2250);
and U2569 (N_2569,N_2238,N_2381);
nor U2570 (N_2570,N_2206,N_2357);
and U2571 (N_2571,N_2316,N_2344);
xnor U2572 (N_2572,N_2220,N_2333);
and U2573 (N_2573,N_2350,N_2326);
xnor U2574 (N_2574,N_2385,N_2378);
nor U2575 (N_2575,N_2275,N_2319);
xnor U2576 (N_2576,N_2302,N_2398);
and U2577 (N_2577,N_2336,N_2266);
nor U2578 (N_2578,N_2203,N_2244);
nor U2579 (N_2579,N_2201,N_2209);
xor U2580 (N_2580,N_2381,N_2201);
and U2581 (N_2581,N_2202,N_2343);
nor U2582 (N_2582,N_2360,N_2330);
nor U2583 (N_2583,N_2375,N_2381);
and U2584 (N_2584,N_2331,N_2277);
xnor U2585 (N_2585,N_2203,N_2390);
xnor U2586 (N_2586,N_2257,N_2309);
and U2587 (N_2587,N_2391,N_2219);
nand U2588 (N_2588,N_2333,N_2381);
and U2589 (N_2589,N_2220,N_2213);
xnor U2590 (N_2590,N_2268,N_2337);
nand U2591 (N_2591,N_2389,N_2387);
or U2592 (N_2592,N_2281,N_2299);
nor U2593 (N_2593,N_2369,N_2371);
xnor U2594 (N_2594,N_2344,N_2392);
nor U2595 (N_2595,N_2375,N_2212);
nor U2596 (N_2596,N_2224,N_2228);
and U2597 (N_2597,N_2365,N_2243);
nand U2598 (N_2598,N_2328,N_2296);
or U2599 (N_2599,N_2202,N_2213);
nand U2600 (N_2600,N_2427,N_2546);
and U2601 (N_2601,N_2491,N_2529);
nand U2602 (N_2602,N_2583,N_2516);
nor U2603 (N_2603,N_2597,N_2480);
or U2604 (N_2604,N_2547,N_2488);
and U2605 (N_2605,N_2543,N_2486);
and U2606 (N_2606,N_2587,N_2420);
or U2607 (N_2607,N_2471,N_2461);
nand U2608 (N_2608,N_2441,N_2492);
or U2609 (N_2609,N_2498,N_2426);
or U2610 (N_2610,N_2533,N_2428);
nor U2611 (N_2611,N_2515,N_2548);
and U2612 (N_2612,N_2410,N_2442);
or U2613 (N_2613,N_2477,N_2481);
nand U2614 (N_2614,N_2447,N_2485);
and U2615 (N_2615,N_2443,N_2556);
nand U2616 (N_2616,N_2408,N_2403);
nor U2617 (N_2617,N_2574,N_2592);
nor U2618 (N_2618,N_2568,N_2484);
or U2619 (N_2619,N_2490,N_2550);
nor U2620 (N_2620,N_2541,N_2584);
xor U2621 (N_2621,N_2431,N_2416);
nand U2622 (N_2622,N_2440,N_2425);
nand U2623 (N_2623,N_2534,N_2499);
nand U2624 (N_2624,N_2494,N_2419);
nand U2625 (N_2625,N_2455,N_2466);
or U2626 (N_2626,N_2538,N_2530);
nand U2627 (N_2627,N_2537,N_2448);
or U2628 (N_2628,N_2478,N_2413);
xnor U2629 (N_2629,N_2472,N_2567);
and U2630 (N_2630,N_2444,N_2565);
and U2631 (N_2631,N_2421,N_2591);
nand U2632 (N_2632,N_2451,N_2470);
or U2633 (N_2633,N_2564,N_2402);
or U2634 (N_2634,N_2532,N_2400);
or U2635 (N_2635,N_2528,N_2454);
nand U2636 (N_2636,N_2405,N_2412);
nor U2637 (N_2637,N_2406,N_2505);
nand U2638 (N_2638,N_2586,N_2446);
xor U2639 (N_2639,N_2489,N_2545);
and U2640 (N_2640,N_2553,N_2424);
or U2641 (N_2641,N_2404,N_2439);
or U2642 (N_2642,N_2409,N_2479);
xnor U2643 (N_2643,N_2525,N_2598);
xor U2644 (N_2644,N_2508,N_2539);
or U2645 (N_2645,N_2435,N_2512);
and U2646 (N_2646,N_2456,N_2473);
xor U2647 (N_2647,N_2522,N_2520);
or U2648 (N_2648,N_2581,N_2589);
xnor U2649 (N_2649,N_2580,N_2555);
or U2650 (N_2650,N_2531,N_2407);
xor U2651 (N_2651,N_2497,N_2493);
xnor U2652 (N_2652,N_2577,N_2569);
nor U2653 (N_2653,N_2436,N_2430);
and U2654 (N_2654,N_2495,N_2571);
and U2655 (N_2655,N_2503,N_2563);
or U2656 (N_2656,N_2562,N_2593);
and U2657 (N_2657,N_2483,N_2596);
or U2658 (N_2658,N_2433,N_2432);
nor U2659 (N_2659,N_2449,N_2573);
and U2660 (N_2660,N_2561,N_2513);
nor U2661 (N_2661,N_2482,N_2507);
and U2662 (N_2662,N_2559,N_2437);
and U2663 (N_2663,N_2509,N_2595);
nand U2664 (N_2664,N_2452,N_2457);
xnor U2665 (N_2665,N_2582,N_2438);
nand U2666 (N_2666,N_2429,N_2572);
nor U2667 (N_2667,N_2434,N_2511);
xor U2668 (N_2668,N_2570,N_2422);
nand U2669 (N_2669,N_2523,N_2557);
nor U2670 (N_2670,N_2536,N_2510);
and U2671 (N_2671,N_2414,N_2459);
or U2672 (N_2672,N_2521,N_2566);
nor U2673 (N_2673,N_2464,N_2423);
nor U2674 (N_2674,N_2467,N_2544);
nand U2675 (N_2675,N_2599,N_2401);
and U2676 (N_2676,N_2458,N_2594);
or U2677 (N_2677,N_2501,N_2535);
or U2678 (N_2678,N_2469,N_2524);
nand U2679 (N_2679,N_2579,N_2411);
xnor U2680 (N_2680,N_2514,N_2453);
nor U2681 (N_2681,N_2474,N_2502);
nand U2682 (N_2682,N_2585,N_2415);
xnor U2683 (N_2683,N_2504,N_2465);
or U2684 (N_2684,N_2588,N_2549);
nand U2685 (N_2685,N_2506,N_2540);
xnor U2686 (N_2686,N_2476,N_2487);
or U2687 (N_2687,N_2518,N_2526);
nand U2688 (N_2688,N_2560,N_2542);
xnor U2689 (N_2689,N_2554,N_2590);
nor U2690 (N_2690,N_2517,N_2496);
xnor U2691 (N_2691,N_2558,N_2527);
nand U2692 (N_2692,N_2450,N_2417);
or U2693 (N_2693,N_2519,N_2552);
nand U2694 (N_2694,N_2463,N_2575);
and U2695 (N_2695,N_2551,N_2578);
or U2696 (N_2696,N_2445,N_2418);
and U2697 (N_2697,N_2500,N_2576);
xnor U2698 (N_2698,N_2462,N_2475);
or U2699 (N_2699,N_2460,N_2468);
nor U2700 (N_2700,N_2461,N_2583);
nor U2701 (N_2701,N_2501,N_2470);
or U2702 (N_2702,N_2483,N_2416);
nor U2703 (N_2703,N_2412,N_2507);
or U2704 (N_2704,N_2471,N_2585);
nand U2705 (N_2705,N_2479,N_2543);
or U2706 (N_2706,N_2541,N_2447);
xor U2707 (N_2707,N_2402,N_2422);
and U2708 (N_2708,N_2562,N_2409);
and U2709 (N_2709,N_2458,N_2429);
nor U2710 (N_2710,N_2589,N_2455);
nand U2711 (N_2711,N_2471,N_2411);
xor U2712 (N_2712,N_2521,N_2527);
nand U2713 (N_2713,N_2400,N_2549);
and U2714 (N_2714,N_2481,N_2507);
nor U2715 (N_2715,N_2402,N_2496);
or U2716 (N_2716,N_2484,N_2520);
nand U2717 (N_2717,N_2533,N_2578);
and U2718 (N_2718,N_2577,N_2420);
and U2719 (N_2719,N_2598,N_2538);
nand U2720 (N_2720,N_2551,N_2408);
or U2721 (N_2721,N_2552,N_2551);
or U2722 (N_2722,N_2424,N_2573);
nor U2723 (N_2723,N_2464,N_2450);
nor U2724 (N_2724,N_2489,N_2587);
and U2725 (N_2725,N_2465,N_2410);
and U2726 (N_2726,N_2568,N_2564);
or U2727 (N_2727,N_2402,N_2490);
nor U2728 (N_2728,N_2547,N_2566);
and U2729 (N_2729,N_2440,N_2542);
nand U2730 (N_2730,N_2595,N_2560);
xnor U2731 (N_2731,N_2487,N_2454);
xor U2732 (N_2732,N_2529,N_2478);
or U2733 (N_2733,N_2418,N_2506);
xnor U2734 (N_2734,N_2440,N_2474);
nor U2735 (N_2735,N_2574,N_2463);
nor U2736 (N_2736,N_2533,N_2539);
xor U2737 (N_2737,N_2554,N_2502);
nand U2738 (N_2738,N_2539,N_2436);
and U2739 (N_2739,N_2543,N_2585);
nand U2740 (N_2740,N_2426,N_2580);
and U2741 (N_2741,N_2460,N_2521);
nand U2742 (N_2742,N_2539,N_2592);
or U2743 (N_2743,N_2579,N_2549);
nand U2744 (N_2744,N_2438,N_2491);
and U2745 (N_2745,N_2498,N_2472);
xor U2746 (N_2746,N_2490,N_2432);
nor U2747 (N_2747,N_2502,N_2574);
nand U2748 (N_2748,N_2489,N_2576);
nand U2749 (N_2749,N_2464,N_2460);
nand U2750 (N_2750,N_2468,N_2502);
or U2751 (N_2751,N_2411,N_2521);
nor U2752 (N_2752,N_2459,N_2437);
and U2753 (N_2753,N_2590,N_2448);
and U2754 (N_2754,N_2534,N_2414);
and U2755 (N_2755,N_2580,N_2417);
and U2756 (N_2756,N_2467,N_2477);
xnor U2757 (N_2757,N_2579,N_2577);
nor U2758 (N_2758,N_2438,N_2432);
or U2759 (N_2759,N_2574,N_2418);
xnor U2760 (N_2760,N_2551,N_2545);
nand U2761 (N_2761,N_2515,N_2420);
and U2762 (N_2762,N_2466,N_2567);
nand U2763 (N_2763,N_2455,N_2543);
xor U2764 (N_2764,N_2571,N_2414);
and U2765 (N_2765,N_2465,N_2554);
xnor U2766 (N_2766,N_2424,N_2554);
xnor U2767 (N_2767,N_2505,N_2529);
xnor U2768 (N_2768,N_2452,N_2535);
and U2769 (N_2769,N_2485,N_2553);
and U2770 (N_2770,N_2468,N_2477);
or U2771 (N_2771,N_2552,N_2466);
xnor U2772 (N_2772,N_2530,N_2472);
or U2773 (N_2773,N_2579,N_2463);
and U2774 (N_2774,N_2546,N_2446);
or U2775 (N_2775,N_2570,N_2582);
nor U2776 (N_2776,N_2492,N_2581);
and U2777 (N_2777,N_2473,N_2524);
or U2778 (N_2778,N_2546,N_2594);
nand U2779 (N_2779,N_2569,N_2537);
and U2780 (N_2780,N_2579,N_2456);
nand U2781 (N_2781,N_2407,N_2456);
nor U2782 (N_2782,N_2465,N_2436);
and U2783 (N_2783,N_2461,N_2469);
or U2784 (N_2784,N_2505,N_2447);
nand U2785 (N_2785,N_2536,N_2446);
or U2786 (N_2786,N_2481,N_2406);
or U2787 (N_2787,N_2413,N_2436);
or U2788 (N_2788,N_2596,N_2514);
or U2789 (N_2789,N_2565,N_2450);
xor U2790 (N_2790,N_2592,N_2465);
nand U2791 (N_2791,N_2420,N_2441);
nor U2792 (N_2792,N_2435,N_2493);
nor U2793 (N_2793,N_2431,N_2450);
nand U2794 (N_2794,N_2568,N_2497);
nand U2795 (N_2795,N_2569,N_2495);
nand U2796 (N_2796,N_2592,N_2521);
nor U2797 (N_2797,N_2427,N_2430);
nor U2798 (N_2798,N_2402,N_2469);
xnor U2799 (N_2799,N_2534,N_2522);
or U2800 (N_2800,N_2792,N_2630);
nor U2801 (N_2801,N_2646,N_2729);
and U2802 (N_2802,N_2657,N_2662);
nor U2803 (N_2803,N_2651,N_2695);
nor U2804 (N_2804,N_2718,N_2690);
nor U2805 (N_2805,N_2764,N_2660);
nand U2806 (N_2806,N_2724,N_2785);
or U2807 (N_2807,N_2756,N_2793);
and U2808 (N_2808,N_2727,N_2674);
or U2809 (N_2809,N_2776,N_2618);
nor U2810 (N_2810,N_2643,N_2687);
xnor U2811 (N_2811,N_2735,N_2711);
nand U2812 (N_2812,N_2613,N_2778);
nor U2813 (N_2813,N_2665,N_2702);
or U2814 (N_2814,N_2721,N_2621);
and U2815 (N_2815,N_2626,N_2753);
nand U2816 (N_2816,N_2611,N_2631);
nand U2817 (N_2817,N_2696,N_2629);
nor U2818 (N_2818,N_2761,N_2606);
and U2819 (N_2819,N_2712,N_2617);
xnor U2820 (N_2820,N_2726,N_2680);
or U2821 (N_2821,N_2710,N_2779);
nor U2822 (N_2822,N_2648,N_2723);
and U2823 (N_2823,N_2732,N_2737);
or U2824 (N_2824,N_2600,N_2786);
xnor U2825 (N_2825,N_2673,N_2628);
or U2826 (N_2826,N_2782,N_2734);
nor U2827 (N_2827,N_2692,N_2689);
xor U2828 (N_2828,N_2610,N_2720);
and U2829 (N_2829,N_2752,N_2766);
nor U2830 (N_2830,N_2619,N_2649);
xor U2831 (N_2831,N_2664,N_2788);
xnor U2832 (N_2832,N_2759,N_2769);
xor U2833 (N_2833,N_2741,N_2627);
or U2834 (N_2834,N_2693,N_2754);
and U2835 (N_2835,N_2671,N_2601);
or U2836 (N_2836,N_2669,N_2795);
nor U2837 (N_2837,N_2659,N_2731);
nor U2838 (N_2838,N_2666,N_2762);
or U2839 (N_2839,N_2738,N_2686);
nand U2840 (N_2840,N_2691,N_2688);
nor U2841 (N_2841,N_2678,N_2796);
xnor U2842 (N_2842,N_2672,N_2768);
nor U2843 (N_2843,N_2638,N_2780);
nor U2844 (N_2844,N_2763,N_2747);
nand U2845 (N_2845,N_2787,N_2767);
or U2846 (N_2846,N_2683,N_2681);
and U2847 (N_2847,N_2700,N_2715);
or U2848 (N_2848,N_2705,N_2789);
or U2849 (N_2849,N_2719,N_2603);
and U2850 (N_2850,N_2765,N_2791);
nor U2851 (N_2851,N_2799,N_2640);
or U2852 (N_2852,N_2623,N_2722);
nand U2853 (N_2853,N_2733,N_2616);
nor U2854 (N_2854,N_2605,N_2633);
nor U2855 (N_2855,N_2717,N_2798);
and U2856 (N_2856,N_2645,N_2676);
nor U2857 (N_2857,N_2708,N_2706);
nand U2858 (N_2858,N_2607,N_2698);
nor U2859 (N_2859,N_2602,N_2663);
and U2860 (N_2860,N_2608,N_2750);
nand U2861 (N_2861,N_2604,N_2771);
nor U2862 (N_2862,N_2755,N_2713);
xor U2863 (N_2863,N_2682,N_2758);
and U2864 (N_2864,N_2642,N_2794);
or U2865 (N_2865,N_2644,N_2736);
nor U2866 (N_2866,N_2728,N_2709);
nand U2867 (N_2867,N_2667,N_2614);
nor U2868 (N_2868,N_2637,N_2745);
nor U2869 (N_2869,N_2632,N_2757);
nand U2870 (N_2870,N_2699,N_2654);
nor U2871 (N_2871,N_2615,N_2668);
nor U2872 (N_2872,N_2636,N_2740);
nand U2873 (N_2873,N_2625,N_2624);
nand U2874 (N_2874,N_2704,N_2748);
or U2875 (N_2875,N_2746,N_2760);
nand U2876 (N_2876,N_2650,N_2661);
nand U2877 (N_2877,N_2697,N_2777);
or U2878 (N_2878,N_2770,N_2656);
or U2879 (N_2879,N_2725,N_2701);
or U2880 (N_2880,N_2653,N_2730);
or U2881 (N_2881,N_2772,N_2783);
nand U2882 (N_2882,N_2773,N_2743);
nand U2883 (N_2883,N_2775,N_2749);
xnor U2884 (N_2884,N_2635,N_2652);
or U2885 (N_2885,N_2658,N_2774);
or U2886 (N_2886,N_2744,N_2675);
nor U2887 (N_2887,N_2742,N_2790);
and U2888 (N_2888,N_2655,N_2784);
xor U2889 (N_2889,N_2639,N_2703);
xnor U2890 (N_2890,N_2714,N_2739);
xnor U2891 (N_2891,N_2612,N_2684);
or U2892 (N_2892,N_2609,N_2622);
xor U2893 (N_2893,N_2751,N_2620);
or U2894 (N_2894,N_2716,N_2707);
or U2895 (N_2895,N_2677,N_2685);
nor U2896 (N_2896,N_2647,N_2641);
or U2897 (N_2897,N_2634,N_2797);
and U2898 (N_2898,N_2781,N_2694);
xnor U2899 (N_2899,N_2670,N_2679);
xor U2900 (N_2900,N_2621,N_2752);
or U2901 (N_2901,N_2670,N_2727);
nand U2902 (N_2902,N_2685,N_2612);
nor U2903 (N_2903,N_2764,N_2794);
nor U2904 (N_2904,N_2632,N_2688);
nor U2905 (N_2905,N_2614,N_2677);
and U2906 (N_2906,N_2704,N_2775);
xor U2907 (N_2907,N_2689,N_2649);
or U2908 (N_2908,N_2773,N_2667);
nand U2909 (N_2909,N_2716,N_2718);
xnor U2910 (N_2910,N_2628,N_2763);
or U2911 (N_2911,N_2614,N_2721);
xor U2912 (N_2912,N_2610,N_2655);
nor U2913 (N_2913,N_2688,N_2631);
and U2914 (N_2914,N_2710,N_2643);
xnor U2915 (N_2915,N_2729,N_2612);
xor U2916 (N_2916,N_2624,N_2695);
or U2917 (N_2917,N_2639,N_2672);
and U2918 (N_2918,N_2615,N_2703);
and U2919 (N_2919,N_2798,N_2669);
nand U2920 (N_2920,N_2708,N_2672);
xor U2921 (N_2921,N_2679,N_2704);
and U2922 (N_2922,N_2794,N_2774);
nand U2923 (N_2923,N_2718,N_2691);
xnor U2924 (N_2924,N_2676,N_2642);
nor U2925 (N_2925,N_2703,N_2675);
or U2926 (N_2926,N_2679,N_2662);
nand U2927 (N_2927,N_2769,N_2780);
nor U2928 (N_2928,N_2748,N_2618);
nand U2929 (N_2929,N_2676,N_2604);
or U2930 (N_2930,N_2724,N_2663);
xor U2931 (N_2931,N_2760,N_2788);
xor U2932 (N_2932,N_2676,N_2660);
xor U2933 (N_2933,N_2753,N_2642);
nand U2934 (N_2934,N_2670,N_2666);
or U2935 (N_2935,N_2700,N_2612);
xor U2936 (N_2936,N_2748,N_2692);
xnor U2937 (N_2937,N_2646,N_2746);
and U2938 (N_2938,N_2676,N_2771);
xor U2939 (N_2939,N_2716,N_2653);
or U2940 (N_2940,N_2696,N_2792);
nor U2941 (N_2941,N_2615,N_2783);
or U2942 (N_2942,N_2709,N_2603);
nand U2943 (N_2943,N_2649,N_2777);
xnor U2944 (N_2944,N_2695,N_2781);
or U2945 (N_2945,N_2713,N_2761);
nand U2946 (N_2946,N_2774,N_2624);
xor U2947 (N_2947,N_2733,N_2754);
xor U2948 (N_2948,N_2663,N_2700);
nor U2949 (N_2949,N_2734,N_2655);
xnor U2950 (N_2950,N_2629,N_2640);
and U2951 (N_2951,N_2606,N_2627);
and U2952 (N_2952,N_2789,N_2781);
or U2953 (N_2953,N_2601,N_2728);
nor U2954 (N_2954,N_2752,N_2694);
xor U2955 (N_2955,N_2654,N_2646);
or U2956 (N_2956,N_2690,N_2681);
nor U2957 (N_2957,N_2755,N_2666);
xor U2958 (N_2958,N_2652,N_2605);
xor U2959 (N_2959,N_2731,N_2692);
or U2960 (N_2960,N_2705,N_2674);
xnor U2961 (N_2961,N_2663,N_2622);
nand U2962 (N_2962,N_2675,N_2705);
nor U2963 (N_2963,N_2786,N_2627);
or U2964 (N_2964,N_2790,N_2700);
nor U2965 (N_2965,N_2764,N_2652);
and U2966 (N_2966,N_2732,N_2795);
nor U2967 (N_2967,N_2745,N_2689);
nand U2968 (N_2968,N_2786,N_2745);
xor U2969 (N_2969,N_2634,N_2785);
xor U2970 (N_2970,N_2655,N_2748);
xor U2971 (N_2971,N_2714,N_2675);
xnor U2972 (N_2972,N_2708,N_2786);
nand U2973 (N_2973,N_2670,N_2765);
nand U2974 (N_2974,N_2632,N_2676);
nand U2975 (N_2975,N_2601,N_2617);
nand U2976 (N_2976,N_2718,N_2673);
and U2977 (N_2977,N_2623,N_2736);
or U2978 (N_2978,N_2659,N_2613);
nor U2979 (N_2979,N_2647,N_2774);
nor U2980 (N_2980,N_2681,N_2670);
xor U2981 (N_2981,N_2604,N_2646);
and U2982 (N_2982,N_2711,N_2744);
and U2983 (N_2983,N_2672,N_2774);
nand U2984 (N_2984,N_2702,N_2640);
xor U2985 (N_2985,N_2668,N_2707);
xnor U2986 (N_2986,N_2782,N_2603);
or U2987 (N_2987,N_2778,N_2728);
xnor U2988 (N_2988,N_2733,N_2643);
and U2989 (N_2989,N_2736,N_2616);
nor U2990 (N_2990,N_2631,N_2773);
or U2991 (N_2991,N_2682,N_2668);
and U2992 (N_2992,N_2635,N_2677);
nor U2993 (N_2993,N_2625,N_2661);
or U2994 (N_2994,N_2784,N_2698);
and U2995 (N_2995,N_2744,N_2664);
or U2996 (N_2996,N_2791,N_2614);
or U2997 (N_2997,N_2777,N_2677);
nor U2998 (N_2998,N_2678,N_2637);
xnor U2999 (N_2999,N_2660,N_2727);
xnor U3000 (N_3000,N_2811,N_2948);
xor U3001 (N_3001,N_2908,N_2968);
nand U3002 (N_3002,N_2856,N_2804);
and U3003 (N_3003,N_2927,N_2983);
xnor U3004 (N_3004,N_2865,N_2870);
xor U3005 (N_3005,N_2985,N_2816);
or U3006 (N_3006,N_2912,N_2885);
or U3007 (N_3007,N_2929,N_2822);
and U3008 (N_3008,N_2916,N_2975);
nand U3009 (N_3009,N_2844,N_2894);
nor U3010 (N_3010,N_2842,N_2861);
nor U3011 (N_3011,N_2841,N_2996);
nand U3012 (N_3012,N_2812,N_2889);
or U3013 (N_3013,N_2805,N_2959);
nand U3014 (N_3014,N_2937,N_2848);
xor U3015 (N_3015,N_2984,N_2864);
nand U3016 (N_3016,N_2827,N_2936);
and U3017 (N_3017,N_2837,N_2880);
nand U3018 (N_3018,N_2866,N_2909);
or U3019 (N_3019,N_2854,N_2886);
xnor U3020 (N_3020,N_2986,N_2823);
nor U3021 (N_3021,N_2891,N_2873);
or U3022 (N_3022,N_2887,N_2839);
and U3023 (N_3023,N_2976,N_2967);
and U3024 (N_3024,N_2925,N_2801);
and U3025 (N_3025,N_2950,N_2900);
xor U3026 (N_3026,N_2896,N_2819);
xnor U3027 (N_3027,N_2846,N_2961);
xnor U3028 (N_3028,N_2851,N_2992);
and U3029 (N_3029,N_2939,N_2809);
nand U3030 (N_3030,N_2833,N_2951);
nor U3031 (N_3031,N_2821,N_2814);
and U3032 (N_3032,N_2935,N_2958);
nor U3033 (N_3033,N_2956,N_2845);
or U3034 (N_3034,N_2834,N_2907);
and U3035 (N_3035,N_2981,N_2957);
nand U3036 (N_3036,N_2982,N_2892);
nor U3037 (N_3037,N_2913,N_2988);
or U3038 (N_3038,N_2843,N_2829);
xnor U3039 (N_3039,N_2836,N_2931);
nor U3040 (N_3040,N_2922,N_2857);
and U3041 (N_3041,N_2847,N_2802);
and U3042 (N_3042,N_2924,N_2852);
and U3043 (N_3043,N_2919,N_2883);
xor U3044 (N_3044,N_2974,N_2820);
xnor U3045 (N_3045,N_2881,N_2989);
nor U3046 (N_3046,N_2944,N_2849);
or U3047 (N_3047,N_2877,N_2990);
nand U3048 (N_3048,N_2914,N_2955);
xnor U3049 (N_3049,N_2902,N_2808);
and U3050 (N_3050,N_2897,N_2998);
xnor U3051 (N_3051,N_2918,N_2835);
or U3052 (N_3052,N_2945,N_2826);
nor U3053 (N_3053,N_2991,N_2930);
or U3054 (N_3054,N_2871,N_2863);
or U3055 (N_3055,N_2932,N_2962);
nand U3056 (N_3056,N_2874,N_2859);
or U3057 (N_3057,N_2824,N_2905);
nor U3058 (N_3058,N_2872,N_2917);
xnor U3059 (N_3059,N_2973,N_2928);
nand U3060 (N_3060,N_2970,N_2999);
and U3061 (N_3061,N_2806,N_2949);
or U3062 (N_3062,N_2964,N_2853);
or U3063 (N_3063,N_2971,N_2828);
and U3064 (N_3064,N_2807,N_2923);
xnor U3065 (N_3065,N_2926,N_2815);
nor U3066 (N_3066,N_2921,N_2893);
and U3067 (N_3067,N_2875,N_2910);
xor U3068 (N_3068,N_2978,N_2888);
or U3069 (N_3069,N_2995,N_2901);
nor U3070 (N_3070,N_2817,N_2832);
nor U3071 (N_3071,N_2941,N_2890);
xor U3072 (N_3072,N_2879,N_2915);
nor U3073 (N_3073,N_2933,N_2800);
xor U3074 (N_3074,N_2947,N_2943);
nor U3075 (N_3075,N_2855,N_2965);
and U3076 (N_3076,N_2966,N_2954);
xor U3077 (N_3077,N_2953,N_2862);
nand U3078 (N_3078,N_2840,N_2997);
nor U3079 (N_3079,N_2940,N_2850);
or U3080 (N_3080,N_2904,N_2938);
or U3081 (N_3081,N_2830,N_2946);
or U3082 (N_3082,N_2963,N_2810);
nor U3083 (N_3083,N_2911,N_2920);
or U3084 (N_3084,N_2903,N_2813);
xnor U3085 (N_3085,N_2979,N_2825);
nand U3086 (N_3086,N_2882,N_2980);
nor U3087 (N_3087,N_2831,N_2867);
and U3088 (N_3088,N_2987,N_2952);
nand U3089 (N_3089,N_2895,N_2869);
or U3090 (N_3090,N_2803,N_2858);
nand U3091 (N_3091,N_2860,N_2960);
or U3092 (N_3092,N_2972,N_2994);
nor U3093 (N_3093,N_2838,N_2868);
nand U3094 (N_3094,N_2977,N_2993);
or U3095 (N_3095,N_2906,N_2818);
nor U3096 (N_3096,N_2969,N_2884);
nand U3097 (N_3097,N_2876,N_2899);
and U3098 (N_3098,N_2878,N_2898);
nand U3099 (N_3099,N_2942,N_2934);
nor U3100 (N_3100,N_2950,N_2882);
nand U3101 (N_3101,N_2855,N_2823);
nand U3102 (N_3102,N_2905,N_2854);
nor U3103 (N_3103,N_2891,N_2992);
nand U3104 (N_3104,N_2911,N_2982);
xor U3105 (N_3105,N_2936,N_2872);
and U3106 (N_3106,N_2803,N_2813);
nand U3107 (N_3107,N_2806,N_2913);
xor U3108 (N_3108,N_2848,N_2857);
nor U3109 (N_3109,N_2999,N_2843);
nor U3110 (N_3110,N_2951,N_2982);
and U3111 (N_3111,N_2900,N_2982);
nor U3112 (N_3112,N_2954,N_2995);
xnor U3113 (N_3113,N_2846,N_2844);
nor U3114 (N_3114,N_2845,N_2919);
nand U3115 (N_3115,N_2853,N_2925);
or U3116 (N_3116,N_2860,N_2935);
xnor U3117 (N_3117,N_2865,N_2826);
xnor U3118 (N_3118,N_2886,N_2939);
and U3119 (N_3119,N_2807,N_2801);
or U3120 (N_3120,N_2986,N_2920);
or U3121 (N_3121,N_2980,N_2886);
and U3122 (N_3122,N_2904,N_2848);
xor U3123 (N_3123,N_2904,N_2934);
nor U3124 (N_3124,N_2975,N_2844);
nor U3125 (N_3125,N_2813,N_2810);
or U3126 (N_3126,N_2886,N_2923);
and U3127 (N_3127,N_2997,N_2892);
nor U3128 (N_3128,N_2960,N_2811);
nand U3129 (N_3129,N_2837,N_2916);
and U3130 (N_3130,N_2995,N_2903);
xnor U3131 (N_3131,N_2946,N_2986);
xnor U3132 (N_3132,N_2968,N_2937);
xnor U3133 (N_3133,N_2818,N_2838);
xor U3134 (N_3134,N_2826,N_2974);
xor U3135 (N_3135,N_2843,N_2972);
or U3136 (N_3136,N_2910,N_2945);
nor U3137 (N_3137,N_2947,N_2921);
or U3138 (N_3138,N_2966,N_2829);
nor U3139 (N_3139,N_2954,N_2880);
xor U3140 (N_3140,N_2817,N_2941);
or U3141 (N_3141,N_2852,N_2895);
nor U3142 (N_3142,N_2867,N_2931);
or U3143 (N_3143,N_2821,N_2898);
and U3144 (N_3144,N_2891,N_2808);
xor U3145 (N_3145,N_2881,N_2927);
and U3146 (N_3146,N_2823,N_2828);
xnor U3147 (N_3147,N_2904,N_2985);
and U3148 (N_3148,N_2854,N_2894);
nand U3149 (N_3149,N_2813,N_2935);
and U3150 (N_3150,N_2902,N_2917);
or U3151 (N_3151,N_2948,N_2966);
or U3152 (N_3152,N_2918,N_2967);
and U3153 (N_3153,N_2859,N_2832);
nor U3154 (N_3154,N_2974,N_2906);
or U3155 (N_3155,N_2846,N_2876);
or U3156 (N_3156,N_2900,N_2807);
nor U3157 (N_3157,N_2804,N_2858);
nor U3158 (N_3158,N_2833,N_2861);
nor U3159 (N_3159,N_2818,N_2809);
or U3160 (N_3160,N_2803,N_2912);
nand U3161 (N_3161,N_2985,N_2915);
and U3162 (N_3162,N_2985,N_2831);
xor U3163 (N_3163,N_2936,N_2996);
or U3164 (N_3164,N_2906,N_2883);
nor U3165 (N_3165,N_2819,N_2942);
nor U3166 (N_3166,N_2904,N_2960);
and U3167 (N_3167,N_2834,N_2999);
xor U3168 (N_3168,N_2860,N_2859);
and U3169 (N_3169,N_2829,N_2800);
nor U3170 (N_3170,N_2999,N_2823);
and U3171 (N_3171,N_2970,N_2865);
xnor U3172 (N_3172,N_2828,N_2811);
and U3173 (N_3173,N_2819,N_2801);
and U3174 (N_3174,N_2808,N_2990);
and U3175 (N_3175,N_2974,N_2997);
nor U3176 (N_3176,N_2968,N_2995);
or U3177 (N_3177,N_2897,N_2867);
or U3178 (N_3178,N_2835,N_2966);
and U3179 (N_3179,N_2880,N_2902);
nor U3180 (N_3180,N_2889,N_2881);
xor U3181 (N_3181,N_2811,N_2918);
nor U3182 (N_3182,N_2966,N_2848);
xnor U3183 (N_3183,N_2836,N_2835);
and U3184 (N_3184,N_2894,N_2908);
and U3185 (N_3185,N_2990,N_2806);
nor U3186 (N_3186,N_2924,N_2962);
and U3187 (N_3187,N_2882,N_2829);
xnor U3188 (N_3188,N_2924,N_2980);
nand U3189 (N_3189,N_2854,N_2824);
or U3190 (N_3190,N_2932,N_2811);
nor U3191 (N_3191,N_2993,N_2941);
and U3192 (N_3192,N_2885,N_2836);
and U3193 (N_3193,N_2933,N_2838);
and U3194 (N_3194,N_2863,N_2911);
or U3195 (N_3195,N_2896,N_2948);
or U3196 (N_3196,N_2936,N_2891);
or U3197 (N_3197,N_2871,N_2827);
nor U3198 (N_3198,N_2920,N_2966);
and U3199 (N_3199,N_2932,N_2884);
nor U3200 (N_3200,N_3020,N_3024);
xnor U3201 (N_3201,N_3062,N_3132);
or U3202 (N_3202,N_3193,N_3156);
nand U3203 (N_3203,N_3185,N_3016);
nor U3204 (N_3204,N_3093,N_3019);
and U3205 (N_3205,N_3060,N_3199);
xor U3206 (N_3206,N_3054,N_3059);
and U3207 (N_3207,N_3142,N_3129);
nor U3208 (N_3208,N_3001,N_3108);
nand U3209 (N_3209,N_3101,N_3047);
xor U3210 (N_3210,N_3168,N_3126);
or U3211 (N_3211,N_3037,N_3086);
or U3212 (N_3212,N_3066,N_3032);
xnor U3213 (N_3213,N_3025,N_3124);
nand U3214 (N_3214,N_3184,N_3096);
and U3215 (N_3215,N_3038,N_3183);
or U3216 (N_3216,N_3084,N_3053);
or U3217 (N_3217,N_3178,N_3153);
and U3218 (N_3218,N_3077,N_3165);
nor U3219 (N_3219,N_3114,N_3048);
nand U3220 (N_3220,N_3118,N_3014);
and U3221 (N_3221,N_3027,N_3041);
xnor U3222 (N_3222,N_3089,N_3011);
or U3223 (N_3223,N_3005,N_3122);
xor U3224 (N_3224,N_3151,N_3069);
nor U3225 (N_3225,N_3198,N_3003);
xnor U3226 (N_3226,N_3070,N_3104);
and U3227 (N_3227,N_3081,N_3051);
or U3228 (N_3228,N_3174,N_3109);
nand U3229 (N_3229,N_3055,N_3026);
xor U3230 (N_3230,N_3128,N_3013);
or U3231 (N_3231,N_3191,N_3067);
nand U3232 (N_3232,N_3082,N_3065);
nand U3233 (N_3233,N_3058,N_3102);
and U3234 (N_3234,N_3111,N_3121);
xnor U3235 (N_3235,N_3036,N_3158);
or U3236 (N_3236,N_3105,N_3177);
xnor U3237 (N_3237,N_3068,N_3149);
or U3238 (N_3238,N_3162,N_3017);
nor U3239 (N_3239,N_3161,N_3103);
xor U3240 (N_3240,N_3004,N_3031);
nand U3241 (N_3241,N_3092,N_3033);
xor U3242 (N_3242,N_3061,N_3099);
or U3243 (N_3243,N_3169,N_3085);
or U3244 (N_3244,N_3190,N_3074);
or U3245 (N_3245,N_3043,N_3006);
nor U3246 (N_3246,N_3091,N_3179);
nand U3247 (N_3247,N_3141,N_3194);
nor U3248 (N_3248,N_3100,N_3147);
nand U3249 (N_3249,N_3052,N_3083);
nor U3250 (N_3250,N_3040,N_3173);
nor U3251 (N_3251,N_3143,N_3073);
and U3252 (N_3252,N_3095,N_3098);
nand U3253 (N_3253,N_3182,N_3189);
and U3254 (N_3254,N_3107,N_3029);
and U3255 (N_3255,N_3002,N_3090);
nor U3256 (N_3256,N_3130,N_3009);
xor U3257 (N_3257,N_3012,N_3018);
or U3258 (N_3258,N_3123,N_3152);
nor U3259 (N_3259,N_3079,N_3030);
or U3260 (N_3260,N_3139,N_3000);
or U3261 (N_3261,N_3140,N_3157);
and U3262 (N_3262,N_3113,N_3164);
xor U3263 (N_3263,N_3166,N_3075);
nor U3264 (N_3264,N_3023,N_3057);
and U3265 (N_3265,N_3137,N_3050);
nor U3266 (N_3266,N_3155,N_3022);
and U3267 (N_3267,N_3035,N_3170);
nand U3268 (N_3268,N_3181,N_3088);
xor U3269 (N_3269,N_3094,N_3167);
or U3270 (N_3270,N_3021,N_3080);
or U3271 (N_3271,N_3138,N_3087);
xor U3272 (N_3272,N_3125,N_3127);
xnor U3273 (N_3273,N_3186,N_3078);
nor U3274 (N_3274,N_3049,N_3097);
and U3275 (N_3275,N_3146,N_3034);
or U3276 (N_3276,N_3044,N_3028);
and U3277 (N_3277,N_3180,N_3175);
xor U3278 (N_3278,N_3131,N_3134);
nand U3279 (N_3279,N_3144,N_3010);
and U3280 (N_3280,N_3171,N_3150);
xnor U3281 (N_3281,N_3159,N_3133);
or U3282 (N_3282,N_3112,N_3172);
or U3283 (N_3283,N_3076,N_3115);
xnor U3284 (N_3284,N_3072,N_3071);
nand U3285 (N_3285,N_3160,N_3042);
nand U3286 (N_3286,N_3196,N_3176);
nand U3287 (N_3287,N_3192,N_3197);
or U3288 (N_3288,N_3187,N_3063);
xnor U3289 (N_3289,N_3039,N_3148);
xnor U3290 (N_3290,N_3145,N_3056);
xor U3291 (N_3291,N_3154,N_3116);
nor U3292 (N_3292,N_3045,N_3015);
nor U3293 (N_3293,N_3008,N_3188);
nand U3294 (N_3294,N_3135,N_3117);
and U3295 (N_3295,N_3064,N_3195);
and U3296 (N_3296,N_3007,N_3106);
and U3297 (N_3297,N_3119,N_3136);
nor U3298 (N_3298,N_3110,N_3046);
xor U3299 (N_3299,N_3163,N_3120);
nand U3300 (N_3300,N_3049,N_3188);
xor U3301 (N_3301,N_3171,N_3006);
nor U3302 (N_3302,N_3004,N_3077);
and U3303 (N_3303,N_3008,N_3132);
nor U3304 (N_3304,N_3192,N_3055);
nand U3305 (N_3305,N_3009,N_3190);
nand U3306 (N_3306,N_3199,N_3075);
and U3307 (N_3307,N_3175,N_3199);
nand U3308 (N_3308,N_3159,N_3197);
nor U3309 (N_3309,N_3056,N_3020);
nor U3310 (N_3310,N_3030,N_3081);
xnor U3311 (N_3311,N_3182,N_3080);
xor U3312 (N_3312,N_3068,N_3021);
nor U3313 (N_3313,N_3080,N_3141);
nor U3314 (N_3314,N_3198,N_3178);
xor U3315 (N_3315,N_3146,N_3013);
and U3316 (N_3316,N_3036,N_3040);
or U3317 (N_3317,N_3141,N_3085);
nand U3318 (N_3318,N_3087,N_3121);
or U3319 (N_3319,N_3093,N_3000);
nor U3320 (N_3320,N_3041,N_3188);
xnor U3321 (N_3321,N_3012,N_3146);
nor U3322 (N_3322,N_3060,N_3109);
nand U3323 (N_3323,N_3114,N_3023);
xnor U3324 (N_3324,N_3058,N_3005);
nand U3325 (N_3325,N_3196,N_3142);
and U3326 (N_3326,N_3193,N_3140);
or U3327 (N_3327,N_3156,N_3034);
and U3328 (N_3328,N_3098,N_3090);
nand U3329 (N_3329,N_3055,N_3007);
or U3330 (N_3330,N_3032,N_3174);
nand U3331 (N_3331,N_3192,N_3079);
or U3332 (N_3332,N_3192,N_3133);
or U3333 (N_3333,N_3003,N_3089);
or U3334 (N_3334,N_3183,N_3128);
nand U3335 (N_3335,N_3009,N_3093);
and U3336 (N_3336,N_3137,N_3169);
and U3337 (N_3337,N_3138,N_3120);
or U3338 (N_3338,N_3011,N_3178);
nand U3339 (N_3339,N_3171,N_3113);
nand U3340 (N_3340,N_3180,N_3052);
xor U3341 (N_3341,N_3159,N_3055);
and U3342 (N_3342,N_3196,N_3080);
nor U3343 (N_3343,N_3074,N_3021);
and U3344 (N_3344,N_3099,N_3196);
nor U3345 (N_3345,N_3126,N_3150);
nand U3346 (N_3346,N_3069,N_3067);
and U3347 (N_3347,N_3040,N_3150);
nor U3348 (N_3348,N_3051,N_3159);
nor U3349 (N_3349,N_3199,N_3111);
nor U3350 (N_3350,N_3197,N_3033);
nor U3351 (N_3351,N_3009,N_3032);
nand U3352 (N_3352,N_3003,N_3130);
and U3353 (N_3353,N_3012,N_3035);
nor U3354 (N_3354,N_3132,N_3002);
nand U3355 (N_3355,N_3143,N_3145);
nand U3356 (N_3356,N_3106,N_3105);
xnor U3357 (N_3357,N_3020,N_3071);
nand U3358 (N_3358,N_3196,N_3066);
nand U3359 (N_3359,N_3062,N_3136);
nand U3360 (N_3360,N_3061,N_3169);
nand U3361 (N_3361,N_3046,N_3053);
or U3362 (N_3362,N_3073,N_3093);
or U3363 (N_3363,N_3094,N_3088);
and U3364 (N_3364,N_3132,N_3057);
and U3365 (N_3365,N_3174,N_3027);
xor U3366 (N_3366,N_3191,N_3044);
nor U3367 (N_3367,N_3057,N_3103);
or U3368 (N_3368,N_3135,N_3034);
nor U3369 (N_3369,N_3120,N_3067);
nor U3370 (N_3370,N_3112,N_3126);
nand U3371 (N_3371,N_3135,N_3187);
xor U3372 (N_3372,N_3125,N_3092);
and U3373 (N_3373,N_3184,N_3018);
nor U3374 (N_3374,N_3026,N_3118);
nand U3375 (N_3375,N_3050,N_3006);
xor U3376 (N_3376,N_3059,N_3189);
and U3377 (N_3377,N_3178,N_3105);
and U3378 (N_3378,N_3062,N_3146);
nor U3379 (N_3379,N_3121,N_3175);
and U3380 (N_3380,N_3046,N_3152);
or U3381 (N_3381,N_3113,N_3186);
nand U3382 (N_3382,N_3169,N_3026);
xor U3383 (N_3383,N_3030,N_3113);
nor U3384 (N_3384,N_3062,N_3155);
or U3385 (N_3385,N_3088,N_3121);
nor U3386 (N_3386,N_3013,N_3098);
and U3387 (N_3387,N_3176,N_3161);
nand U3388 (N_3388,N_3138,N_3139);
or U3389 (N_3389,N_3100,N_3081);
or U3390 (N_3390,N_3049,N_3084);
or U3391 (N_3391,N_3154,N_3082);
xnor U3392 (N_3392,N_3048,N_3108);
nor U3393 (N_3393,N_3037,N_3155);
and U3394 (N_3394,N_3019,N_3049);
nor U3395 (N_3395,N_3180,N_3011);
xnor U3396 (N_3396,N_3144,N_3006);
nand U3397 (N_3397,N_3144,N_3074);
nor U3398 (N_3398,N_3046,N_3075);
nand U3399 (N_3399,N_3094,N_3066);
and U3400 (N_3400,N_3343,N_3354);
or U3401 (N_3401,N_3394,N_3215);
or U3402 (N_3402,N_3264,N_3307);
nand U3403 (N_3403,N_3333,N_3261);
and U3404 (N_3404,N_3204,N_3239);
nor U3405 (N_3405,N_3205,N_3294);
and U3406 (N_3406,N_3260,N_3213);
nor U3407 (N_3407,N_3316,N_3355);
or U3408 (N_3408,N_3393,N_3375);
and U3409 (N_3409,N_3259,N_3310);
xor U3410 (N_3410,N_3225,N_3247);
and U3411 (N_3411,N_3382,N_3278);
and U3412 (N_3412,N_3297,N_3285);
nand U3413 (N_3413,N_3383,N_3207);
or U3414 (N_3414,N_3332,N_3321);
xor U3415 (N_3415,N_3326,N_3371);
nor U3416 (N_3416,N_3399,N_3216);
or U3417 (N_3417,N_3342,N_3234);
xor U3418 (N_3418,N_3346,N_3386);
xnor U3419 (N_3419,N_3398,N_3218);
or U3420 (N_3420,N_3385,N_3363);
nor U3421 (N_3421,N_3317,N_3327);
nor U3422 (N_3422,N_3300,N_3380);
or U3423 (N_3423,N_3286,N_3240);
or U3424 (N_3424,N_3341,N_3389);
nand U3425 (N_3425,N_3373,N_3315);
nand U3426 (N_3426,N_3309,N_3396);
nor U3427 (N_3427,N_3220,N_3311);
or U3428 (N_3428,N_3209,N_3368);
or U3429 (N_3429,N_3219,N_3230);
or U3430 (N_3430,N_3359,N_3356);
xnor U3431 (N_3431,N_3301,N_3267);
nand U3432 (N_3432,N_3338,N_3210);
nor U3433 (N_3433,N_3319,N_3365);
or U3434 (N_3434,N_3206,N_3262);
xnor U3435 (N_3435,N_3306,N_3227);
xor U3436 (N_3436,N_3233,N_3283);
nand U3437 (N_3437,N_3253,N_3387);
or U3438 (N_3438,N_3250,N_3347);
and U3439 (N_3439,N_3296,N_3378);
nand U3440 (N_3440,N_3287,N_3305);
or U3441 (N_3441,N_3256,N_3232);
and U3442 (N_3442,N_3281,N_3243);
or U3443 (N_3443,N_3351,N_3257);
and U3444 (N_3444,N_3397,N_3214);
nand U3445 (N_3445,N_3350,N_3201);
nor U3446 (N_3446,N_3277,N_3254);
nand U3447 (N_3447,N_3302,N_3221);
nand U3448 (N_3448,N_3328,N_3211);
or U3449 (N_3449,N_3345,N_3228);
and U3450 (N_3450,N_3271,N_3231);
or U3451 (N_3451,N_3289,N_3352);
or U3452 (N_3452,N_3392,N_3290);
nand U3453 (N_3453,N_3208,N_3202);
xor U3454 (N_3454,N_3265,N_3335);
and U3455 (N_3455,N_3303,N_3388);
xnor U3456 (N_3456,N_3320,N_3370);
nand U3457 (N_3457,N_3372,N_3249);
nand U3458 (N_3458,N_3272,N_3203);
or U3459 (N_3459,N_3344,N_3299);
or U3460 (N_3460,N_3222,N_3334);
nand U3461 (N_3461,N_3212,N_3376);
and U3462 (N_3462,N_3384,N_3244);
or U3463 (N_3463,N_3298,N_3361);
or U3464 (N_3464,N_3331,N_3241);
nor U3465 (N_3465,N_3273,N_3304);
or U3466 (N_3466,N_3251,N_3377);
or U3467 (N_3467,N_3291,N_3348);
nand U3468 (N_3468,N_3353,N_3324);
xnor U3469 (N_3469,N_3266,N_3366);
and U3470 (N_3470,N_3235,N_3284);
nor U3471 (N_3471,N_3246,N_3282);
xor U3472 (N_3472,N_3280,N_3318);
nor U3473 (N_3473,N_3379,N_3276);
xor U3474 (N_3474,N_3362,N_3248);
xnor U3475 (N_3475,N_3358,N_3312);
xnor U3476 (N_3476,N_3357,N_3274);
and U3477 (N_3477,N_3330,N_3293);
nand U3478 (N_3478,N_3295,N_3263);
xnor U3479 (N_3479,N_3223,N_3242);
nor U3480 (N_3480,N_3374,N_3255);
and U3481 (N_3481,N_3381,N_3229);
nor U3482 (N_3482,N_3236,N_3288);
xor U3483 (N_3483,N_3224,N_3323);
nand U3484 (N_3484,N_3364,N_3270);
and U3485 (N_3485,N_3238,N_3340);
or U3486 (N_3486,N_3325,N_3360);
and U3487 (N_3487,N_3313,N_3258);
xor U3488 (N_3488,N_3245,N_3217);
xnor U3489 (N_3489,N_3395,N_3349);
nor U3490 (N_3490,N_3292,N_3226);
nand U3491 (N_3491,N_3322,N_3390);
nor U3492 (N_3492,N_3339,N_3269);
nor U3493 (N_3493,N_3367,N_3308);
xnor U3494 (N_3494,N_3252,N_3275);
nor U3495 (N_3495,N_3268,N_3279);
nor U3496 (N_3496,N_3314,N_3336);
and U3497 (N_3497,N_3329,N_3237);
nand U3498 (N_3498,N_3391,N_3200);
xor U3499 (N_3499,N_3369,N_3337);
or U3500 (N_3500,N_3220,N_3237);
nor U3501 (N_3501,N_3325,N_3327);
nand U3502 (N_3502,N_3335,N_3327);
nand U3503 (N_3503,N_3288,N_3332);
or U3504 (N_3504,N_3317,N_3286);
xnor U3505 (N_3505,N_3398,N_3322);
xnor U3506 (N_3506,N_3344,N_3282);
nand U3507 (N_3507,N_3288,N_3389);
and U3508 (N_3508,N_3222,N_3391);
or U3509 (N_3509,N_3370,N_3263);
or U3510 (N_3510,N_3336,N_3303);
nor U3511 (N_3511,N_3208,N_3356);
or U3512 (N_3512,N_3269,N_3297);
xnor U3513 (N_3513,N_3296,N_3269);
nor U3514 (N_3514,N_3380,N_3308);
xnor U3515 (N_3515,N_3203,N_3305);
xor U3516 (N_3516,N_3212,N_3397);
xor U3517 (N_3517,N_3304,N_3377);
and U3518 (N_3518,N_3281,N_3307);
or U3519 (N_3519,N_3238,N_3304);
or U3520 (N_3520,N_3204,N_3300);
and U3521 (N_3521,N_3339,N_3396);
and U3522 (N_3522,N_3380,N_3226);
xnor U3523 (N_3523,N_3229,N_3366);
and U3524 (N_3524,N_3282,N_3256);
nand U3525 (N_3525,N_3359,N_3322);
nor U3526 (N_3526,N_3248,N_3328);
or U3527 (N_3527,N_3254,N_3212);
or U3528 (N_3528,N_3313,N_3366);
or U3529 (N_3529,N_3260,N_3289);
nor U3530 (N_3530,N_3345,N_3294);
nand U3531 (N_3531,N_3209,N_3244);
or U3532 (N_3532,N_3301,N_3206);
xor U3533 (N_3533,N_3253,N_3308);
nand U3534 (N_3534,N_3384,N_3315);
or U3535 (N_3535,N_3221,N_3300);
or U3536 (N_3536,N_3319,N_3344);
and U3537 (N_3537,N_3379,N_3265);
and U3538 (N_3538,N_3377,N_3256);
or U3539 (N_3539,N_3388,N_3304);
and U3540 (N_3540,N_3353,N_3329);
xnor U3541 (N_3541,N_3327,N_3261);
nand U3542 (N_3542,N_3368,N_3314);
and U3543 (N_3543,N_3386,N_3293);
nor U3544 (N_3544,N_3273,N_3388);
and U3545 (N_3545,N_3284,N_3268);
and U3546 (N_3546,N_3359,N_3357);
nor U3547 (N_3547,N_3357,N_3239);
or U3548 (N_3548,N_3328,N_3330);
xnor U3549 (N_3549,N_3334,N_3348);
nand U3550 (N_3550,N_3324,N_3230);
nand U3551 (N_3551,N_3278,N_3395);
nor U3552 (N_3552,N_3346,N_3335);
or U3553 (N_3553,N_3375,N_3201);
or U3554 (N_3554,N_3266,N_3209);
nand U3555 (N_3555,N_3304,N_3399);
nand U3556 (N_3556,N_3256,N_3226);
and U3557 (N_3557,N_3204,N_3222);
and U3558 (N_3558,N_3371,N_3277);
nand U3559 (N_3559,N_3244,N_3238);
or U3560 (N_3560,N_3205,N_3267);
nor U3561 (N_3561,N_3394,N_3208);
and U3562 (N_3562,N_3282,N_3284);
and U3563 (N_3563,N_3398,N_3370);
and U3564 (N_3564,N_3361,N_3379);
nand U3565 (N_3565,N_3210,N_3393);
nand U3566 (N_3566,N_3357,N_3269);
nand U3567 (N_3567,N_3270,N_3214);
or U3568 (N_3568,N_3322,N_3318);
nand U3569 (N_3569,N_3228,N_3277);
and U3570 (N_3570,N_3360,N_3237);
or U3571 (N_3571,N_3375,N_3382);
or U3572 (N_3572,N_3258,N_3301);
or U3573 (N_3573,N_3365,N_3310);
nor U3574 (N_3574,N_3354,N_3245);
or U3575 (N_3575,N_3214,N_3274);
and U3576 (N_3576,N_3213,N_3333);
xor U3577 (N_3577,N_3388,N_3263);
or U3578 (N_3578,N_3393,N_3338);
and U3579 (N_3579,N_3282,N_3380);
nor U3580 (N_3580,N_3204,N_3244);
nor U3581 (N_3581,N_3274,N_3247);
xor U3582 (N_3582,N_3328,N_3286);
nor U3583 (N_3583,N_3285,N_3304);
and U3584 (N_3584,N_3367,N_3342);
and U3585 (N_3585,N_3228,N_3266);
nor U3586 (N_3586,N_3213,N_3296);
nand U3587 (N_3587,N_3213,N_3346);
and U3588 (N_3588,N_3211,N_3303);
nor U3589 (N_3589,N_3250,N_3340);
or U3590 (N_3590,N_3220,N_3378);
nand U3591 (N_3591,N_3283,N_3376);
xnor U3592 (N_3592,N_3240,N_3328);
and U3593 (N_3593,N_3275,N_3291);
or U3594 (N_3594,N_3245,N_3314);
xor U3595 (N_3595,N_3378,N_3397);
nand U3596 (N_3596,N_3203,N_3237);
nor U3597 (N_3597,N_3317,N_3234);
and U3598 (N_3598,N_3301,N_3227);
nand U3599 (N_3599,N_3266,N_3346);
nand U3600 (N_3600,N_3494,N_3426);
or U3601 (N_3601,N_3552,N_3567);
xnor U3602 (N_3602,N_3462,N_3525);
or U3603 (N_3603,N_3425,N_3451);
nand U3604 (N_3604,N_3574,N_3515);
or U3605 (N_3605,N_3442,N_3478);
and U3606 (N_3606,N_3437,N_3454);
nand U3607 (N_3607,N_3597,N_3420);
xnor U3608 (N_3608,N_3500,N_3423);
nor U3609 (N_3609,N_3475,N_3592);
nand U3610 (N_3610,N_3460,N_3473);
and U3611 (N_3611,N_3573,N_3471);
and U3612 (N_3612,N_3576,N_3468);
nand U3613 (N_3613,N_3535,N_3529);
or U3614 (N_3614,N_3546,N_3400);
xor U3615 (N_3615,N_3566,N_3541);
xor U3616 (N_3616,N_3418,N_3558);
nand U3617 (N_3617,N_3443,N_3455);
nand U3618 (N_3618,N_3419,N_3452);
nor U3619 (N_3619,N_3410,N_3476);
or U3620 (N_3620,N_3479,N_3467);
and U3621 (N_3621,N_3590,N_3413);
or U3622 (N_3622,N_3445,N_3506);
xnor U3623 (N_3623,N_3596,N_3491);
nor U3624 (N_3624,N_3405,N_3569);
xor U3625 (N_3625,N_3509,N_3415);
xor U3626 (N_3626,N_3516,N_3599);
nor U3627 (N_3627,N_3481,N_3428);
nor U3628 (N_3628,N_3564,N_3524);
and U3629 (N_3629,N_3540,N_3403);
nand U3630 (N_3630,N_3480,N_3430);
or U3631 (N_3631,N_3449,N_3469);
or U3632 (N_3632,N_3549,N_3411);
nor U3633 (N_3633,N_3539,N_3557);
or U3634 (N_3634,N_3448,N_3530);
and U3635 (N_3635,N_3518,N_3434);
xnor U3636 (N_3636,N_3484,N_3458);
nor U3637 (N_3637,N_3501,N_3466);
xnor U3638 (N_3638,N_3595,N_3447);
nand U3639 (N_3639,N_3542,N_3545);
nand U3640 (N_3640,N_3512,N_3538);
nand U3641 (N_3641,N_3589,N_3424);
xnor U3642 (N_3642,N_3562,N_3465);
or U3643 (N_3643,N_3457,N_3526);
nand U3644 (N_3644,N_3474,N_3464);
nand U3645 (N_3645,N_3578,N_3585);
and U3646 (N_3646,N_3586,N_3581);
nand U3647 (N_3647,N_3441,N_3402);
nand U3648 (N_3648,N_3547,N_3528);
or U3649 (N_3649,N_3435,N_3408);
nand U3650 (N_3650,N_3560,N_3587);
and U3651 (N_3651,N_3563,N_3498);
or U3652 (N_3652,N_3488,N_3453);
or U3653 (N_3653,N_3550,N_3461);
nor U3654 (N_3654,N_3470,N_3572);
and U3655 (N_3655,N_3505,N_3598);
or U3656 (N_3656,N_3446,N_3544);
nor U3657 (N_3657,N_3568,N_3427);
or U3658 (N_3658,N_3433,N_3532);
xor U3659 (N_3659,N_3559,N_3438);
xor U3660 (N_3660,N_3561,N_3417);
or U3661 (N_3661,N_3575,N_3502);
nand U3662 (N_3662,N_3444,N_3570);
nand U3663 (N_3663,N_3583,N_3527);
nand U3664 (N_3664,N_3503,N_3522);
or U3665 (N_3665,N_3556,N_3551);
nand U3666 (N_3666,N_3495,N_3450);
nor U3667 (N_3667,N_3490,N_3439);
xor U3668 (N_3668,N_3429,N_3472);
or U3669 (N_3669,N_3507,N_3401);
nand U3670 (N_3670,N_3412,N_3431);
and U3671 (N_3671,N_3519,N_3579);
xnor U3672 (N_3672,N_3492,N_3514);
or U3673 (N_3673,N_3513,N_3520);
and U3674 (N_3674,N_3496,N_3421);
and U3675 (N_3675,N_3432,N_3463);
nand U3676 (N_3676,N_3594,N_3404);
and U3677 (N_3677,N_3485,N_3487);
xnor U3678 (N_3678,N_3591,N_3489);
nand U3679 (N_3679,N_3580,N_3477);
or U3680 (N_3680,N_3577,N_3521);
nand U3681 (N_3681,N_3483,N_3499);
nand U3682 (N_3682,N_3534,N_3504);
or U3683 (N_3683,N_3555,N_3584);
nand U3684 (N_3684,N_3409,N_3493);
or U3685 (N_3685,N_3553,N_3482);
and U3686 (N_3686,N_3531,N_3582);
or U3687 (N_3687,N_3456,N_3554);
or U3688 (N_3688,N_3523,N_3571);
nor U3689 (N_3689,N_3537,N_3533);
xor U3690 (N_3690,N_3543,N_3593);
and U3691 (N_3691,N_3548,N_3510);
or U3692 (N_3692,N_3407,N_3497);
and U3693 (N_3693,N_3422,N_3414);
and U3694 (N_3694,N_3440,N_3436);
nand U3695 (N_3695,N_3508,N_3486);
xor U3696 (N_3696,N_3511,N_3416);
nor U3697 (N_3697,N_3406,N_3517);
and U3698 (N_3698,N_3588,N_3459);
and U3699 (N_3699,N_3565,N_3536);
or U3700 (N_3700,N_3448,N_3474);
nand U3701 (N_3701,N_3514,N_3583);
nor U3702 (N_3702,N_3413,N_3526);
nor U3703 (N_3703,N_3559,N_3549);
nor U3704 (N_3704,N_3503,N_3426);
and U3705 (N_3705,N_3484,N_3434);
xnor U3706 (N_3706,N_3465,N_3595);
and U3707 (N_3707,N_3459,N_3440);
nand U3708 (N_3708,N_3534,N_3555);
xor U3709 (N_3709,N_3524,N_3484);
nor U3710 (N_3710,N_3595,N_3551);
nand U3711 (N_3711,N_3556,N_3576);
nand U3712 (N_3712,N_3464,N_3452);
nand U3713 (N_3713,N_3537,N_3444);
or U3714 (N_3714,N_3400,N_3406);
nand U3715 (N_3715,N_3562,N_3462);
nor U3716 (N_3716,N_3432,N_3443);
or U3717 (N_3717,N_3435,N_3516);
xor U3718 (N_3718,N_3410,N_3477);
nand U3719 (N_3719,N_3479,N_3552);
nand U3720 (N_3720,N_3470,N_3533);
nand U3721 (N_3721,N_3536,N_3538);
nand U3722 (N_3722,N_3489,N_3518);
or U3723 (N_3723,N_3406,N_3506);
nor U3724 (N_3724,N_3419,N_3512);
and U3725 (N_3725,N_3470,N_3515);
or U3726 (N_3726,N_3558,N_3446);
xor U3727 (N_3727,N_3567,N_3558);
xor U3728 (N_3728,N_3590,N_3432);
or U3729 (N_3729,N_3478,N_3413);
or U3730 (N_3730,N_3522,N_3530);
nor U3731 (N_3731,N_3404,N_3434);
xor U3732 (N_3732,N_3517,N_3476);
nor U3733 (N_3733,N_3532,N_3428);
and U3734 (N_3734,N_3539,N_3444);
nor U3735 (N_3735,N_3579,N_3496);
or U3736 (N_3736,N_3598,N_3536);
nor U3737 (N_3737,N_3592,N_3550);
or U3738 (N_3738,N_3498,N_3513);
nand U3739 (N_3739,N_3413,N_3488);
nand U3740 (N_3740,N_3455,N_3547);
xor U3741 (N_3741,N_3477,N_3541);
xnor U3742 (N_3742,N_3408,N_3466);
and U3743 (N_3743,N_3437,N_3425);
xor U3744 (N_3744,N_3479,N_3421);
and U3745 (N_3745,N_3484,N_3541);
xor U3746 (N_3746,N_3503,N_3575);
nor U3747 (N_3747,N_3439,N_3525);
or U3748 (N_3748,N_3424,N_3493);
and U3749 (N_3749,N_3470,N_3479);
xor U3750 (N_3750,N_3449,N_3594);
nor U3751 (N_3751,N_3564,N_3423);
nand U3752 (N_3752,N_3593,N_3549);
xnor U3753 (N_3753,N_3524,N_3585);
nor U3754 (N_3754,N_3488,N_3535);
nor U3755 (N_3755,N_3469,N_3439);
xor U3756 (N_3756,N_3408,N_3503);
or U3757 (N_3757,N_3493,N_3442);
nand U3758 (N_3758,N_3555,N_3592);
nand U3759 (N_3759,N_3574,N_3483);
xor U3760 (N_3760,N_3450,N_3463);
xor U3761 (N_3761,N_3580,N_3405);
and U3762 (N_3762,N_3456,N_3596);
or U3763 (N_3763,N_3492,N_3444);
nor U3764 (N_3764,N_3479,N_3519);
or U3765 (N_3765,N_3524,N_3499);
nand U3766 (N_3766,N_3448,N_3590);
nor U3767 (N_3767,N_3414,N_3421);
nand U3768 (N_3768,N_3579,N_3430);
or U3769 (N_3769,N_3491,N_3518);
nor U3770 (N_3770,N_3521,N_3592);
and U3771 (N_3771,N_3514,N_3413);
or U3772 (N_3772,N_3403,N_3477);
nand U3773 (N_3773,N_3475,N_3487);
xnor U3774 (N_3774,N_3526,N_3561);
and U3775 (N_3775,N_3508,N_3529);
and U3776 (N_3776,N_3526,N_3483);
and U3777 (N_3777,N_3400,N_3402);
and U3778 (N_3778,N_3423,N_3589);
or U3779 (N_3779,N_3533,N_3423);
or U3780 (N_3780,N_3583,N_3436);
or U3781 (N_3781,N_3451,N_3551);
xor U3782 (N_3782,N_3583,N_3550);
or U3783 (N_3783,N_3513,N_3577);
xnor U3784 (N_3784,N_3559,N_3522);
nand U3785 (N_3785,N_3571,N_3485);
nand U3786 (N_3786,N_3457,N_3598);
and U3787 (N_3787,N_3483,N_3475);
and U3788 (N_3788,N_3494,N_3422);
nand U3789 (N_3789,N_3442,N_3587);
and U3790 (N_3790,N_3445,N_3521);
nand U3791 (N_3791,N_3524,N_3459);
nand U3792 (N_3792,N_3496,N_3581);
nand U3793 (N_3793,N_3541,N_3510);
and U3794 (N_3794,N_3524,N_3460);
and U3795 (N_3795,N_3421,N_3528);
nor U3796 (N_3796,N_3496,N_3417);
or U3797 (N_3797,N_3443,N_3465);
and U3798 (N_3798,N_3422,N_3535);
xor U3799 (N_3799,N_3514,N_3566);
or U3800 (N_3800,N_3606,N_3722);
or U3801 (N_3801,N_3608,N_3718);
xnor U3802 (N_3802,N_3648,N_3702);
or U3803 (N_3803,N_3721,N_3689);
nand U3804 (N_3804,N_3677,N_3715);
nand U3805 (N_3805,N_3610,N_3766);
or U3806 (N_3806,N_3651,N_3796);
xnor U3807 (N_3807,N_3773,N_3788);
or U3808 (N_3808,N_3607,N_3734);
nor U3809 (N_3809,N_3764,N_3793);
or U3810 (N_3810,N_3614,N_3641);
or U3811 (N_3811,N_3778,N_3618);
nand U3812 (N_3812,N_3740,N_3629);
nor U3813 (N_3813,N_3631,N_3728);
and U3814 (N_3814,N_3682,N_3753);
nor U3815 (N_3815,N_3635,N_3794);
nand U3816 (N_3816,N_3647,N_3627);
and U3817 (N_3817,N_3643,N_3785);
nor U3818 (N_3818,N_3645,N_3748);
and U3819 (N_3819,N_3638,N_3704);
nor U3820 (N_3820,N_3727,N_3700);
and U3821 (N_3821,N_3665,N_3792);
nor U3822 (N_3822,N_3604,N_3630);
nand U3823 (N_3823,N_3752,N_3768);
nor U3824 (N_3824,N_3632,N_3649);
and U3825 (N_3825,N_3655,N_3725);
xnor U3826 (N_3826,N_3795,N_3737);
nand U3827 (N_3827,N_3771,N_3667);
xor U3828 (N_3828,N_3683,N_3688);
or U3829 (N_3829,N_3776,N_3676);
or U3830 (N_3830,N_3664,N_3690);
and U3831 (N_3831,N_3675,N_3692);
and U3832 (N_3832,N_3733,N_3782);
and U3833 (N_3833,N_3787,N_3637);
nor U3834 (N_3834,N_3626,N_3786);
or U3835 (N_3835,N_3662,N_3747);
or U3836 (N_3836,N_3713,N_3731);
nand U3837 (N_3837,N_3730,N_3741);
xnor U3838 (N_3838,N_3685,N_3745);
nand U3839 (N_3839,N_3628,N_3729);
and U3840 (N_3840,N_3761,N_3777);
nor U3841 (N_3841,N_3671,N_3710);
and U3842 (N_3842,N_3603,N_3661);
nor U3843 (N_3843,N_3652,N_3620);
nor U3844 (N_3844,N_3789,N_3686);
and U3845 (N_3845,N_3640,N_3757);
and U3846 (N_3846,N_3749,N_3624);
nand U3847 (N_3847,N_3611,N_3654);
and U3848 (N_3848,N_3619,N_3657);
nor U3849 (N_3849,N_3775,N_3743);
nand U3850 (N_3850,N_3760,N_3670);
xnor U3851 (N_3851,N_3767,N_3622);
xnor U3852 (N_3852,N_3779,N_3623);
nor U3853 (N_3853,N_3744,N_3724);
xnor U3854 (N_3854,N_3717,N_3696);
xor U3855 (N_3855,N_3668,N_3751);
and U3856 (N_3856,N_3765,N_3798);
or U3857 (N_3857,N_3646,N_3759);
nand U3858 (N_3858,N_3673,N_3781);
nand U3859 (N_3859,N_3780,N_3672);
nand U3860 (N_3860,N_3644,N_3660);
or U3861 (N_3861,N_3625,N_3663);
and U3862 (N_3862,N_3774,N_3684);
or U3863 (N_3863,N_3707,N_3600);
xor U3864 (N_3864,N_3742,N_3754);
nor U3865 (N_3865,N_3732,N_3790);
and U3866 (N_3866,N_3613,N_3612);
or U3867 (N_3867,N_3750,N_3706);
or U3868 (N_3868,N_3634,N_3695);
nor U3869 (N_3869,N_3756,N_3712);
and U3870 (N_3870,N_3615,N_3698);
xnor U3871 (N_3871,N_3714,N_3770);
nand U3872 (N_3872,N_3617,N_3679);
nor U3873 (N_3873,N_3769,N_3758);
nand U3874 (N_3874,N_3658,N_3735);
and U3875 (N_3875,N_3784,N_3659);
nand U3876 (N_3876,N_3797,N_3791);
and U3877 (N_3877,N_3653,N_3697);
nand U3878 (N_3878,N_3726,N_3694);
or U3879 (N_3879,N_3674,N_3738);
and U3880 (N_3880,N_3719,N_3763);
and U3881 (N_3881,N_3709,N_3711);
nor U3882 (N_3882,N_3691,N_3636);
nand U3883 (N_3883,N_3605,N_3783);
xnor U3884 (N_3884,N_3723,N_3687);
and U3885 (N_3885,N_3708,N_3609);
and U3886 (N_3886,N_3746,N_3602);
and U3887 (N_3887,N_3720,N_3703);
nor U3888 (N_3888,N_3701,N_3716);
or U3889 (N_3889,N_3799,N_3699);
nor U3890 (N_3890,N_3633,N_3705);
or U3891 (N_3891,N_3681,N_3736);
nor U3892 (N_3892,N_3669,N_3680);
and U3893 (N_3893,N_3755,N_3616);
xnor U3894 (N_3894,N_3762,N_3601);
nand U3895 (N_3895,N_3678,N_3666);
or U3896 (N_3896,N_3739,N_3772);
or U3897 (N_3897,N_3639,N_3621);
nand U3898 (N_3898,N_3693,N_3642);
nand U3899 (N_3899,N_3650,N_3656);
nand U3900 (N_3900,N_3791,N_3696);
xor U3901 (N_3901,N_3742,N_3757);
nor U3902 (N_3902,N_3724,N_3699);
nor U3903 (N_3903,N_3628,N_3780);
and U3904 (N_3904,N_3763,N_3762);
nor U3905 (N_3905,N_3601,N_3689);
xnor U3906 (N_3906,N_3640,N_3766);
xor U3907 (N_3907,N_3685,N_3699);
xnor U3908 (N_3908,N_3756,N_3656);
and U3909 (N_3909,N_3788,N_3668);
or U3910 (N_3910,N_3791,N_3669);
xnor U3911 (N_3911,N_3647,N_3653);
and U3912 (N_3912,N_3619,N_3780);
nor U3913 (N_3913,N_3717,N_3713);
xor U3914 (N_3914,N_3793,N_3753);
nor U3915 (N_3915,N_3775,N_3794);
xor U3916 (N_3916,N_3774,N_3647);
nand U3917 (N_3917,N_3685,N_3737);
nor U3918 (N_3918,N_3723,N_3758);
xnor U3919 (N_3919,N_3688,N_3643);
nand U3920 (N_3920,N_3702,N_3798);
nand U3921 (N_3921,N_3698,N_3750);
or U3922 (N_3922,N_3753,N_3672);
nand U3923 (N_3923,N_3662,N_3633);
and U3924 (N_3924,N_3779,N_3766);
nand U3925 (N_3925,N_3729,N_3664);
xor U3926 (N_3926,N_3719,N_3762);
and U3927 (N_3927,N_3689,N_3637);
and U3928 (N_3928,N_3700,N_3674);
and U3929 (N_3929,N_3635,N_3649);
or U3930 (N_3930,N_3687,N_3770);
or U3931 (N_3931,N_3797,N_3679);
xnor U3932 (N_3932,N_3730,N_3661);
nor U3933 (N_3933,N_3730,N_3667);
and U3934 (N_3934,N_3717,N_3608);
or U3935 (N_3935,N_3672,N_3707);
and U3936 (N_3936,N_3672,N_3772);
nor U3937 (N_3937,N_3698,N_3681);
or U3938 (N_3938,N_3640,N_3671);
or U3939 (N_3939,N_3707,N_3775);
nor U3940 (N_3940,N_3692,N_3738);
and U3941 (N_3941,N_3789,N_3775);
nand U3942 (N_3942,N_3631,N_3619);
xor U3943 (N_3943,N_3692,N_3772);
nand U3944 (N_3944,N_3692,N_3741);
nand U3945 (N_3945,N_3722,N_3781);
or U3946 (N_3946,N_3635,N_3613);
or U3947 (N_3947,N_3741,N_3645);
nor U3948 (N_3948,N_3636,N_3723);
nand U3949 (N_3949,N_3672,N_3600);
xor U3950 (N_3950,N_3736,N_3749);
nor U3951 (N_3951,N_3753,N_3604);
nand U3952 (N_3952,N_3719,N_3780);
nor U3953 (N_3953,N_3639,N_3739);
or U3954 (N_3954,N_3677,N_3705);
nand U3955 (N_3955,N_3738,N_3605);
and U3956 (N_3956,N_3600,N_3601);
and U3957 (N_3957,N_3673,N_3708);
nor U3958 (N_3958,N_3631,N_3691);
and U3959 (N_3959,N_3798,N_3668);
and U3960 (N_3960,N_3763,N_3720);
nor U3961 (N_3961,N_3714,N_3753);
xor U3962 (N_3962,N_3741,N_3696);
and U3963 (N_3963,N_3604,N_3769);
xor U3964 (N_3964,N_3665,N_3631);
and U3965 (N_3965,N_3793,N_3650);
nand U3966 (N_3966,N_3657,N_3666);
nand U3967 (N_3967,N_3715,N_3618);
and U3968 (N_3968,N_3719,N_3684);
and U3969 (N_3969,N_3668,N_3725);
nand U3970 (N_3970,N_3791,N_3658);
and U3971 (N_3971,N_3664,N_3771);
xor U3972 (N_3972,N_3643,N_3793);
xor U3973 (N_3973,N_3722,N_3649);
nor U3974 (N_3974,N_3684,N_3770);
nor U3975 (N_3975,N_3775,N_3763);
or U3976 (N_3976,N_3767,N_3641);
nand U3977 (N_3977,N_3601,N_3724);
and U3978 (N_3978,N_3785,N_3618);
nor U3979 (N_3979,N_3646,N_3733);
or U3980 (N_3980,N_3675,N_3770);
or U3981 (N_3981,N_3781,N_3798);
nor U3982 (N_3982,N_3792,N_3715);
nor U3983 (N_3983,N_3764,N_3723);
nor U3984 (N_3984,N_3696,N_3706);
nand U3985 (N_3985,N_3643,N_3759);
nand U3986 (N_3986,N_3675,N_3704);
nand U3987 (N_3987,N_3644,N_3782);
or U3988 (N_3988,N_3658,N_3745);
nor U3989 (N_3989,N_3684,N_3611);
nor U3990 (N_3990,N_3761,N_3731);
and U3991 (N_3991,N_3633,N_3669);
nor U3992 (N_3992,N_3737,N_3659);
and U3993 (N_3993,N_3695,N_3664);
and U3994 (N_3994,N_3730,N_3717);
nand U3995 (N_3995,N_3705,N_3616);
xnor U3996 (N_3996,N_3720,N_3710);
nor U3997 (N_3997,N_3658,N_3615);
xor U3998 (N_3998,N_3686,N_3656);
nand U3999 (N_3999,N_3780,N_3730);
xnor U4000 (N_4000,N_3809,N_3868);
nand U4001 (N_4001,N_3811,N_3840);
nor U4002 (N_4002,N_3888,N_3835);
and U4003 (N_4003,N_3997,N_3900);
or U4004 (N_4004,N_3825,N_3837);
nor U4005 (N_4005,N_3947,N_3901);
or U4006 (N_4006,N_3826,N_3818);
or U4007 (N_4007,N_3864,N_3934);
nor U4008 (N_4008,N_3971,N_3824);
and U4009 (N_4009,N_3832,N_3904);
xor U4010 (N_4010,N_3865,N_3965);
or U4011 (N_4011,N_3984,N_3948);
nand U4012 (N_4012,N_3875,N_3960);
xor U4013 (N_4013,N_3909,N_3921);
or U4014 (N_4014,N_3802,N_3863);
and U4015 (N_4015,N_3967,N_3869);
xor U4016 (N_4016,N_3906,N_3895);
nor U4017 (N_4017,N_3988,N_3859);
xnor U4018 (N_4018,N_3985,N_3913);
and U4019 (N_4019,N_3827,N_3970);
xor U4020 (N_4020,N_3949,N_3929);
nand U4021 (N_4021,N_3801,N_3989);
nand U4022 (N_4022,N_3852,N_3890);
xnor U4023 (N_4023,N_3936,N_3963);
or U4024 (N_4024,N_3952,N_3958);
nor U4025 (N_4025,N_3870,N_3871);
xor U4026 (N_4026,N_3814,N_3849);
or U4027 (N_4027,N_3966,N_3907);
xor U4028 (N_4028,N_3816,N_3831);
or U4029 (N_4029,N_3881,N_3896);
nand U4030 (N_4030,N_3830,N_3920);
and U4031 (N_4031,N_3994,N_3819);
nor U4032 (N_4032,N_3919,N_3995);
and U4033 (N_4033,N_3923,N_3918);
or U4034 (N_4034,N_3893,N_3926);
or U4035 (N_4035,N_3854,N_3841);
nor U4036 (N_4036,N_3883,N_3932);
nor U4037 (N_4037,N_3822,N_3861);
xnor U4038 (N_4038,N_3980,N_3823);
xnor U4039 (N_4039,N_3954,N_3815);
nand U4040 (N_4040,N_3806,N_3856);
and U4041 (N_4041,N_3813,N_3891);
xnor U4042 (N_4042,N_3978,N_3858);
xnor U4043 (N_4043,N_3993,N_3999);
or U4044 (N_4044,N_3836,N_3857);
nand U4045 (N_4045,N_3927,N_3817);
nor U4046 (N_4046,N_3944,N_3860);
nand U4047 (N_4047,N_3987,N_3853);
xnor U4048 (N_4048,N_3946,N_3898);
nand U4049 (N_4049,N_3867,N_3940);
and U4050 (N_4050,N_3964,N_3911);
nand U4051 (N_4051,N_3979,N_3962);
nor U4052 (N_4052,N_3955,N_3829);
or U4053 (N_4053,N_3845,N_3957);
or U4054 (N_4054,N_3931,N_3959);
and U4055 (N_4055,N_3945,N_3892);
or U4056 (N_4056,N_3847,N_3937);
nand U4057 (N_4057,N_3807,N_3839);
and U4058 (N_4058,N_3878,N_3848);
or U4059 (N_4059,N_3996,N_3876);
nand U4060 (N_4060,N_3938,N_3922);
nand U4061 (N_4061,N_3976,N_3956);
nand U4062 (N_4062,N_3917,N_3903);
or U4063 (N_4063,N_3973,N_3897);
or U4064 (N_4064,N_3834,N_3866);
nor U4065 (N_4065,N_3975,N_3990);
nand U4066 (N_4066,N_3977,N_3983);
nor U4067 (N_4067,N_3916,N_3969);
nand U4068 (N_4068,N_3981,N_3879);
xor U4069 (N_4069,N_3915,N_3991);
nand U4070 (N_4070,N_3886,N_3808);
or U4071 (N_4071,N_3972,N_3914);
xor U4072 (N_4072,N_3974,N_3910);
or U4073 (N_4073,N_3885,N_3982);
xnor U4074 (N_4074,N_3924,N_3855);
xnor U4075 (N_4075,N_3842,N_3905);
or U4076 (N_4076,N_3874,N_3992);
and U4077 (N_4077,N_3862,N_3908);
xnor U4078 (N_4078,N_3925,N_3850);
nor U4079 (N_4079,N_3912,N_3899);
nor U4080 (N_4080,N_3873,N_3943);
and U4081 (N_4081,N_3953,N_3838);
xor U4082 (N_4082,N_3902,N_3986);
nor U4083 (N_4083,N_3880,N_3803);
xnor U4084 (N_4084,N_3846,N_3805);
and U4085 (N_4085,N_3933,N_3942);
nand U4086 (N_4086,N_3844,N_3887);
and U4087 (N_4087,N_3843,N_3968);
nor U4088 (N_4088,N_3872,N_3882);
nand U4089 (N_4089,N_3930,N_3894);
nand U4090 (N_4090,N_3812,N_3935);
nand U4091 (N_4091,N_3998,N_3928);
and U4092 (N_4092,N_3950,N_3851);
or U4093 (N_4093,N_3889,N_3939);
and U4094 (N_4094,N_3810,N_3800);
or U4095 (N_4095,N_3941,N_3833);
xnor U4096 (N_4096,N_3877,N_3820);
xnor U4097 (N_4097,N_3951,N_3804);
and U4098 (N_4098,N_3821,N_3884);
nand U4099 (N_4099,N_3828,N_3961);
and U4100 (N_4100,N_3892,N_3907);
nor U4101 (N_4101,N_3907,N_3899);
and U4102 (N_4102,N_3840,N_3939);
nor U4103 (N_4103,N_3893,N_3970);
nor U4104 (N_4104,N_3850,N_3858);
or U4105 (N_4105,N_3977,N_3932);
nand U4106 (N_4106,N_3906,N_3863);
xor U4107 (N_4107,N_3916,N_3967);
and U4108 (N_4108,N_3839,N_3909);
nand U4109 (N_4109,N_3823,N_3968);
and U4110 (N_4110,N_3867,N_3903);
nand U4111 (N_4111,N_3867,N_3941);
xor U4112 (N_4112,N_3829,N_3957);
or U4113 (N_4113,N_3921,N_3914);
nor U4114 (N_4114,N_3932,N_3827);
and U4115 (N_4115,N_3906,N_3828);
or U4116 (N_4116,N_3863,N_3853);
or U4117 (N_4117,N_3813,N_3810);
xnor U4118 (N_4118,N_3803,N_3929);
and U4119 (N_4119,N_3896,N_3869);
or U4120 (N_4120,N_3976,N_3932);
and U4121 (N_4121,N_3814,N_3972);
and U4122 (N_4122,N_3963,N_3913);
nand U4123 (N_4123,N_3814,N_3894);
or U4124 (N_4124,N_3996,N_3807);
nand U4125 (N_4125,N_3824,N_3919);
nand U4126 (N_4126,N_3892,N_3820);
xnor U4127 (N_4127,N_3838,N_3907);
nand U4128 (N_4128,N_3876,N_3806);
or U4129 (N_4129,N_3959,N_3900);
or U4130 (N_4130,N_3924,N_3800);
or U4131 (N_4131,N_3915,N_3977);
xnor U4132 (N_4132,N_3948,N_3861);
nor U4133 (N_4133,N_3809,N_3944);
xnor U4134 (N_4134,N_3868,N_3994);
nand U4135 (N_4135,N_3917,N_3939);
or U4136 (N_4136,N_3956,N_3988);
and U4137 (N_4137,N_3846,N_3828);
xor U4138 (N_4138,N_3935,N_3869);
and U4139 (N_4139,N_3870,N_3977);
nand U4140 (N_4140,N_3882,N_3809);
or U4141 (N_4141,N_3807,N_3952);
nand U4142 (N_4142,N_3985,N_3937);
and U4143 (N_4143,N_3978,N_3800);
and U4144 (N_4144,N_3890,N_3936);
and U4145 (N_4145,N_3854,N_3939);
nand U4146 (N_4146,N_3889,N_3927);
xor U4147 (N_4147,N_3888,N_3831);
nor U4148 (N_4148,N_3997,N_3880);
xnor U4149 (N_4149,N_3959,N_3910);
or U4150 (N_4150,N_3833,N_3938);
xnor U4151 (N_4151,N_3836,N_3826);
xor U4152 (N_4152,N_3986,N_3917);
nor U4153 (N_4153,N_3902,N_3953);
or U4154 (N_4154,N_3863,N_3845);
and U4155 (N_4155,N_3860,N_3988);
nor U4156 (N_4156,N_3858,N_3840);
and U4157 (N_4157,N_3939,N_3967);
xnor U4158 (N_4158,N_3968,N_3804);
and U4159 (N_4159,N_3884,N_3957);
and U4160 (N_4160,N_3892,N_3894);
nand U4161 (N_4161,N_3805,N_3815);
or U4162 (N_4162,N_3835,N_3804);
nor U4163 (N_4163,N_3965,N_3906);
nand U4164 (N_4164,N_3858,N_3849);
nand U4165 (N_4165,N_3800,N_3827);
and U4166 (N_4166,N_3949,N_3922);
or U4167 (N_4167,N_3831,N_3913);
or U4168 (N_4168,N_3858,N_3958);
nand U4169 (N_4169,N_3911,N_3991);
or U4170 (N_4170,N_3917,N_3823);
or U4171 (N_4171,N_3868,N_3996);
and U4172 (N_4172,N_3842,N_3901);
or U4173 (N_4173,N_3845,N_3890);
or U4174 (N_4174,N_3936,N_3977);
and U4175 (N_4175,N_3925,N_3878);
or U4176 (N_4176,N_3820,N_3832);
nand U4177 (N_4177,N_3865,N_3832);
nand U4178 (N_4178,N_3849,N_3865);
nor U4179 (N_4179,N_3961,N_3984);
nand U4180 (N_4180,N_3857,N_3889);
nor U4181 (N_4181,N_3854,N_3934);
xor U4182 (N_4182,N_3814,N_3882);
nor U4183 (N_4183,N_3930,N_3836);
or U4184 (N_4184,N_3808,N_3918);
nand U4185 (N_4185,N_3909,N_3803);
and U4186 (N_4186,N_3950,N_3968);
or U4187 (N_4187,N_3856,N_3952);
xnor U4188 (N_4188,N_3873,N_3933);
or U4189 (N_4189,N_3978,N_3817);
and U4190 (N_4190,N_3822,N_3815);
nand U4191 (N_4191,N_3993,N_3868);
or U4192 (N_4192,N_3803,N_3995);
nor U4193 (N_4193,N_3901,N_3827);
or U4194 (N_4194,N_3907,N_3941);
or U4195 (N_4195,N_3871,N_3914);
and U4196 (N_4196,N_3946,N_3800);
nand U4197 (N_4197,N_3827,N_3938);
nor U4198 (N_4198,N_3879,N_3875);
nor U4199 (N_4199,N_3989,N_3955);
xnor U4200 (N_4200,N_4077,N_4144);
nand U4201 (N_4201,N_4161,N_4007);
nor U4202 (N_4202,N_4198,N_4132);
and U4203 (N_4203,N_4047,N_4083);
or U4204 (N_4204,N_4192,N_4041);
and U4205 (N_4205,N_4158,N_4151);
and U4206 (N_4206,N_4062,N_4082);
xnor U4207 (N_4207,N_4130,N_4061);
nand U4208 (N_4208,N_4084,N_4039);
nor U4209 (N_4209,N_4067,N_4168);
nor U4210 (N_4210,N_4054,N_4069);
nand U4211 (N_4211,N_4143,N_4102);
nand U4212 (N_4212,N_4066,N_4169);
and U4213 (N_4213,N_4133,N_4098);
nor U4214 (N_4214,N_4090,N_4197);
or U4215 (N_4215,N_4103,N_4172);
nand U4216 (N_4216,N_4073,N_4194);
nand U4217 (N_4217,N_4121,N_4107);
xnor U4218 (N_4218,N_4049,N_4125);
nor U4219 (N_4219,N_4085,N_4115);
nor U4220 (N_4220,N_4053,N_4150);
nor U4221 (N_4221,N_4068,N_4124);
and U4222 (N_4222,N_4117,N_4114);
and U4223 (N_4223,N_4092,N_4183);
nor U4224 (N_4224,N_4040,N_4142);
nor U4225 (N_4225,N_4081,N_4109);
nor U4226 (N_4226,N_4190,N_4155);
nor U4227 (N_4227,N_4071,N_4187);
and U4228 (N_4228,N_4008,N_4064);
and U4229 (N_4229,N_4112,N_4126);
and U4230 (N_4230,N_4046,N_4023);
and U4231 (N_4231,N_4159,N_4051);
xor U4232 (N_4232,N_4145,N_4036);
xor U4233 (N_4233,N_4113,N_4011);
and U4234 (N_4234,N_4122,N_4178);
and U4235 (N_4235,N_4079,N_4182);
or U4236 (N_4236,N_4184,N_4157);
or U4237 (N_4237,N_4088,N_4152);
xor U4238 (N_4238,N_4119,N_4087);
or U4239 (N_4239,N_4111,N_4170);
nand U4240 (N_4240,N_4013,N_4027);
and U4241 (N_4241,N_4010,N_4193);
nand U4242 (N_4242,N_4163,N_4186);
nand U4243 (N_4243,N_4137,N_4091);
and U4244 (N_4244,N_4162,N_4116);
xnor U4245 (N_4245,N_4086,N_4005);
and U4246 (N_4246,N_4025,N_4056);
nand U4247 (N_4247,N_4100,N_4000);
nand U4248 (N_4248,N_4129,N_4038);
or U4249 (N_4249,N_4120,N_4075);
nor U4250 (N_4250,N_4055,N_4148);
nor U4251 (N_4251,N_4136,N_4188);
nand U4252 (N_4252,N_4195,N_4022);
xor U4253 (N_4253,N_4096,N_4180);
or U4254 (N_4254,N_4065,N_4101);
xnor U4255 (N_4255,N_4089,N_4181);
nor U4256 (N_4256,N_4189,N_4030);
xnor U4257 (N_4257,N_4001,N_4043);
nor U4258 (N_4258,N_4149,N_4108);
or U4259 (N_4259,N_4104,N_4017);
nor U4260 (N_4260,N_4035,N_4072);
and U4261 (N_4261,N_4106,N_4070);
nand U4262 (N_4262,N_4135,N_4174);
xor U4263 (N_4263,N_4019,N_4153);
and U4264 (N_4264,N_4063,N_4110);
xor U4265 (N_4265,N_4080,N_4002);
or U4266 (N_4266,N_4052,N_4097);
xor U4267 (N_4267,N_4050,N_4141);
or U4268 (N_4268,N_4128,N_4015);
or U4269 (N_4269,N_4029,N_4045);
xnor U4270 (N_4270,N_4127,N_4176);
nand U4271 (N_4271,N_4016,N_4026);
nand U4272 (N_4272,N_4160,N_4191);
nand U4273 (N_4273,N_4134,N_4093);
xnor U4274 (N_4274,N_4076,N_4199);
or U4275 (N_4275,N_4164,N_4033);
xor U4276 (N_4276,N_4078,N_4014);
xnor U4277 (N_4277,N_4059,N_4179);
nand U4278 (N_4278,N_4037,N_4118);
and U4279 (N_4279,N_4074,N_4031);
nor U4280 (N_4280,N_4020,N_4154);
or U4281 (N_4281,N_4166,N_4095);
nor U4282 (N_4282,N_4060,N_4139);
xnor U4283 (N_4283,N_4185,N_4028);
nand U4284 (N_4284,N_4003,N_4196);
nor U4285 (N_4285,N_4156,N_4048);
and U4286 (N_4286,N_4099,N_4024);
nor U4287 (N_4287,N_4021,N_4173);
or U4288 (N_4288,N_4044,N_4131);
or U4289 (N_4289,N_4012,N_4034);
xnor U4290 (N_4290,N_4004,N_4171);
xor U4291 (N_4291,N_4140,N_4165);
and U4292 (N_4292,N_4138,N_4009);
nor U4293 (N_4293,N_4123,N_4105);
nor U4294 (N_4294,N_4175,N_4177);
or U4295 (N_4295,N_4032,N_4057);
or U4296 (N_4296,N_4147,N_4094);
or U4297 (N_4297,N_4018,N_4146);
nand U4298 (N_4298,N_4042,N_4167);
and U4299 (N_4299,N_4006,N_4058);
and U4300 (N_4300,N_4009,N_4074);
nand U4301 (N_4301,N_4176,N_4164);
or U4302 (N_4302,N_4158,N_4000);
nor U4303 (N_4303,N_4035,N_4094);
or U4304 (N_4304,N_4162,N_4155);
nor U4305 (N_4305,N_4039,N_4024);
nand U4306 (N_4306,N_4059,N_4001);
and U4307 (N_4307,N_4092,N_4149);
nand U4308 (N_4308,N_4103,N_4011);
xnor U4309 (N_4309,N_4044,N_4169);
or U4310 (N_4310,N_4109,N_4119);
nand U4311 (N_4311,N_4125,N_4071);
nor U4312 (N_4312,N_4051,N_4195);
nor U4313 (N_4313,N_4026,N_4046);
nor U4314 (N_4314,N_4092,N_4011);
nand U4315 (N_4315,N_4127,N_4080);
nor U4316 (N_4316,N_4097,N_4174);
and U4317 (N_4317,N_4177,N_4014);
nor U4318 (N_4318,N_4159,N_4180);
and U4319 (N_4319,N_4133,N_4134);
xnor U4320 (N_4320,N_4031,N_4050);
nor U4321 (N_4321,N_4107,N_4017);
nand U4322 (N_4322,N_4063,N_4038);
nor U4323 (N_4323,N_4085,N_4061);
nand U4324 (N_4324,N_4011,N_4087);
nand U4325 (N_4325,N_4178,N_4044);
or U4326 (N_4326,N_4195,N_4188);
nand U4327 (N_4327,N_4149,N_4095);
and U4328 (N_4328,N_4039,N_4056);
nor U4329 (N_4329,N_4145,N_4124);
nand U4330 (N_4330,N_4154,N_4139);
or U4331 (N_4331,N_4034,N_4110);
xor U4332 (N_4332,N_4049,N_4134);
or U4333 (N_4333,N_4172,N_4050);
or U4334 (N_4334,N_4135,N_4180);
and U4335 (N_4335,N_4115,N_4042);
xnor U4336 (N_4336,N_4113,N_4121);
or U4337 (N_4337,N_4135,N_4178);
xor U4338 (N_4338,N_4049,N_4060);
or U4339 (N_4339,N_4184,N_4102);
or U4340 (N_4340,N_4176,N_4160);
xnor U4341 (N_4341,N_4140,N_4060);
xnor U4342 (N_4342,N_4091,N_4054);
and U4343 (N_4343,N_4021,N_4116);
xor U4344 (N_4344,N_4071,N_4096);
nor U4345 (N_4345,N_4174,N_4033);
nor U4346 (N_4346,N_4061,N_4019);
nand U4347 (N_4347,N_4107,N_4038);
nor U4348 (N_4348,N_4014,N_4082);
and U4349 (N_4349,N_4021,N_4046);
and U4350 (N_4350,N_4087,N_4187);
nor U4351 (N_4351,N_4128,N_4023);
xor U4352 (N_4352,N_4161,N_4149);
or U4353 (N_4353,N_4035,N_4105);
nand U4354 (N_4354,N_4046,N_4095);
xor U4355 (N_4355,N_4159,N_4183);
nand U4356 (N_4356,N_4084,N_4153);
or U4357 (N_4357,N_4027,N_4172);
xor U4358 (N_4358,N_4129,N_4103);
and U4359 (N_4359,N_4080,N_4048);
xnor U4360 (N_4360,N_4171,N_4107);
xnor U4361 (N_4361,N_4020,N_4143);
xnor U4362 (N_4362,N_4157,N_4117);
nand U4363 (N_4363,N_4128,N_4145);
or U4364 (N_4364,N_4009,N_4022);
nor U4365 (N_4365,N_4144,N_4060);
nor U4366 (N_4366,N_4037,N_4082);
and U4367 (N_4367,N_4026,N_4101);
nand U4368 (N_4368,N_4084,N_4149);
nor U4369 (N_4369,N_4143,N_4159);
xnor U4370 (N_4370,N_4020,N_4021);
or U4371 (N_4371,N_4026,N_4065);
nand U4372 (N_4372,N_4053,N_4096);
xor U4373 (N_4373,N_4142,N_4107);
nor U4374 (N_4374,N_4169,N_4128);
nand U4375 (N_4375,N_4096,N_4029);
nand U4376 (N_4376,N_4166,N_4079);
nor U4377 (N_4377,N_4198,N_4117);
nor U4378 (N_4378,N_4124,N_4062);
or U4379 (N_4379,N_4091,N_4093);
nand U4380 (N_4380,N_4044,N_4090);
xor U4381 (N_4381,N_4146,N_4078);
nor U4382 (N_4382,N_4007,N_4160);
xor U4383 (N_4383,N_4164,N_4185);
and U4384 (N_4384,N_4043,N_4106);
xor U4385 (N_4385,N_4043,N_4009);
or U4386 (N_4386,N_4041,N_4107);
xnor U4387 (N_4387,N_4176,N_4130);
xnor U4388 (N_4388,N_4061,N_4107);
or U4389 (N_4389,N_4020,N_4022);
nor U4390 (N_4390,N_4060,N_4013);
nor U4391 (N_4391,N_4110,N_4074);
nand U4392 (N_4392,N_4025,N_4193);
or U4393 (N_4393,N_4069,N_4124);
and U4394 (N_4394,N_4131,N_4046);
nand U4395 (N_4395,N_4182,N_4170);
nor U4396 (N_4396,N_4144,N_4112);
nor U4397 (N_4397,N_4073,N_4172);
or U4398 (N_4398,N_4105,N_4032);
nand U4399 (N_4399,N_4165,N_4087);
and U4400 (N_4400,N_4256,N_4263);
and U4401 (N_4401,N_4227,N_4328);
or U4402 (N_4402,N_4343,N_4281);
or U4403 (N_4403,N_4337,N_4278);
xor U4404 (N_4404,N_4210,N_4232);
nor U4405 (N_4405,N_4384,N_4307);
and U4406 (N_4406,N_4327,N_4303);
or U4407 (N_4407,N_4276,N_4275);
xnor U4408 (N_4408,N_4367,N_4259);
nor U4409 (N_4409,N_4261,N_4368);
or U4410 (N_4410,N_4347,N_4314);
nand U4411 (N_4411,N_4217,N_4308);
and U4412 (N_4412,N_4221,N_4250);
nand U4413 (N_4413,N_4315,N_4224);
xnor U4414 (N_4414,N_4296,N_4331);
and U4415 (N_4415,N_4274,N_4270);
nand U4416 (N_4416,N_4386,N_4234);
or U4417 (N_4417,N_4207,N_4380);
nor U4418 (N_4418,N_4243,N_4372);
xor U4419 (N_4419,N_4216,N_4297);
nor U4420 (N_4420,N_4369,N_4244);
xnor U4421 (N_4421,N_4351,N_4396);
xor U4422 (N_4422,N_4266,N_4313);
nor U4423 (N_4423,N_4371,N_4267);
xor U4424 (N_4424,N_4397,N_4391);
or U4425 (N_4425,N_4346,N_4283);
nand U4426 (N_4426,N_4294,N_4325);
and U4427 (N_4427,N_4302,N_4271);
nor U4428 (N_4428,N_4301,N_4376);
nand U4429 (N_4429,N_4245,N_4357);
nand U4430 (N_4430,N_4335,N_4378);
or U4431 (N_4431,N_4288,N_4203);
xnor U4432 (N_4432,N_4237,N_4353);
nand U4433 (N_4433,N_4280,N_4320);
or U4434 (N_4434,N_4252,N_4238);
and U4435 (N_4435,N_4269,N_4299);
or U4436 (N_4436,N_4338,N_4363);
nand U4437 (N_4437,N_4366,N_4350);
xor U4438 (N_4438,N_4339,N_4392);
and U4439 (N_4439,N_4286,N_4201);
nor U4440 (N_4440,N_4310,N_4390);
nand U4441 (N_4441,N_4379,N_4309);
xor U4442 (N_4442,N_4373,N_4374);
xnor U4443 (N_4443,N_4387,N_4202);
and U4444 (N_4444,N_4300,N_4306);
nor U4445 (N_4445,N_4273,N_4226);
or U4446 (N_4446,N_4362,N_4279);
nand U4447 (N_4447,N_4253,N_4211);
xor U4448 (N_4448,N_4382,N_4388);
nor U4449 (N_4449,N_4355,N_4219);
nand U4450 (N_4450,N_4204,N_4246);
xnor U4451 (N_4451,N_4348,N_4241);
xor U4452 (N_4452,N_4290,N_4289);
nor U4453 (N_4453,N_4236,N_4212);
nor U4454 (N_4454,N_4316,N_4214);
nor U4455 (N_4455,N_4358,N_4282);
and U4456 (N_4456,N_4293,N_4398);
xor U4457 (N_4457,N_4354,N_4342);
and U4458 (N_4458,N_4235,N_4248);
nand U4459 (N_4459,N_4377,N_4240);
or U4460 (N_4460,N_4231,N_4375);
nand U4461 (N_4461,N_4200,N_4319);
or U4462 (N_4462,N_4249,N_4205);
nand U4463 (N_4463,N_4359,N_4260);
xnor U4464 (N_4464,N_4268,N_4361);
nand U4465 (N_4465,N_4365,N_4264);
or U4466 (N_4466,N_4265,N_4277);
nor U4467 (N_4467,N_4364,N_4206);
nor U4468 (N_4468,N_4295,N_4287);
nor U4469 (N_4469,N_4305,N_4333);
xor U4470 (N_4470,N_4330,N_4229);
nand U4471 (N_4471,N_4345,N_4254);
and U4472 (N_4472,N_4218,N_4258);
or U4473 (N_4473,N_4257,N_4322);
and U4474 (N_4474,N_4332,N_4389);
and U4475 (N_4475,N_4208,N_4344);
or U4476 (N_4476,N_4312,N_4399);
and U4477 (N_4477,N_4318,N_4360);
nand U4478 (N_4478,N_4334,N_4213);
xor U4479 (N_4479,N_4395,N_4317);
xor U4480 (N_4480,N_4291,N_4209);
nand U4481 (N_4481,N_4285,N_4341);
xor U4482 (N_4482,N_4215,N_4220);
and U4483 (N_4483,N_4340,N_4222);
nand U4484 (N_4484,N_4394,N_4349);
nor U4485 (N_4485,N_4324,N_4352);
or U4486 (N_4486,N_4304,N_4311);
nor U4487 (N_4487,N_4385,N_4230);
nor U4488 (N_4488,N_4228,N_4272);
xor U4489 (N_4489,N_4242,N_4225);
or U4490 (N_4490,N_4298,N_4255);
or U4491 (N_4491,N_4381,N_4292);
and U4492 (N_4492,N_4262,N_4321);
nor U4493 (N_4493,N_4223,N_4383);
nand U4494 (N_4494,N_4233,N_4326);
nor U4495 (N_4495,N_4329,N_4323);
or U4496 (N_4496,N_4251,N_4247);
nand U4497 (N_4497,N_4370,N_4239);
nor U4498 (N_4498,N_4356,N_4284);
and U4499 (N_4499,N_4393,N_4336);
nand U4500 (N_4500,N_4217,N_4358);
or U4501 (N_4501,N_4242,N_4370);
xnor U4502 (N_4502,N_4320,N_4359);
nor U4503 (N_4503,N_4300,N_4379);
xor U4504 (N_4504,N_4377,N_4243);
and U4505 (N_4505,N_4222,N_4211);
nand U4506 (N_4506,N_4372,N_4310);
xnor U4507 (N_4507,N_4261,N_4353);
nand U4508 (N_4508,N_4350,N_4364);
and U4509 (N_4509,N_4348,N_4336);
xnor U4510 (N_4510,N_4286,N_4397);
or U4511 (N_4511,N_4360,N_4338);
xnor U4512 (N_4512,N_4277,N_4329);
or U4513 (N_4513,N_4366,N_4334);
xor U4514 (N_4514,N_4386,N_4319);
or U4515 (N_4515,N_4315,N_4260);
nor U4516 (N_4516,N_4242,N_4398);
nor U4517 (N_4517,N_4277,N_4261);
nand U4518 (N_4518,N_4210,N_4223);
nor U4519 (N_4519,N_4317,N_4267);
nor U4520 (N_4520,N_4311,N_4367);
nand U4521 (N_4521,N_4316,N_4303);
xnor U4522 (N_4522,N_4311,N_4293);
and U4523 (N_4523,N_4225,N_4343);
xnor U4524 (N_4524,N_4209,N_4207);
nor U4525 (N_4525,N_4241,N_4392);
and U4526 (N_4526,N_4315,N_4261);
or U4527 (N_4527,N_4301,N_4358);
xnor U4528 (N_4528,N_4370,N_4227);
or U4529 (N_4529,N_4227,N_4291);
nand U4530 (N_4530,N_4310,N_4341);
or U4531 (N_4531,N_4365,N_4375);
nand U4532 (N_4532,N_4354,N_4338);
nand U4533 (N_4533,N_4208,N_4336);
or U4534 (N_4534,N_4304,N_4293);
xnor U4535 (N_4535,N_4245,N_4321);
xor U4536 (N_4536,N_4372,N_4327);
or U4537 (N_4537,N_4389,N_4201);
xnor U4538 (N_4538,N_4368,N_4280);
nor U4539 (N_4539,N_4203,N_4222);
and U4540 (N_4540,N_4207,N_4381);
nor U4541 (N_4541,N_4346,N_4251);
or U4542 (N_4542,N_4252,N_4267);
or U4543 (N_4543,N_4266,N_4240);
nor U4544 (N_4544,N_4214,N_4351);
and U4545 (N_4545,N_4256,N_4251);
and U4546 (N_4546,N_4338,N_4234);
or U4547 (N_4547,N_4368,N_4202);
nand U4548 (N_4548,N_4327,N_4398);
nand U4549 (N_4549,N_4216,N_4315);
xnor U4550 (N_4550,N_4255,N_4289);
and U4551 (N_4551,N_4215,N_4244);
nand U4552 (N_4552,N_4383,N_4264);
nor U4553 (N_4553,N_4362,N_4213);
and U4554 (N_4554,N_4264,N_4350);
nand U4555 (N_4555,N_4375,N_4373);
nand U4556 (N_4556,N_4224,N_4387);
xnor U4557 (N_4557,N_4397,N_4268);
nor U4558 (N_4558,N_4284,N_4239);
nor U4559 (N_4559,N_4224,N_4245);
or U4560 (N_4560,N_4396,N_4246);
xnor U4561 (N_4561,N_4213,N_4332);
and U4562 (N_4562,N_4343,N_4243);
or U4563 (N_4563,N_4298,N_4392);
or U4564 (N_4564,N_4286,N_4262);
and U4565 (N_4565,N_4201,N_4203);
and U4566 (N_4566,N_4392,N_4356);
xor U4567 (N_4567,N_4314,N_4359);
and U4568 (N_4568,N_4308,N_4291);
or U4569 (N_4569,N_4311,N_4337);
or U4570 (N_4570,N_4363,N_4221);
xor U4571 (N_4571,N_4377,N_4264);
and U4572 (N_4572,N_4270,N_4338);
nand U4573 (N_4573,N_4311,N_4391);
and U4574 (N_4574,N_4316,N_4339);
and U4575 (N_4575,N_4337,N_4371);
and U4576 (N_4576,N_4286,N_4216);
nand U4577 (N_4577,N_4266,N_4346);
nand U4578 (N_4578,N_4293,N_4240);
nand U4579 (N_4579,N_4394,N_4293);
nor U4580 (N_4580,N_4253,N_4394);
or U4581 (N_4581,N_4260,N_4399);
and U4582 (N_4582,N_4214,N_4296);
nand U4583 (N_4583,N_4355,N_4391);
nor U4584 (N_4584,N_4221,N_4273);
or U4585 (N_4585,N_4202,N_4270);
xnor U4586 (N_4586,N_4397,N_4367);
xnor U4587 (N_4587,N_4322,N_4270);
nor U4588 (N_4588,N_4359,N_4373);
nand U4589 (N_4589,N_4357,N_4356);
xnor U4590 (N_4590,N_4321,N_4388);
nor U4591 (N_4591,N_4284,N_4259);
xor U4592 (N_4592,N_4212,N_4227);
nor U4593 (N_4593,N_4318,N_4335);
nor U4594 (N_4594,N_4358,N_4295);
nor U4595 (N_4595,N_4324,N_4234);
or U4596 (N_4596,N_4250,N_4280);
nand U4597 (N_4597,N_4356,N_4220);
nor U4598 (N_4598,N_4394,N_4371);
nor U4599 (N_4599,N_4362,N_4389);
and U4600 (N_4600,N_4447,N_4489);
and U4601 (N_4601,N_4595,N_4505);
nor U4602 (N_4602,N_4589,N_4484);
nand U4603 (N_4603,N_4526,N_4591);
xor U4604 (N_4604,N_4439,N_4592);
and U4605 (N_4605,N_4535,N_4463);
and U4606 (N_4606,N_4414,N_4593);
and U4607 (N_4607,N_4421,N_4510);
nor U4608 (N_4608,N_4576,N_4423);
nor U4609 (N_4609,N_4415,N_4493);
xnor U4610 (N_4610,N_4467,N_4406);
nand U4611 (N_4611,N_4420,N_4411);
and U4612 (N_4612,N_4405,N_4444);
nor U4613 (N_4613,N_4410,N_4502);
and U4614 (N_4614,N_4494,N_4588);
xor U4615 (N_4615,N_4561,N_4563);
nand U4616 (N_4616,N_4416,N_4582);
and U4617 (N_4617,N_4412,N_4458);
and U4618 (N_4618,N_4516,N_4454);
and U4619 (N_4619,N_4492,N_4441);
xor U4620 (N_4620,N_4513,N_4453);
and U4621 (N_4621,N_4434,N_4557);
or U4622 (N_4622,N_4584,N_4532);
and U4623 (N_4623,N_4597,N_4436);
nor U4624 (N_4624,N_4506,N_4431);
or U4625 (N_4625,N_4417,N_4594);
nand U4626 (N_4626,N_4507,N_4524);
or U4627 (N_4627,N_4586,N_4481);
xnor U4628 (N_4628,N_4583,N_4549);
or U4629 (N_4629,N_4466,N_4459);
xnor U4630 (N_4630,N_4400,N_4501);
nor U4631 (N_4631,N_4473,N_4476);
nor U4632 (N_4632,N_4529,N_4455);
and U4633 (N_4633,N_4518,N_4424);
nor U4634 (N_4634,N_4422,N_4543);
nor U4635 (N_4635,N_4552,N_4512);
nand U4636 (N_4636,N_4440,N_4461);
nand U4637 (N_4637,N_4517,N_4525);
nor U4638 (N_4638,N_4572,N_4490);
or U4639 (N_4639,N_4547,N_4457);
nor U4640 (N_4640,N_4430,N_4475);
nand U4641 (N_4641,N_4564,N_4571);
xor U4642 (N_4642,N_4456,N_4555);
xnor U4643 (N_4643,N_4596,N_4598);
nor U4644 (N_4644,N_4515,N_4565);
nand U4645 (N_4645,N_4465,N_4585);
nor U4646 (N_4646,N_4460,N_4432);
or U4647 (N_4647,N_4581,N_4544);
nand U4648 (N_4648,N_4575,N_4485);
or U4649 (N_4649,N_4504,N_4580);
xnor U4650 (N_4650,N_4542,N_4482);
nor U4651 (N_4651,N_4471,N_4442);
xnor U4652 (N_4652,N_4497,N_4548);
nor U4653 (N_4653,N_4435,N_4537);
and U4654 (N_4654,N_4443,N_4503);
or U4655 (N_4655,N_4401,N_4499);
xor U4656 (N_4656,N_4462,N_4450);
and U4657 (N_4657,N_4578,N_4402);
nand U4658 (N_4658,N_4569,N_4509);
xor U4659 (N_4659,N_4418,N_4469);
and U4660 (N_4660,N_4541,N_4407);
nand U4661 (N_4661,N_4520,N_4496);
or U4662 (N_4662,N_4452,N_4519);
xor U4663 (N_4663,N_4426,N_4464);
xnor U4664 (N_4664,N_4451,N_4546);
or U4665 (N_4665,N_4428,N_4472);
or U4666 (N_4666,N_4508,N_4448);
xor U4667 (N_4667,N_4574,N_4539);
or U4668 (N_4668,N_4403,N_4523);
and U4669 (N_4669,N_4567,N_4545);
nand U4670 (N_4670,N_4533,N_4536);
xnor U4671 (N_4671,N_4554,N_4413);
or U4672 (N_4672,N_4522,N_4570);
xor U4673 (N_4673,N_4553,N_4556);
and U4674 (N_4674,N_4480,N_4425);
nand U4675 (N_4675,N_4573,N_4474);
and U4676 (N_4676,N_4562,N_4551);
nor U4677 (N_4677,N_4478,N_4486);
xor U4678 (N_4678,N_4491,N_4433);
nand U4679 (N_4679,N_4528,N_4540);
and U4680 (N_4680,N_4568,N_4477);
or U4681 (N_4681,N_4579,N_4577);
xnor U4682 (N_4682,N_4483,N_4470);
or U4683 (N_4683,N_4599,N_4498);
nand U4684 (N_4684,N_4419,N_4449);
and U4685 (N_4685,N_4446,N_4495);
nand U4686 (N_4686,N_4429,N_4559);
xnor U4687 (N_4687,N_4511,N_4479);
nand U4688 (N_4688,N_4534,N_4560);
and U4689 (N_4689,N_4500,N_4438);
and U4690 (N_4690,N_4558,N_4404);
and U4691 (N_4691,N_4468,N_4488);
or U4692 (N_4692,N_4550,N_4437);
and U4693 (N_4693,N_4587,N_4566);
nor U4694 (N_4694,N_4445,N_4409);
xor U4695 (N_4695,N_4487,N_4527);
xor U4696 (N_4696,N_4530,N_4427);
xor U4697 (N_4697,N_4538,N_4408);
and U4698 (N_4698,N_4521,N_4590);
xnor U4699 (N_4699,N_4531,N_4514);
and U4700 (N_4700,N_4456,N_4552);
and U4701 (N_4701,N_4491,N_4474);
and U4702 (N_4702,N_4419,N_4496);
or U4703 (N_4703,N_4488,N_4483);
or U4704 (N_4704,N_4467,N_4514);
and U4705 (N_4705,N_4496,N_4483);
and U4706 (N_4706,N_4472,N_4482);
or U4707 (N_4707,N_4445,N_4434);
or U4708 (N_4708,N_4591,N_4521);
or U4709 (N_4709,N_4535,N_4553);
nor U4710 (N_4710,N_4566,N_4408);
and U4711 (N_4711,N_4434,N_4449);
xnor U4712 (N_4712,N_4592,N_4534);
nand U4713 (N_4713,N_4507,N_4572);
xnor U4714 (N_4714,N_4500,N_4528);
nor U4715 (N_4715,N_4479,N_4447);
nand U4716 (N_4716,N_4474,N_4540);
or U4717 (N_4717,N_4458,N_4462);
xor U4718 (N_4718,N_4452,N_4426);
nand U4719 (N_4719,N_4584,N_4540);
and U4720 (N_4720,N_4538,N_4424);
xnor U4721 (N_4721,N_4479,N_4414);
and U4722 (N_4722,N_4479,N_4564);
or U4723 (N_4723,N_4593,N_4503);
and U4724 (N_4724,N_4569,N_4503);
nor U4725 (N_4725,N_4477,N_4472);
or U4726 (N_4726,N_4502,N_4591);
xor U4727 (N_4727,N_4571,N_4497);
nor U4728 (N_4728,N_4486,N_4570);
and U4729 (N_4729,N_4470,N_4445);
or U4730 (N_4730,N_4456,N_4514);
nand U4731 (N_4731,N_4512,N_4513);
xnor U4732 (N_4732,N_4580,N_4573);
nand U4733 (N_4733,N_4537,N_4592);
nand U4734 (N_4734,N_4487,N_4442);
nor U4735 (N_4735,N_4524,N_4578);
or U4736 (N_4736,N_4404,N_4408);
nand U4737 (N_4737,N_4590,N_4498);
or U4738 (N_4738,N_4460,N_4437);
nor U4739 (N_4739,N_4536,N_4514);
nand U4740 (N_4740,N_4424,N_4468);
and U4741 (N_4741,N_4447,N_4557);
nor U4742 (N_4742,N_4591,N_4482);
nor U4743 (N_4743,N_4559,N_4449);
and U4744 (N_4744,N_4574,N_4456);
nor U4745 (N_4745,N_4597,N_4497);
xnor U4746 (N_4746,N_4482,N_4551);
nor U4747 (N_4747,N_4428,N_4547);
nor U4748 (N_4748,N_4582,N_4421);
nand U4749 (N_4749,N_4509,N_4409);
and U4750 (N_4750,N_4502,N_4452);
and U4751 (N_4751,N_4506,N_4590);
nand U4752 (N_4752,N_4514,N_4587);
nand U4753 (N_4753,N_4571,N_4409);
nand U4754 (N_4754,N_4497,N_4577);
or U4755 (N_4755,N_4587,N_4446);
and U4756 (N_4756,N_4578,N_4533);
xnor U4757 (N_4757,N_4596,N_4466);
xnor U4758 (N_4758,N_4588,N_4510);
and U4759 (N_4759,N_4403,N_4483);
xor U4760 (N_4760,N_4496,N_4498);
or U4761 (N_4761,N_4512,N_4547);
nand U4762 (N_4762,N_4488,N_4412);
nand U4763 (N_4763,N_4459,N_4441);
xnor U4764 (N_4764,N_4486,N_4481);
nor U4765 (N_4765,N_4426,N_4502);
nand U4766 (N_4766,N_4537,N_4451);
xnor U4767 (N_4767,N_4472,N_4510);
xor U4768 (N_4768,N_4523,N_4486);
or U4769 (N_4769,N_4421,N_4442);
nor U4770 (N_4770,N_4590,N_4494);
nand U4771 (N_4771,N_4428,N_4457);
nor U4772 (N_4772,N_4420,N_4518);
and U4773 (N_4773,N_4477,N_4474);
nor U4774 (N_4774,N_4433,N_4577);
or U4775 (N_4775,N_4587,N_4584);
or U4776 (N_4776,N_4418,N_4480);
nor U4777 (N_4777,N_4424,N_4559);
nand U4778 (N_4778,N_4555,N_4540);
nand U4779 (N_4779,N_4475,N_4481);
nand U4780 (N_4780,N_4525,N_4425);
or U4781 (N_4781,N_4441,N_4593);
nand U4782 (N_4782,N_4403,N_4515);
and U4783 (N_4783,N_4592,N_4480);
nand U4784 (N_4784,N_4431,N_4503);
xnor U4785 (N_4785,N_4548,N_4479);
xor U4786 (N_4786,N_4550,N_4549);
and U4787 (N_4787,N_4456,N_4587);
xor U4788 (N_4788,N_4431,N_4442);
nand U4789 (N_4789,N_4424,N_4503);
and U4790 (N_4790,N_4530,N_4576);
or U4791 (N_4791,N_4504,N_4447);
nor U4792 (N_4792,N_4559,N_4546);
xnor U4793 (N_4793,N_4551,N_4503);
or U4794 (N_4794,N_4586,N_4550);
xnor U4795 (N_4795,N_4485,N_4583);
and U4796 (N_4796,N_4495,N_4414);
xor U4797 (N_4797,N_4411,N_4462);
or U4798 (N_4798,N_4427,N_4407);
xnor U4799 (N_4799,N_4450,N_4527);
nor U4800 (N_4800,N_4633,N_4614);
xor U4801 (N_4801,N_4716,N_4746);
or U4802 (N_4802,N_4654,N_4753);
xnor U4803 (N_4803,N_4732,N_4605);
xor U4804 (N_4804,N_4659,N_4625);
nand U4805 (N_4805,N_4793,N_4778);
xor U4806 (N_4806,N_4693,N_4734);
and U4807 (N_4807,N_4745,N_4759);
or U4808 (N_4808,N_4738,N_4707);
nor U4809 (N_4809,N_4615,N_4726);
or U4810 (N_4810,N_4660,N_4783);
nand U4811 (N_4811,N_4613,N_4773);
xor U4812 (N_4812,N_4638,N_4607);
or U4813 (N_4813,N_4653,N_4621);
nand U4814 (N_4814,N_4680,N_4733);
or U4815 (N_4815,N_4796,N_4770);
nor U4816 (N_4816,N_4617,N_4658);
nor U4817 (N_4817,N_4708,N_4799);
nor U4818 (N_4818,N_4775,N_4643);
or U4819 (N_4819,N_4720,N_4601);
nor U4820 (N_4820,N_4678,N_4679);
nand U4821 (N_4821,N_4635,N_4692);
xnor U4822 (N_4822,N_4650,N_4785);
or U4823 (N_4823,N_4797,N_4664);
nand U4824 (N_4824,N_4644,N_4705);
nor U4825 (N_4825,N_4767,N_4724);
and U4826 (N_4826,N_4751,N_4616);
or U4827 (N_4827,N_4721,N_4742);
nor U4828 (N_4828,N_4710,N_4730);
nor U4829 (N_4829,N_4694,N_4602);
nand U4830 (N_4830,N_4752,N_4702);
or U4831 (N_4831,N_4631,N_4618);
and U4832 (N_4832,N_4762,N_4784);
and U4833 (N_4833,N_4610,N_4765);
nand U4834 (N_4834,N_4634,N_4626);
or U4835 (N_4835,N_4729,N_4632);
nand U4836 (N_4836,N_4661,N_4737);
and U4837 (N_4837,N_4704,N_4764);
or U4838 (N_4838,N_4624,N_4695);
xnor U4839 (N_4839,N_4779,N_4636);
nor U4840 (N_4840,N_4722,N_4606);
xnor U4841 (N_4841,N_4703,N_4736);
and U4842 (N_4842,N_4788,N_4755);
nor U4843 (N_4843,N_4656,N_4683);
and U4844 (N_4844,N_4671,N_4629);
or U4845 (N_4845,N_4639,N_4665);
or U4846 (N_4846,N_4688,N_4623);
xor U4847 (N_4847,N_4609,N_4646);
or U4848 (N_4848,N_4748,N_4714);
nor U4849 (N_4849,N_4676,N_4677);
xor U4850 (N_4850,N_4630,N_4766);
or U4851 (N_4851,N_4697,N_4603);
and U4852 (N_4852,N_4666,N_4698);
xor U4853 (N_4853,N_4673,N_4608);
nor U4854 (N_4854,N_4675,N_4682);
and U4855 (N_4855,N_4663,N_4685);
nand U4856 (N_4856,N_4648,N_4749);
or U4857 (N_4857,N_4690,N_4647);
nand U4858 (N_4858,N_4781,N_4655);
or U4859 (N_4859,N_4747,N_4754);
xnor U4860 (N_4860,N_4760,N_4798);
or U4861 (N_4861,N_4769,N_4787);
nor U4862 (N_4862,N_4684,N_4645);
or U4863 (N_4863,N_4717,N_4739);
xor U4864 (N_4864,N_4744,N_4670);
and U4865 (N_4865,N_4757,N_4649);
or U4866 (N_4866,N_4622,N_4627);
or U4867 (N_4867,N_4691,N_4709);
or U4868 (N_4868,N_4637,N_4791);
and U4869 (N_4869,N_4604,N_4681);
or U4870 (N_4870,N_4758,N_4761);
nand U4871 (N_4871,N_4689,N_4641);
and U4872 (N_4872,N_4668,N_4768);
nor U4873 (N_4873,N_4686,N_4640);
nor U4874 (N_4874,N_4792,N_4713);
nand U4875 (N_4875,N_4756,N_4750);
nor U4876 (N_4876,N_4612,N_4600);
nor U4877 (N_4877,N_4786,N_4794);
nor U4878 (N_4878,N_4772,N_4672);
nor U4879 (N_4879,N_4725,N_4657);
or U4880 (N_4880,N_4669,N_4628);
nor U4881 (N_4881,N_4667,N_4715);
xnor U4882 (N_4882,N_4771,N_4706);
or U4883 (N_4883,N_4696,N_4662);
or U4884 (N_4884,N_4718,N_4740);
nand U4885 (N_4885,N_4741,N_4700);
and U4886 (N_4886,N_4620,N_4728);
nor U4887 (N_4887,N_4780,N_4712);
or U4888 (N_4888,N_4687,N_4611);
and U4889 (N_4889,N_4723,N_4790);
nor U4890 (N_4890,N_4731,N_4699);
or U4891 (N_4891,N_4795,N_4735);
nor U4892 (N_4892,N_4777,N_4789);
nand U4893 (N_4893,N_4642,N_4674);
nand U4894 (N_4894,N_4619,N_4652);
xnor U4895 (N_4895,N_4782,N_4651);
nor U4896 (N_4896,N_4727,N_4763);
nand U4897 (N_4897,N_4776,N_4701);
or U4898 (N_4898,N_4711,N_4774);
xnor U4899 (N_4899,N_4719,N_4743);
or U4900 (N_4900,N_4684,N_4682);
nand U4901 (N_4901,N_4790,N_4776);
nor U4902 (N_4902,N_4610,N_4783);
xor U4903 (N_4903,N_4647,N_4717);
and U4904 (N_4904,N_4638,N_4780);
xnor U4905 (N_4905,N_4758,N_4661);
xor U4906 (N_4906,N_4768,N_4716);
and U4907 (N_4907,N_4708,N_4772);
or U4908 (N_4908,N_4673,N_4726);
nor U4909 (N_4909,N_4734,N_4706);
xor U4910 (N_4910,N_4654,N_4715);
xnor U4911 (N_4911,N_4698,N_4782);
nor U4912 (N_4912,N_4720,N_4635);
and U4913 (N_4913,N_4635,N_4672);
nor U4914 (N_4914,N_4667,N_4788);
xor U4915 (N_4915,N_4660,N_4633);
nand U4916 (N_4916,N_4736,N_4600);
or U4917 (N_4917,N_4781,N_4720);
nand U4918 (N_4918,N_4784,N_4792);
and U4919 (N_4919,N_4672,N_4707);
xnor U4920 (N_4920,N_4663,N_4634);
nand U4921 (N_4921,N_4664,N_4613);
nand U4922 (N_4922,N_4659,N_4730);
or U4923 (N_4923,N_4718,N_4643);
nand U4924 (N_4924,N_4797,N_4662);
xnor U4925 (N_4925,N_4658,N_4774);
and U4926 (N_4926,N_4763,N_4661);
xnor U4927 (N_4927,N_4721,N_4637);
and U4928 (N_4928,N_4738,N_4767);
xnor U4929 (N_4929,N_4642,N_4661);
nor U4930 (N_4930,N_4627,N_4796);
and U4931 (N_4931,N_4798,N_4732);
and U4932 (N_4932,N_4685,N_4705);
nand U4933 (N_4933,N_4677,N_4617);
xor U4934 (N_4934,N_4626,N_4659);
nor U4935 (N_4935,N_4600,N_4683);
and U4936 (N_4936,N_4793,N_4605);
xnor U4937 (N_4937,N_4608,N_4667);
xor U4938 (N_4938,N_4726,N_4762);
xor U4939 (N_4939,N_4668,N_4705);
or U4940 (N_4940,N_4620,N_4672);
xor U4941 (N_4941,N_4757,N_4797);
or U4942 (N_4942,N_4790,N_4660);
and U4943 (N_4943,N_4744,N_4704);
nand U4944 (N_4944,N_4710,N_4619);
or U4945 (N_4945,N_4648,N_4729);
nand U4946 (N_4946,N_4742,N_4691);
nor U4947 (N_4947,N_4691,N_4673);
nand U4948 (N_4948,N_4706,N_4633);
nand U4949 (N_4949,N_4610,N_4662);
or U4950 (N_4950,N_4650,N_4793);
nor U4951 (N_4951,N_4686,N_4630);
xnor U4952 (N_4952,N_4613,N_4757);
xnor U4953 (N_4953,N_4698,N_4641);
or U4954 (N_4954,N_4791,N_4694);
xor U4955 (N_4955,N_4763,N_4706);
or U4956 (N_4956,N_4795,N_4749);
and U4957 (N_4957,N_4745,N_4656);
or U4958 (N_4958,N_4725,N_4666);
nand U4959 (N_4959,N_4770,N_4637);
nor U4960 (N_4960,N_4666,N_4668);
or U4961 (N_4961,N_4675,N_4756);
or U4962 (N_4962,N_4642,N_4712);
nand U4963 (N_4963,N_4757,N_4667);
or U4964 (N_4964,N_4726,N_4705);
and U4965 (N_4965,N_4731,N_4681);
xnor U4966 (N_4966,N_4728,N_4730);
xnor U4967 (N_4967,N_4715,N_4620);
and U4968 (N_4968,N_4640,N_4741);
and U4969 (N_4969,N_4782,N_4755);
and U4970 (N_4970,N_4748,N_4673);
nand U4971 (N_4971,N_4767,N_4792);
or U4972 (N_4972,N_4721,N_4697);
xor U4973 (N_4973,N_4696,N_4626);
or U4974 (N_4974,N_4708,N_4710);
nand U4975 (N_4975,N_4793,N_4641);
nor U4976 (N_4976,N_4607,N_4673);
or U4977 (N_4977,N_4748,N_4754);
xor U4978 (N_4978,N_4656,N_4719);
nand U4979 (N_4979,N_4727,N_4789);
nand U4980 (N_4980,N_4707,N_4612);
or U4981 (N_4981,N_4724,N_4611);
nand U4982 (N_4982,N_4637,N_4783);
nor U4983 (N_4983,N_4783,N_4695);
or U4984 (N_4984,N_4624,N_4785);
nor U4985 (N_4985,N_4675,N_4731);
and U4986 (N_4986,N_4664,N_4620);
xor U4987 (N_4987,N_4614,N_4757);
or U4988 (N_4988,N_4610,N_4737);
xnor U4989 (N_4989,N_4680,N_4608);
nand U4990 (N_4990,N_4764,N_4602);
xor U4991 (N_4991,N_4735,N_4749);
and U4992 (N_4992,N_4720,N_4650);
xnor U4993 (N_4993,N_4602,N_4670);
nand U4994 (N_4994,N_4773,N_4659);
xor U4995 (N_4995,N_4733,N_4705);
xor U4996 (N_4996,N_4678,N_4662);
nor U4997 (N_4997,N_4732,N_4612);
nor U4998 (N_4998,N_4640,N_4623);
nand U4999 (N_4999,N_4626,N_4766);
nor U5000 (N_5000,N_4838,N_4881);
or U5001 (N_5001,N_4920,N_4817);
or U5002 (N_5002,N_4835,N_4978);
and U5003 (N_5003,N_4968,N_4824);
nand U5004 (N_5004,N_4867,N_4860);
and U5005 (N_5005,N_4868,N_4823);
xnor U5006 (N_5006,N_4861,N_4877);
or U5007 (N_5007,N_4926,N_4895);
and U5008 (N_5008,N_4889,N_4828);
xor U5009 (N_5009,N_4975,N_4939);
and U5010 (N_5010,N_4812,N_4879);
nor U5011 (N_5011,N_4976,N_4891);
or U5012 (N_5012,N_4806,N_4952);
or U5013 (N_5013,N_4992,N_4887);
and U5014 (N_5014,N_4875,N_4837);
and U5015 (N_5015,N_4853,N_4834);
nor U5016 (N_5016,N_4988,N_4847);
or U5017 (N_5017,N_4912,N_4971);
xnor U5018 (N_5018,N_4900,N_4954);
or U5019 (N_5019,N_4878,N_4801);
nand U5020 (N_5020,N_4846,N_4830);
and U5021 (N_5021,N_4808,N_4886);
or U5022 (N_5022,N_4870,N_4928);
nor U5023 (N_5023,N_4977,N_4803);
nand U5024 (N_5024,N_4914,N_4944);
nor U5025 (N_5025,N_4851,N_4854);
nand U5026 (N_5026,N_4951,N_4826);
and U5027 (N_5027,N_4822,N_4913);
xnor U5028 (N_5028,N_4945,N_4898);
xor U5029 (N_5029,N_4862,N_4892);
nand U5030 (N_5030,N_4818,N_4983);
nor U5031 (N_5031,N_4811,N_4940);
or U5032 (N_5032,N_4831,N_4836);
nand U5033 (N_5033,N_4989,N_4972);
nor U5034 (N_5034,N_4963,N_4814);
xor U5035 (N_5035,N_4848,N_4953);
nor U5036 (N_5036,N_4919,N_4894);
or U5037 (N_5037,N_4911,N_4929);
nand U5038 (N_5038,N_4908,N_4902);
xnor U5039 (N_5039,N_4839,N_4950);
or U5040 (N_5040,N_4876,N_4961);
or U5041 (N_5041,N_4857,N_4955);
and U5042 (N_5042,N_4999,N_4987);
or U5043 (N_5043,N_4941,N_4994);
or U5044 (N_5044,N_4804,N_4809);
nand U5045 (N_5045,N_4807,N_4917);
nor U5046 (N_5046,N_4921,N_4903);
nand U5047 (N_5047,N_4872,N_4852);
or U5048 (N_5048,N_4873,N_4905);
nand U5049 (N_5049,N_4985,N_4997);
nand U5050 (N_5050,N_4821,N_4843);
xnor U5051 (N_5051,N_4967,N_4991);
or U5052 (N_5052,N_4958,N_4907);
and U5053 (N_5053,N_4825,N_4864);
nand U5054 (N_5054,N_4943,N_4805);
xnor U5055 (N_5055,N_4841,N_4909);
and U5056 (N_5056,N_4964,N_4930);
xor U5057 (N_5057,N_4934,N_4923);
or U5058 (N_5058,N_4810,N_4910);
or U5059 (N_5059,N_4819,N_4859);
and U5060 (N_5060,N_4842,N_4869);
xnor U5061 (N_5061,N_4959,N_4849);
or U5062 (N_5062,N_4960,N_4936);
and U5063 (N_5063,N_4833,N_4979);
nor U5064 (N_5064,N_4942,N_4965);
and U5065 (N_5065,N_4996,N_4906);
nand U5066 (N_5066,N_4922,N_4924);
and U5067 (N_5067,N_4802,N_4899);
or U5068 (N_5068,N_4884,N_4863);
and U5069 (N_5069,N_4986,N_4829);
xnor U5070 (N_5070,N_4947,N_4915);
nor U5071 (N_5071,N_4970,N_4871);
nor U5072 (N_5072,N_4832,N_4969);
nand U5073 (N_5073,N_4998,N_4827);
nand U5074 (N_5074,N_4933,N_4880);
nor U5075 (N_5075,N_4855,N_4937);
and U5076 (N_5076,N_4845,N_4865);
nand U5077 (N_5077,N_4931,N_4840);
or U5078 (N_5078,N_4890,N_4962);
or U5079 (N_5079,N_4984,N_4813);
xnor U5080 (N_5080,N_4925,N_4966);
and U5081 (N_5081,N_4949,N_4918);
nor U5082 (N_5082,N_4882,N_4874);
nor U5083 (N_5083,N_4885,N_4893);
nor U5084 (N_5084,N_4995,N_4927);
xor U5085 (N_5085,N_4916,N_4866);
and U5086 (N_5086,N_4800,N_4973);
and U5087 (N_5087,N_4888,N_4990);
and U5088 (N_5088,N_4897,N_4938);
and U5089 (N_5089,N_4946,N_4844);
or U5090 (N_5090,N_4901,N_4980);
xnor U5091 (N_5091,N_4858,N_4948);
xnor U5092 (N_5092,N_4856,N_4932);
nand U5093 (N_5093,N_4993,N_4850);
nor U5094 (N_5094,N_4981,N_4816);
and U5095 (N_5095,N_4957,N_4896);
xnor U5096 (N_5096,N_4815,N_4883);
xnor U5097 (N_5097,N_4904,N_4935);
nand U5098 (N_5098,N_4974,N_4820);
or U5099 (N_5099,N_4956,N_4982);
and U5100 (N_5100,N_4974,N_4995);
xor U5101 (N_5101,N_4922,N_4807);
and U5102 (N_5102,N_4998,N_4958);
nand U5103 (N_5103,N_4994,N_4887);
nor U5104 (N_5104,N_4927,N_4839);
nor U5105 (N_5105,N_4872,N_4945);
nor U5106 (N_5106,N_4824,N_4901);
nor U5107 (N_5107,N_4868,N_4830);
or U5108 (N_5108,N_4859,N_4841);
and U5109 (N_5109,N_4877,N_4817);
nor U5110 (N_5110,N_4894,N_4805);
and U5111 (N_5111,N_4860,N_4881);
xor U5112 (N_5112,N_4879,N_4893);
nor U5113 (N_5113,N_4811,N_4896);
and U5114 (N_5114,N_4847,N_4976);
nand U5115 (N_5115,N_4802,N_4806);
and U5116 (N_5116,N_4968,N_4936);
nand U5117 (N_5117,N_4829,N_4980);
or U5118 (N_5118,N_4941,N_4860);
and U5119 (N_5119,N_4900,N_4968);
nor U5120 (N_5120,N_4859,N_4889);
xnor U5121 (N_5121,N_4977,N_4917);
or U5122 (N_5122,N_4831,N_4966);
and U5123 (N_5123,N_4956,N_4889);
xor U5124 (N_5124,N_4853,N_4822);
and U5125 (N_5125,N_4818,N_4846);
nor U5126 (N_5126,N_4902,N_4937);
nor U5127 (N_5127,N_4825,N_4887);
or U5128 (N_5128,N_4839,N_4949);
or U5129 (N_5129,N_4977,N_4826);
nor U5130 (N_5130,N_4975,N_4838);
nand U5131 (N_5131,N_4944,N_4982);
xnor U5132 (N_5132,N_4985,N_4809);
and U5133 (N_5133,N_4811,N_4880);
nor U5134 (N_5134,N_4984,N_4851);
or U5135 (N_5135,N_4810,N_4815);
or U5136 (N_5136,N_4867,N_4943);
and U5137 (N_5137,N_4973,N_4969);
nand U5138 (N_5138,N_4837,N_4874);
nand U5139 (N_5139,N_4818,N_4894);
and U5140 (N_5140,N_4934,N_4930);
nand U5141 (N_5141,N_4875,N_4985);
or U5142 (N_5142,N_4876,N_4837);
nand U5143 (N_5143,N_4969,N_4886);
nand U5144 (N_5144,N_4835,N_4930);
and U5145 (N_5145,N_4847,N_4924);
nor U5146 (N_5146,N_4815,N_4877);
or U5147 (N_5147,N_4906,N_4870);
or U5148 (N_5148,N_4931,N_4997);
xnor U5149 (N_5149,N_4868,N_4869);
and U5150 (N_5150,N_4881,N_4961);
nor U5151 (N_5151,N_4862,N_4986);
xor U5152 (N_5152,N_4856,N_4978);
nand U5153 (N_5153,N_4825,N_4880);
xor U5154 (N_5154,N_4849,N_4878);
or U5155 (N_5155,N_4855,N_4862);
and U5156 (N_5156,N_4997,N_4837);
or U5157 (N_5157,N_4811,N_4991);
nor U5158 (N_5158,N_4916,N_4881);
nand U5159 (N_5159,N_4976,N_4866);
or U5160 (N_5160,N_4858,N_4972);
nand U5161 (N_5161,N_4812,N_4848);
nand U5162 (N_5162,N_4820,N_4811);
and U5163 (N_5163,N_4958,N_4804);
nand U5164 (N_5164,N_4850,N_4870);
or U5165 (N_5165,N_4895,N_4900);
nor U5166 (N_5166,N_4980,N_4864);
or U5167 (N_5167,N_4981,N_4804);
or U5168 (N_5168,N_4943,N_4807);
and U5169 (N_5169,N_4934,N_4843);
and U5170 (N_5170,N_4854,N_4990);
and U5171 (N_5171,N_4872,N_4811);
and U5172 (N_5172,N_4894,N_4821);
and U5173 (N_5173,N_4821,N_4816);
xnor U5174 (N_5174,N_4986,N_4989);
xor U5175 (N_5175,N_4933,N_4908);
nand U5176 (N_5176,N_4857,N_4968);
nor U5177 (N_5177,N_4972,N_4987);
nand U5178 (N_5178,N_4969,N_4927);
nor U5179 (N_5179,N_4923,N_4904);
or U5180 (N_5180,N_4915,N_4849);
xnor U5181 (N_5181,N_4981,N_4882);
nor U5182 (N_5182,N_4847,N_4800);
nand U5183 (N_5183,N_4853,N_4964);
xor U5184 (N_5184,N_4923,N_4819);
or U5185 (N_5185,N_4881,N_4849);
or U5186 (N_5186,N_4833,N_4847);
xor U5187 (N_5187,N_4970,N_4969);
nand U5188 (N_5188,N_4913,N_4942);
and U5189 (N_5189,N_4899,N_4883);
or U5190 (N_5190,N_4911,N_4976);
or U5191 (N_5191,N_4936,N_4846);
xnor U5192 (N_5192,N_4967,N_4892);
or U5193 (N_5193,N_4924,N_4929);
or U5194 (N_5194,N_4903,N_4885);
and U5195 (N_5195,N_4975,N_4969);
xnor U5196 (N_5196,N_4906,N_4995);
or U5197 (N_5197,N_4875,N_4869);
nor U5198 (N_5198,N_4907,N_4818);
xor U5199 (N_5199,N_4831,N_4960);
and U5200 (N_5200,N_5044,N_5100);
nor U5201 (N_5201,N_5039,N_5027);
and U5202 (N_5202,N_5122,N_5180);
nor U5203 (N_5203,N_5120,N_5189);
nor U5204 (N_5204,N_5053,N_5115);
nand U5205 (N_5205,N_5159,N_5192);
nor U5206 (N_5206,N_5194,N_5010);
nand U5207 (N_5207,N_5028,N_5199);
or U5208 (N_5208,N_5009,N_5019);
nand U5209 (N_5209,N_5050,N_5105);
or U5210 (N_5210,N_5131,N_5032);
nand U5211 (N_5211,N_5158,N_5081);
nor U5212 (N_5212,N_5114,N_5049);
and U5213 (N_5213,N_5193,N_5179);
or U5214 (N_5214,N_5030,N_5047);
or U5215 (N_5215,N_5188,N_5056);
nand U5216 (N_5216,N_5134,N_5067);
xnor U5217 (N_5217,N_5026,N_5147);
xnor U5218 (N_5218,N_5137,N_5143);
or U5219 (N_5219,N_5078,N_5161);
and U5220 (N_5220,N_5090,N_5155);
nand U5221 (N_5221,N_5116,N_5111);
nor U5222 (N_5222,N_5172,N_5107);
nor U5223 (N_5223,N_5042,N_5068);
and U5224 (N_5224,N_5185,N_5073);
or U5225 (N_5225,N_5033,N_5003);
xnor U5226 (N_5226,N_5059,N_5173);
nor U5227 (N_5227,N_5025,N_5153);
and U5228 (N_5228,N_5141,N_5076);
and U5229 (N_5229,N_5181,N_5094);
and U5230 (N_5230,N_5096,N_5095);
nor U5231 (N_5231,N_5080,N_5011);
xor U5232 (N_5232,N_5041,N_5029);
xor U5233 (N_5233,N_5110,N_5052);
or U5234 (N_5234,N_5163,N_5121);
nand U5235 (N_5235,N_5182,N_5077);
nand U5236 (N_5236,N_5083,N_5196);
nor U5237 (N_5237,N_5140,N_5171);
or U5238 (N_5238,N_5043,N_5070);
nor U5239 (N_5239,N_5075,N_5015);
nor U5240 (N_5240,N_5035,N_5087);
nand U5241 (N_5241,N_5005,N_5055);
xor U5242 (N_5242,N_5031,N_5136);
xor U5243 (N_5243,N_5169,N_5187);
nand U5244 (N_5244,N_5013,N_5063);
nand U5245 (N_5245,N_5012,N_5069);
nor U5246 (N_5246,N_5119,N_5129);
nand U5247 (N_5247,N_5125,N_5130);
xor U5248 (N_5248,N_5008,N_5071);
or U5249 (N_5249,N_5108,N_5149);
xnor U5250 (N_5250,N_5123,N_5023);
or U5251 (N_5251,N_5138,N_5170);
or U5252 (N_5252,N_5091,N_5154);
and U5253 (N_5253,N_5162,N_5097);
nand U5254 (N_5254,N_5061,N_5133);
nand U5255 (N_5255,N_5024,N_5151);
nand U5256 (N_5256,N_5093,N_5102);
nor U5257 (N_5257,N_5058,N_5152);
nand U5258 (N_5258,N_5062,N_5127);
or U5259 (N_5259,N_5190,N_5020);
nand U5260 (N_5260,N_5002,N_5101);
or U5261 (N_5261,N_5168,N_5166);
nor U5262 (N_5262,N_5040,N_5139);
nor U5263 (N_5263,N_5186,N_5098);
xor U5264 (N_5264,N_5000,N_5178);
xnor U5265 (N_5265,N_5106,N_5165);
or U5266 (N_5266,N_5017,N_5084);
xnor U5267 (N_5267,N_5197,N_5146);
xor U5268 (N_5268,N_5088,N_5034);
xor U5269 (N_5269,N_5086,N_5195);
nand U5270 (N_5270,N_5144,N_5022);
nand U5271 (N_5271,N_5191,N_5079);
xor U5272 (N_5272,N_5184,N_5082);
and U5273 (N_5273,N_5054,N_5176);
nor U5274 (N_5274,N_5085,N_5135);
xnor U5275 (N_5275,N_5174,N_5177);
and U5276 (N_5276,N_5057,N_5113);
and U5277 (N_5277,N_5126,N_5109);
or U5278 (N_5278,N_5048,N_5064);
nand U5279 (N_5279,N_5037,N_5001);
or U5280 (N_5280,N_5036,N_5018);
nand U5281 (N_5281,N_5118,N_5038);
xor U5282 (N_5282,N_5099,N_5112);
xor U5283 (N_5283,N_5092,N_5066);
and U5284 (N_5284,N_5006,N_5060);
xor U5285 (N_5285,N_5065,N_5142);
and U5286 (N_5286,N_5124,N_5132);
nor U5287 (N_5287,N_5145,N_5160);
or U5288 (N_5288,N_5148,N_5089);
nor U5289 (N_5289,N_5167,N_5007);
nor U5290 (N_5290,N_5150,N_5117);
and U5291 (N_5291,N_5004,N_5164);
nor U5292 (N_5292,N_5198,N_5051);
nor U5293 (N_5293,N_5103,N_5183);
and U5294 (N_5294,N_5014,N_5016);
and U5295 (N_5295,N_5074,N_5128);
or U5296 (N_5296,N_5175,N_5046);
xor U5297 (N_5297,N_5072,N_5104);
nor U5298 (N_5298,N_5156,N_5157);
or U5299 (N_5299,N_5021,N_5045);
xor U5300 (N_5300,N_5025,N_5071);
xor U5301 (N_5301,N_5144,N_5055);
nor U5302 (N_5302,N_5019,N_5093);
or U5303 (N_5303,N_5047,N_5120);
or U5304 (N_5304,N_5114,N_5178);
and U5305 (N_5305,N_5003,N_5160);
xnor U5306 (N_5306,N_5070,N_5161);
and U5307 (N_5307,N_5143,N_5023);
or U5308 (N_5308,N_5081,N_5001);
and U5309 (N_5309,N_5139,N_5059);
and U5310 (N_5310,N_5019,N_5195);
or U5311 (N_5311,N_5007,N_5071);
or U5312 (N_5312,N_5106,N_5088);
nand U5313 (N_5313,N_5077,N_5107);
nand U5314 (N_5314,N_5044,N_5170);
nand U5315 (N_5315,N_5018,N_5126);
and U5316 (N_5316,N_5165,N_5148);
nand U5317 (N_5317,N_5044,N_5194);
nor U5318 (N_5318,N_5097,N_5034);
nand U5319 (N_5319,N_5097,N_5025);
or U5320 (N_5320,N_5001,N_5166);
nand U5321 (N_5321,N_5156,N_5048);
and U5322 (N_5322,N_5096,N_5144);
nor U5323 (N_5323,N_5069,N_5083);
or U5324 (N_5324,N_5109,N_5024);
nand U5325 (N_5325,N_5035,N_5186);
nor U5326 (N_5326,N_5184,N_5013);
nand U5327 (N_5327,N_5103,N_5009);
and U5328 (N_5328,N_5080,N_5063);
and U5329 (N_5329,N_5075,N_5161);
nor U5330 (N_5330,N_5005,N_5004);
and U5331 (N_5331,N_5195,N_5133);
xor U5332 (N_5332,N_5182,N_5147);
or U5333 (N_5333,N_5194,N_5086);
nand U5334 (N_5334,N_5008,N_5186);
nor U5335 (N_5335,N_5182,N_5158);
or U5336 (N_5336,N_5173,N_5044);
xor U5337 (N_5337,N_5036,N_5011);
and U5338 (N_5338,N_5008,N_5117);
nand U5339 (N_5339,N_5047,N_5080);
xnor U5340 (N_5340,N_5111,N_5109);
xnor U5341 (N_5341,N_5115,N_5047);
and U5342 (N_5342,N_5048,N_5061);
nand U5343 (N_5343,N_5120,N_5077);
or U5344 (N_5344,N_5035,N_5154);
nand U5345 (N_5345,N_5042,N_5169);
nand U5346 (N_5346,N_5193,N_5019);
xor U5347 (N_5347,N_5185,N_5059);
nor U5348 (N_5348,N_5031,N_5075);
nor U5349 (N_5349,N_5167,N_5097);
nand U5350 (N_5350,N_5099,N_5030);
nand U5351 (N_5351,N_5078,N_5111);
and U5352 (N_5352,N_5078,N_5016);
or U5353 (N_5353,N_5099,N_5013);
and U5354 (N_5354,N_5057,N_5123);
nand U5355 (N_5355,N_5085,N_5157);
xor U5356 (N_5356,N_5197,N_5145);
and U5357 (N_5357,N_5000,N_5128);
xnor U5358 (N_5358,N_5131,N_5162);
and U5359 (N_5359,N_5199,N_5177);
nand U5360 (N_5360,N_5103,N_5028);
xor U5361 (N_5361,N_5125,N_5199);
nor U5362 (N_5362,N_5169,N_5125);
xnor U5363 (N_5363,N_5158,N_5159);
and U5364 (N_5364,N_5041,N_5036);
xnor U5365 (N_5365,N_5003,N_5026);
xnor U5366 (N_5366,N_5004,N_5183);
nand U5367 (N_5367,N_5195,N_5168);
or U5368 (N_5368,N_5106,N_5195);
xor U5369 (N_5369,N_5107,N_5033);
xor U5370 (N_5370,N_5010,N_5119);
nor U5371 (N_5371,N_5105,N_5048);
or U5372 (N_5372,N_5185,N_5117);
xnor U5373 (N_5373,N_5183,N_5056);
or U5374 (N_5374,N_5042,N_5109);
or U5375 (N_5375,N_5029,N_5141);
or U5376 (N_5376,N_5164,N_5162);
xnor U5377 (N_5377,N_5181,N_5175);
or U5378 (N_5378,N_5152,N_5045);
or U5379 (N_5379,N_5100,N_5139);
nand U5380 (N_5380,N_5022,N_5173);
nor U5381 (N_5381,N_5077,N_5006);
xnor U5382 (N_5382,N_5057,N_5072);
nor U5383 (N_5383,N_5015,N_5162);
or U5384 (N_5384,N_5182,N_5083);
xnor U5385 (N_5385,N_5061,N_5155);
xnor U5386 (N_5386,N_5199,N_5051);
nor U5387 (N_5387,N_5170,N_5107);
xnor U5388 (N_5388,N_5093,N_5027);
nand U5389 (N_5389,N_5060,N_5103);
and U5390 (N_5390,N_5041,N_5120);
or U5391 (N_5391,N_5004,N_5000);
and U5392 (N_5392,N_5188,N_5077);
and U5393 (N_5393,N_5070,N_5084);
or U5394 (N_5394,N_5058,N_5176);
nand U5395 (N_5395,N_5194,N_5063);
or U5396 (N_5396,N_5015,N_5146);
or U5397 (N_5397,N_5136,N_5121);
and U5398 (N_5398,N_5013,N_5011);
xnor U5399 (N_5399,N_5121,N_5097);
nand U5400 (N_5400,N_5339,N_5268);
nor U5401 (N_5401,N_5343,N_5272);
or U5402 (N_5402,N_5259,N_5369);
nand U5403 (N_5403,N_5261,N_5356);
or U5404 (N_5404,N_5214,N_5216);
nor U5405 (N_5405,N_5303,N_5364);
or U5406 (N_5406,N_5212,N_5204);
nand U5407 (N_5407,N_5319,N_5320);
nand U5408 (N_5408,N_5340,N_5317);
or U5409 (N_5409,N_5238,N_5371);
or U5410 (N_5410,N_5227,N_5224);
nor U5411 (N_5411,N_5336,N_5219);
nand U5412 (N_5412,N_5300,N_5264);
nand U5413 (N_5413,N_5274,N_5389);
xnor U5414 (N_5414,N_5255,N_5302);
xnor U5415 (N_5415,N_5290,N_5211);
or U5416 (N_5416,N_5246,N_5304);
nor U5417 (N_5417,N_5284,N_5381);
or U5418 (N_5418,N_5269,N_5237);
or U5419 (N_5419,N_5293,N_5361);
nand U5420 (N_5420,N_5251,N_5326);
xor U5421 (N_5421,N_5283,N_5398);
or U5422 (N_5422,N_5257,N_5208);
nand U5423 (N_5423,N_5366,N_5223);
or U5424 (N_5424,N_5393,N_5390);
or U5425 (N_5425,N_5341,N_5279);
nand U5426 (N_5426,N_5351,N_5202);
nand U5427 (N_5427,N_5323,N_5342);
nand U5428 (N_5428,N_5328,N_5265);
nand U5429 (N_5429,N_5225,N_5276);
and U5430 (N_5430,N_5229,N_5350);
and U5431 (N_5431,N_5275,N_5388);
or U5432 (N_5432,N_5365,N_5354);
nor U5433 (N_5433,N_5391,N_5262);
nor U5434 (N_5434,N_5314,N_5235);
or U5435 (N_5435,N_5230,N_5299);
and U5436 (N_5436,N_5392,N_5252);
and U5437 (N_5437,N_5385,N_5220);
nand U5438 (N_5438,N_5209,N_5287);
nor U5439 (N_5439,N_5332,N_5282);
or U5440 (N_5440,N_5294,N_5316);
nand U5441 (N_5441,N_5205,N_5232);
or U5442 (N_5442,N_5241,N_5368);
or U5443 (N_5443,N_5245,N_5318);
nand U5444 (N_5444,N_5396,N_5286);
nand U5445 (N_5445,N_5349,N_5333);
nand U5446 (N_5446,N_5337,N_5308);
and U5447 (N_5447,N_5244,N_5200);
and U5448 (N_5448,N_5222,N_5213);
nor U5449 (N_5449,N_5310,N_5344);
nand U5450 (N_5450,N_5360,N_5267);
nand U5451 (N_5451,N_5215,N_5277);
and U5452 (N_5452,N_5228,N_5285);
nor U5453 (N_5453,N_5297,N_5373);
xor U5454 (N_5454,N_5383,N_5253);
and U5455 (N_5455,N_5309,N_5325);
xnor U5456 (N_5456,N_5270,N_5289);
xor U5457 (N_5457,N_5295,N_5345);
nor U5458 (N_5458,N_5353,N_5311);
nand U5459 (N_5459,N_5370,N_5248);
xnor U5460 (N_5460,N_5394,N_5315);
or U5461 (N_5461,N_5348,N_5327);
nor U5462 (N_5462,N_5242,N_5352);
nand U5463 (N_5463,N_5281,N_5288);
or U5464 (N_5464,N_5263,N_5203);
nor U5465 (N_5465,N_5355,N_5347);
nand U5466 (N_5466,N_5386,N_5379);
nand U5467 (N_5467,N_5243,N_5231);
nor U5468 (N_5468,N_5397,N_5305);
nand U5469 (N_5469,N_5322,N_5359);
nand U5470 (N_5470,N_5292,N_5372);
nand U5471 (N_5471,N_5306,N_5210);
nand U5472 (N_5472,N_5221,N_5218);
nor U5473 (N_5473,N_5378,N_5250);
or U5474 (N_5474,N_5217,N_5387);
or U5475 (N_5475,N_5234,N_5399);
nand U5476 (N_5476,N_5273,N_5247);
or U5477 (N_5477,N_5307,N_5256);
xor U5478 (N_5478,N_5278,N_5240);
or U5479 (N_5479,N_5249,N_5367);
xor U5480 (N_5480,N_5382,N_5254);
or U5481 (N_5481,N_5335,N_5312);
nand U5482 (N_5482,N_5280,N_5329);
and U5483 (N_5483,N_5206,N_5207);
or U5484 (N_5484,N_5260,N_5239);
and U5485 (N_5485,N_5236,N_5346);
or U5486 (N_5486,N_5376,N_5331);
nor U5487 (N_5487,N_5301,N_5201);
xnor U5488 (N_5488,N_5338,N_5258);
nor U5489 (N_5489,N_5271,N_5266);
xor U5490 (N_5490,N_5377,N_5298);
nand U5491 (N_5491,N_5291,N_5384);
or U5492 (N_5492,N_5330,N_5313);
and U5493 (N_5493,N_5358,N_5296);
nor U5494 (N_5494,N_5395,N_5233);
or U5495 (N_5495,N_5334,N_5357);
nand U5496 (N_5496,N_5226,N_5321);
nor U5497 (N_5497,N_5374,N_5362);
nand U5498 (N_5498,N_5380,N_5324);
and U5499 (N_5499,N_5363,N_5375);
nor U5500 (N_5500,N_5243,N_5336);
nand U5501 (N_5501,N_5370,N_5363);
nor U5502 (N_5502,N_5390,N_5330);
nor U5503 (N_5503,N_5221,N_5208);
xor U5504 (N_5504,N_5381,N_5346);
nand U5505 (N_5505,N_5320,N_5251);
nand U5506 (N_5506,N_5324,N_5306);
and U5507 (N_5507,N_5255,N_5315);
nand U5508 (N_5508,N_5297,N_5395);
or U5509 (N_5509,N_5288,N_5348);
or U5510 (N_5510,N_5201,N_5286);
xor U5511 (N_5511,N_5259,N_5247);
or U5512 (N_5512,N_5243,N_5330);
nand U5513 (N_5513,N_5380,N_5256);
nand U5514 (N_5514,N_5306,N_5270);
or U5515 (N_5515,N_5239,N_5202);
nor U5516 (N_5516,N_5230,N_5271);
nor U5517 (N_5517,N_5232,N_5246);
or U5518 (N_5518,N_5218,N_5309);
xor U5519 (N_5519,N_5351,N_5332);
xnor U5520 (N_5520,N_5310,N_5257);
nand U5521 (N_5521,N_5346,N_5215);
nor U5522 (N_5522,N_5206,N_5211);
xnor U5523 (N_5523,N_5383,N_5301);
nand U5524 (N_5524,N_5244,N_5315);
and U5525 (N_5525,N_5385,N_5215);
and U5526 (N_5526,N_5380,N_5296);
nor U5527 (N_5527,N_5377,N_5399);
nor U5528 (N_5528,N_5301,N_5381);
or U5529 (N_5529,N_5263,N_5305);
nand U5530 (N_5530,N_5278,N_5234);
and U5531 (N_5531,N_5292,N_5360);
and U5532 (N_5532,N_5301,N_5203);
nand U5533 (N_5533,N_5230,N_5247);
nor U5534 (N_5534,N_5243,N_5257);
nor U5535 (N_5535,N_5356,N_5236);
xnor U5536 (N_5536,N_5268,N_5373);
and U5537 (N_5537,N_5238,N_5226);
nand U5538 (N_5538,N_5387,N_5215);
xor U5539 (N_5539,N_5327,N_5346);
nor U5540 (N_5540,N_5352,N_5356);
nand U5541 (N_5541,N_5361,N_5399);
nor U5542 (N_5542,N_5307,N_5328);
nand U5543 (N_5543,N_5264,N_5331);
or U5544 (N_5544,N_5239,N_5379);
xnor U5545 (N_5545,N_5278,N_5298);
or U5546 (N_5546,N_5369,N_5362);
or U5547 (N_5547,N_5203,N_5255);
nor U5548 (N_5548,N_5267,N_5220);
nand U5549 (N_5549,N_5358,N_5254);
xnor U5550 (N_5550,N_5384,N_5310);
xor U5551 (N_5551,N_5263,N_5298);
nor U5552 (N_5552,N_5203,N_5307);
nor U5553 (N_5553,N_5220,N_5229);
nand U5554 (N_5554,N_5387,N_5207);
or U5555 (N_5555,N_5361,N_5319);
or U5556 (N_5556,N_5341,N_5296);
nor U5557 (N_5557,N_5357,N_5244);
and U5558 (N_5558,N_5248,N_5237);
xor U5559 (N_5559,N_5352,N_5234);
xnor U5560 (N_5560,N_5395,N_5314);
xor U5561 (N_5561,N_5253,N_5237);
nor U5562 (N_5562,N_5378,N_5356);
or U5563 (N_5563,N_5244,N_5222);
and U5564 (N_5564,N_5275,N_5211);
xnor U5565 (N_5565,N_5270,N_5286);
nor U5566 (N_5566,N_5207,N_5374);
nor U5567 (N_5567,N_5391,N_5377);
or U5568 (N_5568,N_5395,N_5289);
or U5569 (N_5569,N_5366,N_5232);
xor U5570 (N_5570,N_5339,N_5367);
and U5571 (N_5571,N_5217,N_5355);
or U5572 (N_5572,N_5320,N_5285);
xor U5573 (N_5573,N_5319,N_5303);
and U5574 (N_5574,N_5222,N_5323);
or U5575 (N_5575,N_5216,N_5362);
nor U5576 (N_5576,N_5242,N_5208);
and U5577 (N_5577,N_5273,N_5307);
or U5578 (N_5578,N_5261,N_5322);
nor U5579 (N_5579,N_5221,N_5255);
and U5580 (N_5580,N_5258,N_5379);
nor U5581 (N_5581,N_5306,N_5397);
xor U5582 (N_5582,N_5365,N_5355);
and U5583 (N_5583,N_5266,N_5322);
nand U5584 (N_5584,N_5229,N_5275);
or U5585 (N_5585,N_5394,N_5335);
nor U5586 (N_5586,N_5240,N_5359);
xnor U5587 (N_5587,N_5224,N_5259);
nand U5588 (N_5588,N_5282,N_5347);
xnor U5589 (N_5589,N_5318,N_5339);
nor U5590 (N_5590,N_5346,N_5252);
nand U5591 (N_5591,N_5285,N_5367);
and U5592 (N_5592,N_5207,N_5345);
xnor U5593 (N_5593,N_5278,N_5232);
xor U5594 (N_5594,N_5331,N_5260);
nor U5595 (N_5595,N_5286,N_5299);
nand U5596 (N_5596,N_5251,N_5392);
or U5597 (N_5597,N_5303,N_5291);
nand U5598 (N_5598,N_5378,N_5252);
or U5599 (N_5599,N_5240,N_5303);
and U5600 (N_5600,N_5460,N_5536);
and U5601 (N_5601,N_5516,N_5472);
xor U5602 (N_5602,N_5466,N_5586);
nand U5603 (N_5603,N_5535,N_5430);
nor U5604 (N_5604,N_5432,N_5450);
nor U5605 (N_5605,N_5415,N_5493);
nor U5606 (N_5606,N_5537,N_5421);
xnor U5607 (N_5607,N_5514,N_5426);
xnor U5608 (N_5608,N_5562,N_5511);
xor U5609 (N_5609,N_5584,N_5425);
or U5610 (N_5610,N_5594,N_5525);
nor U5611 (N_5611,N_5476,N_5576);
or U5612 (N_5612,N_5458,N_5560);
xor U5613 (N_5613,N_5454,N_5500);
xor U5614 (N_5614,N_5418,N_5527);
nor U5615 (N_5615,N_5484,N_5411);
and U5616 (N_5616,N_5554,N_5461);
nand U5617 (N_5617,N_5565,N_5544);
nand U5618 (N_5618,N_5555,N_5423);
and U5619 (N_5619,N_5459,N_5498);
nor U5620 (N_5620,N_5464,N_5417);
or U5621 (N_5621,N_5446,N_5532);
and U5622 (N_5622,N_5489,N_5409);
or U5623 (N_5623,N_5440,N_5503);
nor U5624 (N_5624,N_5482,N_5568);
nor U5625 (N_5625,N_5595,N_5588);
nor U5626 (N_5626,N_5462,N_5475);
and U5627 (N_5627,N_5422,N_5452);
nand U5628 (N_5628,N_5424,N_5572);
xor U5629 (N_5629,N_5442,N_5505);
nand U5630 (N_5630,N_5542,N_5553);
xnor U5631 (N_5631,N_5551,N_5436);
and U5632 (N_5632,N_5429,N_5491);
or U5633 (N_5633,N_5581,N_5407);
nand U5634 (N_5634,N_5403,N_5577);
nor U5635 (N_5635,N_5502,N_5433);
and U5636 (N_5636,N_5457,N_5413);
nor U5637 (N_5637,N_5412,N_5561);
nor U5638 (N_5638,N_5469,N_5569);
or U5639 (N_5639,N_5596,N_5434);
xor U5640 (N_5640,N_5486,N_5510);
xnor U5641 (N_5641,N_5477,N_5556);
nand U5642 (N_5642,N_5558,N_5419);
and U5643 (N_5643,N_5515,N_5573);
or U5644 (N_5644,N_5571,N_5465);
or U5645 (N_5645,N_5523,N_5517);
nand U5646 (N_5646,N_5490,N_5580);
xor U5647 (N_5647,N_5453,N_5599);
xor U5648 (N_5648,N_5550,N_5541);
xnor U5649 (N_5649,N_5589,N_5445);
xor U5650 (N_5650,N_5471,N_5570);
and U5651 (N_5651,N_5455,N_5534);
nand U5652 (N_5652,N_5410,N_5521);
or U5653 (N_5653,N_5512,N_5531);
nand U5654 (N_5654,N_5435,N_5431);
or U5655 (N_5655,N_5406,N_5408);
xnor U5656 (N_5656,N_5400,N_5590);
xor U5657 (N_5657,N_5528,N_5439);
nor U5658 (N_5658,N_5587,N_5483);
or U5659 (N_5659,N_5591,N_5448);
and U5660 (N_5660,N_5543,N_5427);
or U5661 (N_5661,N_5566,N_5506);
or U5662 (N_5662,N_5478,N_5499);
nor U5663 (N_5663,N_5420,N_5564);
and U5664 (N_5664,N_5593,N_5507);
nand U5665 (N_5665,N_5548,N_5414);
nand U5666 (N_5666,N_5592,N_5547);
nand U5667 (N_5667,N_5492,N_5470);
nor U5668 (N_5668,N_5585,N_5546);
or U5669 (N_5669,N_5451,N_5416);
nand U5670 (N_5670,N_5487,N_5404);
nand U5671 (N_5671,N_5513,N_5549);
nand U5672 (N_5672,N_5467,N_5578);
nand U5673 (N_5673,N_5441,N_5444);
xnor U5674 (N_5674,N_5438,N_5559);
nand U5675 (N_5675,N_5437,N_5563);
or U5676 (N_5676,N_5540,N_5496);
nor U5677 (N_5677,N_5567,N_5402);
and U5678 (N_5678,N_5447,N_5463);
nor U5679 (N_5679,N_5597,N_5474);
or U5680 (N_5680,N_5529,N_5443);
or U5681 (N_5681,N_5526,N_5480);
or U5682 (N_5682,N_5508,N_5519);
or U5683 (N_5683,N_5473,N_5504);
xnor U5684 (N_5684,N_5545,N_5524);
xnor U5685 (N_5685,N_5468,N_5582);
xnor U5686 (N_5686,N_5509,N_5501);
and U5687 (N_5687,N_5479,N_5494);
or U5688 (N_5688,N_5405,N_5522);
and U5689 (N_5689,N_5495,N_5574);
xor U5690 (N_5690,N_5579,N_5539);
nand U5691 (N_5691,N_5485,N_5557);
nor U5692 (N_5692,N_5488,N_5520);
xor U5693 (N_5693,N_5583,N_5575);
and U5694 (N_5694,N_5533,N_5598);
or U5695 (N_5695,N_5497,N_5449);
xnor U5696 (N_5696,N_5530,N_5538);
and U5697 (N_5697,N_5428,N_5401);
nand U5698 (N_5698,N_5456,N_5518);
nor U5699 (N_5699,N_5552,N_5481);
nor U5700 (N_5700,N_5577,N_5492);
nor U5701 (N_5701,N_5474,N_5462);
or U5702 (N_5702,N_5518,N_5438);
nand U5703 (N_5703,N_5570,N_5547);
nand U5704 (N_5704,N_5489,N_5463);
or U5705 (N_5705,N_5557,N_5490);
and U5706 (N_5706,N_5570,N_5486);
and U5707 (N_5707,N_5426,N_5573);
or U5708 (N_5708,N_5556,N_5574);
and U5709 (N_5709,N_5428,N_5555);
nand U5710 (N_5710,N_5485,N_5507);
and U5711 (N_5711,N_5486,N_5515);
nor U5712 (N_5712,N_5439,N_5539);
xor U5713 (N_5713,N_5470,N_5515);
or U5714 (N_5714,N_5518,N_5527);
xor U5715 (N_5715,N_5507,N_5598);
nand U5716 (N_5716,N_5468,N_5414);
nor U5717 (N_5717,N_5590,N_5498);
and U5718 (N_5718,N_5458,N_5595);
nand U5719 (N_5719,N_5537,N_5464);
xnor U5720 (N_5720,N_5458,N_5490);
nand U5721 (N_5721,N_5487,N_5540);
or U5722 (N_5722,N_5438,N_5474);
and U5723 (N_5723,N_5528,N_5589);
nor U5724 (N_5724,N_5414,N_5489);
nand U5725 (N_5725,N_5578,N_5468);
nand U5726 (N_5726,N_5564,N_5540);
xnor U5727 (N_5727,N_5543,N_5544);
nor U5728 (N_5728,N_5562,N_5477);
nand U5729 (N_5729,N_5414,N_5527);
xnor U5730 (N_5730,N_5567,N_5564);
xor U5731 (N_5731,N_5485,N_5414);
nand U5732 (N_5732,N_5432,N_5428);
and U5733 (N_5733,N_5508,N_5590);
xor U5734 (N_5734,N_5481,N_5585);
and U5735 (N_5735,N_5514,N_5458);
nor U5736 (N_5736,N_5535,N_5512);
nand U5737 (N_5737,N_5516,N_5481);
and U5738 (N_5738,N_5541,N_5540);
nand U5739 (N_5739,N_5401,N_5521);
and U5740 (N_5740,N_5552,N_5490);
xor U5741 (N_5741,N_5484,N_5434);
nand U5742 (N_5742,N_5420,N_5451);
xor U5743 (N_5743,N_5556,N_5442);
and U5744 (N_5744,N_5444,N_5516);
nand U5745 (N_5745,N_5568,N_5570);
and U5746 (N_5746,N_5400,N_5544);
nor U5747 (N_5747,N_5412,N_5544);
and U5748 (N_5748,N_5430,N_5556);
nor U5749 (N_5749,N_5571,N_5419);
or U5750 (N_5750,N_5454,N_5570);
nand U5751 (N_5751,N_5537,N_5513);
or U5752 (N_5752,N_5513,N_5521);
nor U5753 (N_5753,N_5449,N_5544);
nand U5754 (N_5754,N_5561,N_5566);
xor U5755 (N_5755,N_5475,N_5502);
nand U5756 (N_5756,N_5505,N_5437);
nand U5757 (N_5757,N_5535,N_5565);
xor U5758 (N_5758,N_5422,N_5590);
and U5759 (N_5759,N_5439,N_5571);
nand U5760 (N_5760,N_5574,N_5541);
xnor U5761 (N_5761,N_5514,N_5478);
xor U5762 (N_5762,N_5566,N_5462);
xor U5763 (N_5763,N_5573,N_5469);
xor U5764 (N_5764,N_5584,N_5580);
and U5765 (N_5765,N_5539,N_5574);
nor U5766 (N_5766,N_5470,N_5504);
nand U5767 (N_5767,N_5497,N_5549);
and U5768 (N_5768,N_5401,N_5455);
nand U5769 (N_5769,N_5400,N_5459);
nor U5770 (N_5770,N_5448,N_5412);
nand U5771 (N_5771,N_5508,N_5460);
and U5772 (N_5772,N_5566,N_5403);
or U5773 (N_5773,N_5568,N_5491);
nand U5774 (N_5774,N_5436,N_5408);
nand U5775 (N_5775,N_5555,N_5479);
and U5776 (N_5776,N_5516,N_5428);
and U5777 (N_5777,N_5401,N_5579);
and U5778 (N_5778,N_5488,N_5489);
xor U5779 (N_5779,N_5566,N_5516);
xnor U5780 (N_5780,N_5573,N_5531);
and U5781 (N_5781,N_5557,N_5507);
xor U5782 (N_5782,N_5530,N_5406);
nand U5783 (N_5783,N_5467,N_5532);
xor U5784 (N_5784,N_5517,N_5456);
or U5785 (N_5785,N_5599,N_5414);
xor U5786 (N_5786,N_5588,N_5584);
or U5787 (N_5787,N_5518,N_5504);
nor U5788 (N_5788,N_5405,N_5465);
and U5789 (N_5789,N_5432,N_5527);
xnor U5790 (N_5790,N_5457,N_5498);
nand U5791 (N_5791,N_5572,N_5533);
nand U5792 (N_5792,N_5401,N_5484);
xor U5793 (N_5793,N_5403,N_5513);
and U5794 (N_5794,N_5548,N_5424);
nor U5795 (N_5795,N_5504,N_5567);
nor U5796 (N_5796,N_5568,N_5412);
or U5797 (N_5797,N_5563,N_5410);
or U5798 (N_5798,N_5473,N_5481);
nor U5799 (N_5799,N_5544,N_5414);
nor U5800 (N_5800,N_5611,N_5715);
nand U5801 (N_5801,N_5739,N_5764);
nor U5802 (N_5802,N_5698,N_5670);
nand U5803 (N_5803,N_5638,N_5693);
nor U5804 (N_5804,N_5709,N_5782);
and U5805 (N_5805,N_5619,N_5726);
and U5806 (N_5806,N_5788,N_5633);
nor U5807 (N_5807,N_5663,N_5692);
nand U5808 (N_5808,N_5718,N_5742);
and U5809 (N_5809,N_5789,N_5736);
nor U5810 (N_5810,N_5706,N_5768);
nor U5811 (N_5811,N_5795,N_5681);
and U5812 (N_5812,N_5760,N_5617);
or U5813 (N_5813,N_5632,N_5705);
nor U5814 (N_5814,N_5635,N_5701);
nor U5815 (N_5815,N_5762,N_5787);
nand U5816 (N_5816,N_5687,N_5647);
or U5817 (N_5817,N_5684,N_5612);
or U5818 (N_5818,N_5748,N_5780);
nand U5819 (N_5819,N_5613,N_5691);
xnor U5820 (N_5820,N_5639,N_5688);
nand U5821 (N_5821,N_5673,N_5771);
or U5822 (N_5822,N_5729,N_5606);
nand U5823 (N_5823,N_5700,N_5625);
and U5824 (N_5824,N_5628,N_5717);
or U5825 (N_5825,N_5744,N_5797);
and U5826 (N_5826,N_5685,N_5724);
nand U5827 (N_5827,N_5620,N_5651);
and U5828 (N_5828,N_5668,N_5624);
and U5829 (N_5829,N_5714,N_5796);
xor U5830 (N_5830,N_5601,N_5786);
nand U5831 (N_5831,N_5773,N_5799);
or U5832 (N_5832,N_5605,N_5740);
xnor U5833 (N_5833,N_5734,N_5677);
and U5834 (N_5834,N_5745,N_5750);
nor U5835 (N_5835,N_5792,N_5636);
nand U5836 (N_5836,N_5607,N_5743);
and U5837 (N_5837,N_5614,N_5656);
nand U5838 (N_5838,N_5728,N_5662);
and U5839 (N_5839,N_5690,N_5712);
and U5840 (N_5840,N_5604,N_5751);
nand U5841 (N_5841,N_5732,N_5770);
nand U5842 (N_5842,N_5618,N_5623);
nor U5843 (N_5843,N_5643,N_5713);
and U5844 (N_5844,N_5682,N_5622);
or U5845 (N_5845,N_5784,N_5689);
xnor U5846 (N_5846,N_5757,N_5737);
nand U5847 (N_5847,N_5735,N_5695);
xor U5848 (N_5848,N_5671,N_5642);
nor U5849 (N_5849,N_5754,N_5730);
xnor U5850 (N_5850,N_5727,N_5704);
nor U5851 (N_5851,N_5758,N_5752);
and U5852 (N_5852,N_5694,N_5697);
nor U5853 (N_5853,N_5763,N_5708);
or U5854 (N_5854,N_5733,N_5666);
nand U5855 (N_5855,N_5753,N_5672);
or U5856 (N_5856,N_5648,N_5678);
xor U5857 (N_5857,N_5608,N_5769);
xor U5858 (N_5858,N_5783,N_5600);
and U5859 (N_5859,N_5602,N_5785);
and U5860 (N_5860,N_5616,N_5657);
nand U5861 (N_5861,N_5634,N_5664);
and U5862 (N_5862,N_5627,N_5603);
nor U5863 (N_5863,N_5675,N_5723);
or U5864 (N_5864,N_5630,N_5667);
or U5865 (N_5865,N_5631,N_5790);
nor U5866 (N_5866,N_5794,N_5756);
and U5867 (N_5867,N_5777,N_5759);
nand U5868 (N_5868,N_5644,N_5680);
nand U5869 (N_5869,N_5721,N_5640);
nand U5870 (N_5870,N_5707,N_5659);
xor U5871 (N_5871,N_5703,N_5749);
or U5872 (N_5872,N_5660,N_5658);
nor U5873 (N_5873,N_5646,N_5779);
xor U5874 (N_5874,N_5615,N_5755);
and U5875 (N_5875,N_5661,N_5665);
xor U5876 (N_5876,N_5626,N_5731);
xor U5877 (N_5877,N_5746,N_5776);
and U5878 (N_5878,N_5650,N_5716);
xnor U5879 (N_5879,N_5621,N_5696);
xor U5880 (N_5880,N_5702,N_5747);
or U5881 (N_5881,N_5798,N_5641);
or U5882 (N_5882,N_5793,N_5674);
xor U5883 (N_5883,N_5791,N_5610);
nand U5884 (N_5884,N_5741,N_5722);
xnor U5885 (N_5885,N_5652,N_5655);
xor U5886 (N_5886,N_5683,N_5774);
nor U5887 (N_5887,N_5649,N_5765);
or U5888 (N_5888,N_5645,N_5629);
nand U5889 (N_5889,N_5767,N_5669);
xor U5890 (N_5890,N_5654,N_5653);
nand U5891 (N_5891,N_5775,N_5778);
and U5892 (N_5892,N_5720,N_5761);
xnor U5893 (N_5893,N_5711,N_5676);
or U5894 (N_5894,N_5766,N_5772);
nor U5895 (N_5895,N_5710,N_5725);
nor U5896 (N_5896,N_5637,N_5679);
nand U5897 (N_5897,N_5699,N_5738);
nand U5898 (N_5898,N_5781,N_5686);
nand U5899 (N_5899,N_5609,N_5719);
xor U5900 (N_5900,N_5688,N_5680);
and U5901 (N_5901,N_5709,N_5794);
and U5902 (N_5902,N_5733,N_5650);
or U5903 (N_5903,N_5601,N_5609);
xnor U5904 (N_5904,N_5738,N_5687);
and U5905 (N_5905,N_5717,N_5680);
and U5906 (N_5906,N_5711,N_5776);
nand U5907 (N_5907,N_5728,N_5671);
or U5908 (N_5908,N_5692,N_5792);
nand U5909 (N_5909,N_5765,N_5754);
or U5910 (N_5910,N_5623,N_5627);
nand U5911 (N_5911,N_5600,N_5774);
or U5912 (N_5912,N_5737,N_5656);
and U5913 (N_5913,N_5794,N_5726);
or U5914 (N_5914,N_5638,N_5776);
nor U5915 (N_5915,N_5730,N_5780);
or U5916 (N_5916,N_5655,N_5744);
and U5917 (N_5917,N_5744,N_5735);
or U5918 (N_5918,N_5714,N_5607);
nor U5919 (N_5919,N_5604,N_5715);
or U5920 (N_5920,N_5678,N_5785);
xor U5921 (N_5921,N_5663,N_5680);
nand U5922 (N_5922,N_5644,N_5695);
nor U5923 (N_5923,N_5750,N_5701);
and U5924 (N_5924,N_5733,N_5608);
and U5925 (N_5925,N_5747,N_5635);
or U5926 (N_5926,N_5762,N_5780);
xnor U5927 (N_5927,N_5666,N_5709);
or U5928 (N_5928,N_5777,N_5744);
and U5929 (N_5929,N_5783,N_5734);
and U5930 (N_5930,N_5741,N_5628);
nand U5931 (N_5931,N_5657,N_5678);
nand U5932 (N_5932,N_5662,N_5776);
nor U5933 (N_5933,N_5664,N_5684);
and U5934 (N_5934,N_5711,N_5643);
nor U5935 (N_5935,N_5613,N_5745);
nor U5936 (N_5936,N_5677,N_5667);
nor U5937 (N_5937,N_5699,N_5779);
xnor U5938 (N_5938,N_5767,N_5788);
nand U5939 (N_5939,N_5717,N_5657);
and U5940 (N_5940,N_5719,N_5768);
or U5941 (N_5941,N_5799,N_5775);
nand U5942 (N_5942,N_5676,N_5708);
and U5943 (N_5943,N_5703,N_5745);
xor U5944 (N_5944,N_5669,N_5783);
xnor U5945 (N_5945,N_5763,N_5694);
nand U5946 (N_5946,N_5663,N_5720);
nor U5947 (N_5947,N_5773,N_5628);
or U5948 (N_5948,N_5762,N_5668);
nor U5949 (N_5949,N_5718,N_5686);
or U5950 (N_5950,N_5733,N_5655);
nand U5951 (N_5951,N_5638,N_5692);
and U5952 (N_5952,N_5699,N_5718);
xor U5953 (N_5953,N_5765,N_5662);
xor U5954 (N_5954,N_5788,N_5618);
nand U5955 (N_5955,N_5657,N_5606);
nand U5956 (N_5956,N_5748,N_5740);
and U5957 (N_5957,N_5691,N_5772);
nor U5958 (N_5958,N_5674,N_5641);
and U5959 (N_5959,N_5752,N_5772);
nand U5960 (N_5960,N_5698,N_5643);
and U5961 (N_5961,N_5762,N_5791);
nor U5962 (N_5962,N_5774,N_5656);
and U5963 (N_5963,N_5729,N_5654);
or U5964 (N_5964,N_5715,N_5727);
nor U5965 (N_5965,N_5644,N_5668);
or U5966 (N_5966,N_5718,N_5663);
nand U5967 (N_5967,N_5700,N_5650);
xor U5968 (N_5968,N_5619,N_5701);
or U5969 (N_5969,N_5761,N_5706);
and U5970 (N_5970,N_5649,N_5724);
xnor U5971 (N_5971,N_5779,N_5771);
nor U5972 (N_5972,N_5754,N_5678);
nand U5973 (N_5973,N_5670,N_5663);
xor U5974 (N_5974,N_5704,N_5792);
xor U5975 (N_5975,N_5719,N_5605);
nand U5976 (N_5976,N_5780,N_5707);
and U5977 (N_5977,N_5776,N_5775);
or U5978 (N_5978,N_5623,N_5784);
nand U5979 (N_5979,N_5655,N_5751);
nor U5980 (N_5980,N_5772,N_5610);
and U5981 (N_5981,N_5657,N_5691);
and U5982 (N_5982,N_5626,N_5676);
nand U5983 (N_5983,N_5606,N_5742);
nor U5984 (N_5984,N_5688,N_5709);
xnor U5985 (N_5985,N_5732,N_5663);
and U5986 (N_5986,N_5722,N_5762);
and U5987 (N_5987,N_5751,N_5629);
xor U5988 (N_5988,N_5628,N_5793);
nor U5989 (N_5989,N_5754,N_5691);
and U5990 (N_5990,N_5755,N_5685);
nor U5991 (N_5991,N_5625,N_5775);
nor U5992 (N_5992,N_5667,N_5776);
xor U5993 (N_5993,N_5774,N_5637);
nand U5994 (N_5994,N_5765,N_5782);
nor U5995 (N_5995,N_5682,N_5628);
and U5996 (N_5996,N_5738,N_5676);
nand U5997 (N_5997,N_5628,N_5727);
xnor U5998 (N_5998,N_5674,N_5693);
xor U5999 (N_5999,N_5629,N_5737);
nor U6000 (N_6000,N_5942,N_5822);
nor U6001 (N_6001,N_5930,N_5975);
nor U6002 (N_6002,N_5964,N_5988);
and U6003 (N_6003,N_5808,N_5998);
nor U6004 (N_6004,N_5961,N_5934);
nand U6005 (N_6005,N_5918,N_5814);
xnor U6006 (N_6006,N_5993,N_5864);
and U6007 (N_6007,N_5804,N_5953);
and U6008 (N_6008,N_5849,N_5928);
or U6009 (N_6009,N_5818,N_5875);
nor U6010 (N_6010,N_5872,N_5938);
or U6011 (N_6011,N_5878,N_5882);
and U6012 (N_6012,N_5974,N_5979);
and U6013 (N_6013,N_5980,N_5807);
xnor U6014 (N_6014,N_5803,N_5880);
and U6015 (N_6015,N_5919,N_5831);
nor U6016 (N_6016,N_5863,N_5970);
and U6017 (N_6017,N_5990,N_5865);
xnor U6018 (N_6018,N_5945,N_5890);
and U6019 (N_6019,N_5892,N_5869);
and U6020 (N_6020,N_5936,N_5944);
nor U6021 (N_6021,N_5940,N_5903);
or U6022 (N_6022,N_5911,N_5985);
or U6023 (N_6023,N_5943,N_5867);
and U6024 (N_6024,N_5810,N_5871);
nand U6025 (N_6025,N_5846,N_5824);
nand U6026 (N_6026,N_5948,N_5819);
and U6027 (N_6027,N_5897,N_5848);
xor U6028 (N_6028,N_5837,N_5922);
nor U6029 (N_6029,N_5832,N_5895);
nand U6030 (N_6030,N_5915,N_5909);
or U6031 (N_6031,N_5853,N_5820);
and U6032 (N_6032,N_5976,N_5874);
xor U6033 (N_6033,N_5830,N_5902);
and U6034 (N_6034,N_5826,N_5941);
nand U6035 (N_6035,N_5883,N_5947);
nor U6036 (N_6036,N_5862,N_5994);
and U6037 (N_6037,N_5933,N_5825);
nor U6038 (N_6038,N_5870,N_5997);
or U6039 (N_6039,N_5885,N_5817);
nor U6040 (N_6040,N_5829,N_5861);
and U6041 (N_6041,N_5811,N_5840);
and U6042 (N_6042,N_5876,N_5937);
xnor U6043 (N_6043,N_5982,N_5821);
or U6044 (N_6044,N_5987,N_5992);
and U6045 (N_6045,N_5801,N_5905);
nand U6046 (N_6046,N_5886,N_5900);
xor U6047 (N_6047,N_5963,N_5884);
xnor U6048 (N_6048,N_5802,N_5910);
or U6049 (N_6049,N_5838,N_5860);
nor U6050 (N_6050,N_5855,N_5908);
or U6051 (N_6051,N_5844,N_5981);
nor U6052 (N_6052,N_5931,N_5839);
or U6053 (N_6053,N_5952,N_5901);
or U6054 (N_6054,N_5923,N_5868);
nand U6055 (N_6055,N_5973,N_5812);
xnor U6056 (N_6056,N_5996,N_5956);
xor U6057 (N_6057,N_5989,N_5881);
and U6058 (N_6058,N_5913,N_5929);
xnor U6059 (N_6059,N_5958,N_5856);
and U6060 (N_6060,N_5894,N_5898);
xnor U6061 (N_6061,N_5806,N_5957);
or U6062 (N_6062,N_5834,N_5916);
nor U6063 (N_6063,N_5950,N_5850);
and U6064 (N_6064,N_5827,N_5984);
xor U6065 (N_6065,N_5800,N_5926);
xor U6066 (N_6066,N_5845,N_5962);
nor U6067 (N_6067,N_5968,N_5967);
nor U6068 (N_6068,N_5907,N_5983);
and U6069 (N_6069,N_5977,N_5912);
nand U6070 (N_6070,N_5888,N_5891);
nand U6071 (N_6071,N_5971,N_5866);
nand U6072 (N_6072,N_5854,N_5935);
xor U6073 (N_6073,N_5966,N_5805);
nor U6074 (N_6074,N_5978,N_5965);
nor U6075 (N_6075,N_5927,N_5960);
nand U6076 (N_6076,N_5925,N_5843);
xnor U6077 (N_6077,N_5921,N_5951);
or U6078 (N_6078,N_5813,N_5924);
xor U6079 (N_6079,N_5842,N_5887);
nand U6080 (N_6080,N_5920,N_5859);
xnor U6081 (N_6081,N_5954,N_5858);
nor U6082 (N_6082,N_5857,N_5816);
nor U6083 (N_6083,N_5893,N_5889);
xnor U6084 (N_6084,N_5946,N_5877);
xor U6085 (N_6085,N_5986,N_5906);
nor U6086 (N_6086,N_5815,N_5939);
and U6087 (N_6087,N_5904,N_5847);
xor U6088 (N_6088,N_5991,N_5969);
and U6089 (N_6089,N_5809,N_5995);
xor U6090 (N_6090,N_5932,N_5959);
xor U6091 (N_6091,N_5896,N_5835);
nor U6092 (N_6092,N_5828,N_5972);
nor U6093 (N_6093,N_5899,N_5949);
xnor U6094 (N_6094,N_5851,N_5879);
or U6095 (N_6095,N_5841,N_5917);
nand U6096 (N_6096,N_5833,N_5852);
nand U6097 (N_6097,N_5999,N_5823);
nand U6098 (N_6098,N_5955,N_5914);
nor U6099 (N_6099,N_5873,N_5836);
and U6100 (N_6100,N_5916,N_5983);
and U6101 (N_6101,N_5903,N_5952);
nor U6102 (N_6102,N_5851,N_5869);
or U6103 (N_6103,N_5829,N_5966);
xnor U6104 (N_6104,N_5945,N_5807);
and U6105 (N_6105,N_5923,N_5853);
nand U6106 (N_6106,N_5932,N_5958);
or U6107 (N_6107,N_5935,N_5967);
xnor U6108 (N_6108,N_5984,N_5964);
or U6109 (N_6109,N_5950,N_5999);
nor U6110 (N_6110,N_5904,N_5851);
xnor U6111 (N_6111,N_5841,N_5830);
nand U6112 (N_6112,N_5825,N_5838);
nor U6113 (N_6113,N_5957,N_5956);
nor U6114 (N_6114,N_5852,N_5953);
and U6115 (N_6115,N_5850,N_5874);
or U6116 (N_6116,N_5997,N_5819);
or U6117 (N_6117,N_5874,N_5982);
nand U6118 (N_6118,N_5965,N_5856);
nand U6119 (N_6119,N_5896,N_5857);
xor U6120 (N_6120,N_5802,N_5988);
nor U6121 (N_6121,N_5928,N_5899);
nand U6122 (N_6122,N_5951,N_5891);
nand U6123 (N_6123,N_5954,N_5821);
and U6124 (N_6124,N_5955,N_5824);
nor U6125 (N_6125,N_5886,N_5802);
xor U6126 (N_6126,N_5869,N_5803);
nand U6127 (N_6127,N_5990,N_5963);
or U6128 (N_6128,N_5886,N_5836);
or U6129 (N_6129,N_5809,N_5931);
xor U6130 (N_6130,N_5902,N_5940);
nand U6131 (N_6131,N_5926,N_5923);
nand U6132 (N_6132,N_5910,N_5861);
xnor U6133 (N_6133,N_5966,N_5819);
nor U6134 (N_6134,N_5911,N_5924);
nor U6135 (N_6135,N_5936,N_5902);
or U6136 (N_6136,N_5975,N_5971);
xnor U6137 (N_6137,N_5860,N_5869);
or U6138 (N_6138,N_5961,N_5885);
nor U6139 (N_6139,N_5942,N_5934);
or U6140 (N_6140,N_5941,N_5972);
or U6141 (N_6141,N_5936,N_5842);
and U6142 (N_6142,N_5832,N_5951);
nand U6143 (N_6143,N_5990,N_5877);
nand U6144 (N_6144,N_5806,N_5866);
xnor U6145 (N_6145,N_5894,N_5991);
and U6146 (N_6146,N_5834,N_5880);
or U6147 (N_6147,N_5855,N_5846);
or U6148 (N_6148,N_5895,N_5948);
and U6149 (N_6149,N_5829,N_5887);
nand U6150 (N_6150,N_5958,N_5867);
nor U6151 (N_6151,N_5904,N_5996);
or U6152 (N_6152,N_5829,N_5925);
xor U6153 (N_6153,N_5914,N_5960);
nand U6154 (N_6154,N_5907,N_5935);
xor U6155 (N_6155,N_5846,N_5987);
nand U6156 (N_6156,N_5878,N_5912);
xor U6157 (N_6157,N_5822,N_5814);
or U6158 (N_6158,N_5820,N_5917);
and U6159 (N_6159,N_5807,N_5888);
xnor U6160 (N_6160,N_5868,N_5817);
nand U6161 (N_6161,N_5944,N_5846);
or U6162 (N_6162,N_5878,N_5942);
nand U6163 (N_6163,N_5817,N_5802);
xnor U6164 (N_6164,N_5915,N_5896);
or U6165 (N_6165,N_5824,N_5800);
and U6166 (N_6166,N_5858,N_5840);
or U6167 (N_6167,N_5860,N_5893);
and U6168 (N_6168,N_5974,N_5859);
nand U6169 (N_6169,N_5950,N_5882);
nor U6170 (N_6170,N_5812,N_5926);
xor U6171 (N_6171,N_5847,N_5874);
or U6172 (N_6172,N_5939,N_5862);
nand U6173 (N_6173,N_5847,N_5828);
or U6174 (N_6174,N_5860,N_5875);
xor U6175 (N_6175,N_5887,N_5803);
or U6176 (N_6176,N_5951,N_5865);
nand U6177 (N_6177,N_5845,N_5999);
nand U6178 (N_6178,N_5831,N_5974);
and U6179 (N_6179,N_5900,N_5924);
nor U6180 (N_6180,N_5931,N_5875);
xor U6181 (N_6181,N_5980,N_5906);
and U6182 (N_6182,N_5895,N_5874);
xnor U6183 (N_6183,N_5899,N_5829);
nor U6184 (N_6184,N_5816,N_5980);
or U6185 (N_6185,N_5954,N_5919);
and U6186 (N_6186,N_5974,N_5962);
xnor U6187 (N_6187,N_5845,N_5953);
nand U6188 (N_6188,N_5927,N_5996);
or U6189 (N_6189,N_5851,N_5846);
nand U6190 (N_6190,N_5928,N_5914);
nor U6191 (N_6191,N_5982,N_5847);
nor U6192 (N_6192,N_5971,N_5988);
and U6193 (N_6193,N_5833,N_5819);
and U6194 (N_6194,N_5949,N_5929);
nand U6195 (N_6195,N_5971,N_5872);
and U6196 (N_6196,N_5885,N_5805);
nor U6197 (N_6197,N_5995,N_5847);
nor U6198 (N_6198,N_5985,N_5810);
xor U6199 (N_6199,N_5919,N_5900);
or U6200 (N_6200,N_6101,N_6147);
nor U6201 (N_6201,N_6180,N_6185);
xor U6202 (N_6202,N_6001,N_6171);
xor U6203 (N_6203,N_6014,N_6030);
and U6204 (N_6204,N_6065,N_6055);
or U6205 (N_6205,N_6051,N_6164);
xnor U6206 (N_6206,N_6034,N_6059);
nor U6207 (N_6207,N_6197,N_6140);
nor U6208 (N_6208,N_6003,N_6125);
nor U6209 (N_6209,N_6150,N_6015);
or U6210 (N_6210,N_6124,N_6033);
nor U6211 (N_6211,N_6190,N_6081);
xnor U6212 (N_6212,N_6174,N_6116);
or U6213 (N_6213,N_6073,N_6079);
xor U6214 (N_6214,N_6069,N_6176);
and U6215 (N_6215,N_6187,N_6144);
xor U6216 (N_6216,N_6184,N_6156);
or U6217 (N_6217,N_6021,N_6026);
nor U6218 (N_6218,N_6017,N_6110);
nand U6219 (N_6219,N_6106,N_6177);
and U6220 (N_6220,N_6158,N_6083);
nor U6221 (N_6221,N_6138,N_6011);
or U6222 (N_6222,N_6092,N_6007);
and U6223 (N_6223,N_6107,N_6086);
or U6224 (N_6224,N_6052,N_6152);
xor U6225 (N_6225,N_6078,N_6148);
nand U6226 (N_6226,N_6044,N_6149);
nor U6227 (N_6227,N_6025,N_6043);
and U6228 (N_6228,N_6120,N_6153);
or U6229 (N_6229,N_6133,N_6159);
and U6230 (N_6230,N_6145,N_6023);
or U6231 (N_6231,N_6090,N_6084);
xor U6232 (N_6232,N_6002,N_6009);
and U6233 (N_6233,N_6006,N_6032);
nand U6234 (N_6234,N_6188,N_6104);
nand U6235 (N_6235,N_6196,N_6024);
nor U6236 (N_6236,N_6022,N_6061);
and U6237 (N_6237,N_6047,N_6020);
xor U6238 (N_6238,N_6045,N_6127);
nand U6239 (N_6239,N_6041,N_6097);
nand U6240 (N_6240,N_6039,N_6082);
and U6241 (N_6241,N_6040,N_6103);
xor U6242 (N_6242,N_6170,N_6042);
or U6243 (N_6243,N_6189,N_6109);
xor U6244 (N_6244,N_6129,N_6013);
xor U6245 (N_6245,N_6178,N_6076);
xnor U6246 (N_6246,N_6058,N_6105);
or U6247 (N_6247,N_6095,N_6010);
and U6248 (N_6248,N_6067,N_6169);
or U6249 (N_6249,N_6191,N_6155);
xor U6250 (N_6250,N_6028,N_6072);
nand U6251 (N_6251,N_6100,N_6050);
and U6252 (N_6252,N_6060,N_6080);
xor U6253 (N_6253,N_6192,N_6165);
nor U6254 (N_6254,N_6122,N_6054);
xor U6255 (N_6255,N_6161,N_6195);
nand U6256 (N_6256,N_6181,N_6099);
or U6257 (N_6257,N_6089,N_6175);
or U6258 (N_6258,N_6085,N_6131);
and U6259 (N_6259,N_6031,N_6114);
and U6260 (N_6260,N_6112,N_6027);
xnor U6261 (N_6261,N_6179,N_6056);
and U6262 (N_6262,N_6005,N_6071);
nand U6263 (N_6263,N_6064,N_6198);
xor U6264 (N_6264,N_6016,N_6193);
and U6265 (N_6265,N_6141,N_6008);
nor U6266 (N_6266,N_6173,N_6019);
and U6267 (N_6267,N_6194,N_6098);
xor U6268 (N_6268,N_6046,N_6121);
nand U6269 (N_6269,N_6000,N_6057);
or U6270 (N_6270,N_6063,N_6018);
nand U6271 (N_6271,N_6162,N_6029);
or U6272 (N_6272,N_6130,N_6111);
nand U6273 (N_6273,N_6137,N_6087);
or U6274 (N_6274,N_6167,N_6183);
or U6275 (N_6275,N_6142,N_6119);
and U6276 (N_6276,N_6038,N_6186);
xor U6277 (N_6277,N_6151,N_6077);
or U6278 (N_6278,N_6126,N_6108);
nor U6279 (N_6279,N_6146,N_6049);
xnor U6280 (N_6280,N_6132,N_6182);
or U6281 (N_6281,N_6136,N_6035);
nand U6282 (N_6282,N_6053,N_6062);
or U6283 (N_6283,N_6115,N_6168);
or U6284 (N_6284,N_6157,N_6066);
or U6285 (N_6285,N_6091,N_6075);
nand U6286 (N_6286,N_6135,N_6093);
or U6287 (N_6287,N_6088,N_6070);
and U6288 (N_6288,N_6134,N_6128);
xnor U6289 (N_6289,N_6163,N_6048);
and U6290 (N_6290,N_6172,N_6118);
nor U6291 (N_6291,N_6102,N_6037);
and U6292 (N_6292,N_6004,N_6012);
or U6293 (N_6293,N_6143,N_6068);
nand U6294 (N_6294,N_6166,N_6074);
xnor U6295 (N_6295,N_6139,N_6113);
or U6296 (N_6296,N_6123,N_6096);
nor U6297 (N_6297,N_6199,N_6094);
or U6298 (N_6298,N_6036,N_6160);
and U6299 (N_6299,N_6117,N_6154);
and U6300 (N_6300,N_6015,N_6047);
nand U6301 (N_6301,N_6143,N_6022);
or U6302 (N_6302,N_6099,N_6084);
nand U6303 (N_6303,N_6170,N_6072);
xnor U6304 (N_6304,N_6109,N_6014);
or U6305 (N_6305,N_6168,N_6079);
nor U6306 (N_6306,N_6129,N_6032);
and U6307 (N_6307,N_6081,N_6030);
xnor U6308 (N_6308,N_6056,N_6072);
xnor U6309 (N_6309,N_6180,N_6162);
xnor U6310 (N_6310,N_6157,N_6006);
nand U6311 (N_6311,N_6126,N_6171);
or U6312 (N_6312,N_6123,N_6164);
nand U6313 (N_6313,N_6023,N_6064);
nor U6314 (N_6314,N_6161,N_6083);
xor U6315 (N_6315,N_6059,N_6088);
nor U6316 (N_6316,N_6068,N_6000);
nand U6317 (N_6317,N_6053,N_6168);
and U6318 (N_6318,N_6113,N_6003);
nor U6319 (N_6319,N_6179,N_6030);
nor U6320 (N_6320,N_6006,N_6101);
xnor U6321 (N_6321,N_6132,N_6056);
nor U6322 (N_6322,N_6171,N_6079);
nor U6323 (N_6323,N_6133,N_6011);
or U6324 (N_6324,N_6015,N_6095);
nand U6325 (N_6325,N_6059,N_6139);
or U6326 (N_6326,N_6125,N_6002);
xor U6327 (N_6327,N_6099,N_6159);
nand U6328 (N_6328,N_6059,N_6119);
xor U6329 (N_6329,N_6149,N_6117);
and U6330 (N_6330,N_6013,N_6119);
and U6331 (N_6331,N_6081,N_6177);
or U6332 (N_6332,N_6127,N_6061);
nor U6333 (N_6333,N_6076,N_6094);
nand U6334 (N_6334,N_6034,N_6126);
or U6335 (N_6335,N_6138,N_6198);
or U6336 (N_6336,N_6062,N_6145);
and U6337 (N_6337,N_6081,N_6181);
nand U6338 (N_6338,N_6082,N_6141);
and U6339 (N_6339,N_6139,N_6101);
nand U6340 (N_6340,N_6137,N_6044);
and U6341 (N_6341,N_6065,N_6185);
or U6342 (N_6342,N_6043,N_6078);
nand U6343 (N_6343,N_6121,N_6079);
xor U6344 (N_6344,N_6180,N_6059);
xor U6345 (N_6345,N_6192,N_6110);
and U6346 (N_6346,N_6150,N_6036);
nor U6347 (N_6347,N_6000,N_6054);
nand U6348 (N_6348,N_6149,N_6081);
nand U6349 (N_6349,N_6128,N_6121);
or U6350 (N_6350,N_6086,N_6072);
xnor U6351 (N_6351,N_6115,N_6160);
xor U6352 (N_6352,N_6165,N_6061);
nand U6353 (N_6353,N_6154,N_6054);
nand U6354 (N_6354,N_6061,N_6107);
xnor U6355 (N_6355,N_6086,N_6082);
nor U6356 (N_6356,N_6137,N_6172);
or U6357 (N_6357,N_6015,N_6193);
and U6358 (N_6358,N_6098,N_6061);
nor U6359 (N_6359,N_6022,N_6157);
and U6360 (N_6360,N_6034,N_6092);
xnor U6361 (N_6361,N_6064,N_6089);
or U6362 (N_6362,N_6138,N_6101);
or U6363 (N_6363,N_6011,N_6179);
nor U6364 (N_6364,N_6094,N_6074);
and U6365 (N_6365,N_6006,N_6154);
xnor U6366 (N_6366,N_6172,N_6034);
and U6367 (N_6367,N_6015,N_6172);
nand U6368 (N_6368,N_6164,N_6139);
xor U6369 (N_6369,N_6083,N_6101);
nor U6370 (N_6370,N_6006,N_6179);
or U6371 (N_6371,N_6093,N_6100);
xor U6372 (N_6372,N_6077,N_6150);
nor U6373 (N_6373,N_6139,N_6086);
and U6374 (N_6374,N_6099,N_6049);
xor U6375 (N_6375,N_6062,N_6052);
xnor U6376 (N_6376,N_6125,N_6182);
and U6377 (N_6377,N_6040,N_6004);
nor U6378 (N_6378,N_6047,N_6036);
and U6379 (N_6379,N_6015,N_6199);
xnor U6380 (N_6380,N_6122,N_6096);
xor U6381 (N_6381,N_6069,N_6091);
nor U6382 (N_6382,N_6020,N_6026);
and U6383 (N_6383,N_6195,N_6096);
xnor U6384 (N_6384,N_6046,N_6107);
nand U6385 (N_6385,N_6105,N_6132);
or U6386 (N_6386,N_6009,N_6100);
and U6387 (N_6387,N_6186,N_6002);
nand U6388 (N_6388,N_6043,N_6115);
nand U6389 (N_6389,N_6007,N_6100);
and U6390 (N_6390,N_6154,N_6030);
xor U6391 (N_6391,N_6119,N_6168);
xnor U6392 (N_6392,N_6065,N_6161);
nor U6393 (N_6393,N_6175,N_6145);
nand U6394 (N_6394,N_6061,N_6136);
nor U6395 (N_6395,N_6124,N_6061);
xnor U6396 (N_6396,N_6024,N_6048);
nor U6397 (N_6397,N_6003,N_6124);
and U6398 (N_6398,N_6039,N_6014);
xnor U6399 (N_6399,N_6060,N_6057);
and U6400 (N_6400,N_6347,N_6246);
nor U6401 (N_6401,N_6330,N_6302);
nor U6402 (N_6402,N_6265,N_6393);
nand U6403 (N_6403,N_6343,N_6375);
xnor U6404 (N_6404,N_6206,N_6267);
or U6405 (N_6405,N_6345,N_6380);
nand U6406 (N_6406,N_6349,N_6276);
or U6407 (N_6407,N_6333,N_6279);
nand U6408 (N_6408,N_6224,N_6309);
xor U6409 (N_6409,N_6369,N_6383);
and U6410 (N_6410,N_6312,N_6386);
nor U6411 (N_6411,N_6325,N_6363);
nand U6412 (N_6412,N_6203,N_6323);
and U6413 (N_6413,N_6376,N_6313);
and U6414 (N_6414,N_6389,N_6213);
nor U6415 (N_6415,N_6377,N_6204);
nor U6416 (N_6416,N_6367,N_6299);
and U6417 (N_6417,N_6354,N_6327);
nand U6418 (N_6418,N_6215,N_6217);
or U6419 (N_6419,N_6227,N_6307);
nand U6420 (N_6420,N_6280,N_6270);
or U6421 (N_6421,N_6301,N_6252);
nor U6422 (N_6422,N_6228,N_6358);
xnor U6423 (N_6423,N_6262,N_6289);
xor U6424 (N_6424,N_6263,N_6306);
nand U6425 (N_6425,N_6310,N_6231);
nand U6426 (N_6426,N_6362,N_6374);
nand U6427 (N_6427,N_6371,N_6253);
and U6428 (N_6428,N_6230,N_6298);
and U6429 (N_6429,N_6281,N_6319);
nor U6430 (N_6430,N_6337,N_6266);
nand U6431 (N_6431,N_6241,N_6212);
nand U6432 (N_6432,N_6214,N_6304);
and U6433 (N_6433,N_6311,N_6248);
nand U6434 (N_6434,N_6342,N_6272);
xor U6435 (N_6435,N_6226,N_6382);
and U6436 (N_6436,N_6392,N_6200);
and U6437 (N_6437,N_6261,N_6300);
nor U6438 (N_6438,N_6317,N_6394);
nand U6439 (N_6439,N_6378,N_6348);
xnor U6440 (N_6440,N_6329,N_6355);
nand U6441 (N_6441,N_6294,N_6297);
nor U6442 (N_6442,N_6372,N_6225);
nand U6443 (N_6443,N_6397,N_6268);
and U6444 (N_6444,N_6336,N_6216);
nand U6445 (N_6445,N_6399,N_6287);
nor U6446 (N_6446,N_6249,N_6277);
xor U6447 (N_6447,N_6210,N_6335);
and U6448 (N_6448,N_6258,N_6219);
nor U6449 (N_6449,N_6364,N_6350);
xnor U6450 (N_6450,N_6283,N_6201);
nand U6451 (N_6451,N_6318,N_6385);
or U6452 (N_6452,N_6396,N_6388);
nor U6453 (N_6453,N_6223,N_6288);
and U6454 (N_6454,N_6292,N_6236);
nand U6455 (N_6455,N_6314,N_6321);
nand U6456 (N_6456,N_6282,N_6361);
or U6457 (N_6457,N_6229,N_6346);
nor U6458 (N_6458,N_6357,N_6290);
nand U6459 (N_6459,N_6332,N_6391);
nand U6460 (N_6460,N_6315,N_6308);
nor U6461 (N_6461,N_6232,N_6243);
and U6462 (N_6462,N_6221,N_6254);
nor U6463 (N_6463,N_6368,N_6260);
and U6464 (N_6464,N_6251,N_6398);
and U6465 (N_6465,N_6275,N_6328);
or U6466 (N_6466,N_6384,N_6295);
xnor U6467 (N_6467,N_6379,N_6285);
nor U6468 (N_6468,N_6341,N_6390);
xor U6469 (N_6469,N_6220,N_6274);
nand U6470 (N_6470,N_6353,N_6365);
or U6471 (N_6471,N_6381,N_6284);
nor U6472 (N_6472,N_6239,N_6247);
or U6473 (N_6473,N_6234,N_6395);
or U6474 (N_6474,N_6334,N_6351);
nor U6475 (N_6475,N_6360,N_6237);
xor U6476 (N_6476,N_6255,N_6240);
nor U6477 (N_6477,N_6244,N_6235);
nand U6478 (N_6478,N_6387,N_6324);
xor U6479 (N_6479,N_6370,N_6245);
nand U6480 (N_6480,N_6259,N_6256);
and U6481 (N_6481,N_6208,N_6242);
xor U6482 (N_6482,N_6233,N_6218);
nand U6483 (N_6483,N_6305,N_6238);
and U6484 (N_6484,N_6269,N_6202);
nand U6485 (N_6485,N_6322,N_6356);
nand U6486 (N_6486,N_6222,N_6273);
nand U6487 (N_6487,N_6340,N_6257);
or U6488 (N_6488,N_6296,N_6278);
nand U6489 (N_6489,N_6264,N_6291);
xor U6490 (N_6490,N_6339,N_6326);
xor U6491 (N_6491,N_6316,N_6293);
nor U6492 (N_6492,N_6211,N_6338);
nor U6493 (N_6493,N_6344,N_6331);
xor U6494 (N_6494,N_6250,N_6359);
or U6495 (N_6495,N_6207,N_6320);
and U6496 (N_6496,N_6205,N_6366);
or U6497 (N_6497,N_6352,N_6303);
xnor U6498 (N_6498,N_6373,N_6209);
nor U6499 (N_6499,N_6271,N_6286);
and U6500 (N_6500,N_6251,N_6385);
nor U6501 (N_6501,N_6322,N_6349);
nand U6502 (N_6502,N_6244,N_6363);
nor U6503 (N_6503,N_6295,N_6290);
nor U6504 (N_6504,N_6390,N_6383);
and U6505 (N_6505,N_6322,N_6378);
and U6506 (N_6506,N_6324,N_6205);
xnor U6507 (N_6507,N_6280,N_6382);
and U6508 (N_6508,N_6318,N_6258);
xnor U6509 (N_6509,N_6285,N_6305);
nand U6510 (N_6510,N_6228,N_6385);
and U6511 (N_6511,N_6289,N_6365);
and U6512 (N_6512,N_6390,N_6258);
nand U6513 (N_6513,N_6387,N_6216);
xnor U6514 (N_6514,N_6261,N_6299);
or U6515 (N_6515,N_6368,N_6206);
and U6516 (N_6516,N_6350,N_6352);
nor U6517 (N_6517,N_6365,N_6249);
and U6518 (N_6518,N_6308,N_6254);
nand U6519 (N_6519,N_6380,N_6315);
and U6520 (N_6520,N_6291,N_6215);
xnor U6521 (N_6521,N_6248,N_6308);
and U6522 (N_6522,N_6333,N_6284);
xor U6523 (N_6523,N_6352,N_6372);
xor U6524 (N_6524,N_6352,N_6323);
or U6525 (N_6525,N_6230,N_6307);
and U6526 (N_6526,N_6333,N_6339);
xnor U6527 (N_6527,N_6379,N_6393);
and U6528 (N_6528,N_6332,N_6324);
nand U6529 (N_6529,N_6234,N_6264);
nand U6530 (N_6530,N_6203,N_6300);
nor U6531 (N_6531,N_6242,N_6233);
or U6532 (N_6532,N_6344,N_6256);
nor U6533 (N_6533,N_6304,N_6356);
nor U6534 (N_6534,N_6270,N_6242);
and U6535 (N_6535,N_6376,N_6253);
nand U6536 (N_6536,N_6289,N_6332);
and U6537 (N_6537,N_6386,N_6317);
nor U6538 (N_6538,N_6216,N_6325);
nand U6539 (N_6539,N_6330,N_6326);
nor U6540 (N_6540,N_6224,N_6366);
or U6541 (N_6541,N_6288,N_6296);
and U6542 (N_6542,N_6277,N_6368);
nand U6543 (N_6543,N_6221,N_6348);
and U6544 (N_6544,N_6269,N_6236);
nand U6545 (N_6545,N_6255,N_6230);
and U6546 (N_6546,N_6330,N_6381);
nor U6547 (N_6547,N_6351,N_6258);
xor U6548 (N_6548,N_6214,N_6203);
nand U6549 (N_6549,N_6297,N_6357);
nor U6550 (N_6550,N_6356,N_6223);
nand U6551 (N_6551,N_6228,N_6314);
nand U6552 (N_6552,N_6342,N_6337);
and U6553 (N_6553,N_6304,N_6207);
or U6554 (N_6554,N_6280,N_6307);
and U6555 (N_6555,N_6363,N_6282);
xnor U6556 (N_6556,N_6286,N_6372);
nand U6557 (N_6557,N_6280,N_6392);
or U6558 (N_6558,N_6319,N_6232);
nor U6559 (N_6559,N_6323,N_6254);
nor U6560 (N_6560,N_6200,N_6365);
nand U6561 (N_6561,N_6345,N_6289);
nor U6562 (N_6562,N_6398,N_6214);
nand U6563 (N_6563,N_6234,N_6299);
xnor U6564 (N_6564,N_6384,N_6263);
or U6565 (N_6565,N_6291,N_6274);
nor U6566 (N_6566,N_6348,N_6330);
xnor U6567 (N_6567,N_6393,N_6285);
nand U6568 (N_6568,N_6200,N_6223);
nand U6569 (N_6569,N_6208,N_6350);
nand U6570 (N_6570,N_6389,N_6362);
xor U6571 (N_6571,N_6254,N_6209);
nand U6572 (N_6572,N_6353,N_6209);
xor U6573 (N_6573,N_6306,N_6385);
nor U6574 (N_6574,N_6201,N_6215);
xor U6575 (N_6575,N_6334,N_6263);
and U6576 (N_6576,N_6340,N_6202);
and U6577 (N_6577,N_6208,N_6201);
or U6578 (N_6578,N_6318,N_6243);
or U6579 (N_6579,N_6318,N_6275);
nand U6580 (N_6580,N_6238,N_6392);
and U6581 (N_6581,N_6357,N_6327);
xnor U6582 (N_6582,N_6309,N_6342);
and U6583 (N_6583,N_6388,N_6343);
xnor U6584 (N_6584,N_6333,N_6254);
nand U6585 (N_6585,N_6286,N_6246);
xor U6586 (N_6586,N_6365,N_6345);
nand U6587 (N_6587,N_6390,N_6326);
and U6588 (N_6588,N_6399,N_6271);
nor U6589 (N_6589,N_6360,N_6379);
nor U6590 (N_6590,N_6296,N_6260);
nor U6591 (N_6591,N_6334,N_6394);
and U6592 (N_6592,N_6364,N_6255);
xor U6593 (N_6593,N_6328,N_6259);
or U6594 (N_6594,N_6395,N_6204);
xnor U6595 (N_6595,N_6212,N_6310);
nand U6596 (N_6596,N_6347,N_6396);
nor U6597 (N_6597,N_6294,N_6310);
and U6598 (N_6598,N_6220,N_6242);
or U6599 (N_6599,N_6328,N_6350);
xor U6600 (N_6600,N_6428,N_6447);
and U6601 (N_6601,N_6480,N_6440);
xor U6602 (N_6602,N_6541,N_6427);
or U6603 (N_6603,N_6414,N_6548);
and U6604 (N_6604,N_6526,N_6423);
and U6605 (N_6605,N_6483,N_6402);
nand U6606 (N_6606,N_6468,N_6433);
nor U6607 (N_6607,N_6566,N_6481);
xnor U6608 (N_6608,N_6530,N_6524);
and U6609 (N_6609,N_6400,N_6422);
or U6610 (N_6610,N_6484,N_6574);
xnor U6611 (N_6611,N_6583,N_6426);
xor U6612 (N_6612,N_6489,N_6552);
xor U6613 (N_6613,N_6490,N_6515);
or U6614 (N_6614,N_6559,N_6417);
nand U6615 (N_6615,N_6505,N_6485);
nor U6616 (N_6616,N_6482,N_6424);
xnor U6617 (N_6617,N_6546,N_6436);
and U6618 (N_6618,N_6555,N_6533);
xnor U6619 (N_6619,N_6598,N_6445);
xor U6620 (N_6620,N_6579,N_6589);
xnor U6621 (N_6621,N_6547,N_6573);
nor U6622 (N_6622,N_6401,N_6560);
nand U6623 (N_6623,N_6487,N_6488);
and U6624 (N_6624,N_6502,N_6593);
or U6625 (N_6625,N_6512,N_6519);
or U6626 (N_6626,N_6495,N_6563);
or U6627 (N_6627,N_6464,N_6461);
nor U6628 (N_6628,N_6569,N_6588);
or U6629 (N_6629,N_6421,N_6458);
nand U6630 (N_6630,N_6514,N_6442);
xor U6631 (N_6631,N_6585,N_6457);
xor U6632 (N_6632,N_6599,N_6581);
and U6633 (N_6633,N_6580,N_6437);
xnor U6634 (N_6634,N_6407,N_6538);
nand U6635 (N_6635,N_6474,N_6439);
nand U6636 (N_6636,N_6410,N_6471);
xor U6637 (N_6637,N_6491,N_6497);
xnor U6638 (N_6638,N_6438,N_6578);
xor U6639 (N_6639,N_6516,N_6539);
nand U6640 (N_6640,N_6494,N_6405);
xnor U6641 (N_6641,N_6556,N_6592);
or U6642 (N_6642,N_6493,N_6465);
xor U6643 (N_6643,N_6492,N_6595);
and U6644 (N_6644,N_6476,N_6521);
nor U6645 (N_6645,N_6561,N_6544);
nor U6646 (N_6646,N_6420,N_6467);
and U6647 (N_6647,N_6527,N_6534);
and U6648 (N_6648,N_6403,N_6475);
nand U6649 (N_6649,N_6553,N_6434);
and U6650 (N_6650,N_6570,N_6511);
nor U6651 (N_6651,N_6411,N_6565);
xor U6652 (N_6652,N_6430,N_6409);
or U6653 (N_6653,N_6523,N_6575);
or U6654 (N_6654,N_6441,N_6562);
and U6655 (N_6655,N_6486,N_6504);
xor U6656 (N_6656,N_6522,N_6429);
or U6657 (N_6657,N_6597,N_6406);
nand U6658 (N_6658,N_6532,N_6454);
and U6659 (N_6659,N_6558,N_6413);
nand U6660 (N_6660,N_6448,N_6435);
xor U6661 (N_6661,N_6450,N_6477);
nand U6662 (N_6662,N_6451,N_6459);
nand U6663 (N_6663,N_6443,N_6517);
nor U6664 (N_6664,N_6528,N_6431);
nor U6665 (N_6665,N_6456,N_6567);
nand U6666 (N_6666,N_6582,N_6472);
xor U6667 (N_6667,N_6554,N_6478);
and U6668 (N_6668,N_6536,N_6463);
nand U6669 (N_6669,N_6576,N_6571);
xor U6670 (N_6670,N_6425,N_6473);
xnor U6671 (N_6671,N_6529,N_6568);
or U6672 (N_6672,N_6509,N_6503);
xor U6673 (N_6673,N_6543,N_6418);
or U6674 (N_6674,N_6594,N_6479);
nand U6675 (N_6675,N_6444,N_6408);
nand U6676 (N_6676,N_6590,N_6551);
and U6677 (N_6677,N_6549,N_6531);
or U6678 (N_6678,N_6577,N_6498);
xnor U6679 (N_6679,N_6542,N_6466);
nand U6680 (N_6680,N_6507,N_6499);
xnor U6681 (N_6681,N_6545,N_6518);
xnor U6682 (N_6682,N_6525,N_6469);
or U6683 (N_6683,N_6415,N_6412);
xnor U6684 (N_6684,N_6572,N_6419);
nor U6685 (N_6685,N_6513,N_6591);
nor U6686 (N_6686,N_6508,N_6596);
nor U6687 (N_6687,N_6537,N_6540);
xnor U6688 (N_6688,N_6455,N_6587);
or U6689 (N_6689,N_6432,N_6510);
xor U6690 (N_6690,N_6550,N_6416);
xnor U6691 (N_6691,N_6470,N_6500);
nor U6692 (N_6692,N_6496,N_6446);
nand U6693 (N_6693,N_6564,N_6535);
nand U6694 (N_6694,N_6506,N_6520);
and U6695 (N_6695,N_6586,N_6557);
nand U6696 (N_6696,N_6584,N_6462);
or U6697 (N_6697,N_6449,N_6452);
and U6698 (N_6698,N_6453,N_6460);
or U6699 (N_6699,N_6404,N_6501);
or U6700 (N_6700,N_6594,N_6580);
xor U6701 (N_6701,N_6569,N_6584);
nand U6702 (N_6702,N_6587,N_6418);
and U6703 (N_6703,N_6422,N_6431);
nand U6704 (N_6704,N_6580,N_6540);
or U6705 (N_6705,N_6545,N_6494);
xnor U6706 (N_6706,N_6450,N_6526);
nor U6707 (N_6707,N_6482,N_6459);
or U6708 (N_6708,N_6585,N_6574);
and U6709 (N_6709,N_6499,N_6401);
or U6710 (N_6710,N_6584,N_6408);
and U6711 (N_6711,N_6421,N_6544);
xnor U6712 (N_6712,N_6577,N_6453);
nand U6713 (N_6713,N_6499,N_6497);
nand U6714 (N_6714,N_6416,N_6415);
or U6715 (N_6715,N_6451,N_6552);
nand U6716 (N_6716,N_6495,N_6546);
or U6717 (N_6717,N_6445,N_6471);
or U6718 (N_6718,N_6588,N_6573);
xnor U6719 (N_6719,N_6414,N_6523);
nor U6720 (N_6720,N_6573,N_6578);
nor U6721 (N_6721,N_6574,N_6529);
or U6722 (N_6722,N_6435,N_6597);
nor U6723 (N_6723,N_6448,N_6436);
xor U6724 (N_6724,N_6591,N_6476);
nand U6725 (N_6725,N_6426,N_6572);
nand U6726 (N_6726,N_6448,N_6572);
and U6727 (N_6727,N_6544,N_6401);
nor U6728 (N_6728,N_6437,N_6574);
xor U6729 (N_6729,N_6400,N_6524);
and U6730 (N_6730,N_6580,N_6592);
nor U6731 (N_6731,N_6439,N_6518);
and U6732 (N_6732,N_6507,N_6588);
or U6733 (N_6733,N_6445,N_6480);
nand U6734 (N_6734,N_6560,N_6594);
and U6735 (N_6735,N_6429,N_6525);
nand U6736 (N_6736,N_6540,N_6464);
nor U6737 (N_6737,N_6430,N_6548);
nor U6738 (N_6738,N_6582,N_6558);
or U6739 (N_6739,N_6424,N_6517);
and U6740 (N_6740,N_6491,N_6461);
or U6741 (N_6741,N_6529,N_6598);
nand U6742 (N_6742,N_6404,N_6402);
and U6743 (N_6743,N_6431,N_6409);
xnor U6744 (N_6744,N_6527,N_6546);
or U6745 (N_6745,N_6516,N_6463);
and U6746 (N_6746,N_6421,N_6411);
or U6747 (N_6747,N_6454,N_6506);
nor U6748 (N_6748,N_6468,N_6449);
xor U6749 (N_6749,N_6479,N_6590);
or U6750 (N_6750,N_6410,N_6595);
xor U6751 (N_6751,N_6523,N_6515);
or U6752 (N_6752,N_6411,N_6446);
or U6753 (N_6753,N_6509,N_6475);
nand U6754 (N_6754,N_6462,N_6505);
xor U6755 (N_6755,N_6578,N_6450);
or U6756 (N_6756,N_6444,N_6474);
xnor U6757 (N_6757,N_6440,N_6463);
or U6758 (N_6758,N_6458,N_6568);
nor U6759 (N_6759,N_6520,N_6497);
nor U6760 (N_6760,N_6464,N_6445);
nand U6761 (N_6761,N_6500,N_6540);
or U6762 (N_6762,N_6462,N_6454);
or U6763 (N_6763,N_6557,N_6573);
xnor U6764 (N_6764,N_6402,N_6592);
or U6765 (N_6765,N_6471,N_6468);
and U6766 (N_6766,N_6539,N_6499);
nor U6767 (N_6767,N_6514,N_6586);
or U6768 (N_6768,N_6519,N_6404);
or U6769 (N_6769,N_6497,N_6432);
or U6770 (N_6770,N_6567,N_6473);
and U6771 (N_6771,N_6580,N_6446);
nand U6772 (N_6772,N_6439,N_6532);
nand U6773 (N_6773,N_6495,N_6433);
xnor U6774 (N_6774,N_6554,N_6564);
and U6775 (N_6775,N_6547,N_6493);
nor U6776 (N_6776,N_6506,N_6411);
nand U6777 (N_6777,N_6431,N_6454);
or U6778 (N_6778,N_6584,N_6507);
xor U6779 (N_6779,N_6534,N_6495);
nor U6780 (N_6780,N_6538,N_6459);
nor U6781 (N_6781,N_6589,N_6539);
nor U6782 (N_6782,N_6513,N_6548);
and U6783 (N_6783,N_6408,N_6526);
xor U6784 (N_6784,N_6407,N_6596);
and U6785 (N_6785,N_6415,N_6406);
nor U6786 (N_6786,N_6563,N_6464);
or U6787 (N_6787,N_6511,N_6451);
nor U6788 (N_6788,N_6494,N_6574);
nand U6789 (N_6789,N_6423,N_6491);
nor U6790 (N_6790,N_6410,N_6414);
nor U6791 (N_6791,N_6565,N_6488);
nor U6792 (N_6792,N_6590,N_6434);
xor U6793 (N_6793,N_6589,N_6534);
and U6794 (N_6794,N_6524,N_6532);
and U6795 (N_6795,N_6466,N_6400);
nor U6796 (N_6796,N_6560,N_6577);
nor U6797 (N_6797,N_6498,N_6431);
nor U6798 (N_6798,N_6410,N_6481);
and U6799 (N_6799,N_6437,N_6482);
nor U6800 (N_6800,N_6671,N_6655);
xnor U6801 (N_6801,N_6788,N_6689);
or U6802 (N_6802,N_6613,N_6694);
or U6803 (N_6803,N_6784,N_6697);
and U6804 (N_6804,N_6639,N_6740);
nand U6805 (N_6805,N_6628,N_6707);
or U6806 (N_6806,N_6736,N_6608);
and U6807 (N_6807,N_6731,N_6747);
nand U6808 (N_6808,N_6760,N_6629);
nor U6809 (N_6809,N_6786,N_6654);
nor U6810 (N_6810,N_6703,N_6710);
xor U6811 (N_6811,N_6781,N_6771);
and U6812 (N_6812,N_6785,N_6797);
and U6813 (N_6813,N_6763,N_6675);
nand U6814 (N_6814,N_6732,N_6657);
nand U6815 (N_6815,N_6630,N_6644);
nor U6816 (N_6816,N_6709,N_6772);
nor U6817 (N_6817,N_6787,N_6706);
xnor U6818 (N_6818,N_6789,N_6717);
nor U6819 (N_6819,N_6605,N_6770);
or U6820 (N_6820,N_6793,N_6688);
and U6821 (N_6821,N_6635,N_6725);
nand U6822 (N_6822,N_6708,N_6743);
nand U6823 (N_6823,N_6746,N_6666);
or U6824 (N_6824,N_6712,N_6691);
and U6825 (N_6825,N_6723,N_6701);
xnor U6826 (N_6826,N_6619,N_6609);
and U6827 (N_6827,N_6711,N_6631);
or U6828 (N_6828,N_6636,N_6659);
nand U6829 (N_6829,N_6751,N_6699);
nand U6830 (N_6830,N_6667,N_6752);
xor U6831 (N_6831,N_6766,N_6750);
nor U6832 (N_6832,N_6737,N_6670);
or U6833 (N_6833,N_6681,N_6662);
nor U6834 (N_6834,N_6791,N_6684);
nor U6835 (N_6835,N_6720,N_6647);
or U6836 (N_6836,N_6741,N_6764);
or U6837 (N_6837,N_6648,N_6674);
or U6838 (N_6838,N_6704,N_6767);
nor U6839 (N_6839,N_6730,N_6624);
or U6840 (N_6840,N_6601,N_6626);
or U6841 (N_6841,N_6738,N_6773);
nand U6842 (N_6842,N_6792,N_6685);
xnor U6843 (N_6843,N_6634,N_6759);
and U6844 (N_6844,N_6649,N_6769);
nand U6845 (N_6845,N_6661,N_6765);
nor U6846 (N_6846,N_6744,N_6753);
nor U6847 (N_6847,N_6627,N_6660);
nand U6848 (N_6848,N_6632,N_6729);
xor U6849 (N_6849,N_6693,N_6620);
or U6850 (N_6850,N_6728,N_6618);
and U6851 (N_6851,N_6762,N_6673);
xor U6852 (N_6852,N_6794,N_6748);
nand U6853 (N_6853,N_6603,N_6656);
xnor U6854 (N_6854,N_6796,N_6780);
nand U6855 (N_6855,N_6749,N_6652);
or U6856 (N_6856,N_6686,N_6611);
or U6857 (N_6857,N_6623,N_6768);
nor U6858 (N_6858,N_6739,N_6602);
xor U6859 (N_6859,N_6776,N_6724);
nand U6860 (N_6860,N_6692,N_6616);
and U6861 (N_6861,N_6641,N_6621);
xnor U6862 (N_6862,N_6690,N_6676);
or U6863 (N_6863,N_6622,N_6698);
or U6864 (N_6864,N_6663,N_6612);
xnor U6865 (N_6865,N_6757,N_6716);
nand U6866 (N_6866,N_6658,N_6735);
or U6867 (N_6867,N_6705,N_6798);
or U6868 (N_6868,N_6782,N_6640);
nand U6869 (N_6869,N_6617,N_6779);
nand U6870 (N_6870,N_6695,N_6680);
nor U6871 (N_6871,N_6715,N_6778);
nor U6872 (N_6872,N_6645,N_6677);
xor U6873 (N_6873,N_6646,N_6678);
nor U6874 (N_6874,N_6713,N_6669);
nand U6875 (N_6875,N_6625,N_6719);
and U6876 (N_6876,N_6718,N_6761);
nor U6877 (N_6877,N_6653,N_6722);
nand U6878 (N_6878,N_6756,N_6687);
and U6879 (N_6879,N_6615,N_6700);
and U6880 (N_6880,N_6643,N_6672);
nand U6881 (N_6881,N_6600,N_6777);
nor U6882 (N_6882,N_6696,N_6745);
xor U6883 (N_6883,N_6755,N_6758);
nand U6884 (N_6884,N_6790,N_6714);
nand U6885 (N_6885,N_6721,N_6650);
and U6886 (N_6886,N_6665,N_6633);
and U6887 (N_6887,N_6774,N_6651);
or U6888 (N_6888,N_6607,N_6642);
nand U6889 (N_6889,N_6799,N_6742);
nand U6890 (N_6890,N_6604,N_6606);
and U6891 (N_6891,N_6702,N_6683);
and U6892 (N_6892,N_6775,N_6783);
xnor U6893 (N_6893,N_6754,N_6727);
xor U6894 (N_6894,N_6614,N_6733);
xor U6895 (N_6895,N_6638,N_6682);
and U6896 (N_6896,N_6668,N_6734);
or U6897 (N_6897,N_6726,N_6795);
or U6898 (N_6898,N_6679,N_6664);
nand U6899 (N_6899,N_6610,N_6637);
nor U6900 (N_6900,N_6629,N_6674);
nand U6901 (N_6901,N_6632,N_6751);
nor U6902 (N_6902,N_6762,N_6704);
xor U6903 (N_6903,N_6639,N_6754);
or U6904 (N_6904,N_6695,N_6652);
nor U6905 (N_6905,N_6635,N_6682);
nor U6906 (N_6906,N_6727,N_6715);
and U6907 (N_6907,N_6645,N_6614);
nor U6908 (N_6908,N_6614,N_6669);
xnor U6909 (N_6909,N_6725,N_6673);
nand U6910 (N_6910,N_6751,N_6660);
nor U6911 (N_6911,N_6662,N_6714);
and U6912 (N_6912,N_6741,N_6690);
xnor U6913 (N_6913,N_6624,N_6620);
or U6914 (N_6914,N_6624,N_6654);
nand U6915 (N_6915,N_6753,N_6622);
and U6916 (N_6916,N_6656,N_6646);
xnor U6917 (N_6917,N_6688,N_6651);
nand U6918 (N_6918,N_6734,N_6765);
or U6919 (N_6919,N_6710,N_6652);
nor U6920 (N_6920,N_6644,N_6779);
nor U6921 (N_6921,N_6716,N_6721);
and U6922 (N_6922,N_6624,N_6670);
or U6923 (N_6923,N_6626,N_6696);
or U6924 (N_6924,N_6735,N_6769);
nor U6925 (N_6925,N_6782,N_6633);
or U6926 (N_6926,N_6710,N_6640);
nand U6927 (N_6927,N_6718,N_6749);
nand U6928 (N_6928,N_6749,N_6782);
nand U6929 (N_6929,N_6637,N_6621);
and U6930 (N_6930,N_6685,N_6627);
nor U6931 (N_6931,N_6628,N_6603);
or U6932 (N_6932,N_6645,N_6752);
nor U6933 (N_6933,N_6759,N_6707);
or U6934 (N_6934,N_6739,N_6601);
nor U6935 (N_6935,N_6718,N_6666);
and U6936 (N_6936,N_6670,N_6767);
xnor U6937 (N_6937,N_6723,N_6748);
and U6938 (N_6938,N_6619,N_6660);
or U6939 (N_6939,N_6755,N_6711);
nand U6940 (N_6940,N_6733,N_6642);
or U6941 (N_6941,N_6734,N_6742);
and U6942 (N_6942,N_6738,N_6618);
or U6943 (N_6943,N_6645,N_6782);
or U6944 (N_6944,N_6671,N_6753);
nand U6945 (N_6945,N_6620,N_6730);
xnor U6946 (N_6946,N_6675,N_6671);
xor U6947 (N_6947,N_6616,N_6752);
nand U6948 (N_6948,N_6605,N_6734);
nand U6949 (N_6949,N_6747,N_6739);
nor U6950 (N_6950,N_6608,N_6754);
nand U6951 (N_6951,N_6697,N_6711);
nor U6952 (N_6952,N_6707,N_6747);
xnor U6953 (N_6953,N_6747,N_6780);
or U6954 (N_6954,N_6792,N_6631);
xor U6955 (N_6955,N_6793,N_6707);
or U6956 (N_6956,N_6799,N_6712);
and U6957 (N_6957,N_6704,N_6659);
or U6958 (N_6958,N_6603,N_6790);
nand U6959 (N_6959,N_6740,N_6757);
xnor U6960 (N_6960,N_6620,N_6629);
xnor U6961 (N_6961,N_6663,N_6775);
or U6962 (N_6962,N_6677,N_6622);
nand U6963 (N_6963,N_6655,N_6710);
or U6964 (N_6964,N_6739,N_6766);
nor U6965 (N_6965,N_6642,N_6697);
nor U6966 (N_6966,N_6766,N_6717);
and U6967 (N_6967,N_6767,N_6797);
and U6968 (N_6968,N_6694,N_6655);
nand U6969 (N_6969,N_6757,N_6722);
nor U6970 (N_6970,N_6681,N_6791);
nand U6971 (N_6971,N_6618,N_6794);
and U6972 (N_6972,N_6741,N_6602);
xor U6973 (N_6973,N_6704,N_6721);
nand U6974 (N_6974,N_6762,N_6612);
or U6975 (N_6975,N_6704,N_6754);
xor U6976 (N_6976,N_6662,N_6744);
nand U6977 (N_6977,N_6647,N_6783);
and U6978 (N_6978,N_6776,N_6710);
or U6979 (N_6979,N_6789,N_6642);
nand U6980 (N_6980,N_6607,N_6623);
nand U6981 (N_6981,N_6713,N_6674);
nor U6982 (N_6982,N_6713,N_6710);
or U6983 (N_6983,N_6757,N_6744);
or U6984 (N_6984,N_6796,N_6639);
and U6985 (N_6985,N_6785,N_6683);
nor U6986 (N_6986,N_6759,N_6672);
nand U6987 (N_6987,N_6681,N_6659);
xor U6988 (N_6988,N_6684,N_6760);
nand U6989 (N_6989,N_6734,N_6769);
xor U6990 (N_6990,N_6610,N_6762);
nor U6991 (N_6991,N_6636,N_6746);
nand U6992 (N_6992,N_6650,N_6687);
and U6993 (N_6993,N_6693,N_6726);
or U6994 (N_6994,N_6625,N_6746);
and U6995 (N_6995,N_6717,N_6600);
xnor U6996 (N_6996,N_6613,N_6737);
nand U6997 (N_6997,N_6777,N_6787);
nand U6998 (N_6998,N_6782,N_6690);
nor U6999 (N_6999,N_6775,N_6794);
nor U7000 (N_7000,N_6908,N_6899);
nor U7001 (N_7001,N_6817,N_6871);
nand U7002 (N_7002,N_6863,N_6806);
nand U7003 (N_7003,N_6903,N_6893);
xnor U7004 (N_7004,N_6983,N_6858);
nor U7005 (N_7005,N_6952,N_6954);
and U7006 (N_7006,N_6913,N_6997);
and U7007 (N_7007,N_6855,N_6854);
nand U7008 (N_7008,N_6868,N_6955);
and U7009 (N_7009,N_6943,N_6818);
nand U7010 (N_7010,N_6852,N_6864);
nor U7011 (N_7011,N_6936,N_6946);
and U7012 (N_7012,N_6883,N_6842);
and U7013 (N_7013,N_6996,N_6870);
xnor U7014 (N_7014,N_6917,N_6982);
nor U7015 (N_7015,N_6987,N_6897);
nand U7016 (N_7016,N_6907,N_6921);
xor U7017 (N_7017,N_6840,N_6935);
or U7018 (N_7018,N_6991,N_6859);
or U7019 (N_7019,N_6999,N_6882);
nand U7020 (N_7020,N_6834,N_6822);
xnor U7021 (N_7021,N_6862,N_6984);
nor U7022 (N_7022,N_6888,N_6826);
nor U7023 (N_7023,N_6835,N_6975);
nor U7024 (N_7024,N_6985,N_6805);
and U7025 (N_7025,N_6986,N_6802);
and U7026 (N_7026,N_6895,N_6894);
and U7027 (N_7027,N_6965,N_6860);
or U7028 (N_7028,N_6973,N_6969);
nand U7029 (N_7029,N_6922,N_6937);
and U7030 (N_7030,N_6816,N_6823);
or U7031 (N_7031,N_6833,N_6953);
and U7032 (N_7032,N_6853,N_6905);
nor U7033 (N_7033,N_6803,N_6938);
or U7034 (N_7034,N_6872,N_6873);
nand U7035 (N_7035,N_6992,N_6876);
xor U7036 (N_7036,N_6980,N_6880);
and U7037 (N_7037,N_6819,N_6960);
xnor U7038 (N_7038,N_6841,N_6962);
and U7039 (N_7039,N_6977,N_6898);
nand U7040 (N_7040,N_6918,N_6912);
or U7041 (N_7041,N_6879,N_6887);
or U7042 (N_7042,N_6933,N_6844);
and U7043 (N_7043,N_6910,N_6845);
or U7044 (N_7044,N_6974,N_6911);
nor U7045 (N_7045,N_6972,N_6824);
and U7046 (N_7046,N_6808,N_6885);
or U7047 (N_7047,N_6837,N_6812);
xnor U7048 (N_7048,N_6990,N_6828);
or U7049 (N_7049,N_6998,N_6814);
nor U7050 (N_7050,N_6830,N_6940);
nor U7051 (N_7051,N_6931,N_6884);
xor U7052 (N_7052,N_6944,N_6861);
or U7053 (N_7053,N_6896,N_6923);
or U7054 (N_7054,N_6900,N_6889);
nand U7055 (N_7055,N_6988,N_6875);
nor U7056 (N_7056,N_6827,N_6971);
and U7057 (N_7057,N_6925,N_6831);
and U7058 (N_7058,N_6866,N_6950);
xor U7059 (N_7059,N_6915,N_6856);
nand U7060 (N_7060,N_6902,N_6949);
or U7061 (N_7061,N_6939,N_6924);
nand U7062 (N_7062,N_6994,N_6966);
nand U7063 (N_7063,N_6967,N_6981);
xor U7064 (N_7064,N_6843,N_6919);
or U7065 (N_7065,N_6820,N_6927);
nand U7066 (N_7066,N_6970,N_6821);
nand U7067 (N_7067,N_6904,N_6838);
and U7068 (N_7068,N_6825,N_6836);
nand U7069 (N_7069,N_6848,N_6813);
nor U7070 (N_7070,N_6959,N_6945);
and U7071 (N_7071,N_6829,N_6847);
nor U7072 (N_7072,N_6947,N_6934);
xnor U7073 (N_7073,N_6909,N_6891);
xor U7074 (N_7074,N_6993,N_6930);
or U7075 (N_7075,N_6914,N_6886);
nor U7076 (N_7076,N_6811,N_6810);
and U7077 (N_7077,N_6979,N_6951);
nand U7078 (N_7078,N_6968,N_6867);
nand U7079 (N_7079,N_6890,N_6874);
nor U7080 (N_7080,N_6932,N_6804);
nor U7081 (N_7081,N_6989,N_6956);
and U7082 (N_7082,N_6857,N_6958);
or U7083 (N_7083,N_6878,N_6839);
nand U7084 (N_7084,N_6941,N_6809);
nor U7085 (N_7085,N_6869,N_6942);
xor U7086 (N_7086,N_6964,N_6800);
nand U7087 (N_7087,N_6865,N_6901);
or U7088 (N_7088,N_6877,N_6928);
nor U7089 (N_7089,N_6892,N_6906);
nand U7090 (N_7090,N_6929,N_6916);
and U7091 (N_7091,N_6957,N_6926);
xor U7092 (N_7092,N_6963,N_6976);
nand U7093 (N_7093,N_6995,N_6961);
or U7094 (N_7094,N_6801,N_6846);
xor U7095 (N_7095,N_6978,N_6948);
nor U7096 (N_7096,N_6850,N_6815);
nand U7097 (N_7097,N_6832,N_6881);
and U7098 (N_7098,N_6920,N_6849);
and U7099 (N_7099,N_6807,N_6851);
nand U7100 (N_7100,N_6877,N_6908);
or U7101 (N_7101,N_6987,N_6894);
nand U7102 (N_7102,N_6961,N_6945);
and U7103 (N_7103,N_6942,N_6867);
nor U7104 (N_7104,N_6890,N_6968);
nor U7105 (N_7105,N_6938,N_6969);
nor U7106 (N_7106,N_6920,N_6800);
xnor U7107 (N_7107,N_6941,N_6909);
xor U7108 (N_7108,N_6984,N_6905);
or U7109 (N_7109,N_6801,N_6818);
nor U7110 (N_7110,N_6809,N_6929);
nand U7111 (N_7111,N_6869,N_6827);
nor U7112 (N_7112,N_6838,N_6837);
or U7113 (N_7113,N_6815,N_6941);
nand U7114 (N_7114,N_6845,N_6974);
or U7115 (N_7115,N_6939,N_6804);
nor U7116 (N_7116,N_6902,N_6983);
nor U7117 (N_7117,N_6977,N_6956);
nor U7118 (N_7118,N_6959,N_6965);
nand U7119 (N_7119,N_6885,N_6882);
nand U7120 (N_7120,N_6966,N_6848);
and U7121 (N_7121,N_6841,N_6824);
nor U7122 (N_7122,N_6925,N_6949);
nor U7123 (N_7123,N_6810,N_6884);
and U7124 (N_7124,N_6929,N_6911);
or U7125 (N_7125,N_6958,N_6943);
and U7126 (N_7126,N_6910,N_6872);
nor U7127 (N_7127,N_6882,N_6942);
xor U7128 (N_7128,N_6995,N_6927);
nor U7129 (N_7129,N_6884,N_6960);
or U7130 (N_7130,N_6834,N_6963);
xor U7131 (N_7131,N_6863,N_6988);
and U7132 (N_7132,N_6978,N_6928);
nand U7133 (N_7133,N_6979,N_6869);
or U7134 (N_7134,N_6993,N_6955);
nor U7135 (N_7135,N_6813,N_6819);
and U7136 (N_7136,N_6882,N_6892);
xnor U7137 (N_7137,N_6963,N_6970);
and U7138 (N_7138,N_6823,N_6869);
nor U7139 (N_7139,N_6956,N_6875);
xor U7140 (N_7140,N_6961,N_6868);
nor U7141 (N_7141,N_6895,N_6960);
nor U7142 (N_7142,N_6819,N_6895);
xnor U7143 (N_7143,N_6990,N_6822);
and U7144 (N_7144,N_6918,N_6882);
or U7145 (N_7145,N_6827,N_6914);
or U7146 (N_7146,N_6989,N_6882);
xnor U7147 (N_7147,N_6865,N_6937);
or U7148 (N_7148,N_6987,N_6862);
nor U7149 (N_7149,N_6993,N_6847);
and U7150 (N_7150,N_6808,N_6818);
nand U7151 (N_7151,N_6954,N_6951);
nor U7152 (N_7152,N_6905,N_6948);
nor U7153 (N_7153,N_6834,N_6978);
xnor U7154 (N_7154,N_6827,N_6979);
xnor U7155 (N_7155,N_6862,N_6824);
xnor U7156 (N_7156,N_6977,N_6856);
or U7157 (N_7157,N_6835,N_6997);
xnor U7158 (N_7158,N_6806,N_6962);
xor U7159 (N_7159,N_6904,N_6945);
or U7160 (N_7160,N_6963,N_6949);
and U7161 (N_7161,N_6916,N_6832);
nand U7162 (N_7162,N_6968,N_6930);
nor U7163 (N_7163,N_6858,N_6810);
nor U7164 (N_7164,N_6940,N_6936);
and U7165 (N_7165,N_6826,N_6825);
xnor U7166 (N_7166,N_6949,N_6828);
nor U7167 (N_7167,N_6950,N_6851);
nand U7168 (N_7168,N_6933,N_6813);
xnor U7169 (N_7169,N_6989,N_6840);
nand U7170 (N_7170,N_6969,N_6891);
xor U7171 (N_7171,N_6905,N_6938);
xor U7172 (N_7172,N_6958,N_6962);
or U7173 (N_7173,N_6858,N_6842);
and U7174 (N_7174,N_6985,N_6825);
xnor U7175 (N_7175,N_6848,N_6820);
nor U7176 (N_7176,N_6982,N_6908);
nand U7177 (N_7177,N_6848,N_6931);
or U7178 (N_7178,N_6837,N_6921);
nand U7179 (N_7179,N_6961,N_6847);
nor U7180 (N_7180,N_6971,N_6991);
nand U7181 (N_7181,N_6902,N_6810);
and U7182 (N_7182,N_6984,N_6854);
or U7183 (N_7183,N_6998,N_6921);
nor U7184 (N_7184,N_6964,N_6914);
nand U7185 (N_7185,N_6835,N_6990);
nor U7186 (N_7186,N_6975,N_6824);
or U7187 (N_7187,N_6960,N_6829);
xor U7188 (N_7188,N_6887,N_6840);
nor U7189 (N_7189,N_6831,N_6845);
or U7190 (N_7190,N_6948,N_6801);
and U7191 (N_7191,N_6832,N_6808);
nand U7192 (N_7192,N_6961,N_6916);
or U7193 (N_7193,N_6802,N_6969);
or U7194 (N_7194,N_6866,N_6836);
nand U7195 (N_7195,N_6934,N_6989);
nor U7196 (N_7196,N_6949,N_6871);
and U7197 (N_7197,N_6806,N_6905);
nor U7198 (N_7198,N_6940,N_6850);
and U7199 (N_7199,N_6805,N_6856);
or U7200 (N_7200,N_7147,N_7075);
or U7201 (N_7201,N_7035,N_7016);
nand U7202 (N_7202,N_7013,N_7025);
xor U7203 (N_7203,N_7173,N_7125);
and U7204 (N_7204,N_7044,N_7076);
nor U7205 (N_7205,N_7057,N_7133);
and U7206 (N_7206,N_7037,N_7071);
nand U7207 (N_7207,N_7169,N_7077);
nor U7208 (N_7208,N_7083,N_7130);
nor U7209 (N_7209,N_7018,N_7186);
and U7210 (N_7210,N_7054,N_7128);
or U7211 (N_7211,N_7010,N_7043);
or U7212 (N_7212,N_7113,N_7156);
nor U7213 (N_7213,N_7074,N_7140);
nand U7214 (N_7214,N_7039,N_7003);
xnor U7215 (N_7215,N_7005,N_7087);
and U7216 (N_7216,N_7150,N_7162);
or U7217 (N_7217,N_7144,N_7029);
xnor U7218 (N_7218,N_7108,N_7123);
nand U7219 (N_7219,N_7103,N_7134);
nor U7220 (N_7220,N_7093,N_7117);
and U7221 (N_7221,N_7024,N_7098);
and U7222 (N_7222,N_7192,N_7052);
nand U7223 (N_7223,N_7167,N_7051);
nor U7224 (N_7224,N_7102,N_7101);
nand U7225 (N_7225,N_7136,N_7143);
nand U7226 (N_7226,N_7197,N_7160);
nor U7227 (N_7227,N_7020,N_7120);
or U7228 (N_7228,N_7171,N_7106);
xor U7229 (N_7229,N_7181,N_7095);
xnor U7230 (N_7230,N_7146,N_7017);
or U7231 (N_7231,N_7032,N_7121);
nor U7232 (N_7232,N_7065,N_7179);
nand U7233 (N_7233,N_7149,N_7023);
nor U7234 (N_7234,N_7008,N_7158);
and U7235 (N_7235,N_7050,N_7176);
nand U7236 (N_7236,N_7124,N_7002);
xor U7237 (N_7237,N_7006,N_7062);
xnor U7238 (N_7238,N_7004,N_7063);
nor U7239 (N_7239,N_7091,N_7155);
and U7240 (N_7240,N_7011,N_7119);
and U7241 (N_7241,N_7079,N_7153);
nand U7242 (N_7242,N_7060,N_7135);
and U7243 (N_7243,N_7099,N_7154);
xnor U7244 (N_7244,N_7081,N_7049);
nand U7245 (N_7245,N_7126,N_7036);
xnor U7246 (N_7246,N_7022,N_7088);
xor U7247 (N_7247,N_7152,N_7067);
or U7248 (N_7248,N_7082,N_7115);
or U7249 (N_7249,N_7177,N_7166);
or U7250 (N_7250,N_7180,N_7058);
or U7251 (N_7251,N_7027,N_7195);
xnor U7252 (N_7252,N_7161,N_7034);
nor U7253 (N_7253,N_7073,N_7178);
nor U7254 (N_7254,N_7092,N_7048);
nor U7255 (N_7255,N_7163,N_7072);
xnor U7256 (N_7256,N_7165,N_7138);
nand U7257 (N_7257,N_7086,N_7183);
nand U7258 (N_7258,N_7198,N_7012);
xor U7259 (N_7259,N_7042,N_7053);
or U7260 (N_7260,N_7038,N_7129);
xor U7261 (N_7261,N_7137,N_7046);
xor U7262 (N_7262,N_7031,N_7187);
nor U7263 (N_7263,N_7116,N_7141);
nor U7264 (N_7264,N_7069,N_7172);
nand U7265 (N_7265,N_7196,N_7194);
and U7266 (N_7266,N_7122,N_7151);
or U7267 (N_7267,N_7068,N_7139);
xor U7268 (N_7268,N_7030,N_7185);
and U7269 (N_7269,N_7055,N_7109);
nand U7270 (N_7270,N_7026,N_7105);
and U7271 (N_7271,N_7170,N_7001);
and U7272 (N_7272,N_7112,N_7059);
nor U7273 (N_7273,N_7007,N_7056);
nand U7274 (N_7274,N_7182,N_7157);
and U7275 (N_7275,N_7191,N_7033);
nand U7276 (N_7276,N_7175,N_7148);
nor U7277 (N_7277,N_7094,N_7064);
or U7278 (N_7278,N_7145,N_7131);
and U7279 (N_7279,N_7090,N_7100);
xnor U7280 (N_7280,N_7000,N_7045);
xnor U7281 (N_7281,N_7009,N_7199);
and U7282 (N_7282,N_7188,N_7061);
or U7283 (N_7283,N_7028,N_7085);
xor U7284 (N_7284,N_7040,N_7110);
xor U7285 (N_7285,N_7014,N_7159);
nand U7286 (N_7286,N_7066,N_7047);
xor U7287 (N_7287,N_7096,N_7168);
nand U7288 (N_7288,N_7111,N_7193);
and U7289 (N_7289,N_7164,N_7041);
and U7290 (N_7290,N_7118,N_7019);
nor U7291 (N_7291,N_7080,N_7127);
nand U7292 (N_7292,N_7189,N_7097);
or U7293 (N_7293,N_7078,N_7021);
and U7294 (N_7294,N_7132,N_7084);
and U7295 (N_7295,N_7114,N_7184);
nor U7296 (N_7296,N_7174,N_7070);
xor U7297 (N_7297,N_7104,N_7107);
xnor U7298 (N_7298,N_7190,N_7015);
nor U7299 (N_7299,N_7089,N_7142);
xnor U7300 (N_7300,N_7003,N_7155);
nand U7301 (N_7301,N_7151,N_7106);
and U7302 (N_7302,N_7102,N_7097);
nand U7303 (N_7303,N_7169,N_7126);
and U7304 (N_7304,N_7157,N_7064);
and U7305 (N_7305,N_7020,N_7167);
xor U7306 (N_7306,N_7145,N_7005);
or U7307 (N_7307,N_7106,N_7094);
and U7308 (N_7308,N_7151,N_7127);
or U7309 (N_7309,N_7036,N_7089);
xor U7310 (N_7310,N_7186,N_7117);
or U7311 (N_7311,N_7084,N_7173);
and U7312 (N_7312,N_7082,N_7091);
and U7313 (N_7313,N_7025,N_7186);
xnor U7314 (N_7314,N_7188,N_7150);
nand U7315 (N_7315,N_7195,N_7018);
nor U7316 (N_7316,N_7009,N_7042);
nor U7317 (N_7317,N_7180,N_7054);
and U7318 (N_7318,N_7122,N_7033);
nor U7319 (N_7319,N_7044,N_7079);
nand U7320 (N_7320,N_7149,N_7087);
nor U7321 (N_7321,N_7173,N_7015);
and U7322 (N_7322,N_7101,N_7026);
nor U7323 (N_7323,N_7031,N_7160);
nor U7324 (N_7324,N_7106,N_7029);
or U7325 (N_7325,N_7079,N_7144);
xnor U7326 (N_7326,N_7114,N_7142);
nand U7327 (N_7327,N_7052,N_7059);
xnor U7328 (N_7328,N_7161,N_7010);
xnor U7329 (N_7329,N_7012,N_7036);
xnor U7330 (N_7330,N_7127,N_7118);
nand U7331 (N_7331,N_7085,N_7053);
nor U7332 (N_7332,N_7194,N_7061);
or U7333 (N_7333,N_7144,N_7138);
nand U7334 (N_7334,N_7099,N_7096);
or U7335 (N_7335,N_7151,N_7041);
and U7336 (N_7336,N_7032,N_7083);
nor U7337 (N_7337,N_7190,N_7023);
xnor U7338 (N_7338,N_7062,N_7034);
nor U7339 (N_7339,N_7100,N_7084);
nand U7340 (N_7340,N_7109,N_7099);
or U7341 (N_7341,N_7111,N_7165);
nand U7342 (N_7342,N_7134,N_7152);
and U7343 (N_7343,N_7063,N_7166);
xnor U7344 (N_7344,N_7030,N_7192);
nand U7345 (N_7345,N_7110,N_7061);
xor U7346 (N_7346,N_7123,N_7192);
or U7347 (N_7347,N_7134,N_7006);
nor U7348 (N_7348,N_7084,N_7122);
and U7349 (N_7349,N_7117,N_7149);
xnor U7350 (N_7350,N_7115,N_7170);
or U7351 (N_7351,N_7186,N_7000);
nor U7352 (N_7352,N_7151,N_7154);
xnor U7353 (N_7353,N_7093,N_7129);
nand U7354 (N_7354,N_7023,N_7117);
xnor U7355 (N_7355,N_7038,N_7027);
and U7356 (N_7356,N_7095,N_7001);
or U7357 (N_7357,N_7106,N_7018);
or U7358 (N_7358,N_7198,N_7045);
xor U7359 (N_7359,N_7125,N_7009);
nor U7360 (N_7360,N_7024,N_7146);
xnor U7361 (N_7361,N_7062,N_7031);
nor U7362 (N_7362,N_7186,N_7056);
or U7363 (N_7363,N_7109,N_7181);
xor U7364 (N_7364,N_7165,N_7172);
nand U7365 (N_7365,N_7144,N_7140);
or U7366 (N_7366,N_7175,N_7039);
and U7367 (N_7367,N_7133,N_7013);
xnor U7368 (N_7368,N_7059,N_7038);
nand U7369 (N_7369,N_7196,N_7108);
xor U7370 (N_7370,N_7177,N_7130);
nand U7371 (N_7371,N_7190,N_7012);
or U7372 (N_7372,N_7024,N_7165);
xor U7373 (N_7373,N_7104,N_7015);
nor U7374 (N_7374,N_7145,N_7040);
xor U7375 (N_7375,N_7138,N_7143);
nand U7376 (N_7376,N_7075,N_7183);
nand U7377 (N_7377,N_7174,N_7050);
nand U7378 (N_7378,N_7189,N_7164);
xor U7379 (N_7379,N_7172,N_7016);
and U7380 (N_7380,N_7105,N_7103);
or U7381 (N_7381,N_7000,N_7073);
nor U7382 (N_7382,N_7013,N_7018);
nand U7383 (N_7383,N_7025,N_7079);
nand U7384 (N_7384,N_7151,N_7145);
nand U7385 (N_7385,N_7086,N_7070);
nor U7386 (N_7386,N_7194,N_7020);
xnor U7387 (N_7387,N_7189,N_7096);
or U7388 (N_7388,N_7069,N_7092);
nand U7389 (N_7389,N_7019,N_7092);
nor U7390 (N_7390,N_7149,N_7129);
and U7391 (N_7391,N_7054,N_7166);
xor U7392 (N_7392,N_7092,N_7188);
or U7393 (N_7393,N_7126,N_7065);
nand U7394 (N_7394,N_7128,N_7006);
xnor U7395 (N_7395,N_7177,N_7169);
nand U7396 (N_7396,N_7105,N_7092);
or U7397 (N_7397,N_7098,N_7188);
nand U7398 (N_7398,N_7099,N_7133);
xnor U7399 (N_7399,N_7195,N_7151);
or U7400 (N_7400,N_7317,N_7290);
or U7401 (N_7401,N_7228,N_7370);
or U7402 (N_7402,N_7301,N_7365);
nand U7403 (N_7403,N_7265,N_7349);
xnor U7404 (N_7404,N_7216,N_7270);
xor U7405 (N_7405,N_7215,N_7350);
and U7406 (N_7406,N_7204,N_7345);
xor U7407 (N_7407,N_7280,N_7236);
or U7408 (N_7408,N_7274,N_7292);
xnor U7409 (N_7409,N_7287,N_7320);
nor U7410 (N_7410,N_7314,N_7336);
and U7411 (N_7411,N_7285,N_7276);
nor U7412 (N_7412,N_7326,N_7267);
xnor U7413 (N_7413,N_7237,N_7227);
nand U7414 (N_7414,N_7311,N_7299);
and U7415 (N_7415,N_7368,N_7347);
nand U7416 (N_7416,N_7353,N_7315);
xor U7417 (N_7417,N_7322,N_7295);
nor U7418 (N_7418,N_7254,N_7214);
nand U7419 (N_7419,N_7217,N_7277);
nor U7420 (N_7420,N_7358,N_7325);
xnor U7421 (N_7421,N_7221,N_7367);
or U7422 (N_7422,N_7324,N_7235);
nand U7423 (N_7423,N_7281,N_7364);
xnor U7424 (N_7424,N_7357,N_7208);
xor U7425 (N_7425,N_7218,N_7256);
xnor U7426 (N_7426,N_7249,N_7327);
and U7427 (N_7427,N_7313,N_7383);
nor U7428 (N_7428,N_7387,N_7306);
xnor U7429 (N_7429,N_7398,N_7262);
nor U7430 (N_7430,N_7219,N_7210);
nor U7431 (N_7431,N_7385,N_7359);
nand U7432 (N_7432,N_7374,N_7294);
and U7433 (N_7433,N_7381,N_7240);
nand U7434 (N_7434,N_7340,N_7307);
and U7435 (N_7435,N_7332,N_7378);
or U7436 (N_7436,N_7375,N_7321);
nor U7437 (N_7437,N_7334,N_7272);
or U7438 (N_7438,N_7373,N_7273);
nand U7439 (N_7439,N_7372,N_7201);
nor U7440 (N_7440,N_7339,N_7233);
nor U7441 (N_7441,N_7377,N_7229);
nor U7442 (N_7442,N_7261,N_7241);
and U7443 (N_7443,N_7275,N_7260);
nor U7444 (N_7444,N_7268,N_7341);
nor U7445 (N_7445,N_7376,N_7386);
nand U7446 (N_7446,N_7369,N_7333);
xor U7447 (N_7447,N_7259,N_7323);
xnor U7448 (N_7448,N_7346,N_7316);
nand U7449 (N_7449,N_7296,N_7384);
nand U7450 (N_7450,N_7366,N_7232);
or U7451 (N_7451,N_7248,N_7211);
or U7452 (N_7452,N_7223,N_7257);
or U7453 (N_7453,N_7250,N_7224);
nand U7454 (N_7454,N_7293,N_7396);
nor U7455 (N_7455,N_7361,N_7278);
and U7456 (N_7456,N_7303,N_7263);
xnor U7457 (N_7457,N_7284,N_7225);
nand U7458 (N_7458,N_7308,N_7264);
and U7459 (N_7459,N_7338,N_7253);
and U7460 (N_7460,N_7343,N_7243);
nand U7461 (N_7461,N_7244,N_7309);
xnor U7462 (N_7462,N_7328,N_7397);
nand U7463 (N_7463,N_7288,N_7202);
xnor U7464 (N_7464,N_7212,N_7391);
and U7465 (N_7465,N_7271,N_7348);
xnor U7466 (N_7466,N_7394,N_7379);
or U7467 (N_7467,N_7239,N_7231);
and U7468 (N_7468,N_7222,N_7344);
nor U7469 (N_7469,N_7393,N_7286);
or U7470 (N_7470,N_7269,N_7312);
nand U7471 (N_7471,N_7251,N_7291);
nand U7472 (N_7472,N_7354,N_7382);
nand U7473 (N_7473,N_7289,N_7363);
and U7474 (N_7474,N_7362,N_7247);
nand U7475 (N_7475,N_7234,N_7330);
or U7476 (N_7476,N_7389,N_7329);
nor U7477 (N_7477,N_7380,N_7356);
nor U7478 (N_7478,N_7304,N_7230);
nor U7479 (N_7479,N_7342,N_7298);
or U7480 (N_7480,N_7238,N_7206);
nand U7481 (N_7481,N_7213,N_7335);
nor U7482 (N_7482,N_7318,N_7297);
nor U7483 (N_7483,N_7390,N_7371);
or U7484 (N_7484,N_7258,N_7255);
or U7485 (N_7485,N_7302,N_7300);
nand U7486 (N_7486,N_7392,N_7266);
nor U7487 (N_7487,N_7319,N_7279);
or U7488 (N_7488,N_7282,N_7246);
and U7489 (N_7489,N_7200,N_7220);
or U7490 (N_7490,N_7209,N_7360);
nand U7491 (N_7491,N_7245,N_7283);
and U7492 (N_7492,N_7226,N_7352);
nand U7493 (N_7493,N_7252,N_7355);
xor U7494 (N_7494,N_7395,N_7351);
nor U7495 (N_7495,N_7331,N_7399);
and U7496 (N_7496,N_7242,N_7388);
nand U7497 (N_7497,N_7203,N_7310);
xnor U7498 (N_7498,N_7305,N_7337);
and U7499 (N_7499,N_7207,N_7205);
nand U7500 (N_7500,N_7316,N_7387);
and U7501 (N_7501,N_7311,N_7284);
or U7502 (N_7502,N_7237,N_7364);
nor U7503 (N_7503,N_7204,N_7358);
and U7504 (N_7504,N_7325,N_7305);
or U7505 (N_7505,N_7346,N_7303);
or U7506 (N_7506,N_7394,N_7325);
nand U7507 (N_7507,N_7360,N_7366);
or U7508 (N_7508,N_7267,N_7235);
nor U7509 (N_7509,N_7207,N_7267);
or U7510 (N_7510,N_7225,N_7282);
and U7511 (N_7511,N_7221,N_7378);
xor U7512 (N_7512,N_7357,N_7268);
nor U7513 (N_7513,N_7299,N_7266);
or U7514 (N_7514,N_7340,N_7326);
and U7515 (N_7515,N_7352,N_7379);
and U7516 (N_7516,N_7241,N_7288);
nand U7517 (N_7517,N_7280,N_7242);
and U7518 (N_7518,N_7351,N_7334);
and U7519 (N_7519,N_7355,N_7278);
or U7520 (N_7520,N_7311,N_7347);
nor U7521 (N_7521,N_7258,N_7289);
and U7522 (N_7522,N_7356,N_7371);
or U7523 (N_7523,N_7343,N_7389);
nand U7524 (N_7524,N_7391,N_7225);
nor U7525 (N_7525,N_7247,N_7296);
or U7526 (N_7526,N_7367,N_7218);
xor U7527 (N_7527,N_7351,N_7331);
xnor U7528 (N_7528,N_7269,N_7256);
xnor U7529 (N_7529,N_7318,N_7219);
xor U7530 (N_7530,N_7240,N_7331);
and U7531 (N_7531,N_7264,N_7276);
or U7532 (N_7532,N_7381,N_7348);
and U7533 (N_7533,N_7333,N_7277);
nor U7534 (N_7534,N_7390,N_7381);
and U7535 (N_7535,N_7375,N_7280);
nor U7536 (N_7536,N_7228,N_7322);
or U7537 (N_7537,N_7221,N_7354);
nor U7538 (N_7538,N_7214,N_7358);
xnor U7539 (N_7539,N_7210,N_7201);
or U7540 (N_7540,N_7204,N_7201);
xnor U7541 (N_7541,N_7339,N_7390);
and U7542 (N_7542,N_7264,N_7317);
nor U7543 (N_7543,N_7240,N_7362);
nand U7544 (N_7544,N_7391,N_7368);
and U7545 (N_7545,N_7225,N_7311);
nor U7546 (N_7546,N_7216,N_7306);
and U7547 (N_7547,N_7342,N_7336);
nand U7548 (N_7548,N_7265,N_7269);
or U7549 (N_7549,N_7209,N_7254);
xnor U7550 (N_7550,N_7313,N_7252);
or U7551 (N_7551,N_7253,N_7220);
and U7552 (N_7552,N_7327,N_7373);
xor U7553 (N_7553,N_7384,N_7388);
and U7554 (N_7554,N_7216,N_7390);
or U7555 (N_7555,N_7212,N_7392);
nor U7556 (N_7556,N_7251,N_7329);
nand U7557 (N_7557,N_7234,N_7297);
nor U7558 (N_7558,N_7359,N_7240);
and U7559 (N_7559,N_7397,N_7281);
xnor U7560 (N_7560,N_7362,N_7344);
nand U7561 (N_7561,N_7295,N_7225);
or U7562 (N_7562,N_7326,N_7296);
and U7563 (N_7563,N_7272,N_7370);
nand U7564 (N_7564,N_7287,N_7341);
nand U7565 (N_7565,N_7387,N_7204);
and U7566 (N_7566,N_7353,N_7268);
nor U7567 (N_7567,N_7201,N_7290);
nor U7568 (N_7568,N_7226,N_7332);
nor U7569 (N_7569,N_7366,N_7379);
nor U7570 (N_7570,N_7380,N_7287);
nand U7571 (N_7571,N_7310,N_7335);
nor U7572 (N_7572,N_7397,N_7353);
nor U7573 (N_7573,N_7377,N_7372);
nand U7574 (N_7574,N_7259,N_7344);
xor U7575 (N_7575,N_7227,N_7205);
nand U7576 (N_7576,N_7230,N_7205);
xor U7577 (N_7577,N_7387,N_7324);
nor U7578 (N_7578,N_7313,N_7254);
nor U7579 (N_7579,N_7341,N_7326);
xnor U7580 (N_7580,N_7388,N_7320);
and U7581 (N_7581,N_7222,N_7328);
nor U7582 (N_7582,N_7323,N_7298);
nand U7583 (N_7583,N_7256,N_7362);
nand U7584 (N_7584,N_7224,N_7206);
nor U7585 (N_7585,N_7328,N_7213);
and U7586 (N_7586,N_7272,N_7244);
nand U7587 (N_7587,N_7280,N_7249);
nand U7588 (N_7588,N_7360,N_7283);
and U7589 (N_7589,N_7325,N_7329);
nor U7590 (N_7590,N_7381,N_7323);
and U7591 (N_7591,N_7372,N_7279);
nand U7592 (N_7592,N_7242,N_7337);
and U7593 (N_7593,N_7390,N_7277);
or U7594 (N_7594,N_7237,N_7200);
or U7595 (N_7595,N_7223,N_7387);
xor U7596 (N_7596,N_7316,N_7376);
nor U7597 (N_7597,N_7296,N_7379);
or U7598 (N_7598,N_7349,N_7342);
or U7599 (N_7599,N_7276,N_7302);
nand U7600 (N_7600,N_7428,N_7592);
nor U7601 (N_7601,N_7581,N_7552);
or U7602 (N_7602,N_7598,N_7591);
and U7603 (N_7603,N_7473,N_7437);
xnor U7604 (N_7604,N_7596,N_7541);
nor U7605 (N_7605,N_7432,N_7443);
nor U7606 (N_7606,N_7416,N_7410);
and U7607 (N_7607,N_7498,N_7565);
or U7608 (N_7608,N_7535,N_7524);
nor U7609 (N_7609,N_7457,N_7433);
or U7610 (N_7610,N_7442,N_7465);
xnor U7611 (N_7611,N_7403,N_7463);
nor U7612 (N_7612,N_7427,N_7475);
xor U7613 (N_7613,N_7519,N_7454);
xor U7614 (N_7614,N_7587,N_7435);
and U7615 (N_7615,N_7446,N_7597);
or U7616 (N_7616,N_7499,N_7488);
xnor U7617 (N_7617,N_7570,N_7513);
or U7618 (N_7618,N_7599,N_7583);
nor U7619 (N_7619,N_7422,N_7474);
or U7620 (N_7620,N_7400,N_7530);
or U7621 (N_7621,N_7531,N_7559);
nor U7622 (N_7622,N_7436,N_7471);
nor U7623 (N_7623,N_7525,N_7464);
nand U7624 (N_7624,N_7506,N_7508);
nor U7625 (N_7625,N_7555,N_7423);
nor U7626 (N_7626,N_7569,N_7568);
and U7627 (N_7627,N_7572,N_7549);
or U7628 (N_7628,N_7538,N_7448);
nand U7629 (N_7629,N_7571,N_7495);
or U7630 (N_7630,N_7574,N_7479);
and U7631 (N_7631,N_7487,N_7523);
xor U7632 (N_7632,N_7467,N_7551);
or U7633 (N_7633,N_7539,N_7540);
nor U7634 (N_7634,N_7589,N_7418);
and U7635 (N_7635,N_7485,N_7480);
or U7636 (N_7636,N_7470,N_7478);
or U7637 (N_7637,N_7514,N_7411);
nand U7638 (N_7638,N_7586,N_7483);
nor U7639 (N_7639,N_7404,N_7438);
nand U7640 (N_7640,N_7577,N_7505);
and U7641 (N_7641,N_7558,N_7567);
xnor U7642 (N_7642,N_7526,N_7430);
or U7643 (N_7643,N_7460,N_7462);
nand U7644 (N_7644,N_7492,N_7500);
nor U7645 (N_7645,N_7595,N_7566);
xor U7646 (N_7646,N_7494,N_7439);
and U7647 (N_7647,N_7580,N_7413);
xnor U7648 (N_7648,N_7431,N_7578);
xnor U7649 (N_7649,N_7515,N_7518);
nand U7650 (N_7650,N_7489,N_7554);
xnor U7651 (N_7651,N_7590,N_7501);
xor U7652 (N_7652,N_7409,N_7517);
xnor U7653 (N_7653,N_7461,N_7405);
nand U7654 (N_7654,N_7502,N_7544);
and U7655 (N_7655,N_7575,N_7579);
xnor U7656 (N_7656,N_7553,N_7455);
nand U7657 (N_7657,N_7545,N_7496);
xnor U7658 (N_7658,N_7532,N_7550);
nand U7659 (N_7659,N_7481,N_7447);
xor U7660 (N_7660,N_7415,N_7419);
nand U7661 (N_7661,N_7516,N_7491);
or U7662 (N_7662,N_7407,N_7588);
and U7663 (N_7663,N_7561,N_7563);
xnor U7664 (N_7664,N_7584,N_7412);
xor U7665 (N_7665,N_7456,N_7420);
nand U7666 (N_7666,N_7414,N_7458);
or U7667 (N_7667,N_7468,N_7445);
and U7668 (N_7668,N_7426,N_7421);
and U7669 (N_7669,N_7406,N_7594);
nor U7670 (N_7670,N_7451,N_7522);
nand U7671 (N_7671,N_7477,N_7476);
nor U7672 (N_7672,N_7512,N_7441);
nor U7673 (N_7673,N_7576,N_7425);
and U7674 (N_7674,N_7520,N_7450);
nand U7675 (N_7675,N_7434,N_7452);
nand U7676 (N_7676,N_7585,N_7529);
or U7677 (N_7677,N_7548,N_7453);
nand U7678 (N_7678,N_7593,N_7507);
nand U7679 (N_7679,N_7503,N_7486);
nor U7680 (N_7680,N_7534,N_7497);
nand U7681 (N_7681,N_7573,N_7493);
xor U7682 (N_7682,N_7582,N_7449);
xnor U7683 (N_7683,N_7429,N_7560);
or U7684 (N_7684,N_7511,N_7444);
xnor U7685 (N_7685,N_7536,N_7417);
nor U7686 (N_7686,N_7402,N_7547);
nor U7687 (N_7687,N_7466,N_7472);
nand U7688 (N_7688,N_7543,N_7459);
nand U7689 (N_7689,N_7527,N_7504);
xnor U7690 (N_7690,N_7546,N_7484);
xor U7691 (N_7691,N_7482,N_7509);
nor U7692 (N_7692,N_7528,N_7557);
nor U7693 (N_7693,N_7521,N_7440);
xor U7694 (N_7694,N_7564,N_7469);
xnor U7695 (N_7695,N_7490,N_7408);
nand U7696 (N_7696,N_7556,N_7533);
xor U7697 (N_7697,N_7562,N_7510);
and U7698 (N_7698,N_7424,N_7542);
xor U7699 (N_7699,N_7537,N_7401);
nand U7700 (N_7700,N_7462,N_7546);
xnor U7701 (N_7701,N_7400,N_7407);
nor U7702 (N_7702,N_7421,N_7509);
xnor U7703 (N_7703,N_7496,N_7585);
nor U7704 (N_7704,N_7404,N_7449);
and U7705 (N_7705,N_7535,N_7561);
and U7706 (N_7706,N_7587,N_7414);
or U7707 (N_7707,N_7446,N_7542);
and U7708 (N_7708,N_7470,N_7408);
nor U7709 (N_7709,N_7560,N_7541);
or U7710 (N_7710,N_7479,N_7417);
xnor U7711 (N_7711,N_7569,N_7488);
nand U7712 (N_7712,N_7504,N_7559);
xnor U7713 (N_7713,N_7544,N_7546);
nor U7714 (N_7714,N_7580,N_7516);
nand U7715 (N_7715,N_7577,N_7467);
or U7716 (N_7716,N_7497,N_7513);
or U7717 (N_7717,N_7421,N_7557);
nor U7718 (N_7718,N_7580,N_7421);
or U7719 (N_7719,N_7537,N_7512);
nand U7720 (N_7720,N_7425,N_7445);
nand U7721 (N_7721,N_7435,N_7406);
xnor U7722 (N_7722,N_7553,N_7546);
or U7723 (N_7723,N_7501,N_7564);
and U7724 (N_7724,N_7566,N_7487);
xor U7725 (N_7725,N_7458,N_7599);
or U7726 (N_7726,N_7484,N_7590);
xor U7727 (N_7727,N_7555,N_7475);
nor U7728 (N_7728,N_7514,N_7423);
nor U7729 (N_7729,N_7486,N_7447);
or U7730 (N_7730,N_7491,N_7460);
nand U7731 (N_7731,N_7478,N_7518);
or U7732 (N_7732,N_7519,N_7530);
nand U7733 (N_7733,N_7570,N_7522);
nor U7734 (N_7734,N_7461,N_7530);
and U7735 (N_7735,N_7534,N_7530);
nor U7736 (N_7736,N_7434,N_7492);
nand U7737 (N_7737,N_7454,N_7404);
or U7738 (N_7738,N_7584,N_7498);
and U7739 (N_7739,N_7528,N_7412);
xnor U7740 (N_7740,N_7504,N_7580);
nand U7741 (N_7741,N_7592,N_7401);
nor U7742 (N_7742,N_7434,N_7442);
and U7743 (N_7743,N_7473,N_7589);
or U7744 (N_7744,N_7454,N_7447);
nor U7745 (N_7745,N_7598,N_7525);
and U7746 (N_7746,N_7401,N_7585);
xor U7747 (N_7747,N_7451,N_7440);
and U7748 (N_7748,N_7525,N_7597);
nand U7749 (N_7749,N_7405,N_7566);
and U7750 (N_7750,N_7561,N_7449);
or U7751 (N_7751,N_7484,N_7462);
or U7752 (N_7752,N_7575,N_7494);
xnor U7753 (N_7753,N_7597,N_7414);
nor U7754 (N_7754,N_7535,N_7581);
nor U7755 (N_7755,N_7466,N_7507);
nor U7756 (N_7756,N_7558,N_7547);
and U7757 (N_7757,N_7426,N_7461);
xnor U7758 (N_7758,N_7426,N_7413);
nor U7759 (N_7759,N_7578,N_7406);
xnor U7760 (N_7760,N_7422,N_7492);
nand U7761 (N_7761,N_7474,N_7540);
and U7762 (N_7762,N_7568,N_7401);
nor U7763 (N_7763,N_7572,N_7551);
or U7764 (N_7764,N_7407,N_7578);
xnor U7765 (N_7765,N_7547,N_7550);
and U7766 (N_7766,N_7557,N_7494);
nor U7767 (N_7767,N_7447,N_7475);
or U7768 (N_7768,N_7416,N_7435);
nor U7769 (N_7769,N_7585,N_7508);
and U7770 (N_7770,N_7466,N_7568);
xnor U7771 (N_7771,N_7574,N_7522);
or U7772 (N_7772,N_7539,N_7430);
nand U7773 (N_7773,N_7594,N_7497);
xnor U7774 (N_7774,N_7465,N_7597);
nor U7775 (N_7775,N_7593,N_7465);
xnor U7776 (N_7776,N_7511,N_7485);
nor U7777 (N_7777,N_7578,N_7489);
xor U7778 (N_7778,N_7479,N_7596);
nand U7779 (N_7779,N_7464,N_7531);
nand U7780 (N_7780,N_7478,N_7461);
nand U7781 (N_7781,N_7514,N_7441);
xnor U7782 (N_7782,N_7464,N_7553);
xnor U7783 (N_7783,N_7555,N_7589);
and U7784 (N_7784,N_7496,N_7587);
xor U7785 (N_7785,N_7444,N_7572);
xor U7786 (N_7786,N_7558,N_7440);
xor U7787 (N_7787,N_7540,N_7459);
nor U7788 (N_7788,N_7425,N_7459);
or U7789 (N_7789,N_7577,N_7527);
nand U7790 (N_7790,N_7495,N_7407);
nand U7791 (N_7791,N_7559,N_7576);
or U7792 (N_7792,N_7498,N_7425);
and U7793 (N_7793,N_7516,N_7444);
nor U7794 (N_7794,N_7442,N_7549);
nor U7795 (N_7795,N_7478,N_7487);
and U7796 (N_7796,N_7516,N_7543);
xnor U7797 (N_7797,N_7518,N_7556);
xor U7798 (N_7798,N_7506,N_7446);
or U7799 (N_7799,N_7586,N_7431);
xnor U7800 (N_7800,N_7689,N_7756);
nor U7801 (N_7801,N_7739,N_7754);
or U7802 (N_7802,N_7637,N_7791);
nor U7803 (N_7803,N_7798,N_7606);
nor U7804 (N_7804,N_7679,N_7686);
xnor U7805 (N_7805,N_7788,N_7603);
nor U7806 (N_7806,N_7675,N_7766);
nor U7807 (N_7807,N_7671,N_7668);
or U7808 (N_7808,N_7629,N_7619);
or U7809 (N_7809,N_7647,N_7748);
and U7810 (N_7810,N_7630,N_7690);
nor U7811 (N_7811,N_7666,N_7734);
and U7812 (N_7812,N_7627,N_7626);
nand U7813 (N_7813,N_7718,N_7698);
and U7814 (N_7814,N_7692,N_7765);
nor U7815 (N_7815,N_7747,N_7681);
xnor U7816 (N_7816,N_7760,N_7741);
nor U7817 (N_7817,N_7772,N_7638);
nor U7818 (N_7818,N_7608,N_7743);
and U7819 (N_7819,N_7759,N_7701);
xor U7820 (N_7820,N_7727,N_7688);
nand U7821 (N_7821,N_7649,N_7613);
and U7822 (N_7822,N_7716,N_7687);
or U7823 (N_7823,N_7790,N_7665);
nor U7824 (N_7824,N_7601,N_7634);
nor U7825 (N_7825,N_7709,N_7669);
xnor U7826 (N_7826,N_7758,N_7632);
and U7827 (N_7827,N_7725,N_7731);
or U7828 (N_7828,N_7616,N_7643);
and U7829 (N_7829,N_7721,N_7642);
or U7830 (N_7830,N_7658,N_7706);
and U7831 (N_7831,N_7635,N_7719);
xnor U7832 (N_7832,N_7787,N_7663);
nand U7833 (N_7833,N_7715,N_7612);
nand U7834 (N_7834,N_7652,N_7636);
and U7835 (N_7835,N_7742,N_7710);
xnor U7836 (N_7836,N_7746,N_7789);
xnor U7837 (N_7837,N_7785,N_7783);
nor U7838 (N_7838,N_7620,N_7653);
xor U7839 (N_7839,N_7685,N_7720);
nand U7840 (N_7840,N_7763,N_7662);
or U7841 (N_7841,N_7661,N_7769);
nand U7842 (N_7842,N_7796,N_7778);
nand U7843 (N_7843,N_7728,N_7757);
nand U7844 (N_7844,N_7729,N_7610);
nor U7845 (N_7845,N_7693,N_7707);
and U7846 (N_7846,N_7604,N_7781);
xor U7847 (N_7847,N_7792,N_7767);
xnor U7848 (N_7848,N_7624,N_7700);
nand U7849 (N_7849,N_7705,N_7695);
xor U7850 (N_7850,N_7622,N_7777);
or U7851 (N_7851,N_7625,N_7646);
nand U7852 (N_7852,N_7618,N_7672);
nand U7853 (N_7853,N_7628,N_7771);
and U7854 (N_7854,N_7793,N_7670);
xnor U7855 (N_7855,N_7645,N_7696);
and U7856 (N_7856,N_7656,N_7752);
or U7857 (N_7857,N_7703,N_7744);
and U7858 (N_7858,N_7684,N_7722);
and U7859 (N_7859,N_7664,N_7699);
xor U7860 (N_7860,N_7673,N_7770);
and U7861 (N_7861,N_7768,N_7786);
nand U7862 (N_7862,N_7654,N_7733);
nor U7863 (N_7863,N_7762,N_7615);
and U7864 (N_7864,N_7680,N_7730);
or U7865 (N_7865,N_7797,N_7683);
and U7866 (N_7866,N_7753,N_7761);
or U7867 (N_7867,N_7650,N_7740);
nor U7868 (N_7868,N_7614,N_7773);
xor U7869 (N_7869,N_7732,N_7776);
xnor U7870 (N_7870,N_7648,N_7697);
and U7871 (N_7871,N_7600,N_7712);
xor U7872 (N_7872,N_7726,N_7711);
nand U7873 (N_7873,N_7644,N_7659);
or U7874 (N_7874,N_7702,N_7736);
and U7875 (N_7875,N_7602,N_7674);
or U7876 (N_7876,N_7691,N_7633);
and U7877 (N_7877,N_7779,N_7640);
nand U7878 (N_7878,N_7751,N_7651);
nor U7879 (N_7879,N_7631,N_7704);
nor U7880 (N_7880,N_7795,N_7782);
xor U7881 (N_7881,N_7641,N_7639);
nor U7882 (N_7882,N_7623,N_7714);
and U7883 (N_7883,N_7667,N_7713);
nor U7884 (N_7884,N_7738,N_7660);
xnor U7885 (N_7885,N_7745,N_7724);
nor U7886 (N_7886,N_7755,N_7737);
or U7887 (N_7887,N_7774,N_7717);
nor U7888 (N_7888,N_7775,N_7621);
xnor U7889 (N_7889,N_7723,N_7607);
and U7890 (N_7890,N_7708,N_7678);
xnor U7891 (N_7891,N_7676,N_7605);
xnor U7892 (N_7892,N_7682,N_7657);
or U7893 (N_7893,N_7764,N_7735);
and U7894 (N_7894,N_7611,N_7794);
nor U7895 (N_7895,N_7694,N_7799);
xnor U7896 (N_7896,N_7609,N_7677);
xnor U7897 (N_7897,N_7749,N_7655);
and U7898 (N_7898,N_7780,N_7784);
nor U7899 (N_7899,N_7617,N_7750);
and U7900 (N_7900,N_7729,N_7787);
nand U7901 (N_7901,N_7613,N_7754);
or U7902 (N_7902,N_7683,N_7736);
or U7903 (N_7903,N_7684,N_7708);
and U7904 (N_7904,N_7649,N_7688);
nor U7905 (N_7905,N_7782,N_7758);
nor U7906 (N_7906,N_7676,N_7678);
or U7907 (N_7907,N_7607,N_7761);
nor U7908 (N_7908,N_7772,N_7661);
and U7909 (N_7909,N_7609,N_7730);
xnor U7910 (N_7910,N_7783,N_7660);
nor U7911 (N_7911,N_7712,N_7739);
nor U7912 (N_7912,N_7747,N_7732);
or U7913 (N_7913,N_7755,N_7601);
xnor U7914 (N_7914,N_7706,N_7742);
nand U7915 (N_7915,N_7667,N_7761);
nor U7916 (N_7916,N_7608,N_7716);
xnor U7917 (N_7917,N_7732,N_7647);
xor U7918 (N_7918,N_7702,N_7771);
and U7919 (N_7919,N_7787,N_7760);
nor U7920 (N_7920,N_7676,N_7789);
or U7921 (N_7921,N_7758,N_7655);
and U7922 (N_7922,N_7746,N_7727);
nor U7923 (N_7923,N_7719,N_7782);
nor U7924 (N_7924,N_7734,N_7669);
and U7925 (N_7925,N_7704,N_7789);
xor U7926 (N_7926,N_7742,N_7727);
and U7927 (N_7927,N_7665,N_7705);
xor U7928 (N_7928,N_7644,N_7628);
or U7929 (N_7929,N_7611,N_7607);
xor U7930 (N_7930,N_7724,N_7708);
xor U7931 (N_7931,N_7630,N_7786);
or U7932 (N_7932,N_7635,N_7704);
and U7933 (N_7933,N_7775,N_7721);
nor U7934 (N_7934,N_7733,N_7618);
and U7935 (N_7935,N_7682,N_7797);
nor U7936 (N_7936,N_7765,N_7794);
xnor U7937 (N_7937,N_7716,N_7674);
xnor U7938 (N_7938,N_7650,N_7711);
nand U7939 (N_7939,N_7743,N_7781);
or U7940 (N_7940,N_7742,N_7760);
xnor U7941 (N_7941,N_7787,N_7659);
xor U7942 (N_7942,N_7628,N_7723);
nand U7943 (N_7943,N_7664,N_7767);
xnor U7944 (N_7944,N_7783,N_7727);
nand U7945 (N_7945,N_7672,N_7609);
and U7946 (N_7946,N_7690,N_7700);
xnor U7947 (N_7947,N_7799,N_7730);
nand U7948 (N_7948,N_7750,N_7687);
nor U7949 (N_7949,N_7612,N_7664);
nor U7950 (N_7950,N_7758,N_7722);
xnor U7951 (N_7951,N_7616,N_7625);
and U7952 (N_7952,N_7797,N_7752);
or U7953 (N_7953,N_7652,N_7606);
nand U7954 (N_7954,N_7658,N_7760);
nand U7955 (N_7955,N_7719,N_7756);
nand U7956 (N_7956,N_7778,N_7703);
or U7957 (N_7957,N_7795,N_7778);
and U7958 (N_7958,N_7639,N_7636);
nand U7959 (N_7959,N_7686,N_7668);
xor U7960 (N_7960,N_7727,N_7710);
xnor U7961 (N_7961,N_7610,N_7759);
or U7962 (N_7962,N_7787,N_7670);
or U7963 (N_7963,N_7698,N_7756);
or U7964 (N_7964,N_7638,N_7682);
or U7965 (N_7965,N_7747,N_7627);
nand U7966 (N_7966,N_7784,N_7709);
or U7967 (N_7967,N_7710,N_7619);
nor U7968 (N_7968,N_7680,N_7770);
nand U7969 (N_7969,N_7653,N_7604);
and U7970 (N_7970,N_7609,N_7693);
or U7971 (N_7971,N_7792,N_7682);
xor U7972 (N_7972,N_7659,N_7641);
nor U7973 (N_7973,N_7732,N_7799);
or U7974 (N_7974,N_7685,N_7631);
and U7975 (N_7975,N_7689,N_7675);
nand U7976 (N_7976,N_7640,N_7794);
nand U7977 (N_7977,N_7795,N_7713);
or U7978 (N_7978,N_7731,N_7616);
nand U7979 (N_7979,N_7744,N_7736);
xor U7980 (N_7980,N_7655,N_7600);
xor U7981 (N_7981,N_7653,N_7768);
nor U7982 (N_7982,N_7651,N_7750);
and U7983 (N_7983,N_7773,N_7675);
or U7984 (N_7984,N_7693,N_7601);
xor U7985 (N_7985,N_7644,N_7759);
and U7986 (N_7986,N_7689,N_7719);
xnor U7987 (N_7987,N_7659,N_7695);
nor U7988 (N_7988,N_7605,N_7664);
and U7989 (N_7989,N_7684,N_7679);
and U7990 (N_7990,N_7786,N_7783);
or U7991 (N_7991,N_7781,N_7633);
nor U7992 (N_7992,N_7608,N_7672);
nand U7993 (N_7993,N_7771,N_7674);
nand U7994 (N_7994,N_7754,N_7690);
nand U7995 (N_7995,N_7654,N_7792);
and U7996 (N_7996,N_7626,N_7616);
nand U7997 (N_7997,N_7762,N_7795);
xor U7998 (N_7998,N_7729,N_7683);
nor U7999 (N_7999,N_7717,N_7639);
or U8000 (N_8000,N_7897,N_7956);
xnor U8001 (N_8001,N_7953,N_7921);
xnor U8002 (N_8002,N_7967,N_7927);
or U8003 (N_8003,N_7876,N_7841);
and U8004 (N_8004,N_7842,N_7835);
or U8005 (N_8005,N_7895,N_7874);
nor U8006 (N_8006,N_7922,N_7930);
nor U8007 (N_8007,N_7866,N_7906);
and U8008 (N_8008,N_7825,N_7857);
or U8009 (N_8009,N_7908,N_7988);
nor U8010 (N_8010,N_7870,N_7802);
and U8011 (N_8011,N_7965,N_7821);
or U8012 (N_8012,N_7845,N_7884);
xnor U8013 (N_8013,N_7947,N_7997);
nor U8014 (N_8014,N_7992,N_7892);
nor U8015 (N_8015,N_7812,N_7971);
and U8016 (N_8016,N_7826,N_7887);
and U8017 (N_8017,N_7915,N_7989);
xnor U8018 (N_8018,N_7970,N_7869);
nand U8019 (N_8019,N_7804,N_7871);
and U8020 (N_8020,N_7873,N_7838);
or U8021 (N_8021,N_7941,N_7924);
and U8022 (N_8022,N_7942,N_7879);
xor U8023 (N_8023,N_7911,N_7963);
or U8024 (N_8024,N_7945,N_7902);
and U8025 (N_8025,N_7834,N_7889);
or U8026 (N_8026,N_7976,N_7803);
xor U8027 (N_8027,N_7916,N_7934);
nor U8028 (N_8028,N_7846,N_7894);
and U8029 (N_8029,N_7805,N_7984);
or U8030 (N_8030,N_7943,N_7909);
xnor U8031 (N_8031,N_7914,N_7961);
nand U8032 (N_8032,N_7928,N_7861);
nor U8033 (N_8033,N_7983,N_7831);
xor U8034 (N_8034,N_7926,N_7837);
or U8035 (N_8035,N_7810,N_7840);
nor U8036 (N_8036,N_7951,N_7912);
nor U8037 (N_8037,N_7907,N_7990);
nand U8038 (N_8038,N_7815,N_7998);
xor U8039 (N_8039,N_7813,N_7852);
xor U8040 (N_8040,N_7981,N_7940);
nand U8041 (N_8041,N_7962,N_7935);
nor U8042 (N_8042,N_7929,N_7939);
nand U8043 (N_8043,N_7944,N_7800);
or U8044 (N_8044,N_7882,N_7985);
and U8045 (N_8045,N_7823,N_7822);
and U8046 (N_8046,N_7888,N_7844);
nor U8047 (N_8047,N_7905,N_7959);
and U8048 (N_8048,N_7807,N_7955);
nor U8049 (N_8049,N_7923,N_7918);
or U8050 (N_8050,N_7860,N_7999);
nor U8051 (N_8051,N_7966,N_7901);
nor U8052 (N_8052,N_7855,N_7913);
or U8053 (N_8053,N_7991,N_7903);
xor U8054 (N_8054,N_7817,N_7858);
nor U8055 (N_8055,N_7853,N_7919);
nand U8056 (N_8056,N_7925,N_7896);
nand U8057 (N_8057,N_7865,N_7931);
nor U8058 (N_8058,N_7859,N_7964);
nor U8059 (N_8059,N_7849,N_7885);
xnor U8060 (N_8060,N_7832,N_7877);
and U8061 (N_8061,N_7973,N_7946);
and U8062 (N_8062,N_7878,N_7890);
or U8063 (N_8063,N_7818,N_7995);
or U8064 (N_8064,N_7972,N_7868);
and U8065 (N_8065,N_7904,N_7886);
xor U8066 (N_8066,N_7979,N_7854);
nand U8067 (N_8067,N_7977,N_7987);
nor U8068 (N_8068,N_7872,N_7862);
nor U8069 (N_8069,N_7856,N_7829);
nand U8070 (N_8070,N_7996,N_7938);
nand U8071 (N_8071,N_7816,N_7899);
nand U8072 (N_8072,N_7883,N_7801);
nand U8073 (N_8073,N_7936,N_7917);
nor U8074 (N_8074,N_7833,N_7828);
xor U8075 (N_8075,N_7948,N_7986);
nor U8076 (N_8076,N_7820,N_7900);
nor U8077 (N_8077,N_7827,N_7824);
nor U8078 (N_8078,N_7937,N_7968);
and U8079 (N_8079,N_7819,N_7809);
nand U8080 (N_8080,N_7814,N_7954);
nand U8081 (N_8081,N_7875,N_7974);
nand U8082 (N_8082,N_7848,N_7958);
xor U8083 (N_8083,N_7994,N_7952);
or U8084 (N_8084,N_7864,N_7949);
or U8085 (N_8085,N_7933,N_7850);
and U8086 (N_8086,N_7843,N_7982);
and U8087 (N_8087,N_7830,N_7808);
or U8088 (N_8088,N_7898,N_7893);
xnor U8089 (N_8089,N_7969,N_7806);
nand U8090 (N_8090,N_7881,N_7920);
nor U8091 (N_8091,N_7847,N_7980);
nand U8092 (N_8092,N_7957,N_7993);
xor U8093 (N_8093,N_7851,N_7863);
nor U8094 (N_8094,N_7880,N_7975);
and U8095 (N_8095,N_7910,N_7950);
nand U8096 (N_8096,N_7960,N_7836);
or U8097 (N_8097,N_7839,N_7891);
and U8098 (N_8098,N_7932,N_7867);
and U8099 (N_8099,N_7811,N_7978);
nand U8100 (N_8100,N_7860,N_7908);
xor U8101 (N_8101,N_7863,N_7905);
xnor U8102 (N_8102,N_7857,N_7971);
xor U8103 (N_8103,N_7901,N_7813);
and U8104 (N_8104,N_7994,N_7937);
and U8105 (N_8105,N_7860,N_7892);
nand U8106 (N_8106,N_7864,N_7883);
nand U8107 (N_8107,N_7880,N_7813);
nor U8108 (N_8108,N_7999,N_7959);
xor U8109 (N_8109,N_7910,N_7938);
or U8110 (N_8110,N_7921,N_7881);
nand U8111 (N_8111,N_7913,N_7922);
and U8112 (N_8112,N_7833,N_7868);
nor U8113 (N_8113,N_7839,N_7821);
nor U8114 (N_8114,N_7883,N_7893);
nor U8115 (N_8115,N_7920,N_7915);
xnor U8116 (N_8116,N_7811,N_7938);
xor U8117 (N_8117,N_7876,N_7836);
or U8118 (N_8118,N_7971,N_7924);
xnor U8119 (N_8119,N_7900,N_7938);
or U8120 (N_8120,N_7969,N_7867);
and U8121 (N_8121,N_7892,N_7972);
and U8122 (N_8122,N_7816,N_7836);
nor U8123 (N_8123,N_7812,N_7843);
xnor U8124 (N_8124,N_7901,N_7982);
xor U8125 (N_8125,N_7899,N_7835);
nor U8126 (N_8126,N_7888,N_7808);
or U8127 (N_8127,N_7909,N_7886);
nor U8128 (N_8128,N_7943,N_7871);
nand U8129 (N_8129,N_7880,N_7887);
nand U8130 (N_8130,N_7889,N_7844);
nor U8131 (N_8131,N_7998,N_7968);
nand U8132 (N_8132,N_7821,N_7977);
or U8133 (N_8133,N_7961,N_7909);
or U8134 (N_8134,N_7831,N_7938);
xor U8135 (N_8135,N_7952,N_7897);
xnor U8136 (N_8136,N_7974,N_7827);
and U8137 (N_8137,N_7940,N_7859);
or U8138 (N_8138,N_7989,N_7818);
or U8139 (N_8139,N_7962,N_7972);
xor U8140 (N_8140,N_7862,N_7913);
nor U8141 (N_8141,N_7810,N_7884);
nand U8142 (N_8142,N_7829,N_7870);
nand U8143 (N_8143,N_7949,N_7811);
xor U8144 (N_8144,N_7812,N_7826);
nand U8145 (N_8145,N_7961,N_7956);
nor U8146 (N_8146,N_7801,N_7815);
xnor U8147 (N_8147,N_7938,N_7987);
nor U8148 (N_8148,N_7940,N_7967);
xor U8149 (N_8149,N_7969,N_7883);
nor U8150 (N_8150,N_7815,N_7908);
or U8151 (N_8151,N_7932,N_7911);
and U8152 (N_8152,N_7802,N_7959);
and U8153 (N_8153,N_7893,N_7930);
nor U8154 (N_8154,N_7973,N_7834);
nand U8155 (N_8155,N_7827,N_7806);
and U8156 (N_8156,N_7948,N_7877);
or U8157 (N_8157,N_7826,N_7913);
xor U8158 (N_8158,N_7910,N_7842);
or U8159 (N_8159,N_7947,N_7939);
and U8160 (N_8160,N_7879,N_7880);
xor U8161 (N_8161,N_7805,N_7960);
xor U8162 (N_8162,N_7925,N_7999);
nand U8163 (N_8163,N_7980,N_7904);
and U8164 (N_8164,N_7978,N_7810);
nor U8165 (N_8165,N_7845,N_7943);
nand U8166 (N_8166,N_7896,N_7857);
or U8167 (N_8167,N_7821,N_7868);
xor U8168 (N_8168,N_7876,N_7981);
and U8169 (N_8169,N_7964,N_7898);
or U8170 (N_8170,N_7933,N_7945);
nand U8171 (N_8171,N_7974,N_7958);
xnor U8172 (N_8172,N_7873,N_7889);
and U8173 (N_8173,N_7828,N_7854);
nand U8174 (N_8174,N_7853,N_7818);
nand U8175 (N_8175,N_7832,N_7860);
xnor U8176 (N_8176,N_7880,N_7804);
nor U8177 (N_8177,N_7893,N_7921);
nand U8178 (N_8178,N_7846,N_7850);
xor U8179 (N_8179,N_7832,N_7833);
nand U8180 (N_8180,N_7818,N_7883);
xnor U8181 (N_8181,N_7933,N_7872);
xor U8182 (N_8182,N_7840,N_7888);
or U8183 (N_8183,N_7899,N_7960);
xor U8184 (N_8184,N_7971,N_7962);
nor U8185 (N_8185,N_7902,N_7839);
xor U8186 (N_8186,N_7978,N_7835);
nand U8187 (N_8187,N_7959,N_7997);
nor U8188 (N_8188,N_7959,N_7817);
or U8189 (N_8189,N_7932,N_7994);
nor U8190 (N_8190,N_7917,N_7902);
nand U8191 (N_8191,N_7978,N_7821);
nand U8192 (N_8192,N_7980,N_7935);
nor U8193 (N_8193,N_7809,N_7811);
and U8194 (N_8194,N_7829,N_7986);
nor U8195 (N_8195,N_7870,N_7941);
nand U8196 (N_8196,N_7936,N_7906);
nor U8197 (N_8197,N_7843,N_7827);
nor U8198 (N_8198,N_7985,N_7892);
or U8199 (N_8199,N_7845,N_7830);
and U8200 (N_8200,N_8056,N_8089);
xor U8201 (N_8201,N_8193,N_8020);
nand U8202 (N_8202,N_8021,N_8081);
nand U8203 (N_8203,N_8151,N_8189);
and U8204 (N_8204,N_8185,N_8179);
nand U8205 (N_8205,N_8054,N_8107);
and U8206 (N_8206,N_8044,N_8190);
and U8207 (N_8207,N_8194,N_8113);
and U8208 (N_8208,N_8159,N_8146);
and U8209 (N_8209,N_8143,N_8086);
nand U8210 (N_8210,N_8162,N_8039);
xor U8211 (N_8211,N_8040,N_8172);
and U8212 (N_8212,N_8095,N_8037);
xor U8213 (N_8213,N_8002,N_8060);
nor U8214 (N_8214,N_8186,N_8170);
or U8215 (N_8215,N_8097,N_8191);
or U8216 (N_8216,N_8177,N_8150);
or U8217 (N_8217,N_8154,N_8041);
nand U8218 (N_8218,N_8199,N_8094);
nor U8219 (N_8219,N_8168,N_8031);
xor U8220 (N_8220,N_8050,N_8069);
xnor U8221 (N_8221,N_8182,N_8018);
nand U8222 (N_8222,N_8001,N_8132);
xnor U8223 (N_8223,N_8167,N_8008);
nor U8224 (N_8224,N_8016,N_8131);
or U8225 (N_8225,N_8005,N_8128);
and U8226 (N_8226,N_8022,N_8165);
and U8227 (N_8227,N_8063,N_8100);
nor U8228 (N_8228,N_8102,N_8080);
nor U8229 (N_8229,N_8048,N_8171);
nor U8230 (N_8230,N_8047,N_8114);
or U8231 (N_8231,N_8026,N_8030);
nand U8232 (N_8232,N_8071,N_8155);
or U8233 (N_8233,N_8135,N_8073);
nor U8234 (N_8234,N_8157,N_8042);
or U8235 (N_8235,N_8079,N_8015);
or U8236 (N_8236,N_8121,N_8043);
nand U8237 (N_8237,N_8108,N_8127);
nand U8238 (N_8238,N_8125,N_8096);
xnor U8239 (N_8239,N_8084,N_8090);
xnor U8240 (N_8240,N_8126,N_8198);
and U8241 (N_8241,N_8023,N_8136);
and U8242 (N_8242,N_8025,N_8130);
and U8243 (N_8243,N_8176,N_8116);
nor U8244 (N_8244,N_8046,N_8109);
or U8245 (N_8245,N_8085,N_8049);
nand U8246 (N_8246,N_8087,N_8051);
nor U8247 (N_8247,N_8187,N_8078);
and U8248 (N_8248,N_8012,N_8158);
nand U8249 (N_8249,N_8068,N_8153);
and U8250 (N_8250,N_8184,N_8076);
or U8251 (N_8251,N_8028,N_8075);
and U8252 (N_8252,N_8148,N_8163);
xor U8253 (N_8253,N_8098,N_8061);
nor U8254 (N_8254,N_8035,N_8007);
nand U8255 (N_8255,N_8059,N_8117);
nand U8256 (N_8256,N_8106,N_8034);
or U8257 (N_8257,N_8093,N_8147);
nand U8258 (N_8258,N_8149,N_8092);
nor U8259 (N_8259,N_8101,N_8142);
or U8260 (N_8260,N_8055,N_8104);
and U8261 (N_8261,N_8072,N_8169);
or U8262 (N_8262,N_8105,N_8160);
and U8263 (N_8263,N_8137,N_8120);
xor U8264 (N_8264,N_8141,N_8118);
xor U8265 (N_8265,N_8009,N_8111);
nand U8266 (N_8266,N_8175,N_8077);
or U8267 (N_8267,N_8122,N_8197);
or U8268 (N_8268,N_8112,N_8161);
nor U8269 (N_8269,N_8134,N_8027);
nand U8270 (N_8270,N_8013,N_8083);
or U8271 (N_8271,N_8010,N_8006);
nand U8272 (N_8272,N_8195,N_8057);
xnor U8273 (N_8273,N_8053,N_8032);
xnor U8274 (N_8274,N_8192,N_8064);
and U8275 (N_8275,N_8033,N_8166);
or U8276 (N_8276,N_8052,N_8183);
nand U8277 (N_8277,N_8088,N_8145);
and U8278 (N_8278,N_8173,N_8099);
nor U8279 (N_8279,N_8066,N_8152);
xor U8280 (N_8280,N_8004,N_8139);
xor U8281 (N_8281,N_8133,N_8038);
nand U8282 (N_8282,N_8011,N_8017);
and U8283 (N_8283,N_8019,N_8058);
or U8284 (N_8284,N_8014,N_8180);
nor U8285 (N_8285,N_8164,N_8036);
and U8286 (N_8286,N_8178,N_8045);
xor U8287 (N_8287,N_8074,N_8174);
and U8288 (N_8288,N_8140,N_8029);
and U8289 (N_8289,N_8181,N_8065);
xnor U8290 (N_8290,N_8067,N_8196);
nand U8291 (N_8291,N_8062,N_8070);
nand U8292 (N_8292,N_8188,N_8082);
and U8293 (N_8293,N_8156,N_8000);
and U8294 (N_8294,N_8123,N_8115);
or U8295 (N_8295,N_8119,N_8144);
nand U8296 (N_8296,N_8003,N_8103);
nand U8297 (N_8297,N_8138,N_8091);
nor U8298 (N_8298,N_8024,N_8110);
xor U8299 (N_8299,N_8129,N_8124);
or U8300 (N_8300,N_8056,N_8050);
xnor U8301 (N_8301,N_8101,N_8077);
nor U8302 (N_8302,N_8125,N_8196);
and U8303 (N_8303,N_8137,N_8016);
and U8304 (N_8304,N_8109,N_8093);
or U8305 (N_8305,N_8132,N_8069);
or U8306 (N_8306,N_8038,N_8193);
nor U8307 (N_8307,N_8194,N_8030);
nand U8308 (N_8308,N_8056,N_8111);
xor U8309 (N_8309,N_8017,N_8152);
and U8310 (N_8310,N_8057,N_8029);
or U8311 (N_8311,N_8026,N_8002);
nor U8312 (N_8312,N_8185,N_8176);
nor U8313 (N_8313,N_8050,N_8017);
and U8314 (N_8314,N_8142,N_8009);
nor U8315 (N_8315,N_8139,N_8061);
and U8316 (N_8316,N_8148,N_8080);
and U8317 (N_8317,N_8173,N_8062);
and U8318 (N_8318,N_8117,N_8022);
xor U8319 (N_8319,N_8097,N_8062);
nor U8320 (N_8320,N_8028,N_8115);
nor U8321 (N_8321,N_8074,N_8064);
xor U8322 (N_8322,N_8122,N_8056);
and U8323 (N_8323,N_8160,N_8195);
and U8324 (N_8324,N_8167,N_8187);
xor U8325 (N_8325,N_8033,N_8055);
nor U8326 (N_8326,N_8059,N_8187);
or U8327 (N_8327,N_8157,N_8041);
nand U8328 (N_8328,N_8016,N_8157);
and U8329 (N_8329,N_8105,N_8076);
nor U8330 (N_8330,N_8031,N_8000);
nor U8331 (N_8331,N_8004,N_8153);
or U8332 (N_8332,N_8058,N_8105);
or U8333 (N_8333,N_8188,N_8134);
nand U8334 (N_8334,N_8034,N_8064);
nand U8335 (N_8335,N_8199,N_8055);
and U8336 (N_8336,N_8057,N_8177);
and U8337 (N_8337,N_8113,N_8019);
and U8338 (N_8338,N_8167,N_8006);
nand U8339 (N_8339,N_8153,N_8121);
or U8340 (N_8340,N_8000,N_8146);
and U8341 (N_8341,N_8105,N_8060);
and U8342 (N_8342,N_8153,N_8198);
xnor U8343 (N_8343,N_8091,N_8128);
or U8344 (N_8344,N_8047,N_8036);
nor U8345 (N_8345,N_8002,N_8059);
or U8346 (N_8346,N_8091,N_8144);
xor U8347 (N_8347,N_8036,N_8003);
nor U8348 (N_8348,N_8190,N_8143);
xor U8349 (N_8349,N_8107,N_8099);
xnor U8350 (N_8350,N_8150,N_8057);
nor U8351 (N_8351,N_8142,N_8083);
or U8352 (N_8352,N_8142,N_8155);
and U8353 (N_8353,N_8060,N_8038);
nand U8354 (N_8354,N_8187,N_8106);
or U8355 (N_8355,N_8104,N_8059);
nand U8356 (N_8356,N_8118,N_8148);
nor U8357 (N_8357,N_8186,N_8104);
or U8358 (N_8358,N_8177,N_8160);
and U8359 (N_8359,N_8010,N_8116);
xor U8360 (N_8360,N_8193,N_8150);
nand U8361 (N_8361,N_8070,N_8034);
or U8362 (N_8362,N_8043,N_8128);
and U8363 (N_8363,N_8111,N_8052);
nor U8364 (N_8364,N_8121,N_8165);
nor U8365 (N_8365,N_8017,N_8142);
nor U8366 (N_8366,N_8167,N_8180);
or U8367 (N_8367,N_8004,N_8109);
or U8368 (N_8368,N_8168,N_8160);
nand U8369 (N_8369,N_8192,N_8039);
and U8370 (N_8370,N_8047,N_8115);
nor U8371 (N_8371,N_8045,N_8181);
nand U8372 (N_8372,N_8105,N_8099);
xnor U8373 (N_8373,N_8010,N_8079);
and U8374 (N_8374,N_8179,N_8041);
or U8375 (N_8375,N_8104,N_8151);
nand U8376 (N_8376,N_8091,N_8092);
xnor U8377 (N_8377,N_8000,N_8078);
nand U8378 (N_8378,N_8067,N_8085);
nand U8379 (N_8379,N_8154,N_8057);
xor U8380 (N_8380,N_8134,N_8164);
nand U8381 (N_8381,N_8015,N_8115);
nand U8382 (N_8382,N_8137,N_8034);
nor U8383 (N_8383,N_8050,N_8139);
and U8384 (N_8384,N_8072,N_8143);
nor U8385 (N_8385,N_8137,N_8004);
and U8386 (N_8386,N_8159,N_8079);
xor U8387 (N_8387,N_8144,N_8056);
or U8388 (N_8388,N_8041,N_8021);
nand U8389 (N_8389,N_8075,N_8080);
and U8390 (N_8390,N_8152,N_8159);
nand U8391 (N_8391,N_8166,N_8091);
nand U8392 (N_8392,N_8050,N_8104);
nand U8393 (N_8393,N_8045,N_8183);
xor U8394 (N_8394,N_8175,N_8040);
and U8395 (N_8395,N_8000,N_8013);
or U8396 (N_8396,N_8165,N_8010);
xnor U8397 (N_8397,N_8178,N_8023);
xor U8398 (N_8398,N_8152,N_8117);
and U8399 (N_8399,N_8158,N_8102);
or U8400 (N_8400,N_8389,N_8278);
xnor U8401 (N_8401,N_8321,N_8260);
and U8402 (N_8402,N_8391,N_8345);
nand U8403 (N_8403,N_8315,N_8398);
nand U8404 (N_8404,N_8336,N_8230);
xor U8405 (N_8405,N_8271,N_8262);
nand U8406 (N_8406,N_8352,N_8340);
and U8407 (N_8407,N_8320,N_8232);
or U8408 (N_8408,N_8395,N_8225);
nand U8409 (N_8409,N_8314,N_8331);
nand U8410 (N_8410,N_8293,N_8229);
and U8411 (N_8411,N_8339,N_8241);
nor U8412 (N_8412,N_8373,N_8233);
xnor U8413 (N_8413,N_8329,N_8354);
or U8414 (N_8414,N_8223,N_8282);
nor U8415 (N_8415,N_8246,N_8256);
and U8416 (N_8416,N_8379,N_8203);
and U8417 (N_8417,N_8372,N_8251);
nand U8418 (N_8418,N_8390,N_8239);
or U8419 (N_8419,N_8328,N_8351);
xnor U8420 (N_8420,N_8384,N_8310);
nor U8421 (N_8421,N_8344,N_8243);
and U8422 (N_8422,N_8356,N_8371);
or U8423 (N_8423,N_8333,N_8220);
xor U8424 (N_8424,N_8376,N_8215);
or U8425 (N_8425,N_8304,N_8349);
nor U8426 (N_8426,N_8252,N_8366);
nor U8427 (N_8427,N_8202,N_8322);
nand U8428 (N_8428,N_8264,N_8298);
xnor U8429 (N_8429,N_8394,N_8270);
nor U8430 (N_8430,N_8267,N_8327);
and U8431 (N_8431,N_8334,N_8347);
nor U8432 (N_8432,N_8295,N_8231);
nor U8433 (N_8433,N_8318,N_8288);
or U8434 (N_8434,N_8272,N_8388);
nor U8435 (N_8435,N_8253,N_8244);
nor U8436 (N_8436,N_8346,N_8248);
and U8437 (N_8437,N_8381,N_8259);
nor U8438 (N_8438,N_8365,N_8257);
or U8439 (N_8439,N_8383,N_8317);
xor U8440 (N_8440,N_8399,N_8330);
xor U8441 (N_8441,N_8361,N_8364);
or U8442 (N_8442,N_8305,N_8222);
nand U8443 (N_8443,N_8221,N_8268);
xnor U8444 (N_8444,N_8374,N_8338);
or U8445 (N_8445,N_8206,N_8357);
or U8446 (N_8446,N_8228,N_8286);
or U8447 (N_8447,N_8387,N_8393);
or U8448 (N_8448,N_8316,N_8217);
or U8449 (N_8449,N_8378,N_8312);
or U8450 (N_8450,N_8324,N_8363);
nand U8451 (N_8451,N_8290,N_8358);
and U8452 (N_8452,N_8367,N_8258);
nand U8453 (N_8453,N_8307,N_8210);
or U8454 (N_8454,N_8309,N_8227);
nor U8455 (N_8455,N_8237,N_8303);
nand U8456 (N_8456,N_8208,N_8294);
nor U8457 (N_8457,N_8200,N_8275);
and U8458 (N_8458,N_8302,N_8283);
and U8459 (N_8459,N_8289,N_8359);
nor U8460 (N_8460,N_8311,N_8204);
xnor U8461 (N_8461,N_8287,N_8226);
xnor U8462 (N_8462,N_8261,N_8235);
or U8463 (N_8463,N_8284,N_8254);
nor U8464 (N_8464,N_8385,N_8301);
nand U8465 (N_8465,N_8273,N_8313);
nand U8466 (N_8466,N_8296,N_8380);
nand U8467 (N_8467,N_8355,N_8396);
nor U8468 (N_8468,N_8280,N_8250);
xnor U8469 (N_8469,N_8285,N_8360);
nand U8470 (N_8470,N_8245,N_8274);
and U8471 (N_8471,N_8375,N_8214);
and U8472 (N_8472,N_8277,N_8319);
nand U8473 (N_8473,N_8218,N_8279);
or U8474 (N_8474,N_8234,N_8350);
xnor U8475 (N_8475,N_8397,N_8269);
nor U8476 (N_8476,N_8297,N_8219);
and U8477 (N_8477,N_8242,N_8323);
nor U8478 (N_8478,N_8209,N_8332);
or U8479 (N_8479,N_8348,N_8201);
and U8480 (N_8480,N_8353,N_8249);
nand U8481 (N_8481,N_8292,N_8335);
nand U8482 (N_8482,N_8276,N_8205);
nand U8483 (N_8483,N_8266,N_8216);
nand U8484 (N_8484,N_8369,N_8240);
xor U8485 (N_8485,N_8337,N_8236);
and U8486 (N_8486,N_8362,N_8212);
nor U8487 (N_8487,N_8207,N_8247);
nor U8488 (N_8488,N_8281,N_8341);
and U8489 (N_8489,N_8291,N_8306);
xor U8490 (N_8490,N_8325,N_8343);
or U8491 (N_8491,N_8299,N_8342);
xor U8492 (N_8492,N_8382,N_8308);
xnor U8493 (N_8493,N_8238,N_8368);
xnor U8494 (N_8494,N_8386,N_8377);
or U8495 (N_8495,N_8263,N_8392);
or U8496 (N_8496,N_8326,N_8224);
and U8497 (N_8497,N_8255,N_8370);
xor U8498 (N_8498,N_8211,N_8265);
and U8499 (N_8499,N_8213,N_8300);
nor U8500 (N_8500,N_8364,N_8396);
nand U8501 (N_8501,N_8391,N_8378);
and U8502 (N_8502,N_8355,N_8237);
nand U8503 (N_8503,N_8270,N_8245);
nand U8504 (N_8504,N_8372,N_8310);
or U8505 (N_8505,N_8230,N_8256);
or U8506 (N_8506,N_8290,N_8264);
nor U8507 (N_8507,N_8336,N_8369);
nor U8508 (N_8508,N_8210,N_8208);
or U8509 (N_8509,N_8289,N_8355);
or U8510 (N_8510,N_8346,N_8245);
nor U8511 (N_8511,N_8302,N_8349);
or U8512 (N_8512,N_8370,N_8304);
or U8513 (N_8513,N_8228,N_8202);
nor U8514 (N_8514,N_8312,N_8209);
nand U8515 (N_8515,N_8305,N_8337);
nand U8516 (N_8516,N_8272,N_8242);
or U8517 (N_8517,N_8243,N_8339);
xor U8518 (N_8518,N_8217,N_8363);
nor U8519 (N_8519,N_8217,N_8294);
xor U8520 (N_8520,N_8251,N_8392);
nand U8521 (N_8521,N_8307,N_8225);
xor U8522 (N_8522,N_8205,N_8330);
xnor U8523 (N_8523,N_8345,N_8283);
xor U8524 (N_8524,N_8328,N_8369);
and U8525 (N_8525,N_8238,N_8272);
nand U8526 (N_8526,N_8374,N_8254);
and U8527 (N_8527,N_8282,N_8344);
xor U8528 (N_8528,N_8332,N_8295);
nor U8529 (N_8529,N_8341,N_8292);
nand U8530 (N_8530,N_8267,N_8308);
nand U8531 (N_8531,N_8326,N_8381);
or U8532 (N_8532,N_8208,N_8284);
xnor U8533 (N_8533,N_8340,N_8249);
nand U8534 (N_8534,N_8272,N_8243);
nand U8535 (N_8535,N_8396,N_8377);
nor U8536 (N_8536,N_8295,N_8321);
nand U8537 (N_8537,N_8356,N_8324);
and U8538 (N_8538,N_8214,N_8246);
xnor U8539 (N_8539,N_8330,N_8216);
xor U8540 (N_8540,N_8310,N_8353);
xnor U8541 (N_8541,N_8232,N_8381);
nand U8542 (N_8542,N_8329,N_8226);
or U8543 (N_8543,N_8236,N_8220);
xor U8544 (N_8544,N_8319,N_8347);
or U8545 (N_8545,N_8261,N_8365);
xnor U8546 (N_8546,N_8360,N_8228);
xor U8547 (N_8547,N_8232,N_8332);
nor U8548 (N_8548,N_8370,N_8371);
and U8549 (N_8549,N_8395,N_8351);
nand U8550 (N_8550,N_8273,N_8281);
nand U8551 (N_8551,N_8327,N_8393);
and U8552 (N_8552,N_8316,N_8227);
xnor U8553 (N_8553,N_8209,N_8204);
nor U8554 (N_8554,N_8308,N_8344);
and U8555 (N_8555,N_8205,N_8306);
or U8556 (N_8556,N_8245,N_8361);
nor U8557 (N_8557,N_8344,N_8229);
nor U8558 (N_8558,N_8238,N_8258);
xor U8559 (N_8559,N_8362,N_8233);
or U8560 (N_8560,N_8350,N_8354);
or U8561 (N_8561,N_8335,N_8358);
nor U8562 (N_8562,N_8296,N_8207);
and U8563 (N_8563,N_8314,N_8350);
xnor U8564 (N_8564,N_8323,N_8386);
nor U8565 (N_8565,N_8278,N_8293);
or U8566 (N_8566,N_8398,N_8236);
and U8567 (N_8567,N_8307,N_8329);
and U8568 (N_8568,N_8312,N_8393);
or U8569 (N_8569,N_8241,N_8273);
nor U8570 (N_8570,N_8311,N_8340);
and U8571 (N_8571,N_8226,N_8318);
or U8572 (N_8572,N_8395,N_8388);
or U8573 (N_8573,N_8365,N_8378);
nand U8574 (N_8574,N_8325,N_8202);
and U8575 (N_8575,N_8390,N_8290);
xor U8576 (N_8576,N_8310,N_8267);
or U8577 (N_8577,N_8387,N_8273);
nand U8578 (N_8578,N_8385,N_8270);
and U8579 (N_8579,N_8311,N_8367);
or U8580 (N_8580,N_8298,N_8216);
nor U8581 (N_8581,N_8200,N_8386);
and U8582 (N_8582,N_8394,N_8235);
or U8583 (N_8583,N_8285,N_8294);
nor U8584 (N_8584,N_8335,N_8295);
or U8585 (N_8585,N_8321,N_8239);
or U8586 (N_8586,N_8231,N_8314);
or U8587 (N_8587,N_8313,N_8390);
and U8588 (N_8588,N_8391,N_8204);
and U8589 (N_8589,N_8374,N_8200);
or U8590 (N_8590,N_8368,N_8325);
nor U8591 (N_8591,N_8213,N_8273);
nand U8592 (N_8592,N_8279,N_8226);
nor U8593 (N_8593,N_8210,N_8386);
and U8594 (N_8594,N_8215,N_8315);
nor U8595 (N_8595,N_8369,N_8278);
nand U8596 (N_8596,N_8287,N_8367);
xnor U8597 (N_8597,N_8208,N_8256);
and U8598 (N_8598,N_8260,N_8349);
xnor U8599 (N_8599,N_8332,N_8208);
nand U8600 (N_8600,N_8476,N_8591);
xnor U8601 (N_8601,N_8452,N_8487);
nand U8602 (N_8602,N_8593,N_8561);
xor U8603 (N_8603,N_8510,N_8535);
xnor U8604 (N_8604,N_8483,N_8433);
or U8605 (N_8605,N_8599,N_8400);
or U8606 (N_8606,N_8477,N_8435);
nor U8607 (N_8607,N_8588,N_8563);
nor U8608 (N_8608,N_8598,N_8580);
nand U8609 (N_8609,N_8542,N_8576);
nor U8610 (N_8610,N_8564,N_8578);
and U8611 (N_8611,N_8557,N_8532);
or U8612 (N_8612,N_8421,N_8437);
nor U8613 (N_8613,N_8402,N_8526);
and U8614 (N_8614,N_8486,N_8566);
nor U8615 (N_8615,N_8468,N_8499);
or U8616 (N_8616,N_8527,N_8597);
nand U8617 (N_8617,N_8469,N_8443);
nand U8618 (N_8618,N_8592,N_8520);
nand U8619 (N_8619,N_8451,N_8497);
or U8620 (N_8620,N_8423,N_8569);
nand U8621 (N_8621,N_8460,N_8506);
and U8622 (N_8622,N_8467,N_8472);
and U8623 (N_8623,N_8466,N_8533);
or U8624 (N_8624,N_8428,N_8485);
nor U8625 (N_8625,N_8560,N_8595);
and U8626 (N_8626,N_8571,N_8447);
nor U8627 (N_8627,N_8517,N_8482);
and U8628 (N_8628,N_8550,N_8463);
xnor U8629 (N_8629,N_8551,N_8543);
nand U8630 (N_8630,N_8409,N_8465);
or U8631 (N_8631,N_8556,N_8496);
nand U8632 (N_8632,N_8410,N_8538);
nand U8633 (N_8633,N_8449,N_8459);
or U8634 (N_8634,N_8500,N_8586);
xnor U8635 (N_8635,N_8453,N_8417);
nor U8636 (N_8636,N_8504,N_8445);
nand U8637 (N_8637,N_8408,N_8440);
or U8638 (N_8638,N_8583,N_8577);
xnor U8639 (N_8639,N_8521,N_8462);
xor U8640 (N_8640,N_8559,N_8479);
nand U8641 (N_8641,N_8587,N_8478);
nor U8642 (N_8642,N_8581,N_8407);
nor U8643 (N_8643,N_8574,N_8488);
nor U8644 (N_8644,N_8411,N_8495);
nor U8645 (N_8645,N_8596,N_8457);
nand U8646 (N_8646,N_8544,N_8420);
nor U8647 (N_8647,N_8531,N_8562);
xnor U8648 (N_8648,N_8515,N_8425);
and U8649 (N_8649,N_8512,N_8590);
and U8650 (N_8650,N_8464,N_8528);
nor U8651 (N_8651,N_8429,N_8511);
nand U8652 (N_8652,N_8492,N_8436);
xor U8653 (N_8653,N_8481,N_8427);
xor U8654 (N_8654,N_8442,N_8455);
or U8655 (N_8655,N_8518,N_8432);
nand U8656 (N_8656,N_8524,N_8575);
xor U8657 (N_8657,N_8415,N_8529);
xor U8658 (N_8658,N_8547,N_8404);
nand U8659 (N_8659,N_8414,N_8490);
and U8660 (N_8660,N_8461,N_8419);
or U8661 (N_8661,N_8505,N_8507);
and U8662 (N_8662,N_8567,N_8545);
nor U8663 (N_8663,N_8554,N_8502);
nor U8664 (N_8664,N_8434,N_8474);
or U8665 (N_8665,N_8491,N_8484);
and U8666 (N_8666,N_8480,N_8458);
nor U8667 (N_8667,N_8475,N_8406);
nand U8668 (N_8668,N_8431,N_8509);
nand U8669 (N_8669,N_8541,N_8446);
nand U8670 (N_8670,N_8585,N_8470);
or U8671 (N_8671,N_8498,N_8413);
xor U8672 (N_8672,N_8536,N_8513);
xor U8673 (N_8673,N_8438,N_8448);
or U8674 (N_8674,N_8534,N_8555);
nand U8675 (N_8675,N_8401,N_8424);
nand U8676 (N_8676,N_8489,N_8405);
and U8677 (N_8677,N_8426,N_8471);
nand U8678 (N_8678,N_8549,N_8539);
nand U8679 (N_8679,N_8589,N_8552);
xor U8680 (N_8680,N_8522,N_8444);
nor U8681 (N_8681,N_8546,N_8558);
xnor U8682 (N_8682,N_8594,N_8441);
nor U8683 (N_8683,N_8422,N_8403);
xor U8684 (N_8684,N_8579,N_8418);
nor U8685 (N_8685,N_8540,N_8503);
and U8686 (N_8686,N_8573,N_8439);
and U8687 (N_8687,N_8508,N_8501);
or U8688 (N_8688,N_8519,N_8582);
or U8689 (N_8689,N_8584,N_8523);
or U8690 (N_8690,N_8568,N_8430);
nor U8691 (N_8691,N_8456,N_8416);
nand U8692 (N_8692,N_8450,N_8565);
nand U8693 (N_8693,N_8454,N_8514);
xnor U8694 (N_8694,N_8412,N_8548);
nor U8695 (N_8695,N_8516,N_8493);
or U8696 (N_8696,N_8473,N_8572);
and U8697 (N_8697,N_8530,N_8553);
and U8698 (N_8698,N_8537,N_8570);
xor U8699 (N_8699,N_8494,N_8525);
xor U8700 (N_8700,N_8477,N_8586);
and U8701 (N_8701,N_8487,N_8565);
nand U8702 (N_8702,N_8475,N_8519);
nand U8703 (N_8703,N_8441,N_8533);
nand U8704 (N_8704,N_8424,N_8494);
nand U8705 (N_8705,N_8550,N_8425);
nor U8706 (N_8706,N_8528,N_8560);
or U8707 (N_8707,N_8584,N_8532);
xnor U8708 (N_8708,N_8517,N_8579);
nand U8709 (N_8709,N_8417,N_8525);
nor U8710 (N_8710,N_8527,N_8584);
and U8711 (N_8711,N_8555,N_8443);
nor U8712 (N_8712,N_8451,N_8486);
and U8713 (N_8713,N_8476,N_8500);
and U8714 (N_8714,N_8564,N_8519);
nand U8715 (N_8715,N_8571,N_8545);
nor U8716 (N_8716,N_8576,N_8547);
xor U8717 (N_8717,N_8595,N_8552);
xnor U8718 (N_8718,N_8539,N_8450);
nor U8719 (N_8719,N_8460,N_8529);
and U8720 (N_8720,N_8532,N_8486);
or U8721 (N_8721,N_8447,N_8465);
nor U8722 (N_8722,N_8529,N_8419);
nor U8723 (N_8723,N_8500,N_8480);
and U8724 (N_8724,N_8513,N_8456);
or U8725 (N_8725,N_8546,N_8532);
and U8726 (N_8726,N_8477,N_8549);
nor U8727 (N_8727,N_8555,N_8581);
xnor U8728 (N_8728,N_8568,N_8425);
or U8729 (N_8729,N_8499,N_8461);
nand U8730 (N_8730,N_8547,N_8416);
or U8731 (N_8731,N_8546,N_8544);
or U8732 (N_8732,N_8562,N_8428);
and U8733 (N_8733,N_8435,N_8572);
or U8734 (N_8734,N_8540,N_8487);
or U8735 (N_8735,N_8417,N_8437);
xnor U8736 (N_8736,N_8445,N_8465);
nand U8737 (N_8737,N_8564,N_8403);
nand U8738 (N_8738,N_8494,N_8540);
and U8739 (N_8739,N_8439,N_8507);
xor U8740 (N_8740,N_8599,N_8476);
nor U8741 (N_8741,N_8449,N_8575);
or U8742 (N_8742,N_8446,N_8578);
nand U8743 (N_8743,N_8580,N_8406);
or U8744 (N_8744,N_8533,N_8569);
nor U8745 (N_8745,N_8546,N_8520);
nor U8746 (N_8746,N_8545,N_8419);
nand U8747 (N_8747,N_8593,N_8427);
and U8748 (N_8748,N_8487,N_8543);
and U8749 (N_8749,N_8513,N_8576);
xor U8750 (N_8750,N_8485,N_8535);
xor U8751 (N_8751,N_8467,N_8474);
and U8752 (N_8752,N_8423,N_8587);
xnor U8753 (N_8753,N_8568,N_8588);
xor U8754 (N_8754,N_8423,N_8482);
or U8755 (N_8755,N_8536,N_8573);
or U8756 (N_8756,N_8551,N_8529);
or U8757 (N_8757,N_8452,N_8468);
nor U8758 (N_8758,N_8535,N_8410);
nor U8759 (N_8759,N_8454,N_8571);
nand U8760 (N_8760,N_8473,N_8477);
nor U8761 (N_8761,N_8443,N_8542);
nand U8762 (N_8762,N_8505,N_8502);
and U8763 (N_8763,N_8562,N_8570);
xor U8764 (N_8764,N_8585,N_8414);
nand U8765 (N_8765,N_8540,N_8410);
nor U8766 (N_8766,N_8540,N_8595);
nand U8767 (N_8767,N_8401,N_8590);
nor U8768 (N_8768,N_8425,N_8421);
and U8769 (N_8769,N_8568,N_8491);
nor U8770 (N_8770,N_8521,N_8592);
nor U8771 (N_8771,N_8405,N_8462);
xor U8772 (N_8772,N_8528,N_8530);
and U8773 (N_8773,N_8402,N_8563);
and U8774 (N_8774,N_8440,N_8497);
and U8775 (N_8775,N_8594,N_8499);
or U8776 (N_8776,N_8595,N_8503);
and U8777 (N_8777,N_8430,N_8401);
or U8778 (N_8778,N_8564,N_8521);
nor U8779 (N_8779,N_8515,N_8546);
nand U8780 (N_8780,N_8425,N_8434);
and U8781 (N_8781,N_8580,N_8420);
xor U8782 (N_8782,N_8448,N_8479);
nor U8783 (N_8783,N_8511,N_8553);
and U8784 (N_8784,N_8446,N_8447);
xnor U8785 (N_8785,N_8485,N_8462);
and U8786 (N_8786,N_8449,N_8406);
xnor U8787 (N_8787,N_8540,N_8425);
or U8788 (N_8788,N_8463,N_8512);
or U8789 (N_8789,N_8570,N_8549);
nor U8790 (N_8790,N_8487,N_8495);
xnor U8791 (N_8791,N_8496,N_8578);
or U8792 (N_8792,N_8597,N_8456);
xnor U8793 (N_8793,N_8548,N_8431);
and U8794 (N_8794,N_8416,N_8534);
or U8795 (N_8795,N_8400,N_8597);
xor U8796 (N_8796,N_8557,N_8558);
or U8797 (N_8797,N_8432,N_8529);
xor U8798 (N_8798,N_8515,N_8568);
nand U8799 (N_8799,N_8549,N_8453);
and U8800 (N_8800,N_8761,N_8728);
xnor U8801 (N_8801,N_8682,N_8645);
nand U8802 (N_8802,N_8743,N_8685);
nand U8803 (N_8803,N_8746,N_8749);
xnor U8804 (N_8804,N_8631,N_8620);
or U8805 (N_8805,N_8748,N_8683);
nand U8806 (N_8806,N_8677,N_8687);
nor U8807 (N_8807,N_8666,N_8633);
nand U8808 (N_8808,N_8635,N_8625);
or U8809 (N_8809,N_8793,N_8655);
or U8810 (N_8810,N_8726,N_8660);
or U8811 (N_8811,N_8626,N_8763);
or U8812 (N_8812,N_8698,N_8667);
xnor U8813 (N_8813,N_8730,N_8676);
nand U8814 (N_8814,N_8795,N_8637);
or U8815 (N_8815,N_8721,N_8799);
xor U8816 (N_8816,N_8711,N_8638);
and U8817 (N_8817,N_8784,N_8605);
nor U8818 (N_8818,N_8782,N_8767);
and U8819 (N_8819,N_8670,N_8719);
nor U8820 (N_8820,N_8790,N_8702);
nand U8821 (N_8821,N_8715,N_8641);
nor U8822 (N_8822,N_8706,N_8756);
or U8823 (N_8823,N_8610,N_8770);
nand U8824 (N_8824,N_8658,N_8663);
and U8825 (N_8825,N_8695,N_8759);
or U8826 (N_8826,N_8603,N_8752);
nor U8827 (N_8827,N_8762,N_8733);
nor U8828 (N_8828,N_8785,N_8742);
xor U8829 (N_8829,N_8704,N_8639);
nor U8830 (N_8830,N_8741,N_8656);
nor U8831 (N_8831,N_8773,N_8652);
xnor U8832 (N_8832,N_8700,N_8640);
nand U8833 (N_8833,N_8707,N_8727);
or U8834 (N_8834,N_8643,N_8750);
nor U8835 (N_8835,N_8751,N_8632);
xnor U8836 (N_8836,N_8613,N_8703);
nor U8837 (N_8837,N_8681,N_8654);
nor U8838 (N_8838,N_8604,N_8771);
and U8839 (N_8839,N_8772,N_8601);
or U8840 (N_8840,N_8732,N_8757);
or U8841 (N_8841,N_8674,N_8648);
xor U8842 (N_8842,N_8754,N_8650);
or U8843 (N_8843,N_8705,N_8708);
and U8844 (N_8844,N_8686,N_8787);
and U8845 (N_8845,N_8636,N_8680);
or U8846 (N_8846,N_8780,N_8775);
nand U8847 (N_8847,N_8789,N_8788);
xor U8848 (N_8848,N_8628,N_8724);
nand U8849 (N_8849,N_8664,N_8768);
and U8850 (N_8850,N_8622,N_8614);
nand U8851 (N_8851,N_8618,N_8689);
nand U8852 (N_8852,N_8747,N_8778);
nor U8853 (N_8853,N_8769,N_8649);
and U8854 (N_8854,N_8671,N_8621);
nand U8855 (N_8855,N_8745,N_8607);
nor U8856 (N_8856,N_8600,N_8616);
xor U8857 (N_8857,N_8647,N_8723);
nand U8858 (N_8858,N_8735,N_8764);
nand U8859 (N_8859,N_8634,N_8714);
nor U8860 (N_8860,N_8672,N_8684);
xnor U8861 (N_8861,N_8692,N_8678);
xor U8862 (N_8862,N_8669,N_8697);
nor U8863 (N_8863,N_8694,N_8675);
nand U8864 (N_8864,N_8783,N_8661);
nor U8865 (N_8865,N_8786,N_8738);
and U8866 (N_8866,N_8796,N_8792);
nor U8867 (N_8867,N_8624,N_8798);
nand U8868 (N_8868,N_8779,N_8797);
nor U8869 (N_8869,N_8615,N_8606);
nor U8870 (N_8870,N_8731,N_8794);
nor U8871 (N_8871,N_8617,N_8611);
and U8872 (N_8872,N_8791,N_8710);
nor U8873 (N_8873,N_8716,N_8665);
and U8874 (N_8874,N_8740,N_8668);
nand U8875 (N_8875,N_8623,N_8651);
nor U8876 (N_8876,N_8696,N_8644);
xnor U8877 (N_8877,N_8602,N_8758);
nand U8878 (N_8878,N_8699,N_8729);
xnor U8879 (N_8879,N_8646,N_8627);
nand U8880 (N_8880,N_8739,N_8720);
nor U8881 (N_8881,N_8713,N_8679);
nand U8882 (N_8882,N_8659,N_8642);
xnor U8883 (N_8883,N_8765,N_8766);
xnor U8884 (N_8884,N_8718,N_8609);
and U8885 (N_8885,N_8736,N_8608);
xnor U8886 (N_8886,N_8760,N_8612);
nand U8887 (N_8887,N_8657,N_8734);
nor U8888 (N_8888,N_8690,N_8722);
or U8889 (N_8889,N_8688,N_8709);
xnor U8890 (N_8890,N_8776,N_8662);
or U8891 (N_8891,N_8725,N_8744);
and U8892 (N_8892,N_8755,N_8630);
nand U8893 (N_8893,N_8774,N_8673);
or U8894 (N_8894,N_8619,N_8693);
nor U8895 (N_8895,N_8777,N_8753);
nand U8896 (N_8896,N_8691,N_8717);
nor U8897 (N_8897,N_8712,N_8653);
or U8898 (N_8898,N_8629,N_8737);
or U8899 (N_8899,N_8701,N_8781);
nand U8900 (N_8900,N_8644,N_8772);
xor U8901 (N_8901,N_8611,N_8660);
nand U8902 (N_8902,N_8721,N_8600);
and U8903 (N_8903,N_8678,N_8706);
nand U8904 (N_8904,N_8724,N_8693);
nand U8905 (N_8905,N_8675,N_8772);
and U8906 (N_8906,N_8642,N_8614);
nand U8907 (N_8907,N_8637,N_8702);
xnor U8908 (N_8908,N_8653,N_8742);
or U8909 (N_8909,N_8674,N_8732);
and U8910 (N_8910,N_8634,N_8739);
or U8911 (N_8911,N_8678,N_8752);
or U8912 (N_8912,N_8623,N_8703);
nor U8913 (N_8913,N_8654,N_8723);
and U8914 (N_8914,N_8762,N_8697);
or U8915 (N_8915,N_8647,N_8750);
nor U8916 (N_8916,N_8620,N_8714);
and U8917 (N_8917,N_8700,N_8605);
nor U8918 (N_8918,N_8605,N_8747);
and U8919 (N_8919,N_8705,N_8787);
or U8920 (N_8920,N_8689,N_8690);
nand U8921 (N_8921,N_8739,N_8662);
nand U8922 (N_8922,N_8613,N_8676);
nor U8923 (N_8923,N_8629,N_8709);
nand U8924 (N_8924,N_8761,N_8781);
and U8925 (N_8925,N_8651,N_8693);
xor U8926 (N_8926,N_8731,N_8789);
and U8927 (N_8927,N_8634,N_8732);
or U8928 (N_8928,N_8799,N_8647);
or U8929 (N_8929,N_8764,N_8603);
and U8930 (N_8930,N_8712,N_8640);
nor U8931 (N_8931,N_8779,N_8766);
and U8932 (N_8932,N_8693,N_8744);
and U8933 (N_8933,N_8789,N_8726);
nor U8934 (N_8934,N_8794,N_8606);
or U8935 (N_8935,N_8747,N_8612);
and U8936 (N_8936,N_8619,N_8695);
and U8937 (N_8937,N_8783,N_8789);
and U8938 (N_8938,N_8712,N_8756);
and U8939 (N_8939,N_8742,N_8694);
nand U8940 (N_8940,N_8628,N_8614);
nor U8941 (N_8941,N_8721,N_8657);
or U8942 (N_8942,N_8637,N_8777);
nand U8943 (N_8943,N_8634,N_8773);
xor U8944 (N_8944,N_8711,N_8608);
or U8945 (N_8945,N_8628,N_8795);
xnor U8946 (N_8946,N_8761,N_8681);
and U8947 (N_8947,N_8776,N_8724);
xor U8948 (N_8948,N_8761,N_8670);
and U8949 (N_8949,N_8758,N_8683);
and U8950 (N_8950,N_8617,N_8637);
or U8951 (N_8951,N_8617,N_8710);
nand U8952 (N_8952,N_8616,N_8694);
and U8953 (N_8953,N_8632,N_8701);
nor U8954 (N_8954,N_8718,N_8679);
and U8955 (N_8955,N_8679,N_8750);
xnor U8956 (N_8956,N_8707,N_8616);
or U8957 (N_8957,N_8618,N_8721);
nor U8958 (N_8958,N_8673,N_8633);
nor U8959 (N_8959,N_8699,N_8708);
and U8960 (N_8960,N_8616,N_8793);
xor U8961 (N_8961,N_8748,N_8618);
and U8962 (N_8962,N_8705,N_8788);
or U8963 (N_8963,N_8654,N_8682);
nor U8964 (N_8964,N_8633,N_8782);
nor U8965 (N_8965,N_8771,N_8672);
and U8966 (N_8966,N_8721,N_8793);
xnor U8967 (N_8967,N_8681,N_8694);
nand U8968 (N_8968,N_8615,N_8656);
and U8969 (N_8969,N_8770,N_8731);
nand U8970 (N_8970,N_8647,N_8664);
nor U8971 (N_8971,N_8658,N_8702);
nor U8972 (N_8972,N_8648,N_8770);
xor U8973 (N_8973,N_8724,N_8631);
nor U8974 (N_8974,N_8620,N_8603);
nor U8975 (N_8975,N_8761,N_8764);
or U8976 (N_8976,N_8732,N_8755);
or U8977 (N_8977,N_8696,N_8618);
or U8978 (N_8978,N_8739,N_8729);
nor U8979 (N_8979,N_8776,N_8686);
xor U8980 (N_8980,N_8690,N_8625);
xor U8981 (N_8981,N_8767,N_8702);
xnor U8982 (N_8982,N_8774,N_8634);
nand U8983 (N_8983,N_8716,N_8655);
or U8984 (N_8984,N_8695,N_8763);
nor U8985 (N_8985,N_8690,N_8644);
nand U8986 (N_8986,N_8777,N_8664);
nor U8987 (N_8987,N_8661,N_8780);
xnor U8988 (N_8988,N_8648,N_8633);
or U8989 (N_8989,N_8725,N_8674);
or U8990 (N_8990,N_8630,N_8691);
nand U8991 (N_8991,N_8654,N_8649);
or U8992 (N_8992,N_8691,N_8690);
nor U8993 (N_8993,N_8671,N_8715);
nor U8994 (N_8994,N_8761,N_8672);
or U8995 (N_8995,N_8736,N_8745);
and U8996 (N_8996,N_8707,N_8673);
xor U8997 (N_8997,N_8778,N_8739);
nor U8998 (N_8998,N_8761,N_8705);
nand U8999 (N_8999,N_8787,N_8646);
or U9000 (N_9000,N_8814,N_8823);
and U9001 (N_9001,N_8898,N_8981);
nand U9002 (N_9002,N_8888,N_8881);
or U9003 (N_9003,N_8963,N_8987);
nor U9004 (N_9004,N_8970,N_8844);
nand U9005 (N_9005,N_8942,N_8926);
and U9006 (N_9006,N_8890,N_8800);
or U9007 (N_9007,N_8977,N_8990);
and U9008 (N_9008,N_8849,N_8955);
nor U9009 (N_9009,N_8916,N_8870);
and U9010 (N_9010,N_8818,N_8828);
and U9011 (N_9011,N_8880,N_8991);
and U9012 (N_9012,N_8997,N_8982);
xor U9013 (N_9013,N_8819,N_8868);
xor U9014 (N_9014,N_8901,N_8899);
or U9015 (N_9015,N_8809,N_8873);
nor U9016 (N_9016,N_8937,N_8989);
nor U9017 (N_9017,N_8863,N_8968);
nor U9018 (N_9018,N_8872,N_8962);
nor U9019 (N_9019,N_8978,N_8948);
nor U9020 (N_9020,N_8815,N_8920);
and U9021 (N_9021,N_8998,N_8886);
or U9022 (N_9022,N_8864,N_8851);
or U9023 (N_9023,N_8858,N_8904);
xor U9024 (N_9024,N_8971,N_8893);
or U9025 (N_9025,N_8935,N_8914);
or U9026 (N_9026,N_8999,N_8902);
or U9027 (N_9027,N_8887,N_8835);
nand U9028 (N_9028,N_8950,N_8833);
nand U9029 (N_9029,N_8891,N_8974);
xor U9030 (N_9030,N_8976,N_8923);
nand U9031 (N_9031,N_8985,N_8945);
nor U9032 (N_9032,N_8909,N_8846);
xor U9033 (N_9033,N_8918,N_8944);
nor U9034 (N_9034,N_8878,N_8958);
and U9035 (N_9035,N_8939,N_8894);
nand U9036 (N_9036,N_8861,N_8842);
and U9037 (N_9037,N_8884,N_8946);
xor U9038 (N_9038,N_8951,N_8984);
xor U9039 (N_9039,N_8869,N_8836);
or U9040 (N_9040,N_8889,N_8829);
nor U9041 (N_9041,N_8988,N_8841);
nand U9042 (N_9042,N_8956,N_8949);
or U9043 (N_9043,N_8822,N_8912);
nor U9044 (N_9044,N_8930,N_8847);
and U9045 (N_9045,N_8850,N_8871);
nand U9046 (N_9046,N_8805,N_8996);
xnor U9047 (N_9047,N_8854,N_8804);
and U9048 (N_9048,N_8906,N_8897);
nor U9049 (N_9049,N_8883,N_8853);
nor U9050 (N_9050,N_8866,N_8860);
nor U9051 (N_9051,N_8924,N_8919);
and U9052 (N_9052,N_8964,N_8816);
and U9053 (N_9053,N_8807,N_8936);
and U9054 (N_9054,N_8925,N_8839);
or U9055 (N_9055,N_8986,N_8938);
and U9056 (N_9056,N_8859,N_8845);
nand U9057 (N_9057,N_8905,N_8972);
or U9058 (N_9058,N_8855,N_8813);
or U9059 (N_9059,N_8862,N_8910);
or U9060 (N_9060,N_8913,N_8911);
or U9061 (N_9061,N_8952,N_8852);
nand U9062 (N_9062,N_8874,N_8900);
nor U9063 (N_9063,N_8895,N_8801);
or U9064 (N_9064,N_8826,N_8803);
and U9065 (N_9065,N_8940,N_8980);
or U9066 (N_9066,N_8885,N_8933);
nand U9067 (N_9067,N_8879,N_8843);
or U9068 (N_9068,N_8832,N_8865);
nand U9069 (N_9069,N_8825,N_8932);
nor U9070 (N_9070,N_8907,N_8966);
nor U9071 (N_9071,N_8867,N_8953);
nand U9072 (N_9072,N_8928,N_8983);
nor U9073 (N_9073,N_8973,N_8959);
xor U9074 (N_9074,N_8967,N_8875);
nor U9075 (N_9075,N_8838,N_8993);
nand U9076 (N_9076,N_8929,N_8957);
xnor U9077 (N_9077,N_8975,N_8947);
nand U9078 (N_9078,N_8915,N_8848);
nor U9079 (N_9079,N_8943,N_8820);
or U9080 (N_9080,N_8837,N_8812);
nand U9081 (N_9081,N_8994,N_8931);
nand U9082 (N_9082,N_8830,N_8960);
nor U9083 (N_9083,N_8965,N_8969);
or U9084 (N_9084,N_8877,N_8831);
nor U9085 (N_9085,N_8810,N_8892);
and U9086 (N_9086,N_8954,N_8995);
nor U9087 (N_9087,N_8827,N_8857);
or U9088 (N_9088,N_8922,N_8896);
nand U9089 (N_9089,N_8808,N_8811);
xnor U9090 (N_9090,N_8806,N_8856);
or U9091 (N_9091,N_8834,N_8934);
and U9092 (N_9092,N_8979,N_8908);
nor U9093 (N_9093,N_8876,N_8802);
nand U9094 (N_9094,N_8961,N_8927);
nand U9095 (N_9095,N_8840,N_8903);
and U9096 (N_9096,N_8824,N_8941);
or U9097 (N_9097,N_8821,N_8882);
xor U9098 (N_9098,N_8921,N_8917);
and U9099 (N_9099,N_8992,N_8817);
xnor U9100 (N_9100,N_8807,N_8868);
nand U9101 (N_9101,N_8831,N_8930);
nand U9102 (N_9102,N_8862,N_8958);
xor U9103 (N_9103,N_8939,N_8919);
nor U9104 (N_9104,N_8880,N_8954);
nor U9105 (N_9105,N_8915,N_8893);
xor U9106 (N_9106,N_8864,N_8926);
xor U9107 (N_9107,N_8897,N_8934);
nand U9108 (N_9108,N_8823,N_8917);
xor U9109 (N_9109,N_8890,N_8980);
nor U9110 (N_9110,N_8858,N_8859);
or U9111 (N_9111,N_8856,N_8910);
xnor U9112 (N_9112,N_8871,N_8909);
nand U9113 (N_9113,N_8842,N_8992);
and U9114 (N_9114,N_8983,N_8860);
nand U9115 (N_9115,N_8852,N_8956);
nor U9116 (N_9116,N_8878,N_8804);
nand U9117 (N_9117,N_8903,N_8832);
nand U9118 (N_9118,N_8949,N_8808);
nor U9119 (N_9119,N_8994,N_8941);
nor U9120 (N_9120,N_8962,N_8828);
nand U9121 (N_9121,N_8811,N_8959);
xor U9122 (N_9122,N_8962,N_8944);
nor U9123 (N_9123,N_8863,N_8896);
nor U9124 (N_9124,N_8947,N_8914);
nand U9125 (N_9125,N_8972,N_8934);
nand U9126 (N_9126,N_8910,N_8903);
and U9127 (N_9127,N_8935,N_8973);
or U9128 (N_9128,N_8829,N_8918);
and U9129 (N_9129,N_8889,N_8819);
and U9130 (N_9130,N_8814,N_8817);
and U9131 (N_9131,N_8974,N_8863);
nor U9132 (N_9132,N_8886,N_8823);
nand U9133 (N_9133,N_8921,N_8816);
or U9134 (N_9134,N_8888,N_8914);
xor U9135 (N_9135,N_8827,N_8878);
nor U9136 (N_9136,N_8841,N_8999);
or U9137 (N_9137,N_8922,N_8937);
nor U9138 (N_9138,N_8875,N_8887);
nor U9139 (N_9139,N_8816,N_8918);
nor U9140 (N_9140,N_8932,N_8891);
nand U9141 (N_9141,N_8811,N_8826);
nor U9142 (N_9142,N_8886,N_8997);
or U9143 (N_9143,N_8811,N_8810);
and U9144 (N_9144,N_8935,N_8974);
and U9145 (N_9145,N_8860,N_8870);
nand U9146 (N_9146,N_8906,N_8973);
nor U9147 (N_9147,N_8910,N_8966);
xor U9148 (N_9148,N_8916,N_8803);
nor U9149 (N_9149,N_8831,N_8946);
or U9150 (N_9150,N_8856,N_8817);
and U9151 (N_9151,N_8957,N_8944);
nand U9152 (N_9152,N_8945,N_8857);
nor U9153 (N_9153,N_8826,N_8819);
xor U9154 (N_9154,N_8831,N_8830);
nor U9155 (N_9155,N_8959,N_8837);
nand U9156 (N_9156,N_8920,N_8888);
nand U9157 (N_9157,N_8993,N_8881);
xor U9158 (N_9158,N_8873,N_8886);
and U9159 (N_9159,N_8882,N_8851);
and U9160 (N_9160,N_8802,N_8928);
xnor U9161 (N_9161,N_8903,N_8827);
and U9162 (N_9162,N_8957,N_8844);
xnor U9163 (N_9163,N_8974,N_8909);
nor U9164 (N_9164,N_8925,N_8927);
xnor U9165 (N_9165,N_8900,N_8956);
or U9166 (N_9166,N_8931,N_8961);
nor U9167 (N_9167,N_8872,N_8806);
xnor U9168 (N_9168,N_8946,N_8812);
nand U9169 (N_9169,N_8956,N_8961);
xnor U9170 (N_9170,N_8876,N_8974);
or U9171 (N_9171,N_8936,N_8990);
or U9172 (N_9172,N_8901,N_8964);
or U9173 (N_9173,N_8881,N_8875);
and U9174 (N_9174,N_8839,N_8985);
and U9175 (N_9175,N_8925,N_8867);
xor U9176 (N_9176,N_8900,N_8870);
or U9177 (N_9177,N_8889,N_8924);
nor U9178 (N_9178,N_8874,N_8836);
and U9179 (N_9179,N_8868,N_8829);
xnor U9180 (N_9180,N_8844,N_8833);
or U9181 (N_9181,N_8883,N_8932);
nand U9182 (N_9182,N_8916,N_8958);
and U9183 (N_9183,N_8879,N_8877);
nor U9184 (N_9184,N_8831,N_8817);
nand U9185 (N_9185,N_8909,N_8895);
nand U9186 (N_9186,N_8897,N_8983);
nand U9187 (N_9187,N_8871,N_8856);
nand U9188 (N_9188,N_8813,N_8843);
nand U9189 (N_9189,N_8916,N_8938);
and U9190 (N_9190,N_8997,N_8884);
and U9191 (N_9191,N_8879,N_8948);
nor U9192 (N_9192,N_8986,N_8959);
and U9193 (N_9193,N_8925,N_8905);
and U9194 (N_9194,N_8978,N_8891);
or U9195 (N_9195,N_8808,N_8868);
nor U9196 (N_9196,N_8884,N_8848);
and U9197 (N_9197,N_8875,N_8894);
nor U9198 (N_9198,N_8814,N_8985);
nand U9199 (N_9199,N_8862,N_8809);
xnor U9200 (N_9200,N_9074,N_9140);
or U9201 (N_9201,N_9141,N_9165);
nand U9202 (N_9202,N_9090,N_9171);
and U9203 (N_9203,N_9180,N_9115);
nor U9204 (N_9204,N_9096,N_9143);
nor U9205 (N_9205,N_9101,N_9131);
and U9206 (N_9206,N_9052,N_9142);
and U9207 (N_9207,N_9166,N_9072);
and U9208 (N_9208,N_9054,N_9087);
and U9209 (N_9209,N_9123,N_9167);
nor U9210 (N_9210,N_9037,N_9047);
nor U9211 (N_9211,N_9153,N_9110);
and U9212 (N_9212,N_9125,N_9026);
or U9213 (N_9213,N_9084,N_9192);
xor U9214 (N_9214,N_9092,N_9046);
nand U9215 (N_9215,N_9000,N_9124);
and U9216 (N_9216,N_9158,N_9055);
and U9217 (N_9217,N_9027,N_9029);
nand U9218 (N_9218,N_9011,N_9107);
nand U9219 (N_9219,N_9059,N_9042);
xnor U9220 (N_9220,N_9195,N_9088);
or U9221 (N_9221,N_9068,N_9015);
and U9222 (N_9222,N_9089,N_9028);
xnor U9223 (N_9223,N_9170,N_9062);
or U9224 (N_9224,N_9024,N_9145);
and U9225 (N_9225,N_9113,N_9160);
and U9226 (N_9226,N_9112,N_9019);
or U9227 (N_9227,N_9130,N_9183);
nand U9228 (N_9228,N_9187,N_9091);
xnor U9229 (N_9229,N_9001,N_9151);
and U9230 (N_9230,N_9128,N_9106);
and U9231 (N_9231,N_9191,N_9005);
nand U9232 (N_9232,N_9033,N_9109);
nor U9233 (N_9233,N_9023,N_9117);
or U9234 (N_9234,N_9133,N_9134);
nand U9235 (N_9235,N_9061,N_9045);
nor U9236 (N_9236,N_9039,N_9032);
nand U9237 (N_9237,N_9065,N_9083);
xnor U9238 (N_9238,N_9149,N_9058);
nor U9239 (N_9239,N_9014,N_9021);
xnor U9240 (N_9240,N_9198,N_9002);
nor U9241 (N_9241,N_9114,N_9199);
nand U9242 (N_9242,N_9111,N_9067);
nand U9243 (N_9243,N_9152,N_9146);
nand U9244 (N_9244,N_9157,N_9012);
nor U9245 (N_9245,N_9094,N_9136);
xnor U9246 (N_9246,N_9186,N_9116);
nor U9247 (N_9247,N_9178,N_9020);
nand U9248 (N_9248,N_9138,N_9030);
nor U9249 (N_9249,N_9079,N_9105);
or U9250 (N_9250,N_9078,N_9036);
and U9251 (N_9251,N_9008,N_9098);
xor U9252 (N_9252,N_9189,N_9044);
nor U9253 (N_9253,N_9135,N_9075);
and U9254 (N_9254,N_9003,N_9102);
nand U9255 (N_9255,N_9070,N_9048);
and U9256 (N_9256,N_9077,N_9172);
xor U9257 (N_9257,N_9051,N_9161);
nand U9258 (N_9258,N_9095,N_9173);
nor U9259 (N_9259,N_9007,N_9154);
nand U9260 (N_9260,N_9038,N_9139);
nor U9261 (N_9261,N_9069,N_9184);
xnor U9262 (N_9262,N_9168,N_9179);
or U9263 (N_9263,N_9035,N_9018);
and U9264 (N_9264,N_9164,N_9085);
and U9265 (N_9265,N_9147,N_9022);
xnor U9266 (N_9266,N_9155,N_9043);
and U9267 (N_9267,N_9176,N_9122);
and U9268 (N_9268,N_9006,N_9196);
and U9269 (N_9269,N_9132,N_9063);
xor U9270 (N_9270,N_9159,N_9056);
nand U9271 (N_9271,N_9190,N_9119);
and U9272 (N_9272,N_9076,N_9148);
nand U9273 (N_9273,N_9057,N_9004);
nor U9274 (N_9274,N_9082,N_9041);
nor U9275 (N_9275,N_9193,N_9129);
nand U9276 (N_9276,N_9103,N_9118);
or U9277 (N_9277,N_9031,N_9093);
xnor U9278 (N_9278,N_9182,N_9144);
xnor U9279 (N_9279,N_9064,N_9169);
and U9280 (N_9280,N_9177,N_9013);
or U9281 (N_9281,N_9126,N_9066);
xnor U9282 (N_9282,N_9181,N_9034);
nand U9283 (N_9283,N_9025,N_9053);
nor U9284 (N_9284,N_9009,N_9081);
nand U9285 (N_9285,N_9097,N_9071);
and U9286 (N_9286,N_9121,N_9100);
nor U9287 (N_9287,N_9049,N_9197);
nand U9288 (N_9288,N_9185,N_9174);
nand U9289 (N_9289,N_9163,N_9080);
or U9290 (N_9290,N_9175,N_9127);
xnor U9291 (N_9291,N_9099,N_9150);
nand U9292 (N_9292,N_9188,N_9050);
and U9293 (N_9293,N_9017,N_9194);
nor U9294 (N_9294,N_9010,N_9086);
xnor U9295 (N_9295,N_9073,N_9156);
and U9296 (N_9296,N_9016,N_9120);
and U9297 (N_9297,N_9162,N_9108);
or U9298 (N_9298,N_9104,N_9060);
nor U9299 (N_9299,N_9040,N_9137);
and U9300 (N_9300,N_9106,N_9192);
nand U9301 (N_9301,N_9152,N_9057);
and U9302 (N_9302,N_9180,N_9098);
xnor U9303 (N_9303,N_9073,N_9152);
nand U9304 (N_9304,N_9008,N_9147);
nand U9305 (N_9305,N_9189,N_9160);
xnor U9306 (N_9306,N_9160,N_9192);
and U9307 (N_9307,N_9171,N_9102);
xnor U9308 (N_9308,N_9171,N_9189);
and U9309 (N_9309,N_9079,N_9025);
xnor U9310 (N_9310,N_9119,N_9088);
or U9311 (N_9311,N_9164,N_9017);
or U9312 (N_9312,N_9154,N_9079);
nor U9313 (N_9313,N_9149,N_9156);
nor U9314 (N_9314,N_9145,N_9118);
xnor U9315 (N_9315,N_9120,N_9107);
or U9316 (N_9316,N_9138,N_9018);
nand U9317 (N_9317,N_9180,N_9005);
or U9318 (N_9318,N_9007,N_9088);
nand U9319 (N_9319,N_9153,N_9048);
nand U9320 (N_9320,N_9088,N_9115);
xor U9321 (N_9321,N_9120,N_9005);
nand U9322 (N_9322,N_9124,N_9143);
or U9323 (N_9323,N_9020,N_9062);
or U9324 (N_9324,N_9164,N_9070);
or U9325 (N_9325,N_9185,N_9007);
nand U9326 (N_9326,N_9056,N_9193);
or U9327 (N_9327,N_9195,N_9166);
and U9328 (N_9328,N_9079,N_9126);
xor U9329 (N_9329,N_9167,N_9066);
nand U9330 (N_9330,N_9190,N_9168);
xnor U9331 (N_9331,N_9108,N_9016);
xor U9332 (N_9332,N_9009,N_9194);
nand U9333 (N_9333,N_9022,N_9084);
xnor U9334 (N_9334,N_9160,N_9012);
or U9335 (N_9335,N_9195,N_9121);
nor U9336 (N_9336,N_9186,N_9141);
and U9337 (N_9337,N_9025,N_9196);
or U9338 (N_9338,N_9159,N_9153);
xnor U9339 (N_9339,N_9135,N_9020);
or U9340 (N_9340,N_9188,N_9107);
and U9341 (N_9341,N_9185,N_9043);
or U9342 (N_9342,N_9108,N_9068);
nand U9343 (N_9343,N_9118,N_9018);
or U9344 (N_9344,N_9164,N_9097);
xor U9345 (N_9345,N_9003,N_9142);
nand U9346 (N_9346,N_9026,N_9190);
nor U9347 (N_9347,N_9066,N_9113);
xnor U9348 (N_9348,N_9005,N_9156);
nor U9349 (N_9349,N_9011,N_9109);
nand U9350 (N_9350,N_9139,N_9078);
and U9351 (N_9351,N_9011,N_9140);
nor U9352 (N_9352,N_9175,N_9079);
and U9353 (N_9353,N_9074,N_9053);
and U9354 (N_9354,N_9159,N_9112);
nand U9355 (N_9355,N_9107,N_9191);
xnor U9356 (N_9356,N_9006,N_9063);
nor U9357 (N_9357,N_9139,N_9150);
nor U9358 (N_9358,N_9199,N_9023);
or U9359 (N_9359,N_9143,N_9024);
and U9360 (N_9360,N_9127,N_9015);
or U9361 (N_9361,N_9005,N_9117);
xnor U9362 (N_9362,N_9098,N_9071);
or U9363 (N_9363,N_9109,N_9019);
nand U9364 (N_9364,N_9168,N_9098);
nand U9365 (N_9365,N_9012,N_9072);
nor U9366 (N_9366,N_9188,N_9143);
or U9367 (N_9367,N_9059,N_9007);
nand U9368 (N_9368,N_9089,N_9098);
nor U9369 (N_9369,N_9015,N_9162);
nand U9370 (N_9370,N_9086,N_9058);
and U9371 (N_9371,N_9145,N_9172);
nand U9372 (N_9372,N_9094,N_9112);
nor U9373 (N_9373,N_9151,N_9179);
xor U9374 (N_9374,N_9128,N_9114);
nor U9375 (N_9375,N_9135,N_9157);
nand U9376 (N_9376,N_9158,N_9155);
and U9377 (N_9377,N_9040,N_9078);
or U9378 (N_9378,N_9002,N_9167);
or U9379 (N_9379,N_9183,N_9053);
xor U9380 (N_9380,N_9176,N_9160);
nor U9381 (N_9381,N_9000,N_9184);
and U9382 (N_9382,N_9044,N_9048);
and U9383 (N_9383,N_9038,N_9123);
xnor U9384 (N_9384,N_9036,N_9147);
nor U9385 (N_9385,N_9016,N_9156);
nor U9386 (N_9386,N_9102,N_9145);
xnor U9387 (N_9387,N_9091,N_9095);
and U9388 (N_9388,N_9184,N_9005);
nor U9389 (N_9389,N_9133,N_9086);
or U9390 (N_9390,N_9101,N_9106);
nor U9391 (N_9391,N_9090,N_9130);
nor U9392 (N_9392,N_9031,N_9111);
xnor U9393 (N_9393,N_9003,N_9083);
nor U9394 (N_9394,N_9049,N_9196);
nand U9395 (N_9395,N_9034,N_9087);
nor U9396 (N_9396,N_9194,N_9175);
xnor U9397 (N_9397,N_9101,N_9147);
or U9398 (N_9398,N_9050,N_9015);
and U9399 (N_9399,N_9048,N_9049);
nor U9400 (N_9400,N_9247,N_9278);
or U9401 (N_9401,N_9392,N_9394);
nand U9402 (N_9402,N_9255,N_9375);
or U9403 (N_9403,N_9315,N_9213);
nand U9404 (N_9404,N_9296,N_9271);
and U9405 (N_9405,N_9306,N_9364);
nand U9406 (N_9406,N_9303,N_9376);
and U9407 (N_9407,N_9265,N_9219);
xor U9408 (N_9408,N_9372,N_9244);
or U9409 (N_9409,N_9206,N_9241);
nand U9410 (N_9410,N_9357,N_9359);
and U9411 (N_9411,N_9331,N_9277);
xor U9412 (N_9412,N_9238,N_9338);
nand U9413 (N_9413,N_9339,N_9388);
xor U9414 (N_9414,N_9363,N_9262);
and U9415 (N_9415,N_9371,N_9288);
xor U9416 (N_9416,N_9253,N_9208);
xnor U9417 (N_9417,N_9217,N_9270);
and U9418 (N_9418,N_9382,N_9209);
xnor U9419 (N_9419,N_9389,N_9378);
nand U9420 (N_9420,N_9311,N_9314);
nor U9421 (N_9421,N_9239,N_9292);
nand U9422 (N_9422,N_9350,N_9325);
nand U9423 (N_9423,N_9243,N_9283);
nor U9424 (N_9424,N_9286,N_9345);
and U9425 (N_9425,N_9301,N_9201);
nor U9426 (N_9426,N_9231,N_9294);
xor U9427 (N_9427,N_9398,N_9276);
nor U9428 (N_9428,N_9362,N_9387);
nand U9429 (N_9429,N_9220,N_9399);
xnor U9430 (N_9430,N_9366,N_9282);
xnor U9431 (N_9431,N_9384,N_9313);
nor U9432 (N_9432,N_9369,N_9302);
xor U9433 (N_9433,N_9308,N_9321);
and U9434 (N_9434,N_9335,N_9386);
nand U9435 (N_9435,N_9344,N_9305);
nor U9436 (N_9436,N_9379,N_9377);
xor U9437 (N_9437,N_9307,N_9237);
xnor U9438 (N_9438,N_9360,N_9333);
nor U9439 (N_9439,N_9367,N_9267);
xor U9440 (N_9440,N_9356,N_9273);
nand U9441 (N_9441,N_9318,N_9340);
and U9442 (N_9442,N_9353,N_9229);
and U9443 (N_9443,N_9210,N_9395);
nor U9444 (N_9444,N_9279,N_9355);
and U9445 (N_9445,N_9365,N_9212);
and U9446 (N_9446,N_9261,N_9290);
xnor U9447 (N_9447,N_9248,N_9274);
and U9448 (N_9448,N_9380,N_9312);
or U9449 (N_9449,N_9397,N_9242);
nand U9450 (N_9450,N_9250,N_9256);
or U9451 (N_9451,N_9245,N_9249);
xnor U9452 (N_9452,N_9200,N_9348);
xor U9453 (N_9453,N_9383,N_9309);
xor U9454 (N_9454,N_9260,N_9352);
nand U9455 (N_9455,N_9346,N_9203);
and U9456 (N_9456,N_9343,N_9205);
nand U9457 (N_9457,N_9299,N_9337);
and U9458 (N_9458,N_9264,N_9234);
nor U9459 (N_9459,N_9232,N_9204);
nand U9460 (N_9460,N_9287,N_9235);
xnor U9461 (N_9461,N_9396,N_9323);
xnor U9462 (N_9462,N_9289,N_9226);
xor U9463 (N_9463,N_9342,N_9297);
nor U9464 (N_9464,N_9324,N_9221);
nor U9465 (N_9465,N_9233,N_9224);
or U9466 (N_9466,N_9254,N_9216);
or U9467 (N_9467,N_9218,N_9317);
nor U9468 (N_9468,N_9257,N_9215);
nor U9469 (N_9469,N_9351,N_9284);
xor U9470 (N_9470,N_9236,N_9230);
xor U9471 (N_9471,N_9334,N_9223);
xnor U9472 (N_9472,N_9329,N_9298);
xnor U9473 (N_9473,N_9246,N_9272);
or U9474 (N_9474,N_9361,N_9295);
and U9475 (N_9475,N_9390,N_9370);
and U9476 (N_9476,N_9281,N_9381);
nor U9477 (N_9477,N_9251,N_9341);
or U9478 (N_9478,N_9358,N_9275);
nand U9479 (N_9479,N_9202,N_9300);
nor U9480 (N_9480,N_9336,N_9368);
or U9481 (N_9481,N_9316,N_9263);
xor U9482 (N_9482,N_9207,N_9328);
xnor U9483 (N_9483,N_9373,N_9259);
nor U9484 (N_9484,N_9293,N_9330);
or U9485 (N_9485,N_9332,N_9240);
nand U9486 (N_9486,N_9354,N_9211);
and U9487 (N_9487,N_9322,N_9326);
xnor U9488 (N_9488,N_9214,N_9349);
nand U9489 (N_9489,N_9310,N_9266);
xnor U9490 (N_9490,N_9393,N_9347);
xor U9491 (N_9491,N_9225,N_9319);
and U9492 (N_9492,N_9304,N_9252);
or U9493 (N_9493,N_9222,N_9228);
and U9494 (N_9494,N_9269,N_9285);
xnor U9495 (N_9495,N_9391,N_9280);
xor U9496 (N_9496,N_9374,N_9291);
xor U9497 (N_9497,N_9327,N_9268);
or U9498 (N_9498,N_9258,N_9320);
or U9499 (N_9499,N_9227,N_9385);
nor U9500 (N_9500,N_9368,N_9249);
nor U9501 (N_9501,N_9299,N_9378);
xnor U9502 (N_9502,N_9208,N_9320);
nor U9503 (N_9503,N_9235,N_9358);
nand U9504 (N_9504,N_9376,N_9248);
nand U9505 (N_9505,N_9325,N_9377);
and U9506 (N_9506,N_9282,N_9229);
and U9507 (N_9507,N_9254,N_9223);
xnor U9508 (N_9508,N_9308,N_9364);
nand U9509 (N_9509,N_9363,N_9204);
and U9510 (N_9510,N_9267,N_9217);
nand U9511 (N_9511,N_9368,N_9292);
or U9512 (N_9512,N_9396,N_9346);
xor U9513 (N_9513,N_9300,N_9377);
or U9514 (N_9514,N_9206,N_9369);
or U9515 (N_9515,N_9302,N_9392);
nand U9516 (N_9516,N_9394,N_9375);
nand U9517 (N_9517,N_9352,N_9218);
nor U9518 (N_9518,N_9305,N_9382);
xnor U9519 (N_9519,N_9270,N_9299);
nor U9520 (N_9520,N_9302,N_9269);
or U9521 (N_9521,N_9251,N_9384);
or U9522 (N_9522,N_9373,N_9287);
nor U9523 (N_9523,N_9359,N_9275);
xnor U9524 (N_9524,N_9320,N_9345);
and U9525 (N_9525,N_9349,N_9289);
xnor U9526 (N_9526,N_9367,N_9371);
and U9527 (N_9527,N_9273,N_9256);
or U9528 (N_9528,N_9326,N_9215);
or U9529 (N_9529,N_9341,N_9213);
or U9530 (N_9530,N_9386,N_9288);
xor U9531 (N_9531,N_9376,N_9334);
or U9532 (N_9532,N_9283,N_9240);
nor U9533 (N_9533,N_9211,N_9312);
and U9534 (N_9534,N_9399,N_9293);
nor U9535 (N_9535,N_9398,N_9355);
or U9536 (N_9536,N_9233,N_9226);
or U9537 (N_9537,N_9381,N_9303);
or U9538 (N_9538,N_9268,N_9386);
nor U9539 (N_9539,N_9306,N_9255);
or U9540 (N_9540,N_9301,N_9343);
nand U9541 (N_9541,N_9244,N_9373);
nand U9542 (N_9542,N_9346,N_9320);
nand U9543 (N_9543,N_9334,N_9383);
or U9544 (N_9544,N_9273,N_9274);
or U9545 (N_9545,N_9300,N_9299);
nand U9546 (N_9546,N_9207,N_9331);
or U9547 (N_9547,N_9338,N_9369);
or U9548 (N_9548,N_9280,N_9389);
nor U9549 (N_9549,N_9279,N_9370);
nand U9550 (N_9550,N_9357,N_9240);
and U9551 (N_9551,N_9312,N_9242);
nand U9552 (N_9552,N_9204,N_9371);
nor U9553 (N_9553,N_9205,N_9301);
xor U9554 (N_9554,N_9241,N_9248);
nor U9555 (N_9555,N_9239,N_9334);
or U9556 (N_9556,N_9325,N_9324);
or U9557 (N_9557,N_9330,N_9228);
and U9558 (N_9558,N_9374,N_9250);
nand U9559 (N_9559,N_9239,N_9349);
nand U9560 (N_9560,N_9239,N_9275);
xnor U9561 (N_9561,N_9289,N_9301);
xnor U9562 (N_9562,N_9305,N_9357);
or U9563 (N_9563,N_9209,N_9254);
or U9564 (N_9564,N_9353,N_9349);
and U9565 (N_9565,N_9281,N_9396);
xnor U9566 (N_9566,N_9248,N_9279);
and U9567 (N_9567,N_9357,N_9386);
or U9568 (N_9568,N_9332,N_9255);
nor U9569 (N_9569,N_9384,N_9204);
nand U9570 (N_9570,N_9257,N_9237);
xor U9571 (N_9571,N_9389,N_9226);
nor U9572 (N_9572,N_9374,N_9394);
xor U9573 (N_9573,N_9332,N_9362);
or U9574 (N_9574,N_9212,N_9231);
nor U9575 (N_9575,N_9277,N_9295);
nand U9576 (N_9576,N_9323,N_9249);
xor U9577 (N_9577,N_9253,N_9284);
nand U9578 (N_9578,N_9320,N_9268);
nand U9579 (N_9579,N_9207,N_9266);
and U9580 (N_9580,N_9238,N_9350);
and U9581 (N_9581,N_9261,N_9388);
xor U9582 (N_9582,N_9384,N_9390);
or U9583 (N_9583,N_9263,N_9393);
nand U9584 (N_9584,N_9328,N_9320);
xor U9585 (N_9585,N_9383,N_9277);
and U9586 (N_9586,N_9274,N_9332);
or U9587 (N_9587,N_9322,N_9370);
xor U9588 (N_9588,N_9323,N_9324);
nand U9589 (N_9589,N_9289,N_9205);
nor U9590 (N_9590,N_9249,N_9374);
xnor U9591 (N_9591,N_9348,N_9208);
and U9592 (N_9592,N_9367,N_9212);
nand U9593 (N_9593,N_9284,N_9208);
xor U9594 (N_9594,N_9383,N_9236);
nor U9595 (N_9595,N_9337,N_9350);
xor U9596 (N_9596,N_9386,N_9253);
and U9597 (N_9597,N_9219,N_9247);
xnor U9598 (N_9598,N_9292,N_9311);
and U9599 (N_9599,N_9321,N_9255);
and U9600 (N_9600,N_9581,N_9569);
nand U9601 (N_9601,N_9563,N_9475);
nor U9602 (N_9602,N_9440,N_9429);
or U9603 (N_9603,N_9519,N_9560);
and U9604 (N_9604,N_9520,N_9532);
nand U9605 (N_9605,N_9423,N_9461);
nor U9606 (N_9606,N_9593,N_9524);
nand U9607 (N_9607,N_9452,N_9506);
nand U9608 (N_9608,N_9580,N_9402);
nor U9609 (N_9609,N_9512,N_9582);
xor U9610 (N_9610,N_9443,N_9557);
nand U9611 (N_9611,N_9472,N_9533);
and U9612 (N_9612,N_9430,N_9568);
or U9613 (N_9613,N_9528,N_9553);
xor U9614 (N_9614,N_9438,N_9449);
and U9615 (N_9615,N_9482,N_9459);
xor U9616 (N_9616,N_9477,N_9505);
and U9617 (N_9617,N_9487,N_9561);
and U9618 (N_9618,N_9471,N_9501);
nand U9619 (N_9619,N_9525,N_9485);
nand U9620 (N_9620,N_9515,N_9473);
nor U9621 (N_9621,N_9474,N_9586);
nor U9622 (N_9622,N_9454,N_9433);
or U9623 (N_9623,N_9464,N_9518);
nor U9624 (N_9624,N_9543,N_9457);
or U9625 (N_9625,N_9508,N_9489);
xnor U9626 (N_9626,N_9427,N_9573);
xnor U9627 (N_9627,N_9495,N_9496);
nor U9628 (N_9628,N_9546,N_9597);
and U9629 (N_9629,N_9585,N_9534);
or U9630 (N_9630,N_9444,N_9539);
xor U9631 (N_9631,N_9535,N_9523);
nand U9632 (N_9632,N_9583,N_9577);
or U9633 (N_9633,N_9400,N_9590);
and U9634 (N_9634,N_9484,N_9432);
nand U9635 (N_9635,N_9467,N_9480);
nor U9636 (N_9636,N_9456,N_9510);
nand U9637 (N_9637,N_9572,N_9566);
nand U9638 (N_9638,N_9405,N_9556);
or U9639 (N_9639,N_9447,N_9504);
or U9640 (N_9640,N_9576,N_9409);
and U9641 (N_9641,N_9530,N_9536);
nand U9642 (N_9642,N_9413,N_9578);
or U9643 (N_9643,N_9542,N_9458);
or U9644 (N_9644,N_9417,N_9403);
or U9645 (N_9645,N_9550,N_9404);
or U9646 (N_9646,N_9595,N_9552);
nor U9647 (N_9647,N_9425,N_9559);
nor U9648 (N_9648,N_9493,N_9468);
nand U9649 (N_9649,N_9410,N_9579);
or U9650 (N_9650,N_9488,N_9416);
and U9651 (N_9651,N_9481,N_9509);
and U9652 (N_9652,N_9503,N_9526);
nor U9653 (N_9653,N_9406,N_9574);
nor U9654 (N_9654,N_9531,N_9465);
xor U9655 (N_9655,N_9497,N_9414);
xnor U9656 (N_9656,N_9599,N_9588);
xnor U9657 (N_9657,N_9537,N_9478);
nor U9658 (N_9658,N_9421,N_9470);
xor U9659 (N_9659,N_9411,N_9511);
and U9660 (N_9660,N_9451,N_9469);
xnor U9661 (N_9661,N_9426,N_9502);
nor U9662 (N_9662,N_9567,N_9545);
nor U9663 (N_9663,N_9492,N_9548);
and U9664 (N_9664,N_9446,N_9462);
xor U9665 (N_9665,N_9596,N_9419);
nor U9666 (N_9666,N_9538,N_9522);
nand U9667 (N_9667,N_9453,N_9460);
nand U9668 (N_9668,N_9499,N_9435);
nand U9669 (N_9669,N_9521,N_9500);
and U9670 (N_9670,N_9514,N_9491);
nand U9671 (N_9671,N_9558,N_9434);
or U9672 (N_9672,N_9476,N_9562);
nand U9673 (N_9673,N_9565,N_9439);
nand U9674 (N_9674,N_9494,N_9431);
xor U9675 (N_9675,N_9592,N_9437);
nand U9676 (N_9676,N_9415,N_9441);
or U9677 (N_9677,N_9541,N_9442);
nor U9678 (N_9678,N_9575,N_9455);
or U9679 (N_9679,N_9448,N_9450);
nand U9680 (N_9680,N_9570,N_9418);
or U9681 (N_9681,N_9479,N_9498);
xnor U9682 (N_9682,N_9540,N_9420);
or U9683 (N_9683,N_9555,N_9466);
or U9684 (N_9684,N_9428,N_9587);
nor U9685 (N_9685,N_9513,N_9571);
nor U9686 (N_9686,N_9554,N_9517);
nor U9687 (N_9687,N_9422,N_9412);
xnor U9688 (N_9688,N_9486,N_9527);
or U9689 (N_9689,N_9445,N_9490);
xnor U9690 (N_9690,N_9401,N_9544);
xnor U9691 (N_9691,N_9551,N_9591);
nand U9692 (N_9692,N_9407,N_9424);
nand U9693 (N_9693,N_9516,N_9436);
or U9694 (N_9694,N_9598,N_9483);
nor U9695 (N_9695,N_9584,N_9408);
and U9696 (N_9696,N_9589,N_9549);
xor U9697 (N_9697,N_9507,N_9594);
nor U9698 (N_9698,N_9529,N_9564);
or U9699 (N_9699,N_9463,N_9547);
and U9700 (N_9700,N_9496,N_9576);
and U9701 (N_9701,N_9491,N_9472);
and U9702 (N_9702,N_9546,N_9453);
xor U9703 (N_9703,N_9426,N_9561);
nor U9704 (N_9704,N_9552,N_9597);
and U9705 (N_9705,N_9518,N_9513);
nor U9706 (N_9706,N_9497,N_9565);
nand U9707 (N_9707,N_9474,N_9549);
or U9708 (N_9708,N_9494,N_9562);
nor U9709 (N_9709,N_9523,N_9441);
or U9710 (N_9710,N_9408,N_9583);
nor U9711 (N_9711,N_9498,N_9574);
and U9712 (N_9712,N_9520,N_9516);
nand U9713 (N_9713,N_9404,N_9496);
xnor U9714 (N_9714,N_9527,N_9430);
nor U9715 (N_9715,N_9471,N_9599);
or U9716 (N_9716,N_9507,N_9450);
nor U9717 (N_9717,N_9407,N_9587);
nand U9718 (N_9718,N_9526,N_9443);
xnor U9719 (N_9719,N_9518,N_9463);
xnor U9720 (N_9720,N_9532,N_9592);
xnor U9721 (N_9721,N_9417,N_9565);
xnor U9722 (N_9722,N_9586,N_9498);
xor U9723 (N_9723,N_9465,N_9479);
xor U9724 (N_9724,N_9415,N_9584);
nand U9725 (N_9725,N_9433,N_9578);
and U9726 (N_9726,N_9518,N_9563);
or U9727 (N_9727,N_9408,N_9483);
and U9728 (N_9728,N_9569,N_9478);
nor U9729 (N_9729,N_9441,N_9521);
xnor U9730 (N_9730,N_9588,N_9446);
or U9731 (N_9731,N_9515,N_9467);
nor U9732 (N_9732,N_9421,N_9413);
and U9733 (N_9733,N_9594,N_9501);
nor U9734 (N_9734,N_9526,N_9516);
or U9735 (N_9735,N_9519,N_9523);
or U9736 (N_9736,N_9485,N_9460);
nor U9737 (N_9737,N_9484,N_9588);
or U9738 (N_9738,N_9569,N_9423);
or U9739 (N_9739,N_9536,N_9551);
and U9740 (N_9740,N_9495,N_9593);
nand U9741 (N_9741,N_9538,N_9596);
and U9742 (N_9742,N_9471,N_9586);
nand U9743 (N_9743,N_9491,N_9419);
and U9744 (N_9744,N_9519,N_9593);
xor U9745 (N_9745,N_9486,N_9423);
nor U9746 (N_9746,N_9505,N_9524);
and U9747 (N_9747,N_9492,N_9443);
xor U9748 (N_9748,N_9472,N_9450);
xnor U9749 (N_9749,N_9529,N_9448);
or U9750 (N_9750,N_9514,N_9525);
xnor U9751 (N_9751,N_9493,N_9480);
nand U9752 (N_9752,N_9593,N_9477);
xor U9753 (N_9753,N_9583,N_9442);
or U9754 (N_9754,N_9452,N_9425);
or U9755 (N_9755,N_9493,N_9522);
nand U9756 (N_9756,N_9429,N_9521);
xnor U9757 (N_9757,N_9497,N_9581);
or U9758 (N_9758,N_9568,N_9556);
xnor U9759 (N_9759,N_9533,N_9515);
or U9760 (N_9760,N_9482,N_9514);
nand U9761 (N_9761,N_9519,N_9489);
nor U9762 (N_9762,N_9564,N_9434);
and U9763 (N_9763,N_9401,N_9554);
or U9764 (N_9764,N_9423,N_9538);
nor U9765 (N_9765,N_9430,N_9411);
or U9766 (N_9766,N_9522,N_9446);
nor U9767 (N_9767,N_9538,N_9572);
xor U9768 (N_9768,N_9594,N_9431);
nor U9769 (N_9769,N_9573,N_9403);
or U9770 (N_9770,N_9488,N_9571);
or U9771 (N_9771,N_9571,N_9529);
nand U9772 (N_9772,N_9443,N_9530);
nand U9773 (N_9773,N_9441,N_9503);
and U9774 (N_9774,N_9497,N_9433);
xor U9775 (N_9775,N_9573,N_9537);
and U9776 (N_9776,N_9442,N_9524);
or U9777 (N_9777,N_9484,N_9586);
xnor U9778 (N_9778,N_9426,N_9568);
or U9779 (N_9779,N_9499,N_9528);
nor U9780 (N_9780,N_9574,N_9562);
nand U9781 (N_9781,N_9497,N_9501);
xor U9782 (N_9782,N_9407,N_9414);
and U9783 (N_9783,N_9457,N_9563);
nand U9784 (N_9784,N_9412,N_9565);
nand U9785 (N_9785,N_9475,N_9513);
nor U9786 (N_9786,N_9479,N_9530);
and U9787 (N_9787,N_9465,N_9411);
and U9788 (N_9788,N_9540,N_9495);
xor U9789 (N_9789,N_9402,N_9512);
and U9790 (N_9790,N_9567,N_9556);
nand U9791 (N_9791,N_9591,N_9575);
nor U9792 (N_9792,N_9442,N_9469);
or U9793 (N_9793,N_9520,N_9556);
nor U9794 (N_9794,N_9598,N_9500);
xnor U9795 (N_9795,N_9407,N_9543);
nand U9796 (N_9796,N_9553,N_9505);
xor U9797 (N_9797,N_9429,N_9557);
or U9798 (N_9798,N_9425,N_9429);
nor U9799 (N_9799,N_9479,N_9421);
and U9800 (N_9800,N_9655,N_9754);
nor U9801 (N_9801,N_9631,N_9791);
or U9802 (N_9802,N_9710,N_9740);
or U9803 (N_9803,N_9693,N_9780);
xor U9804 (N_9804,N_9797,N_9739);
xnor U9805 (N_9805,N_9604,N_9657);
nor U9806 (N_9806,N_9783,N_9672);
nor U9807 (N_9807,N_9744,N_9666);
and U9808 (N_9808,N_9768,N_9728);
xor U9809 (N_9809,N_9712,N_9733);
xnor U9810 (N_9810,N_9701,N_9749);
nor U9811 (N_9811,N_9608,N_9772);
nand U9812 (N_9812,N_9775,N_9784);
xnor U9813 (N_9813,N_9626,N_9747);
or U9814 (N_9814,N_9792,N_9602);
xnor U9815 (N_9815,N_9796,N_9702);
and U9816 (N_9816,N_9774,N_9600);
xor U9817 (N_9817,N_9676,N_9644);
xnor U9818 (N_9818,N_9659,N_9715);
or U9819 (N_9819,N_9789,N_9724);
nor U9820 (N_9820,N_9759,N_9748);
xnor U9821 (N_9821,N_9786,N_9645);
nand U9822 (N_9822,N_9623,N_9713);
or U9823 (N_9823,N_9764,N_9723);
nand U9824 (N_9824,N_9656,N_9681);
nand U9825 (N_9825,N_9790,N_9781);
nor U9826 (N_9826,N_9741,N_9606);
xnor U9827 (N_9827,N_9738,N_9716);
nand U9828 (N_9828,N_9782,N_9660);
or U9829 (N_9829,N_9650,N_9665);
nand U9830 (N_9830,N_9717,N_9767);
nor U9831 (N_9831,N_9758,N_9615);
and U9832 (N_9832,N_9787,N_9755);
or U9833 (N_9833,N_9640,N_9722);
nor U9834 (N_9834,N_9674,N_9621);
or U9835 (N_9835,N_9699,N_9680);
xor U9836 (N_9836,N_9779,N_9730);
or U9837 (N_9837,N_9620,N_9647);
nand U9838 (N_9838,N_9751,N_9766);
nor U9839 (N_9839,N_9703,N_9669);
and U9840 (N_9840,N_9698,N_9601);
nor U9841 (N_9841,N_9616,N_9641);
xor U9842 (N_9842,N_9663,N_9605);
or U9843 (N_9843,N_9736,N_9709);
nand U9844 (N_9844,N_9675,N_9682);
and U9845 (N_9845,N_9707,N_9765);
and U9846 (N_9846,N_9607,N_9636);
and U9847 (N_9847,N_9706,N_9750);
xor U9848 (N_9848,N_9731,N_9684);
xnor U9849 (N_9849,N_9637,N_9757);
or U9850 (N_9850,N_9688,N_9726);
xor U9851 (N_9851,N_9756,N_9610);
or U9852 (N_9852,N_9795,N_9668);
xnor U9853 (N_9853,N_9687,N_9760);
or U9854 (N_9854,N_9671,N_9737);
nor U9855 (N_9855,N_9634,N_9617);
nor U9856 (N_9856,N_9679,N_9695);
nor U9857 (N_9857,N_9727,N_9611);
or U9858 (N_9858,N_9619,N_9633);
nor U9859 (N_9859,N_9705,N_9742);
or U9860 (N_9860,N_9670,N_9649);
nand U9861 (N_9861,N_9714,N_9643);
and U9862 (N_9862,N_9799,N_9652);
nand U9863 (N_9863,N_9720,N_9735);
or U9864 (N_9864,N_9694,N_9614);
nand U9865 (N_9865,N_9662,N_9632);
xnor U9866 (N_9866,N_9794,N_9721);
and U9867 (N_9867,N_9770,N_9776);
nor U9868 (N_9868,N_9661,N_9685);
and U9869 (N_9869,N_9769,N_9648);
or U9870 (N_9870,N_9704,N_9651);
nand U9871 (N_9871,N_9628,N_9683);
nand U9872 (N_9872,N_9708,N_9778);
or U9873 (N_9873,N_9732,N_9658);
xor U9874 (N_9874,N_9788,N_9677);
or U9875 (N_9875,N_9696,N_9725);
xnor U9876 (N_9876,N_9734,N_9664);
or U9877 (N_9877,N_9771,N_9653);
nor U9878 (N_9878,N_9654,N_9603);
nor U9879 (N_9879,N_9686,N_9678);
nor U9880 (N_9880,N_9793,N_9773);
xor U9881 (N_9881,N_9743,N_9746);
nor U9882 (N_9882,N_9612,N_9763);
and U9883 (N_9883,N_9642,N_9798);
or U9884 (N_9884,N_9618,N_9785);
and U9885 (N_9885,N_9625,N_9635);
nor U9886 (N_9886,N_9718,N_9752);
or U9887 (N_9887,N_9624,N_9700);
or U9888 (N_9888,N_9630,N_9691);
and U9889 (N_9889,N_9673,N_9762);
or U9890 (N_9890,N_9646,N_9711);
xor U9891 (N_9891,N_9777,N_9719);
nor U9892 (N_9892,N_9690,N_9627);
xor U9893 (N_9893,N_9638,N_9692);
nor U9894 (N_9894,N_9629,N_9745);
nand U9895 (N_9895,N_9697,N_9753);
or U9896 (N_9896,N_9761,N_9667);
nand U9897 (N_9897,N_9613,N_9729);
or U9898 (N_9898,N_9639,N_9622);
nor U9899 (N_9899,N_9609,N_9689);
nand U9900 (N_9900,N_9707,N_9795);
or U9901 (N_9901,N_9703,N_9605);
or U9902 (N_9902,N_9657,N_9684);
and U9903 (N_9903,N_9697,N_9716);
and U9904 (N_9904,N_9663,N_9741);
or U9905 (N_9905,N_9627,N_9705);
xnor U9906 (N_9906,N_9697,N_9653);
nor U9907 (N_9907,N_9626,N_9678);
xnor U9908 (N_9908,N_9766,N_9626);
nand U9909 (N_9909,N_9757,N_9755);
nor U9910 (N_9910,N_9686,N_9734);
xnor U9911 (N_9911,N_9793,N_9681);
or U9912 (N_9912,N_9696,N_9636);
nand U9913 (N_9913,N_9631,N_9735);
xnor U9914 (N_9914,N_9758,N_9683);
nor U9915 (N_9915,N_9718,N_9630);
xor U9916 (N_9916,N_9602,N_9638);
xor U9917 (N_9917,N_9629,N_9618);
and U9918 (N_9918,N_9649,N_9728);
nand U9919 (N_9919,N_9654,N_9661);
or U9920 (N_9920,N_9655,N_9639);
and U9921 (N_9921,N_9778,N_9632);
and U9922 (N_9922,N_9771,N_9674);
xnor U9923 (N_9923,N_9711,N_9657);
nand U9924 (N_9924,N_9736,N_9612);
or U9925 (N_9925,N_9623,N_9647);
nand U9926 (N_9926,N_9666,N_9648);
or U9927 (N_9927,N_9695,N_9757);
and U9928 (N_9928,N_9755,N_9768);
xor U9929 (N_9929,N_9759,N_9715);
nand U9930 (N_9930,N_9762,N_9674);
and U9931 (N_9931,N_9783,N_9606);
nor U9932 (N_9932,N_9765,N_9612);
and U9933 (N_9933,N_9616,N_9734);
nor U9934 (N_9934,N_9606,N_9610);
nor U9935 (N_9935,N_9699,N_9647);
nand U9936 (N_9936,N_9756,N_9722);
nor U9937 (N_9937,N_9683,N_9611);
or U9938 (N_9938,N_9678,N_9643);
nand U9939 (N_9939,N_9620,N_9663);
or U9940 (N_9940,N_9604,N_9612);
nand U9941 (N_9941,N_9653,N_9794);
nor U9942 (N_9942,N_9742,N_9712);
xor U9943 (N_9943,N_9727,N_9632);
xor U9944 (N_9944,N_9771,N_9602);
xnor U9945 (N_9945,N_9777,N_9754);
or U9946 (N_9946,N_9666,N_9682);
xnor U9947 (N_9947,N_9717,N_9708);
nor U9948 (N_9948,N_9617,N_9776);
nor U9949 (N_9949,N_9744,N_9752);
nand U9950 (N_9950,N_9643,N_9737);
nand U9951 (N_9951,N_9784,N_9712);
xor U9952 (N_9952,N_9614,N_9775);
or U9953 (N_9953,N_9709,N_9793);
nand U9954 (N_9954,N_9733,N_9754);
xnor U9955 (N_9955,N_9671,N_9672);
xnor U9956 (N_9956,N_9667,N_9705);
and U9957 (N_9957,N_9768,N_9622);
or U9958 (N_9958,N_9706,N_9703);
nor U9959 (N_9959,N_9632,N_9658);
xor U9960 (N_9960,N_9743,N_9646);
nand U9961 (N_9961,N_9729,N_9601);
nor U9962 (N_9962,N_9713,N_9683);
xnor U9963 (N_9963,N_9774,N_9658);
xor U9964 (N_9964,N_9770,N_9768);
or U9965 (N_9965,N_9739,N_9708);
xnor U9966 (N_9966,N_9791,N_9758);
xor U9967 (N_9967,N_9792,N_9629);
nand U9968 (N_9968,N_9789,N_9732);
or U9969 (N_9969,N_9789,N_9609);
nand U9970 (N_9970,N_9798,N_9609);
xor U9971 (N_9971,N_9735,N_9788);
nor U9972 (N_9972,N_9635,N_9791);
nand U9973 (N_9973,N_9610,N_9755);
nor U9974 (N_9974,N_9783,N_9762);
xnor U9975 (N_9975,N_9769,N_9612);
nand U9976 (N_9976,N_9738,N_9786);
nor U9977 (N_9977,N_9770,N_9662);
and U9978 (N_9978,N_9716,N_9731);
or U9979 (N_9979,N_9713,N_9644);
xor U9980 (N_9980,N_9706,N_9660);
xnor U9981 (N_9981,N_9773,N_9769);
nor U9982 (N_9982,N_9624,N_9602);
nor U9983 (N_9983,N_9719,N_9713);
xor U9984 (N_9984,N_9772,N_9744);
nand U9985 (N_9985,N_9718,N_9607);
and U9986 (N_9986,N_9674,N_9778);
nor U9987 (N_9987,N_9767,N_9686);
xor U9988 (N_9988,N_9613,N_9703);
and U9989 (N_9989,N_9698,N_9715);
nor U9990 (N_9990,N_9622,N_9643);
nor U9991 (N_9991,N_9644,N_9650);
nand U9992 (N_9992,N_9756,N_9693);
nor U9993 (N_9993,N_9734,N_9707);
and U9994 (N_9994,N_9685,N_9614);
or U9995 (N_9995,N_9706,N_9761);
nand U9996 (N_9996,N_9776,N_9769);
or U9997 (N_9997,N_9677,N_9790);
xor U9998 (N_9998,N_9694,N_9792);
xnor U9999 (N_9999,N_9684,N_9633);
nor U10000 (N_10000,N_9954,N_9967);
and U10001 (N_10001,N_9816,N_9956);
nor U10002 (N_10002,N_9952,N_9811);
nand U10003 (N_10003,N_9986,N_9812);
nor U10004 (N_10004,N_9961,N_9910);
nand U10005 (N_10005,N_9832,N_9942);
and U10006 (N_10006,N_9810,N_9899);
xor U10007 (N_10007,N_9980,N_9839);
and U10008 (N_10008,N_9851,N_9886);
nand U10009 (N_10009,N_9997,N_9809);
and U10010 (N_10010,N_9999,N_9892);
xnor U10011 (N_10011,N_9978,N_9893);
nand U10012 (N_10012,N_9920,N_9820);
or U10013 (N_10013,N_9857,N_9911);
nand U10014 (N_10014,N_9891,N_9938);
nor U10015 (N_10015,N_9968,N_9971);
nor U10016 (N_10016,N_9885,N_9991);
xnor U10017 (N_10017,N_9840,N_9951);
or U10018 (N_10018,N_9982,N_9960);
and U10019 (N_10019,N_9950,N_9970);
nor U10020 (N_10020,N_9888,N_9930);
xnor U10021 (N_10021,N_9932,N_9922);
xnor U10022 (N_10022,N_9824,N_9829);
or U10023 (N_10023,N_9965,N_9807);
nand U10024 (N_10024,N_9963,N_9936);
and U10025 (N_10025,N_9831,N_9800);
and U10026 (N_10026,N_9988,N_9926);
nor U10027 (N_10027,N_9958,N_9803);
and U10028 (N_10028,N_9858,N_9947);
nand U10029 (N_10029,N_9868,N_9901);
and U10030 (N_10030,N_9924,N_9828);
and U10031 (N_10031,N_9964,N_9996);
and U10032 (N_10032,N_9909,N_9976);
and U10033 (N_10033,N_9802,N_9877);
xor U10034 (N_10034,N_9849,N_9940);
xor U10035 (N_10035,N_9833,N_9902);
xnor U10036 (N_10036,N_9973,N_9869);
and U10037 (N_10037,N_9846,N_9850);
and U10038 (N_10038,N_9896,N_9919);
xnor U10039 (N_10039,N_9863,N_9908);
nor U10040 (N_10040,N_9992,N_9962);
and U10041 (N_10041,N_9998,N_9881);
or U10042 (N_10042,N_9853,N_9972);
xnor U10043 (N_10043,N_9925,N_9861);
or U10044 (N_10044,N_9979,N_9990);
nand U10045 (N_10045,N_9921,N_9887);
xnor U10046 (N_10046,N_9981,N_9854);
nor U10047 (N_10047,N_9928,N_9834);
nand U10048 (N_10048,N_9989,N_9934);
nand U10049 (N_10049,N_9848,N_9856);
and U10050 (N_10050,N_9826,N_9819);
and U10051 (N_10051,N_9917,N_9873);
and U10052 (N_10052,N_9813,N_9953);
xor U10053 (N_10053,N_9955,N_9859);
or U10054 (N_10054,N_9895,N_9927);
or U10055 (N_10055,N_9801,N_9935);
or U10056 (N_10056,N_9984,N_9879);
nor U10057 (N_10057,N_9823,N_9852);
nand U10058 (N_10058,N_9949,N_9866);
nor U10059 (N_10059,N_9845,N_9843);
or U10060 (N_10060,N_9876,N_9874);
nand U10061 (N_10061,N_9941,N_9870);
or U10062 (N_10062,N_9966,N_9806);
nand U10063 (N_10063,N_9903,N_9842);
or U10064 (N_10064,N_9918,N_9841);
nand U10065 (N_10065,N_9975,N_9864);
nand U10066 (N_10066,N_9844,N_9983);
xnor U10067 (N_10067,N_9860,N_9937);
nor U10068 (N_10068,N_9957,N_9916);
xor U10069 (N_10069,N_9945,N_9946);
nand U10070 (N_10070,N_9987,N_9822);
and U10071 (N_10071,N_9974,N_9808);
xor U10072 (N_10072,N_9875,N_9900);
or U10073 (N_10073,N_9871,N_9929);
xnor U10074 (N_10074,N_9818,N_9906);
or U10075 (N_10075,N_9867,N_9884);
xnor U10076 (N_10076,N_9931,N_9865);
and U10077 (N_10077,N_9855,N_9872);
or U10078 (N_10078,N_9883,N_9835);
and U10079 (N_10079,N_9830,N_9804);
nand U10080 (N_10080,N_9993,N_9894);
nor U10081 (N_10081,N_9969,N_9821);
xnor U10082 (N_10082,N_9890,N_9862);
nand U10083 (N_10083,N_9815,N_9837);
nor U10084 (N_10084,N_9913,N_9880);
and U10085 (N_10085,N_9905,N_9944);
or U10086 (N_10086,N_9817,N_9897);
xor U10087 (N_10087,N_9939,N_9814);
or U10088 (N_10088,N_9827,N_9878);
nand U10089 (N_10089,N_9882,N_9912);
nor U10090 (N_10090,N_9995,N_9915);
or U10091 (N_10091,N_9985,N_9923);
or U10092 (N_10092,N_9889,N_9836);
xnor U10093 (N_10093,N_9948,N_9805);
nor U10094 (N_10094,N_9959,N_9994);
xnor U10095 (N_10095,N_9907,N_9898);
and U10096 (N_10096,N_9825,N_9838);
nand U10097 (N_10097,N_9943,N_9904);
nor U10098 (N_10098,N_9977,N_9933);
or U10099 (N_10099,N_9914,N_9847);
or U10100 (N_10100,N_9973,N_9876);
nor U10101 (N_10101,N_9914,N_9954);
xnor U10102 (N_10102,N_9959,N_9891);
xnor U10103 (N_10103,N_9979,N_9811);
and U10104 (N_10104,N_9866,N_9962);
xor U10105 (N_10105,N_9961,N_9852);
xor U10106 (N_10106,N_9921,N_9822);
xnor U10107 (N_10107,N_9814,N_9810);
xnor U10108 (N_10108,N_9842,N_9965);
or U10109 (N_10109,N_9878,N_9931);
nand U10110 (N_10110,N_9940,N_9802);
xor U10111 (N_10111,N_9988,N_9985);
and U10112 (N_10112,N_9907,N_9934);
or U10113 (N_10113,N_9960,N_9946);
xor U10114 (N_10114,N_9901,N_9824);
xnor U10115 (N_10115,N_9982,N_9921);
nand U10116 (N_10116,N_9864,N_9945);
and U10117 (N_10117,N_9828,N_9897);
and U10118 (N_10118,N_9831,N_9897);
nor U10119 (N_10119,N_9848,N_9996);
xor U10120 (N_10120,N_9979,N_9946);
nand U10121 (N_10121,N_9823,N_9834);
xnor U10122 (N_10122,N_9928,N_9818);
nor U10123 (N_10123,N_9958,N_9998);
or U10124 (N_10124,N_9940,N_9838);
and U10125 (N_10125,N_9810,N_9857);
and U10126 (N_10126,N_9818,N_9859);
xor U10127 (N_10127,N_9838,N_9986);
nand U10128 (N_10128,N_9873,N_9913);
nand U10129 (N_10129,N_9906,N_9845);
nor U10130 (N_10130,N_9803,N_9994);
xor U10131 (N_10131,N_9963,N_9849);
and U10132 (N_10132,N_9897,N_9852);
nor U10133 (N_10133,N_9859,N_9867);
nor U10134 (N_10134,N_9884,N_9871);
xor U10135 (N_10135,N_9970,N_9869);
xor U10136 (N_10136,N_9988,N_9827);
nor U10137 (N_10137,N_9833,N_9856);
and U10138 (N_10138,N_9852,N_9870);
and U10139 (N_10139,N_9939,N_9810);
nand U10140 (N_10140,N_9842,N_9953);
or U10141 (N_10141,N_9982,N_9803);
nand U10142 (N_10142,N_9924,N_9807);
and U10143 (N_10143,N_9846,N_9885);
xor U10144 (N_10144,N_9967,N_9869);
nand U10145 (N_10145,N_9940,N_9878);
nand U10146 (N_10146,N_9961,N_9829);
nor U10147 (N_10147,N_9816,N_9950);
xnor U10148 (N_10148,N_9876,N_9864);
nand U10149 (N_10149,N_9989,N_9889);
nor U10150 (N_10150,N_9845,N_9820);
or U10151 (N_10151,N_9939,N_9986);
nor U10152 (N_10152,N_9925,N_9877);
or U10153 (N_10153,N_9895,N_9958);
nand U10154 (N_10154,N_9999,N_9828);
and U10155 (N_10155,N_9878,N_9986);
nand U10156 (N_10156,N_9812,N_9895);
or U10157 (N_10157,N_9851,N_9949);
nand U10158 (N_10158,N_9867,N_9985);
nor U10159 (N_10159,N_9899,N_9873);
and U10160 (N_10160,N_9963,N_9944);
or U10161 (N_10161,N_9977,N_9900);
nand U10162 (N_10162,N_9842,N_9827);
or U10163 (N_10163,N_9935,N_9838);
or U10164 (N_10164,N_9934,N_9890);
nor U10165 (N_10165,N_9964,N_9919);
or U10166 (N_10166,N_9950,N_9903);
xor U10167 (N_10167,N_9986,N_9993);
or U10168 (N_10168,N_9863,N_9915);
nor U10169 (N_10169,N_9947,N_9843);
and U10170 (N_10170,N_9819,N_9882);
xor U10171 (N_10171,N_9923,N_9895);
xnor U10172 (N_10172,N_9830,N_9941);
xnor U10173 (N_10173,N_9877,N_9904);
or U10174 (N_10174,N_9963,N_9965);
nand U10175 (N_10175,N_9821,N_9939);
and U10176 (N_10176,N_9927,N_9963);
xor U10177 (N_10177,N_9802,N_9932);
and U10178 (N_10178,N_9966,N_9999);
xnor U10179 (N_10179,N_9838,N_9949);
and U10180 (N_10180,N_9972,N_9808);
nor U10181 (N_10181,N_9806,N_9935);
xor U10182 (N_10182,N_9943,N_9853);
xor U10183 (N_10183,N_9809,N_9990);
and U10184 (N_10184,N_9824,N_9935);
nor U10185 (N_10185,N_9875,N_9881);
or U10186 (N_10186,N_9815,N_9810);
nor U10187 (N_10187,N_9980,N_9835);
or U10188 (N_10188,N_9815,N_9955);
or U10189 (N_10189,N_9996,N_9805);
nand U10190 (N_10190,N_9822,N_9979);
nand U10191 (N_10191,N_9962,N_9855);
nand U10192 (N_10192,N_9968,N_9918);
and U10193 (N_10193,N_9965,N_9992);
or U10194 (N_10194,N_9822,N_9841);
or U10195 (N_10195,N_9943,N_9989);
xor U10196 (N_10196,N_9950,N_9854);
nor U10197 (N_10197,N_9938,N_9955);
nand U10198 (N_10198,N_9803,N_9948);
xnor U10199 (N_10199,N_9847,N_9835);
nor U10200 (N_10200,N_10010,N_10030);
or U10201 (N_10201,N_10199,N_10162);
nand U10202 (N_10202,N_10111,N_10123);
and U10203 (N_10203,N_10044,N_10128);
or U10204 (N_10204,N_10102,N_10143);
and U10205 (N_10205,N_10029,N_10095);
nand U10206 (N_10206,N_10194,N_10121);
nor U10207 (N_10207,N_10116,N_10184);
nor U10208 (N_10208,N_10087,N_10060);
and U10209 (N_10209,N_10131,N_10022);
nand U10210 (N_10210,N_10046,N_10100);
nand U10211 (N_10211,N_10141,N_10070);
xor U10212 (N_10212,N_10172,N_10105);
and U10213 (N_10213,N_10197,N_10097);
nor U10214 (N_10214,N_10024,N_10084);
nor U10215 (N_10215,N_10074,N_10021);
or U10216 (N_10216,N_10023,N_10055);
and U10217 (N_10217,N_10049,N_10138);
nand U10218 (N_10218,N_10176,N_10028);
xor U10219 (N_10219,N_10135,N_10004);
nor U10220 (N_10220,N_10040,N_10114);
nand U10221 (N_10221,N_10191,N_10025);
and U10222 (N_10222,N_10042,N_10003);
nor U10223 (N_10223,N_10034,N_10056);
and U10224 (N_10224,N_10079,N_10092);
or U10225 (N_10225,N_10149,N_10071);
and U10226 (N_10226,N_10190,N_10112);
xnor U10227 (N_10227,N_10122,N_10140);
or U10228 (N_10228,N_10125,N_10072);
nor U10229 (N_10229,N_10158,N_10189);
xor U10230 (N_10230,N_10136,N_10053);
nor U10231 (N_10231,N_10065,N_10075);
xnor U10232 (N_10232,N_10057,N_10059);
and U10233 (N_10233,N_10076,N_10089);
or U10234 (N_10234,N_10082,N_10148);
and U10235 (N_10235,N_10073,N_10164);
nor U10236 (N_10236,N_10093,N_10129);
or U10237 (N_10237,N_10033,N_10038);
nand U10238 (N_10238,N_10110,N_10007);
nand U10239 (N_10239,N_10005,N_10167);
or U10240 (N_10240,N_10163,N_10181);
xor U10241 (N_10241,N_10147,N_10168);
and U10242 (N_10242,N_10054,N_10026);
or U10243 (N_10243,N_10017,N_10002);
nor U10244 (N_10244,N_10118,N_10179);
or U10245 (N_10245,N_10193,N_10088);
nor U10246 (N_10246,N_10186,N_10183);
and U10247 (N_10247,N_10098,N_10000);
nor U10248 (N_10248,N_10083,N_10019);
nand U10249 (N_10249,N_10165,N_10146);
or U10250 (N_10250,N_10012,N_10036);
nor U10251 (N_10251,N_10177,N_10144);
or U10252 (N_10252,N_10182,N_10086);
and U10253 (N_10253,N_10081,N_10117);
xnor U10254 (N_10254,N_10159,N_10015);
xor U10255 (N_10255,N_10067,N_10134);
nor U10256 (N_10256,N_10156,N_10068);
or U10257 (N_10257,N_10062,N_10139);
or U10258 (N_10258,N_10103,N_10195);
nand U10259 (N_10259,N_10152,N_10187);
nand U10260 (N_10260,N_10009,N_10064);
xor U10261 (N_10261,N_10014,N_10047);
xnor U10262 (N_10262,N_10192,N_10185);
xor U10263 (N_10263,N_10085,N_10171);
or U10264 (N_10264,N_10066,N_10126);
or U10265 (N_10265,N_10150,N_10006);
nand U10266 (N_10266,N_10178,N_10101);
nand U10267 (N_10267,N_10013,N_10018);
nor U10268 (N_10268,N_10173,N_10106);
or U10269 (N_10269,N_10142,N_10127);
nand U10270 (N_10270,N_10174,N_10096);
xnor U10271 (N_10271,N_10050,N_10069);
nor U10272 (N_10272,N_10031,N_10032);
or U10273 (N_10273,N_10137,N_10035);
and U10274 (N_10274,N_10052,N_10107);
or U10275 (N_10275,N_10115,N_10094);
nor U10276 (N_10276,N_10166,N_10154);
nand U10277 (N_10277,N_10037,N_10169);
xor U10278 (N_10278,N_10020,N_10161);
and U10279 (N_10279,N_10188,N_10043);
xor U10280 (N_10280,N_10153,N_10051);
nand U10281 (N_10281,N_10124,N_10198);
xnor U10282 (N_10282,N_10109,N_10080);
nor U10283 (N_10283,N_10011,N_10077);
and U10284 (N_10284,N_10099,N_10090);
xor U10285 (N_10285,N_10145,N_10008);
and U10286 (N_10286,N_10170,N_10157);
and U10287 (N_10287,N_10119,N_10196);
and U10288 (N_10288,N_10133,N_10151);
nor U10289 (N_10289,N_10061,N_10132);
nor U10290 (N_10290,N_10039,N_10113);
nor U10291 (N_10291,N_10155,N_10180);
and U10292 (N_10292,N_10108,N_10048);
xor U10293 (N_10293,N_10058,N_10078);
nor U10294 (N_10294,N_10130,N_10027);
or U10295 (N_10295,N_10001,N_10175);
nand U10296 (N_10296,N_10091,N_10104);
nor U10297 (N_10297,N_10120,N_10016);
or U10298 (N_10298,N_10063,N_10045);
or U10299 (N_10299,N_10041,N_10160);
or U10300 (N_10300,N_10080,N_10041);
xnor U10301 (N_10301,N_10153,N_10093);
and U10302 (N_10302,N_10084,N_10078);
nor U10303 (N_10303,N_10096,N_10132);
and U10304 (N_10304,N_10089,N_10040);
nor U10305 (N_10305,N_10176,N_10046);
nor U10306 (N_10306,N_10058,N_10153);
and U10307 (N_10307,N_10047,N_10088);
nor U10308 (N_10308,N_10071,N_10059);
xnor U10309 (N_10309,N_10018,N_10032);
nand U10310 (N_10310,N_10138,N_10161);
nand U10311 (N_10311,N_10143,N_10008);
or U10312 (N_10312,N_10007,N_10178);
and U10313 (N_10313,N_10117,N_10075);
xnor U10314 (N_10314,N_10162,N_10072);
and U10315 (N_10315,N_10087,N_10059);
nand U10316 (N_10316,N_10069,N_10058);
xor U10317 (N_10317,N_10075,N_10181);
nand U10318 (N_10318,N_10033,N_10120);
and U10319 (N_10319,N_10102,N_10016);
nand U10320 (N_10320,N_10173,N_10125);
nor U10321 (N_10321,N_10072,N_10083);
nand U10322 (N_10322,N_10180,N_10083);
nand U10323 (N_10323,N_10047,N_10050);
xor U10324 (N_10324,N_10136,N_10009);
or U10325 (N_10325,N_10017,N_10025);
xor U10326 (N_10326,N_10116,N_10198);
nor U10327 (N_10327,N_10138,N_10137);
or U10328 (N_10328,N_10109,N_10166);
or U10329 (N_10329,N_10142,N_10123);
and U10330 (N_10330,N_10089,N_10077);
or U10331 (N_10331,N_10021,N_10105);
nor U10332 (N_10332,N_10130,N_10141);
and U10333 (N_10333,N_10157,N_10061);
or U10334 (N_10334,N_10170,N_10058);
nand U10335 (N_10335,N_10120,N_10161);
and U10336 (N_10336,N_10144,N_10011);
and U10337 (N_10337,N_10186,N_10156);
xnor U10338 (N_10338,N_10036,N_10042);
and U10339 (N_10339,N_10000,N_10198);
xor U10340 (N_10340,N_10001,N_10148);
nor U10341 (N_10341,N_10015,N_10004);
and U10342 (N_10342,N_10119,N_10116);
and U10343 (N_10343,N_10024,N_10156);
or U10344 (N_10344,N_10149,N_10098);
xor U10345 (N_10345,N_10082,N_10018);
or U10346 (N_10346,N_10153,N_10122);
or U10347 (N_10347,N_10186,N_10122);
xor U10348 (N_10348,N_10055,N_10030);
xor U10349 (N_10349,N_10008,N_10014);
and U10350 (N_10350,N_10199,N_10108);
and U10351 (N_10351,N_10031,N_10035);
nor U10352 (N_10352,N_10146,N_10198);
nand U10353 (N_10353,N_10134,N_10174);
and U10354 (N_10354,N_10087,N_10064);
nor U10355 (N_10355,N_10133,N_10071);
and U10356 (N_10356,N_10133,N_10088);
nor U10357 (N_10357,N_10159,N_10003);
nand U10358 (N_10358,N_10069,N_10183);
nand U10359 (N_10359,N_10190,N_10028);
nor U10360 (N_10360,N_10174,N_10197);
nor U10361 (N_10361,N_10186,N_10039);
nand U10362 (N_10362,N_10136,N_10170);
and U10363 (N_10363,N_10114,N_10095);
or U10364 (N_10364,N_10056,N_10062);
or U10365 (N_10365,N_10163,N_10064);
nor U10366 (N_10366,N_10041,N_10103);
nand U10367 (N_10367,N_10084,N_10199);
xor U10368 (N_10368,N_10014,N_10154);
xor U10369 (N_10369,N_10132,N_10146);
and U10370 (N_10370,N_10116,N_10064);
xnor U10371 (N_10371,N_10098,N_10143);
nor U10372 (N_10372,N_10118,N_10084);
or U10373 (N_10373,N_10008,N_10081);
xor U10374 (N_10374,N_10002,N_10027);
or U10375 (N_10375,N_10068,N_10021);
nor U10376 (N_10376,N_10055,N_10147);
or U10377 (N_10377,N_10068,N_10029);
nand U10378 (N_10378,N_10186,N_10133);
nor U10379 (N_10379,N_10047,N_10086);
nand U10380 (N_10380,N_10190,N_10120);
and U10381 (N_10381,N_10183,N_10001);
xnor U10382 (N_10382,N_10147,N_10068);
xnor U10383 (N_10383,N_10010,N_10051);
nor U10384 (N_10384,N_10047,N_10040);
xor U10385 (N_10385,N_10124,N_10117);
xnor U10386 (N_10386,N_10092,N_10191);
or U10387 (N_10387,N_10034,N_10163);
or U10388 (N_10388,N_10016,N_10155);
and U10389 (N_10389,N_10028,N_10183);
xor U10390 (N_10390,N_10193,N_10187);
or U10391 (N_10391,N_10130,N_10163);
nor U10392 (N_10392,N_10098,N_10030);
nand U10393 (N_10393,N_10136,N_10035);
nand U10394 (N_10394,N_10045,N_10113);
and U10395 (N_10395,N_10135,N_10143);
nand U10396 (N_10396,N_10086,N_10009);
and U10397 (N_10397,N_10022,N_10090);
or U10398 (N_10398,N_10150,N_10035);
and U10399 (N_10399,N_10119,N_10088);
nor U10400 (N_10400,N_10251,N_10329);
or U10401 (N_10401,N_10342,N_10341);
nor U10402 (N_10402,N_10252,N_10356);
nor U10403 (N_10403,N_10264,N_10316);
nand U10404 (N_10404,N_10302,N_10399);
nor U10405 (N_10405,N_10398,N_10333);
and U10406 (N_10406,N_10358,N_10366);
and U10407 (N_10407,N_10339,N_10325);
nor U10408 (N_10408,N_10204,N_10234);
nand U10409 (N_10409,N_10269,N_10337);
or U10410 (N_10410,N_10382,N_10393);
xnor U10411 (N_10411,N_10321,N_10216);
and U10412 (N_10412,N_10267,N_10281);
and U10413 (N_10413,N_10298,N_10351);
nand U10414 (N_10414,N_10312,N_10215);
nand U10415 (N_10415,N_10219,N_10328);
or U10416 (N_10416,N_10282,N_10392);
xor U10417 (N_10417,N_10353,N_10305);
and U10418 (N_10418,N_10364,N_10313);
xor U10419 (N_10419,N_10306,N_10285);
nor U10420 (N_10420,N_10370,N_10209);
and U10421 (N_10421,N_10287,N_10304);
xnor U10422 (N_10422,N_10248,N_10318);
xor U10423 (N_10423,N_10231,N_10297);
nand U10424 (N_10424,N_10327,N_10268);
and U10425 (N_10425,N_10319,N_10386);
or U10426 (N_10426,N_10324,N_10389);
xnor U10427 (N_10427,N_10273,N_10322);
and U10428 (N_10428,N_10228,N_10238);
or U10429 (N_10429,N_10368,N_10373);
nor U10430 (N_10430,N_10288,N_10348);
xor U10431 (N_10431,N_10245,N_10291);
or U10432 (N_10432,N_10253,N_10380);
or U10433 (N_10433,N_10246,N_10263);
or U10434 (N_10434,N_10222,N_10289);
nand U10435 (N_10435,N_10229,N_10378);
and U10436 (N_10436,N_10295,N_10284);
nand U10437 (N_10437,N_10354,N_10256);
xor U10438 (N_10438,N_10210,N_10332);
and U10439 (N_10439,N_10331,N_10375);
nor U10440 (N_10440,N_10343,N_10395);
and U10441 (N_10441,N_10236,N_10275);
and U10442 (N_10442,N_10286,N_10349);
nor U10443 (N_10443,N_10235,N_10243);
nor U10444 (N_10444,N_10292,N_10227);
and U10445 (N_10445,N_10369,N_10213);
nand U10446 (N_10446,N_10359,N_10385);
and U10447 (N_10447,N_10315,N_10277);
or U10448 (N_10448,N_10218,N_10326);
and U10449 (N_10449,N_10266,N_10347);
or U10450 (N_10450,N_10272,N_10224);
nand U10451 (N_10451,N_10360,N_10207);
nor U10452 (N_10452,N_10240,N_10361);
and U10453 (N_10453,N_10221,N_10350);
nor U10454 (N_10454,N_10271,N_10390);
xor U10455 (N_10455,N_10241,N_10377);
or U10456 (N_10456,N_10344,N_10391);
and U10457 (N_10457,N_10239,N_10371);
nand U10458 (N_10458,N_10244,N_10279);
xor U10459 (N_10459,N_10363,N_10340);
xnor U10460 (N_10460,N_10345,N_10294);
or U10461 (N_10461,N_10293,N_10346);
or U10462 (N_10462,N_10396,N_10205);
and U10463 (N_10463,N_10320,N_10250);
xnor U10464 (N_10464,N_10365,N_10274);
and U10465 (N_10465,N_10230,N_10307);
and U10466 (N_10466,N_10372,N_10379);
or U10467 (N_10467,N_10384,N_10257);
nor U10468 (N_10468,N_10362,N_10374);
and U10469 (N_10469,N_10311,N_10352);
xnor U10470 (N_10470,N_10381,N_10397);
nand U10471 (N_10471,N_10336,N_10265);
and U10472 (N_10472,N_10330,N_10203);
xor U10473 (N_10473,N_10283,N_10309);
nor U10474 (N_10474,N_10208,N_10367);
nor U10475 (N_10475,N_10255,N_10262);
and U10476 (N_10476,N_10394,N_10220);
xnor U10477 (N_10477,N_10387,N_10290);
xor U10478 (N_10478,N_10254,N_10299);
nand U10479 (N_10479,N_10383,N_10249);
and U10480 (N_10480,N_10357,N_10301);
nand U10481 (N_10481,N_10226,N_10376);
or U10482 (N_10482,N_10247,N_10261);
nor U10483 (N_10483,N_10237,N_10300);
nand U10484 (N_10484,N_10323,N_10296);
and U10485 (N_10485,N_10278,N_10260);
and U10486 (N_10486,N_10334,N_10314);
nand U10487 (N_10487,N_10225,N_10388);
nor U10488 (N_10488,N_10310,N_10233);
nand U10489 (N_10489,N_10338,N_10280);
nor U10490 (N_10490,N_10355,N_10223);
and U10491 (N_10491,N_10214,N_10200);
xnor U10492 (N_10492,N_10212,N_10317);
nand U10493 (N_10493,N_10206,N_10259);
xnor U10494 (N_10494,N_10211,N_10270);
nand U10495 (N_10495,N_10242,N_10232);
and U10496 (N_10496,N_10258,N_10335);
xor U10497 (N_10497,N_10202,N_10276);
nand U10498 (N_10498,N_10308,N_10201);
or U10499 (N_10499,N_10303,N_10217);
nor U10500 (N_10500,N_10209,N_10376);
or U10501 (N_10501,N_10300,N_10251);
and U10502 (N_10502,N_10394,N_10313);
nand U10503 (N_10503,N_10304,N_10316);
nand U10504 (N_10504,N_10210,N_10253);
nor U10505 (N_10505,N_10331,N_10275);
nand U10506 (N_10506,N_10274,N_10251);
xnor U10507 (N_10507,N_10212,N_10260);
nor U10508 (N_10508,N_10362,N_10213);
nand U10509 (N_10509,N_10359,N_10290);
or U10510 (N_10510,N_10258,N_10251);
or U10511 (N_10511,N_10298,N_10311);
xor U10512 (N_10512,N_10381,N_10309);
and U10513 (N_10513,N_10247,N_10370);
or U10514 (N_10514,N_10268,N_10394);
and U10515 (N_10515,N_10309,N_10322);
or U10516 (N_10516,N_10394,N_10281);
nand U10517 (N_10517,N_10332,N_10279);
nand U10518 (N_10518,N_10222,N_10298);
or U10519 (N_10519,N_10359,N_10238);
xnor U10520 (N_10520,N_10356,N_10390);
and U10521 (N_10521,N_10350,N_10342);
xnor U10522 (N_10522,N_10289,N_10309);
or U10523 (N_10523,N_10336,N_10235);
nor U10524 (N_10524,N_10377,N_10293);
xor U10525 (N_10525,N_10201,N_10206);
and U10526 (N_10526,N_10265,N_10219);
and U10527 (N_10527,N_10223,N_10314);
nor U10528 (N_10528,N_10306,N_10329);
or U10529 (N_10529,N_10258,N_10294);
or U10530 (N_10530,N_10326,N_10288);
xor U10531 (N_10531,N_10322,N_10372);
nand U10532 (N_10532,N_10398,N_10355);
nand U10533 (N_10533,N_10377,N_10267);
nor U10534 (N_10534,N_10339,N_10368);
nor U10535 (N_10535,N_10335,N_10257);
xnor U10536 (N_10536,N_10344,N_10225);
or U10537 (N_10537,N_10390,N_10398);
nand U10538 (N_10538,N_10378,N_10367);
xor U10539 (N_10539,N_10397,N_10331);
and U10540 (N_10540,N_10288,N_10223);
nand U10541 (N_10541,N_10349,N_10206);
nor U10542 (N_10542,N_10326,N_10327);
xnor U10543 (N_10543,N_10302,N_10348);
xor U10544 (N_10544,N_10389,N_10298);
and U10545 (N_10545,N_10355,N_10245);
nor U10546 (N_10546,N_10316,N_10393);
or U10547 (N_10547,N_10377,N_10341);
or U10548 (N_10548,N_10386,N_10331);
xor U10549 (N_10549,N_10393,N_10360);
xnor U10550 (N_10550,N_10307,N_10272);
xnor U10551 (N_10551,N_10235,N_10329);
nor U10552 (N_10552,N_10226,N_10389);
xor U10553 (N_10553,N_10322,N_10304);
or U10554 (N_10554,N_10277,N_10302);
or U10555 (N_10555,N_10340,N_10202);
xnor U10556 (N_10556,N_10270,N_10210);
nor U10557 (N_10557,N_10368,N_10388);
nor U10558 (N_10558,N_10233,N_10313);
or U10559 (N_10559,N_10287,N_10319);
nand U10560 (N_10560,N_10306,N_10294);
nand U10561 (N_10561,N_10203,N_10219);
nand U10562 (N_10562,N_10338,N_10347);
or U10563 (N_10563,N_10213,N_10251);
or U10564 (N_10564,N_10245,N_10304);
or U10565 (N_10565,N_10260,N_10344);
nor U10566 (N_10566,N_10365,N_10347);
nor U10567 (N_10567,N_10339,N_10343);
nor U10568 (N_10568,N_10242,N_10323);
xnor U10569 (N_10569,N_10357,N_10370);
xnor U10570 (N_10570,N_10354,N_10297);
nand U10571 (N_10571,N_10303,N_10293);
or U10572 (N_10572,N_10350,N_10232);
nand U10573 (N_10573,N_10219,N_10271);
and U10574 (N_10574,N_10242,N_10259);
and U10575 (N_10575,N_10205,N_10258);
nand U10576 (N_10576,N_10388,N_10362);
and U10577 (N_10577,N_10380,N_10262);
and U10578 (N_10578,N_10237,N_10259);
and U10579 (N_10579,N_10356,N_10318);
nand U10580 (N_10580,N_10248,N_10252);
xnor U10581 (N_10581,N_10280,N_10383);
and U10582 (N_10582,N_10362,N_10346);
nand U10583 (N_10583,N_10259,N_10240);
nor U10584 (N_10584,N_10221,N_10228);
or U10585 (N_10585,N_10300,N_10293);
and U10586 (N_10586,N_10396,N_10296);
and U10587 (N_10587,N_10277,N_10259);
nor U10588 (N_10588,N_10311,N_10354);
or U10589 (N_10589,N_10293,N_10399);
and U10590 (N_10590,N_10227,N_10276);
or U10591 (N_10591,N_10300,N_10232);
and U10592 (N_10592,N_10279,N_10371);
and U10593 (N_10593,N_10242,N_10251);
and U10594 (N_10594,N_10201,N_10383);
nor U10595 (N_10595,N_10256,N_10319);
nor U10596 (N_10596,N_10345,N_10334);
nand U10597 (N_10597,N_10391,N_10357);
nand U10598 (N_10598,N_10373,N_10248);
nor U10599 (N_10599,N_10218,N_10250);
nor U10600 (N_10600,N_10460,N_10523);
xor U10601 (N_10601,N_10595,N_10445);
xnor U10602 (N_10602,N_10512,N_10453);
nand U10603 (N_10603,N_10454,N_10412);
xor U10604 (N_10604,N_10480,N_10591);
or U10605 (N_10605,N_10559,N_10515);
or U10606 (N_10606,N_10543,N_10463);
nor U10607 (N_10607,N_10528,N_10501);
or U10608 (N_10608,N_10420,N_10503);
and U10609 (N_10609,N_10549,N_10527);
nand U10610 (N_10610,N_10592,N_10487);
xnor U10611 (N_10611,N_10500,N_10536);
xor U10612 (N_10612,N_10579,N_10430);
nand U10613 (N_10613,N_10552,N_10587);
and U10614 (N_10614,N_10581,N_10423);
nand U10615 (N_10615,N_10493,N_10477);
and U10616 (N_10616,N_10535,N_10583);
or U10617 (N_10617,N_10472,N_10404);
xor U10618 (N_10618,N_10498,N_10400);
or U10619 (N_10619,N_10529,N_10506);
nor U10620 (N_10620,N_10599,N_10433);
nor U10621 (N_10621,N_10418,N_10458);
nand U10622 (N_10622,N_10546,N_10469);
xor U10623 (N_10623,N_10538,N_10462);
nor U10624 (N_10624,N_10438,N_10588);
xnor U10625 (N_10625,N_10491,N_10516);
xnor U10626 (N_10626,N_10513,N_10473);
xnor U10627 (N_10627,N_10571,N_10451);
xnor U10628 (N_10628,N_10570,N_10428);
xnor U10629 (N_10629,N_10402,N_10470);
xor U10630 (N_10630,N_10578,N_10439);
nand U10631 (N_10631,N_10505,N_10432);
nand U10632 (N_10632,N_10422,N_10408);
nor U10633 (N_10633,N_10490,N_10568);
and U10634 (N_10634,N_10586,N_10457);
xnor U10635 (N_10635,N_10403,N_10514);
or U10636 (N_10636,N_10424,N_10577);
xnor U10637 (N_10637,N_10496,N_10449);
or U10638 (N_10638,N_10455,N_10524);
and U10639 (N_10639,N_10476,N_10541);
and U10640 (N_10640,N_10589,N_10479);
nand U10641 (N_10641,N_10532,N_10431);
nand U10642 (N_10642,N_10556,N_10567);
or U10643 (N_10643,N_10485,N_10413);
or U10644 (N_10644,N_10450,N_10427);
nand U10645 (N_10645,N_10594,N_10533);
xnor U10646 (N_10646,N_10411,N_10415);
nor U10647 (N_10647,N_10585,N_10459);
nor U10648 (N_10648,N_10560,N_10444);
and U10649 (N_10649,N_10530,N_10509);
or U10650 (N_10650,N_10573,N_10526);
nor U10651 (N_10651,N_10522,N_10426);
nor U10652 (N_10652,N_10537,N_10575);
or U10653 (N_10653,N_10484,N_10547);
nor U10654 (N_10654,N_10558,N_10507);
or U10655 (N_10655,N_10414,N_10421);
or U10656 (N_10656,N_10553,N_10405);
and U10657 (N_10657,N_10499,N_10434);
nor U10658 (N_10658,N_10483,N_10443);
xnor U10659 (N_10659,N_10566,N_10584);
nand U10660 (N_10660,N_10486,N_10540);
and U10661 (N_10661,N_10417,N_10401);
and U10662 (N_10662,N_10545,N_10593);
or U10663 (N_10663,N_10442,N_10429);
and U10664 (N_10664,N_10466,N_10569);
nand U10665 (N_10665,N_10416,N_10474);
nand U10666 (N_10666,N_10576,N_10539);
and U10667 (N_10667,N_10557,N_10452);
nand U10668 (N_10668,N_10517,N_10468);
and U10669 (N_10669,N_10489,N_10488);
and U10670 (N_10670,N_10520,N_10465);
and U10671 (N_10671,N_10437,N_10531);
or U10672 (N_10672,N_10521,N_10436);
nand U10673 (N_10673,N_10448,N_10598);
and U10674 (N_10674,N_10542,N_10482);
and U10675 (N_10675,N_10525,N_10582);
nand U10676 (N_10676,N_10502,N_10478);
or U10677 (N_10677,N_10572,N_10441);
or U10678 (N_10678,N_10406,N_10467);
and U10679 (N_10679,N_10511,N_10596);
xor U10680 (N_10680,N_10407,N_10504);
nand U10681 (N_10681,N_10508,N_10446);
xor U10682 (N_10682,N_10492,N_10475);
or U10683 (N_10683,N_10534,N_10456);
and U10684 (N_10684,N_10561,N_10554);
xnor U10685 (N_10685,N_10574,N_10580);
xnor U10686 (N_10686,N_10564,N_10519);
and U10687 (N_10687,N_10435,N_10481);
nand U10688 (N_10688,N_10471,N_10440);
nor U10689 (N_10689,N_10425,N_10447);
and U10690 (N_10690,N_10464,N_10518);
or U10691 (N_10691,N_10562,N_10497);
xor U10692 (N_10692,N_10409,N_10555);
nand U10693 (N_10693,N_10551,N_10565);
or U10694 (N_10694,N_10494,N_10597);
xnor U10695 (N_10695,N_10544,N_10550);
nand U10696 (N_10696,N_10510,N_10590);
nor U10697 (N_10697,N_10410,N_10461);
or U10698 (N_10698,N_10548,N_10419);
nand U10699 (N_10699,N_10495,N_10563);
nand U10700 (N_10700,N_10452,N_10422);
nand U10701 (N_10701,N_10489,N_10490);
xnor U10702 (N_10702,N_10491,N_10441);
xor U10703 (N_10703,N_10532,N_10569);
and U10704 (N_10704,N_10420,N_10501);
and U10705 (N_10705,N_10524,N_10492);
xor U10706 (N_10706,N_10407,N_10400);
and U10707 (N_10707,N_10413,N_10534);
xor U10708 (N_10708,N_10581,N_10430);
xor U10709 (N_10709,N_10590,N_10453);
and U10710 (N_10710,N_10414,N_10571);
xnor U10711 (N_10711,N_10482,N_10551);
or U10712 (N_10712,N_10471,N_10595);
nand U10713 (N_10713,N_10481,N_10528);
nor U10714 (N_10714,N_10591,N_10438);
nand U10715 (N_10715,N_10519,N_10572);
nand U10716 (N_10716,N_10411,N_10524);
nand U10717 (N_10717,N_10446,N_10443);
and U10718 (N_10718,N_10409,N_10576);
nor U10719 (N_10719,N_10586,N_10598);
nand U10720 (N_10720,N_10522,N_10525);
xor U10721 (N_10721,N_10577,N_10440);
and U10722 (N_10722,N_10502,N_10578);
nor U10723 (N_10723,N_10483,N_10409);
nor U10724 (N_10724,N_10568,N_10558);
or U10725 (N_10725,N_10491,N_10592);
or U10726 (N_10726,N_10457,N_10517);
and U10727 (N_10727,N_10533,N_10402);
nand U10728 (N_10728,N_10515,N_10528);
nor U10729 (N_10729,N_10532,N_10544);
xnor U10730 (N_10730,N_10515,N_10436);
or U10731 (N_10731,N_10451,N_10412);
and U10732 (N_10732,N_10430,N_10471);
and U10733 (N_10733,N_10454,N_10522);
nor U10734 (N_10734,N_10522,N_10533);
nor U10735 (N_10735,N_10514,N_10578);
and U10736 (N_10736,N_10522,N_10591);
nand U10737 (N_10737,N_10518,N_10489);
and U10738 (N_10738,N_10542,N_10585);
xor U10739 (N_10739,N_10498,N_10444);
xnor U10740 (N_10740,N_10582,N_10581);
and U10741 (N_10741,N_10471,N_10433);
xnor U10742 (N_10742,N_10463,N_10534);
xor U10743 (N_10743,N_10479,N_10410);
or U10744 (N_10744,N_10538,N_10490);
nand U10745 (N_10745,N_10448,N_10460);
and U10746 (N_10746,N_10403,N_10568);
or U10747 (N_10747,N_10464,N_10402);
nor U10748 (N_10748,N_10597,N_10421);
nand U10749 (N_10749,N_10546,N_10427);
nand U10750 (N_10750,N_10448,N_10455);
and U10751 (N_10751,N_10458,N_10467);
nand U10752 (N_10752,N_10442,N_10577);
nand U10753 (N_10753,N_10584,N_10535);
nor U10754 (N_10754,N_10507,N_10486);
and U10755 (N_10755,N_10466,N_10482);
and U10756 (N_10756,N_10577,N_10584);
nand U10757 (N_10757,N_10402,N_10510);
or U10758 (N_10758,N_10565,N_10486);
or U10759 (N_10759,N_10405,N_10429);
nand U10760 (N_10760,N_10461,N_10508);
and U10761 (N_10761,N_10407,N_10415);
and U10762 (N_10762,N_10564,N_10433);
xor U10763 (N_10763,N_10443,N_10547);
nand U10764 (N_10764,N_10467,N_10429);
nand U10765 (N_10765,N_10545,N_10436);
nand U10766 (N_10766,N_10594,N_10437);
xnor U10767 (N_10767,N_10560,N_10506);
nor U10768 (N_10768,N_10587,N_10499);
or U10769 (N_10769,N_10475,N_10409);
and U10770 (N_10770,N_10516,N_10465);
and U10771 (N_10771,N_10428,N_10542);
nor U10772 (N_10772,N_10560,N_10525);
nand U10773 (N_10773,N_10593,N_10462);
xor U10774 (N_10774,N_10504,N_10564);
and U10775 (N_10775,N_10490,N_10414);
or U10776 (N_10776,N_10528,N_10525);
or U10777 (N_10777,N_10558,N_10531);
or U10778 (N_10778,N_10583,N_10450);
or U10779 (N_10779,N_10488,N_10507);
or U10780 (N_10780,N_10414,N_10483);
or U10781 (N_10781,N_10520,N_10515);
xnor U10782 (N_10782,N_10445,N_10493);
or U10783 (N_10783,N_10570,N_10592);
nand U10784 (N_10784,N_10483,N_10570);
xnor U10785 (N_10785,N_10581,N_10537);
or U10786 (N_10786,N_10581,N_10431);
nand U10787 (N_10787,N_10541,N_10557);
nand U10788 (N_10788,N_10554,N_10541);
or U10789 (N_10789,N_10520,N_10564);
nor U10790 (N_10790,N_10467,N_10522);
nand U10791 (N_10791,N_10559,N_10581);
xnor U10792 (N_10792,N_10510,N_10447);
xnor U10793 (N_10793,N_10560,N_10546);
and U10794 (N_10794,N_10486,N_10525);
nand U10795 (N_10795,N_10587,N_10415);
nand U10796 (N_10796,N_10438,N_10472);
xnor U10797 (N_10797,N_10470,N_10443);
nor U10798 (N_10798,N_10567,N_10584);
nor U10799 (N_10799,N_10570,N_10400);
or U10800 (N_10800,N_10723,N_10604);
or U10801 (N_10801,N_10707,N_10748);
xor U10802 (N_10802,N_10743,N_10606);
nor U10803 (N_10803,N_10769,N_10720);
nand U10804 (N_10804,N_10662,N_10643);
nor U10805 (N_10805,N_10616,N_10760);
or U10806 (N_10806,N_10629,N_10749);
nor U10807 (N_10807,N_10763,N_10747);
xnor U10808 (N_10808,N_10703,N_10781);
xnor U10809 (N_10809,N_10766,N_10730);
xor U10810 (N_10810,N_10757,N_10799);
or U10811 (N_10811,N_10620,N_10729);
xor U10812 (N_10812,N_10665,N_10787);
or U10813 (N_10813,N_10671,N_10732);
and U10814 (N_10814,N_10696,N_10634);
nor U10815 (N_10815,N_10624,N_10704);
nor U10816 (N_10816,N_10794,N_10735);
nand U10817 (N_10817,N_10790,N_10608);
nor U10818 (N_10818,N_10652,N_10712);
nand U10819 (N_10819,N_10626,N_10650);
xnor U10820 (N_10820,N_10780,N_10728);
nand U10821 (N_10821,N_10654,N_10702);
or U10822 (N_10822,N_10685,N_10711);
or U10823 (N_10823,N_10689,N_10791);
nor U10824 (N_10824,N_10625,N_10687);
and U10825 (N_10825,N_10674,N_10614);
and U10826 (N_10826,N_10755,N_10644);
and U10827 (N_10827,N_10676,N_10758);
or U10828 (N_10828,N_10738,N_10611);
xor U10829 (N_10829,N_10661,N_10726);
nand U10830 (N_10830,N_10683,N_10772);
nand U10831 (N_10831,N_10601,N_10693);
or U10832 (N_10832,N_10713,N_10646);
nand U10833 (N_10833,N_10784,N_10767);
or U10834 (N_10834,N_10768,N_10668);
or U10835 (N_10835,N_10690,N_10754);
nand U10836 (N_10836,N_10714,N_10691);
xor U10837 (N_10837,N_10716,N_10797);
nand U10838 (N_10838,N_10649,N_10633);
or U10839 (N_10839,N_10778,N_10786);
xnor U10840 (N_10840,N_10655,N_10706);
nor U10841 (N_10841,N_10751,N_10752);
or U10842 (N_10842,N_10721,N_10637);
nor U10843 (N_10843,N_10621,N_10724);
nor U10844 (N_10844,N_10789,N_10619);
nand U10845 (N_10845,N_10651,N_10719);
xor U10846 (N_10846,N_10670,N_10793);
and U10847 (N_10847,N_10739,N_10648);
and U10848 (N_10848,N_10666,N_10770);
nand U10849 (N_10849,N_10737,N_10761);
nand U10850 (N_10850,N_10694,N_10656);
or U10851 (N_10851,N_10622,N_10605);
and U10852 (N_10852,N_10630,N_10672);
nand U10853 (N_10853,N_10765,N_10771);
nor U10854 (N_10854,N_10708,N_10725);
or U10855 (N_10855,N_10613,N_10684);
nand U10856 (N_10856,N_10779,N_10635);
nand U10857 (N_10857,N_10764,N_10612);
nor U10858 (N_10858,N_10653,N_10785);
xnor U10859 (N_10859,N_10688,N_10657);
and U10860 (N_10860,N_10618,N_10776);
xor U10861 (N_10861,N_10680,N_10673);
nand U10862 (N_10862,N_10627,N_10734);
or U10863 (N_10863,N_10699,N_10698);
or U10864 (N_10864,N_10742,N_10681);
or U10865 (N_10865,N_10715,N_10664);
nand U10866 (N_10866,N_10669,N_10609);
nand U10867 (N_10867,N_10733,N_10647);
and U10868 (N_10868,N_10756,N_10600);
or U10869 (N_10869,N_10659,N_10610);
nand U10870 (N_10870,N_10774,N_10603);
nor U10871 (N_10871,N_10745,N_10798);
xor U10872 (N_10872,N_10718,N_10727);
xor U10873 (N_10873,N_10640,N_10641);
xnor U10874 (N_10874,N_10788,N_10602);
or U10875 (N_10875,N_10692,N_10795);
nand U10876 (N_10876,N_10658,N_10638);
or U10877 (N_10877,N_10783,N_10645);
or U10878 (N_10878,N_10628,N_10736);
nand U10879 (N_10879,N_10660,N_10796);
nand U10880 (N_10880,N_10775,N_10678);
and U10881 (N_10881,N_10677,N_10617);
or U10882 (N_10882,N_10679,N_10615);
and U10883 (N_10883,N_10667,N_10762);
or U10884 (N_10884,N_10722,N_10695);
xor U10885 (N_10885,N_10682,N_10773);
xor U10886 (N_10886,N_10639,N_10709);
or U10887 (N_10887,N_10746,N_10686);
and U10888 (N_10888,N_10700,N_10675);
nand U10889 (N_10889,N_10753,N_10632);
and U10890 (N_10890,N_10782,N_10705);
xor U10891 (N_10891,N_10740,N_10642);
nor U10892 (N_10892,N_10744,N_10792);
and U10893 (N_10893,N_10741,N_10636);
nand U10894 (N_10894,N_10623,N_10701);
and U10895 (N_10895,N_10697,N_10777);
or U10896 (N_10896,N_10607,N_10631);
xnor U10897 (N_10897,N_10731,N_10710);
and U10898 (N_10898,N_10750,N_10759);
xor U10899 (N_10899,N_10717,N_10663);
and U10900 (N_10900,N_10752,N_10784);
nor U10901 (N_10901,N_10788,N_10622);
and U10902 (N_10902,N_10692,N_10617);
nor U10903 (N_10903,N_10731,N_10651);
xnor U10904 (N_10904,N_10788,N_10701);
xnor U10905 (N_10905,N_10792,N_10643);
nand U10906 (N_10906,N_10748,N_10776);
or U10907 (N_10907,N_10798,N_10722);
and U10908 (N_10908,N_10633,N_10756);
xor U10909 (N_10909,N_10689,N_10764);
nor U10910 (N_10910,N_10676,N_10631);
nor U10911 (N_10911,N_10695,N_10713);
or U10912 (N_10912,N_10683,N_10773);
nor U10913 (N_10913,N_10714,N_10737);
nand U10914 (N_10914,N_10796,N_10661);
or U10915 (N_10915,N_10783,N_10632);
nand U10916 (N_10916,N_10792,N_10630);
and U10917 (N_10917,N_10690,N_10654);
nand U10918 (N_10918,N_10666,N_10773);
nor U10919 (N_10919,N_10681,N_10787);
nand U10920 (N_10920,N_10646,N_10783);
or U10921 (N_10921,N_10637,N_10713);
nor U10922 (N_10922,N_10655,N_10686);
xnor U10923 (N_10923,N_10646,N_10679);
and U10924 (N_10924,N_10790,N_10687);
nor U10925 (N_10925,N_10693,N_10706);
or U10926 (N_10926,N_10632,N_10674);
xnor U10927 (N_10927,N_10731,N_10742);
nor U10928 (N_10928,N_10662,N_10741);
and U10929 (N_10929,N_10716,N_10625);
or U10930 (N_10930,N_10714,N_10634);
nor U10931 (N_10931,N_10653,N_10793);
nor U10932 (N_10932,N_10707,N_10703);
nand U10933 (N_10933,N_10651,N_10638);
and U10934 (N_10934,N_10712,N_10670);
and U10935 (N_10935,N_10621,N_10722);
xor U10936 (N_10936,N_10718,N_10659);
and U10937 (N_10937,N_10695,N_10778);
nor U10938 (N_10938,N_10603,N_10756);
xnor U10939 (N_10939,N_10627,N_10669);
nor U10940 (N_10940,N_10655,N_10737);
and U10941 (N_10941,N_10710,N_10691);
nand U10942 (N_10942,N_10607,N_10641);
and U10943 (N_10943,N_10677,N_10611);
or U10944 (N_10944,N_10653,N_10716);
or U10945 (N_10945,N_10674,N_10685);
and U10946 (N_10946,N_10637,N_10630);
and U10947 (N_10947,N_10782,N_10677);
or U10948 (N_10948,N_10796,N_10743);
xnor U10949 (N_10949,N_10636,N_10734);
or U10950 (N_10950,N_10694,N_10739);
nor U10951 (N_10951,N_10663,N_10724);
and U10952 (N_10952,N_10706,N_10617);
xnor U10953 (N_10953,N_10606,N_10755);
and U10954 (N_10954,N_10733,N_10627);
and U10955 (N_10955,N_10731,N_10627);
nor U10956 (N_10956,N_10757,N_10653);
or U10957 (N_10957,N_10667,N_10760);
xor U10958 (N_10958,N_10600,N_10617);
nor U10959 (N_10959,N_10653,N_10639);
nand U10960 (N_10960,N_10706,N_10699);
nand U10961 (N_10961,N_10609,N_10715);
and U10962 (N_10962,N_10603,N_10612);
nand U10963 (N_10963,N_10651,N_10771);
nor U10964 (N_10964,N_10649,N_10757);
xnor U10965 (N_10965,N_10713,N_10724);
nor U10966 (N_10966,N_10797,N_10719);
or U10967 (N_10967,N_10735,N_10722);
xor U10968 (N_10968,N_10655,N_10751);
nand U10969 (N_10969,N_10608,N_10709);
nand U10970 (N_10970,N_10784,N_10771);
nand U10971 (N_10971,N_10620,N_10635);
xnor U10972 (N_10972,N_10717,N_10675);
or U10973 (N_10973,N_10764,N_10659);
and U10974 (N_10974,N_10618,N_10777);
xnor U10975 (N_10975,N_10669,N_10780);
and U10976 (N_10976,N_10620,N_10709);
or U10977 (N_10977,N_10743,N_10626);
nor U10978 (N_10978,N_10786,N_10774);
xnor U10979 (N_10979,N_10797,N_10661);
nor U10980 (N_10980,N_10690,N_10731);
xnor U10981 (N_10981,N_10682,N_10701);
and U10982 (N_10982,N_10651,N_10637);
nor U10983 (N_10983,N_10762,N_10710);
nor U10984 (N_10984,N_10668,N_10649);
nand U10985 (N_10985,N_10691,N_10740);
and U10986 (N_10986,N_10603,N_10666);
or U10987 (N_10987,N_10778,N_10661);
or U10988 (N_10988,N_10648,N_10632);
xor U10989 (N_10989,N_10696,N_10742);
or U10990 (N_10990,N_10742,N_10734);
xor U10991 (N_10991,N_10771,N_10643);
and U10992 (N_10992,N_10731,N_10780);
nand U10993 (N_10993,N_10651,N_10799);
nor U10994 (N_10994,N_10663,N_10764);
and U10995 (N_10995,N_10637,N_10638);
xor U10996 (N_10996,N_10649,N_10752);
xor U10997 (N_10997,N_10652,N_10656);
or U10998 (N_10998,N_10621,N_10639);
xnor U10999 (N_10999,N_10697,N_10723);
xnor U11000 (N_11000,N_10823,N_10910);
nor U11001 (N_11001,N_10946,N_10940);
xnor U11002 (N_11002,N_10907,N_10949);
and U11003 (N_11003,N_10812,N_10869);
xnor U11004 (N_11004,N_10942,N_10830);
and U11005 (N_11005,N_10937,N_10825);
nor U11006 (N_11006,N_10847,N_10820);
nand U11007 (N_11007,N_10968,N_10906);
and U11008 (N_11008,N_10965,N_10880);
xor U11009 (N_11009,N_10894,N_10974);
and U11010 (N_11010,N_10809,N_10989);
or U11011 (N_11011,N_10994,N_10886);
xnor U11012 (N_11012,N_10851,N_10838);
or U11013 (N_11013,N_10859,N_10826);
and U11014 (N_11014,N_10842,N_10955);
and U11015 (N_11015,N_10899,N_10829);
and U11016 (N_11016,N_10996,N_10803);
and U11017 (N_11017,N_10818,N_10879);
or U11018 (N_11018,N_10944,N_10991);
or U11019 (N_11019,N_10952,N_10973);
nand U11020 (N_11020,N_10972,N_10885);
xnor U11021 (N_11021,N_10975,N_10927);
nor U11022 (N_11022,N_10961,N_10800);
nor U11023 (N_11023,N_10925,N_10987);
nand U11024 (N_11024,N_10922,N_10959);
or U11025 (N_11025,N_10941,N_10846);
or U11026 (N_11026,N_10900,N_10871);
and U11027 (N_11027,N_10856,N_10878);
and U11028 (N_11028,N_10870,N_10914);
nand U11029 (N_11029,N_10862,N_10898);
nand U11030 (N_11030,N_10836,N_10984);
and U11031 (N_11031,N_10930,N_10860);
or U11032 (N_11032,N_10837,N_10909);
nand U11033 (N_11033,N_10857,N_10916);
and U11034 (N_11034,N_10917,N_10971);
xnor U11035 (N_11035,N_10893,N_10938);
or U11036 (N_11036,N_10913,N_10883);
nand U11037 (N_11037,N_10806,N_10835);
nand U11038 (N_11038,N_10817,N_10978);
nand U11039 (N_11039,N_10892,N_10969);
and U11040 (N_11040,N_10874,N_10918);
or U11041 (N_11041,N_10924,N_10819);
nand U11042 (N_11042,N_10982,N_10811);
and U11043 (N_11043,N_10861,N_10936);
nand U11044 (N_11044,N_10888,N_10957);
or U11045 (N_11045,N_10902,N_10901);
or U11046 (N_11046,N_10866,N_10849);
or U11047 (N_11047,N_10943,N_10875);
or U11048 (N_11048,N_10889,N_10998);
nand U11049 (N_11049,N_10995,N_10802);
nor U11050 (N_11050,N_10990,N_10897);
nand U11051 (N_11051,N_10993,N_10980);
nand U11052 (N_11052,N_10976,N_10884);
nor U11053 (N_11053,N_10915,N_10841);
and U11054 (N_11054,N_10852,N_10945);
and U11055 (N_11055,N_10905,N_10810);
nand U11056 (N_11056,N_10853,N_10986);
and U11057 (N_11057,N_10815,N_10967);
nand U11058 (N_11058,N_10981,N_10950);
or U11059 (N_11059,N_10960,N_10822);
and U11060 (N_11060,N_10948,N_10843);
nor U11061 (N_11061,N_10921,N_10896);
nor U11062 (N_11062,N_10804,N_10963);
or U11063 (N_11063,N_10876,N_10992);
nand U11064 (N_11064,N_10887,N_10821);
and U11065 (N_11065,N_10947,N_10912);
nand U11066 (N_11066,N_10926,N_10813);
nor U11067 (N_11067,N_10904,N_10839);
or U11068 (N_11068,N_10873,N_10872);
or U11069 (N_11069,N_10816,N_10868);
or U11070 (N_11070,N_10919,N_10882);
and U11071 (N_11071,N_10855,N_10966);
and U11072 (N_11072,N_10833,N_10890);
xnor U11073 (N_11073,N_10977,N_10954);
nor U11074 (N_11074,N_10979,N_10958);
and U11075 (N_11075,N_10931,N_10805);
and U11076 (N_11076,N_10911,N_10848);
and U11077 (N_11077,N_10923,N_10863);
and U11078 (N_11078,N_10824,N_10908);
nor U11079 (N_11079,N_10932,N_10997);
nor U11080 (N_11080,N_10827,N_10985);
and U11081 (N_11081,N_10903,N_10939);
nor U11082 (N_11082,N_10934,N_10814);
nor U11083 (N_11083,N_10845,N_10970);
nor U11084 (N_11084,N_10867,N_10807);
and U11085 (N_11085,N_10850,N_10808);
nand U11086 (N_11086,N_10928,N_10832);
xnor U11087 (N_11087,N_10834,N_10999);
and U11088 (N_11088,N_10895,N_10854);
and U11089 (N_11089,N_10891,N_10844);
or U11090 (N_11090,N_10956,N_10831);
and U11091 (N_11091,N_10983,N_10935);
nand U11092 (N_11092,N_10964,N_10865);
or U11093 (N_11093,N_10951,N_10877);
xor U11094 (N_11094,N_10840,N_10929);
nand U11095 (N_11095,N_10953,N_10864);
or U11096 (N_11096,N_10933,N_10920);
nor U11097 (N_11097,N_10828,N_10881);
nor U11098 (N_11098,N_10858,N_10801);
and U11099 (N_11099,N_10962,N_10988);
xnor U11100 (N_11100,N_10926,N_10819);
and U11101 (N_11101,N_10944,N_10829);
nor U11102 (N_11102,N_10971,N_10842);
nor U11103 (N_11103,N_10834,N_10860);
or U11104 (N_11104,N_10834,N_10858);
nor U11105 (N_11105,N_10871,N_10844);
xor U11106 (N_11106,N_10814,N_10856);
and U11107 (N_11107,N_10878,N_10872);
nor U11108 (N_11108,N_10872,N_10809);
xnor U11109 (N_11109,N_10982,N_10997);
nor U11110 (N_11110,N_10859,N_10810);
nor U11111 (N_11111,N_10903,N_10857);
xor U11112 (N_11112,N_10840,N_10995);
and U11113 (N_11113,N_10948,N_10830);
and U11114 (N_11114,N_10922,N_10900);
nand U11115 (N_11115,N_10896,N_10855);
or U11116 (N_11116,N_10991,N_10970);
and U11117 (N_11117,N_10961,N_10938);
nand U11118 (N_11118,N_10904,N_10997);
xor U11119 (N_11119,N_10855,N_10882);
or U11120 (N_11120,N_10994,N_10893);
and U11121 (N_11121,N_10825,N_10987);
xnor U11122 (N_11122,N_10972,N_10822);
nor U11123 (N_11123,N_10993,N_10901);
xor U11124 (N_11124,N_10979,N_10977);
xor U11125 (N_11125,N_10966,N_10990);
and U11126 (N_11126,N_10810,N_10904);
nand U11127 (N_11127,N_10845,N_10899);
xor U11128 (N_11128,N_10952,N_10827);
and U11129 (N_11129,N_10835,N_10818);
and U11130 (N_11130,N_10844,N_10925);
nor U11131 (N_11131,N_10809,N_10833);
nor U11132 (N_11132,N_10875,N_10895);
xor U11133 (N_11133,N_10857,N_10806);
and U11134 (N_11134,N_10964,N_10950);
and U11135 (N_11135,N_10950,N_10958);
or U11136 (N_11136,N_10929,N_10879);
or U11137 (N_11137,N_10832,N_10950);
nand U11138 (N_11138,N_10843,N_10908);
xnor U11139 (N_11139,N_10805,N_10831);
or U11140 (N_11140,N_10831,N_10940);
nand U11141 (N_11141,N_10938,N_10937);
xor U11142 (N_11142,N_10898,N_10912);
and U11143 (N_11143,N_10959,N_10990);
nor U11144 (N_11144,N_10876,N_10849);
and U11145 (N_11145,N_10896,N_10895);
nand U11146 (N_11146,N_10887,N_10986);
nand U11147 (N_11147,N_10983,N_10976);
or U11148 (N_11148,N_10819,N_10822);
and U11149 (N_11149,N_10930,N_10919);
and U11150 (N_11150,N_10963,N_10885);
nor U11151 (N_11151,N_10869,N_10856);
or U11152 (N_11152,N_10963,N_10934);
or U11153 (N_11153,N_10971,N_10862);
and U11154 (N_11154,N_10844,N_10956);
nor U11155 (N_11155,N_10866,N_10938);
xor U11156 (N_11156,N_10898,N_10945);
or U11157 (N_11157,N_10899,N_10906);
xnor U11158 (N_11158,N_10952,N_10988);
and U11159 (N_11159,N_10971,N_10927);
and U11160 (N_11160,N_10993,N_10900);
or U11161 (N_11161,N_10874,N_10961);
nor U11162 (N_11162,N_10944,N_10900);
nor U11163 (N_11163,N_10976,N_10923);
nand U11164 (N_11164,N_10892,N_10902);
xor U11165 (N_11165,N_10908,N_10930);
nor U11166 (N_11166,N_10925,N_10941);
and U11167 (N_11167,N_10854,N_10945);
and U11168 (N_11168,N_10878,N_10933);
nand U11169 (N_11169,N_10949,N_10936);
xnor U11170 (N_11170,N_10884,N_10975);
or U11171 (N_11171,N_10911,N_10912);
nor U11172 (N_11172,N_10890,N_10845);
and U11173 (N_11173,N_10897,N_10931);
nor U11174 (N_11174,N_10971,N_10980);
nand U11175 (N_11175,N_10938,N_10843);
nor U11176 (N_11176,N_10806,N_10866);
xnor U11177 (N_11177,N_10837,N_10919);
or U11178 (N_11178,N_10811,N_10909);
xor U11179 (N_11179,N_10946,N_10927);
and U11180 (N_11180,N_10948,N_10803);
or U11181 (N_11181,N_10995,N_10870);
or U11182 (N_11182,N_10943,N_10919);
and U11183 (N_11183,N_10948,N_10847);
nor U11184 (N_11184,N_10831,N_10907);
and U11185 (N_11185,N_10924,N_10860);
nor U11186 (N_11186,N_10930,N_10986);
and U11187 (N_11187,N_10828,N_10818);
and U11188 (N_11188,N_10872,N_10835);
and U11189 (N_11189,N_10959,N_10901);
and U11190 (N_11190,N_10891,N_10883);
and U11191 (N_11191,N_10987,N_10947);
xnor U11192 (N_11192,N_10916,N_10930);
nand U11193 (N_11193,N_10815,N_10888);
xnor U11194 (N_11194,N_10966,N_10875);
nor U11195 (N_11195,N_10963,N_10959);
nand U11196 (N_11196,N_10924,N_10961);
and U11197 (N_11197,N_10935,N_10826);
or U11198 (N_11198,N_10868,N_10911);
xor U11199 (N_11199,N_10941,N_10994);
or U11200 (N_11200,N_11173,N_11144);
and U11201 (N_11201,N_11057,N_11160);
nand U11202 (N_11202,N_11053,N_11073);
and U11203 (N_11203,N_11190,N_11185);
nand U11204 (N_11204,N_11157,N_11016);
nand U11205 (N_11205,N_11197,N_11076);
nand U11206 (N_11206,N_11028,N_11067);
xnor U11207 (N_11207,N_11043,N_11049);
nor U11208 (N_11208,N_11129,N_11145);
or U11209 (N_11209,N_11105,N_11100);
nand U11210 (N_11210,N_11163,N_11079);
xor U11211 (N_11211,N_11065,N_11095);
nor U11212 (N_11212,N_11027,N_11121);
xor U11213 (N_11213,N_11114,N_11112);
and U11214 (N_11214,N_11050,N_11060);
nand U11215 (N_11215,N_11153,N_11124);
nor U11216 (N_11216,N_11137,N_11098);
xnor U11217 (N_11217,N_11007,N_11178);
or U11218 (N_11218,N_11054,N_11110);
and U11219 (N_11219,N_11139,N_11142);
nand U11220 (N_11220,N_11196,N_11046);
or U11221 (N_11221,N_11063,N_11096);
and U11222 (N_11222,N_11059,N_11188);
or U11223 (N_11223,N_11187,N_11193);
xor U11224 (N_11224,N_11039,N_11094);
and U11225 (N_11225,N_11198,N_11044);
nand U11226 (N_11226,N_11015,N_11131);
nor U11227 (N_11227,N_11146,N_11074);
or U11228 (N_11228,N_11170,N_11070);
and U11229 (N_11229,N_11075,N_11014);
xnor U11230 (N_11230,N_11152,N_11017);
nor U11231 (N_11231,N_11162,N_11036);
nand U11232 (N_11232,N_11001,N_11056);
nand U11233 (N_11233,N_11021,N_11080);
nand U11234 (N_11234,N_11109,N_11026);
xor U11235 (N_11235,N_11130,N_11104);
nand U11236 (N_11236,N_11072,N_11004);
nand U11237 (N_11237,N_11180,N_11090);
or U11238 (N_11238,N_11133,N_11179);
xnor U11239 (N_11239,N_11011,N_11003);
nor U11240 (N_11240,N_11199,N_11089);
nor U11241 (N_11241,N_11158,N_11033);
or U11242 (N_11242,N_11102,N_11009);
nand U11243 (N_11243,N_11052,N_11078);
and U11244 (N_11244,N_11062,N_11136);
nand U11245 (N_11245,N_11000,N_11111);
or U11246 (N_11246,N_11022,N_11002);
xnor U11247 (N_11247,N_11058,N_11183);
or U11248 (N_11248,N_11025,N_11101);
nor U11249 (N_11249,N_11154,N_11168);
and U11250 (N_11250,N_11127,N_11055);
and U11251 (N_11251,N_11172,N_11051);
xnor U11252 (N_11252,N_11176,N_11149);
and U11253 (N_11253,N_11069,N_11126);
and U11254 (N_11254,N_11135,N_11161);
xor U11255 (N_11255,N_11119,N_11181);
and U11256 (N_11256,N_11010,N_11138);
xnor U11257 (N_11257,N_11159,N_11174);
and U11258 (N_11258,N_11038,N_11165);
or U11259 (N_11259,N_11031,N_11115);
nor U11260 (N_11260,N_11045,N_11141);
nand U11261 (N_11261,N_11186,N_11113);
nor U11262 (N_11262,N_11128,N_11191);
nor U11263 (N_11263,N_11156,N_11164);
xnor U11264 (N_11264,N_11171,N_11082);
xnor U11265 (N_11265,N_11061,N_11013);
nor U11266 (N_11266,N_11192,N_11019);
nand U11267 (N_11267,N_11194,N_11150);
nor U11268 (N_11268,N_11106,N_11143);
nor U11269 (N_11269,N_11108,N_11118);
xor U11270 (N_11270,N_11068,N_11008);
and U11271 (N_11271,N_11132,N_11099);
nor U11272 (N_11272,N_11122,N_11120);
nand U11273 (N_11273,N_11084,N_11117);
xor U11274 (N_11274,N_11155,N_11103);
nor U11275 (N_11275,N_11125,N_11047);
nand U11276 (N_11276,N_11035,N_11097);
and U11277 (N_11277,N_11184,N_11140);
or U11278 (N_11278,N_11085,N_11147);
or U11279 (N_11279,N_11029,N_11048);
or U11280 (N_11280,N_11189,N_11166);
nand U11281 (N_11281,N_11169,N_11081);
and U11282 (N_11282,N_11123,N_11195);
or U11283 (N_11283,N_11034,N_11182);
and U11284 (N_11284,N_11091,N_11037);
nor U11285 (N_11285,N_11167,N_11148);
or U11286 (N_11286,N_11071,N_11116);
and U11287 (N_11287,N_11107,N_11151);
nor U11288 (N_11288,N_11066,N_11020);
nor U11289 (N_11289,N_11024,N_11093);
xnor U11290 (N_11290,N_11042,N_11040);
nor U11291 (N_11291,N_11064,N_11012);
nor U11292 (N_11292,N_11041,N_11087);
and U11293 (N_11293,N_11018,N_11032);
nand U11294 (N_11294,N_11086,N_11177);
nor U11295 (N_11295,N_11088,N_11083);
nand U11296 (N_11296,N_11134,N_11092);
xnor U11297 (N_11297,N_11175,N_11006);
nor U11298 (N_11298,N_11023,N_11077);
nor U11299 (N_11299,N_11005,N_11030);
or U11300 (N_11300,N_11194,N_11055);
xor U11301 (N_11301,N_11037,N_11157);
nand U11302 (N_11302,N_11088,N_11102);
xnor U11303 (N_11303,N_11187,N_11111);
and U11304 (N_11304,N_11125,N_11166);
or U11305 (N_11305,N_11007,N_11106);
and U11306 (N_11306,N_11005,N_11089);
nand U11307 (N_11307,N_11118,N_11138);
nor U11308 (N_11308,N_11058,N_11087);
or U11309 (N_11309,N_11049,N_11009);
and U11310 (N_11310,N_11174,N_11005);
nand U11311 (N_11311,N_11055,N_11145);
or U11312 (N_11312,N_11138,N_11107);
nor U11313 (N_11313,N_11113,N_11059);
nor U11314 (N_11314,N_11107,N_11124);
xor U11315 (N_11315,N_11025,N_11008);
or U11316 (N_11316,N_11039,N_11020);
or U11317 (N_11317,N_11166,N_11080);
nor U11318 (N_11318,N_11161,N_11192);
xor U11319 (N_11319,N_11139,N_11065);
xnor U11320 (N_11320,N_11034,N_11097);
xor U11321 (N_11321,N_11045,N_11136);
or U11322 (N_11322,N_11192,N_11024);
nor U11323 (N_11323,N_11179,N_11074);
or U11324 (N_11324,N_11052,N_11174);
nand U11325 (N_11325,N_11119,N_11040);
nand U11326 (N_11326,N_11129,N_11037);
nand U11327 (N_11327,N_11049,N_11013);
nand U11328 (N_11328,N_11079,N_11106);
xor U11329 (N_11329,N_11190,N_11064);
or U11330 (N_11330,N_11180,N_11171);
xor U11331 (N_11331,N_11186,N_11011);
nand U11332 (N_11332,N_11055,N_11071);
nand U11333 (N_11333,N_11011,N_11064);
nor U11334 (N_11334,N_11006,N_11043);
xnor U11335 (N_11335,N_11014,N_11104);
and U11336 (N_11336,N_11040,N_11070);
xor U11337 (N_11337,N_11028,N_11188);
nand U11338 (N_11338,N_11085,N_11053);
xor U11339 (N_11339,N_11108,N_11138);
and U11340 (N_11340,N_11097,N_11124);
nand U11341 (N_11341,N_11068,N_11090);
nand U11342 (N_11342,N_11188,N_11021);
or U11343 (N_11343,N_11135,N_11079);
and U11344 (N_11344,N_11063,N_11113);
and U11345 (N_11345,N_11043,N_11130);
nor U11346 (N_11346,N_11072,N_11011);
xnor U11347 (N_11347,N_11158,N_11130);
nand U11348 (N_11348,N_11040,N_11000);
or U11349 (N_11349,N_11026,N_11040);
or U11350 (N_11350,N_11074,N_11080);
nand U11351 (N_11351,N_11041,N_11098);
and U11352 (N_11352,N_11011,N_11078);
nand U11353 (N_11353,N_11058,N_11191);
xnor U11354 (N_11354,N_11079,N_11174);
or U11355 (N_11355,N_11018,N_11111);
or U11356 (N_11356,N_11011,N_11034);
or U11357 (N_11357,N_11157,N_11008);
nand U11358 (N_11358,N_11117,N_11157);
or U11359 (N_11359,N_11123,N_11103);
xnor U11360 (N_11360,N_11054,N_11049);
nor U11361 (N_11361,N_11130,N_11049);
nand U11362 (N_11362,N_11147,N_11162);
xor U11363 (N_11363,N_11028,N_11135);
and U11364 (N_11364,N_11042,N_11060);
or U11365 (N_11365,N_11006,N_11170);
nand U11366 (N_11366,N_11104,N_11043);
nor U11367 (N_11367,N_11133,N_11079);
nand U11368 (N_11368,N_11110,N_11108);
nor U11369 (N_11369,N_11192,N_11132);
and U11370 (N_11370,N_11170,N_11048);
or U11371 (N_11371,N_11069,N_11188);
and U11372 (N_11372,N_11126,N_11005);
or U11373 (N_11373,N_11053,N_11117);
nor U11374 (N_11374,N_11123,N_11128);
nor U11375 (N_11375,N_11043,N_11176);
nor U11376 (N_11376,N_11062,N_11031);
and U11377 (N_11377,N_11016,N_11044);
nand U11378 (N_11378,N_11183,N_11129);
and U11379 (N_11379,N_11177,N_11026);
and U11380 (N_11380,N_11136,N_11170);
nand U11381 (N_11381,N_11109,N_11039);
nand U11382 (N_11382,N_11096,N_11076);
nor U11383 (N_11383,N_11079,N_11142);
xnor U11384 (N_11384,N_11040,N_11085);
xor U11385 (N_11385,N_11173,N_11193);
nand U11386 (N_11386,N_11097,N_11165);
nor U11387 (N_11387,N_11106,N_11048);
nor U11388 (N_11388,N_11199,N_11110);
nor U11389 (N_11389,N_11125,N_11004);
or U11390 (N_11390,N_11133,N_11145);
nor U11391 (N_11391,N_11064,N_11172);
xnor U11392 (N_11392,N_11134,N_11020);
nand U11393 (N_11393,N_11199,N_11132);
nand U11394 (N_11394,N_11060,N_11002);
nor U11395 (N_11395,N_11120,N_11102);
nand U11396 (N_11396,N_11057,N_11002);
nand U11397 (N_11397,N_11066,N_11100);
or U11398 (N_11398,N_11126,N_11115);
or U11399 (N_11399,N_11035,N_11183);
and U11400 (N_11400,N_11264,N_11281);
xor U11401 (N_11401,N_11262,N_11345);
nor U11402 (N_11402,N_11321,N_11295);
and U11403 (N_11403,N_11308,N_11356);
nand U11404 (N_11404,N_11296,N_11238);
xnor U11405 (N_11405,N_11395,N_11343);
and U11406 (N_11406,N_11387,N_11313);
nand U11407 (N_11407,N_11361,N_11302);
or U11408 (N_11408,N_11366,N_11273);
nand U11409 (N_11409,N_11344,N_11334);
and U11410 (N_11410,N_11222,N_11215);
nor U11411 (N_11411,N_11248,N_11367);
and U11412 (N_11412,N_11223,N_11319);
nor U11413 (N_11413,N_11329,N_11201);
or U11414 (N_11414,N_11259,N_11340);
and U11415 (N_11415,N_11290,N_11202);
or U11416 (N_11416,N_11205,N_11265);
nand U11417 (N_11417,N_11375,N_11324);
xnor U11418 (N_11418,N_11224,N_11261);
nand U11419 (N_11419,N_11227,N_11271);
or U11420 (N_11420,N_11346,N_11278);
nor U11421 (N_11421,N_11210,N_11245);
nand U11422 (N_11422,N_11256,N_11228);
nand U11423 (N_11423,N_11276,N_11233);
and U11424 (N_11424,N_11355,N_11235);
or U11425 (N_11425,N_11305,N_11301);
xnor U11426 (N_11426,N_11326,N_11330);
or U11427 (N_11427,N_11286,N_11275);
nand U11428 (N_11428,N_11268,N_11328);
xnor U11429 (N_11429,N_11325,N_11337);
nor U11430 (N_11430,N_11255,N_11378);
or U11431 (N_11431,N_11382,N_11293);
and U11432 (N_11432,N_11311,N_11317);
nor U11433 (N_11433,N_11348,N_11254);
nand U11434 (N_11434,N_11388,N_11243);
xor U11435 (N_11435,N_11280,N_11251);
nand U11436 (N_11436,N_11269,N_11320);
nor U11437 (N_11437,N_11307,N_11209);
and U11438 (N_11438,N_11327,N_11270);
nand U11439 (N_11439,N_11285,N_11391);
nor U11440 (N_11440,N_11381,N_11394);
nor U11441 (N_11441,N_11252,N_11212);
nand U11442 (N_11442,N_11314,N_11284);
xor U11443 (N_11443,N_11369,N_11208);
nand U11444 (N_11444,N_11266,N_11289);
and U11445 (N_11445,N_11257,N_11300);
and U11446 (N_11446,N_11229,N_11341);
nor U11447 (N_11447,N_11225,N_11246);
nand U11448 (N_11448,N_11312,N_11333);
xnor U11449 (N_11449,N_11203,N_11379);
xor U11450 (N_11450,N_11332,N_11309);
xor U11451 (N_11451,N_11318,N_11230);
xor U11452 (N_11452,N_11216,N_11376);
or U11453 (N_11453,N_11338,N_11383);
or U11454 (N_11454,N_11304,N_11297);
nor U11455 (N_11455,N_11374,N_11206);
and U11456 (N_11456,N_11213,N_11279);
and U11457 (N_11457,N_11299,N_11342);
and U11458 (N_11458,N_11358,N_11385);
and U11459 (N_11459,N_11370,N_11336);
xor U11460 (N_11460,N_11204,N_11260);
xor U11461 (N_11461,N_11352,N_11277);
nor U11462 (N_11462,N_11322,N_11214);
nor U11463 (N_11463,N_11221,N_11372);
nand U11464 (N_11464,N_11219,N_11303);
xor U11465 (N_11465,N_11310,N_11207);
nor U11466 (N_11466,N_11350,N_11390);
or U11467 (N_11467,N_11315,N_11398);
nand U11468 (N_11468,N_11294,N_11283);
or U11469 (N_11469,N_11234,N_11335);
xor U11470 (N_11470,N_11392,N_11247);
or U11471 (N_11471,N_11349,N_11220);
or U11472 (N_11472,N_11298,N_11389);
nand U11473 (N_11473,N_11244,N_11291);
nor U11474 (N_11474,N_11360,N_11339);
nor U11475 (N_11475,N_11347,N_11365);
and U11476 (N_11476,N_11292,N_11288);
and U11477 (N_11477,N_11354,N_11218);
nand U11478 (N_11478,N_11217,N_11263);
nor U11479 (N_11479,N_11272,N_11231);
and U11480 (N_11480,N_11240,N_11237);
and U11481 (N_11481,N_11306,N_11242);
or U11482 (N_11482,N_11386,N_11353);
xnor U11483 (N_11483,N_11351,N_11380);
and U11484 (N_11484,N_11363,N_11371);
xnor U11485 (N_11485,N_11211,N_11377);
xnor U11486 (N_11486,N_11267,N_11226);
or U11487 (N_11487,N_11239,N_11249);
and U11488 (N_11488,N_11258,N_11384);
nand U11489 (N_11489,N_11323,N_11331);
nor U11490 (N_11490,N_11397,N_11357);
or U11491 (N_11491,N_11396,N_11200);
xnor U11492 (N_11492,N_11241,N_11362);
xor U11493 (N_11493,N_11274,N_11236);
xnor U11494 (N_11494,N_11393,N_11232);
nor U11495 (N_11495,N_11316,N_11282);
and U11496 (N_11496,N_11250,N_11364);
nand U11497 (N_11497,N_11253,N_11399);
xnor U11498 (N_11498,N_11368,N_11373);
nor U11499 (N_11499,N_11359,N_11287);
or U11500 (N_11500,N_11280,N_11309);
or U11501 (N_11501,N_11312,N_11286);
nor U11502 (N_11502,N_11342,N_11378);
xnor U11503 (N_11503,N_11339,N_11249);
nor U11504 (N_11504,N_11390,N_11201);
xnor U11505 (N_11505,N_11372,N_11241);
or U11506 (N_11506,N_11263,N_11271);
xnor U11507 (N_11507,N_11209,N_11204);
and U11508 (N_11508,N_11309,N_11256);
and U11509 (N_11509,N_11332,N_11300);
or U11510 (N_11510,N_11399,N_11324);
and U11511 (N_11511,N_11316,N_11312);
or U11512 (N_11512,N_11368,N_11298);
nor U11513 (N_11513,N_11371,N_11385);
nand U11514 (N_11514,N_11284,N_11226);
nand U11515 (N_11515,N_11346,N_11204);
nand U11516 (N_11516,N_11201,N_11373);
nor U11517 (N_11517,N_11381,N_11296);
nand U11518 (N_11518,N_11362,N_11398);
nor U11519 (N_11519,N_11208,N_11341);
and U11520 (N_11520,N_11249,N_11307);
nor U11521 (N_11521,N_11212,N_11388);
xnor U11522 (N_11522,N_11319,N_11263);
and U11523 (N_11523,N_11256,N_11214);
nand U11524 (N_11524,N_11261,N_11275);
nor U11525 (N_11525,N_11214,N_11388);
or U11526 (N_11526,N_11386,N_11318);
and U11527 (N_11527,N_11239,N_11235);
nor U11528 (N_11528,N_11362,N_11214);
nand U11529 (N_11529,N_11392,N_11399);
nand U11530 (N_11530,N_11384,N_11317);
and U11531 (N_11531,N_11333,N_11291);
nand U11532 (N_11532,N_11312,N_11299);
and U11533 (N_11533,N_11360,N_11355);
nand U11534 (N_11534,N_11287,N_11364);
xnor U11535 (N_11535,N_11225,N_11321);
or U11536 (N_11536,N_11302,N_11270);
or U11537 (N_11537,N_11365,N_11396);
xor U11538 (N_11538,N_11294,N_11344);
nand U11539 (N_11539,N_11309,N_11318);
xnor U11540 (N_11540,N_11344,N_11244);
and U11541 (N_11541,N_11389,N_11374);
and U11542 (N_11542,N_11343,N_11285);
nor U11543 (N_11543,N_11396,N_11262);
nand U11544 (N_11544,N_11242,N_11399);
and U11545 (N_11545,N_11205,N_11337);
xor U11546 (N_11546,N_11336,N_11354);
nand U11547 (N_11547,N_11226,N_11258);
and U11548 (N_11548,N_11309,N_11251);
nand U11549 (N_11549,N_11233,N_11346);
xnor U11550 (N_11550,N_11375,N_11376);
xnor U11551 (N_11551,N_11274,N_11309);
nand U11552 (N_11552,N_11216,N_11221);
and U11553 (N_11553,N_11337,N_11242);
nor U11554 (N_11554,N_11263,N_11399);
nor U11555 (N_11555,N_11290,N_11254);
or U11556 (N_11556,N_11213,N_11375);
and U11557 (N_11557,N_11213,N_11356);
xnor U11558 (N_11558,N_11240,N_11234);
or U11559 (N_11559,N_11328,N_11388);
xnor U11560 (N_11560,N_11347,N_11224);
xor U11561 (N_11561,N_11337,N_11314);
nor U11562 (N_11562,N_11240,N_11344);
nand U11563 (N_11563,N_11323,N_11233);
nand U11564 (N_11564,N_11391,N_11396);
nand U11565 (N_11565,N_11244,N_11279);
xnor U11566 (N_11566,N_11308,N_11236);
xor U11567 (N_11567,N_11325,N_11375);
or U11568 (N_11568,N_11267,N_11297);
or U11569 (N_11569,N_11325,N_11263);
or U11570 (N_11570,N_11325,N_11232);
or U11571 (N_11571,N_11345,N_11361);
xnor U11572 (N_11572,N_11352,N_11254);
xor U11573 (N_11573,N_11250,N_11239);
and U11574 (N_11574,N_11286,N_11333);
and U11575 (N_11575,N_11206,N_11341);
nor U11576 (N_11576,N_11257,N_11329);
nor U11577 (N_11577,N_11230,N_11337);
nand U11578 (N_11578,N_11376,N_11345);
and U11579 (N_11579,N_11306,N_11381);
and U11580 (N_11580,N_11293,N_11295);
and U11581 (N_11581,N_11210,N_11349);
and U11582 (N_11582,N_11343,N_11227);
xor U11583 (N_11583,N_11235,N_11203);
nand U11584 (N_11584,N_11228,N_11277);
and U11585 (N_11585,N_11306,N_11378);
nand U11586 (N_11586,N_11239,N_11248);
and U11587 (N_11587,N_11220,N_11330);
xnor U11588 (N_11588,N_11302,N_11380);
or U11589 (N_11589,N_11301,N_11280);
nand U11590 (N_11590,N_11362,N_11319);
nand U11591 (N_11591,N_11211,N_11313);
or U11592 (N_11592,N_11292,N_11283);
and U11593 (N_11593,N_11234,N_11261);
and U11594 (N_11594,N_11269,N_11294);
nor U11595 (N_11595,N_11252,N_11352);
and U11596 (N_11596,N_11209,N_11384);
xor U11597 (N_11597,N_11368,N_11348);
nand U11598 (N_11598,N_11361,N_11237);
and U11599 (N_11599,N_11328,N_11307);
or U11600 (N_11600,N_11572,N_11548);
and U11601 (N_11601,N_11568,N_11528);
nand U11602 (N_11602,N_11431,N_11566);
nand U11603 (N_11603,N_11487,N_11460);
or U11604 (N_11604,N_11511,N_11493);
and U11605 (N_11605,N_11442,N_11541);
or U11606 (N_11606,N_11443,N_11481);
nor U11607 (N_11607,N_11419,N_11588);
and U11608 (N_11608,N_11582,N_11410);
nand U11609 (N_11609,N_11427,N_11547);
nor U11610 (N_11610,N_11455,N_11423);
or U11611 (N_11611,N_11407,N_11584);
nand U11612 (N_11612,N_11537,N_11474);
and U11613 (N_11613,N_11482,N_11401);
and U11614 (N_11614,N_11497,N_11492);
nand U11615 (N_11615,N_11479,N_11424);
or U11616 (N_11616,N_11596,N_11494);
xor U11617 (N_11617,N_11552,N_11430);
nor U11618 (N_11618,N_11496,N_11435);
nand U11619 (N_11619,N_11565,N_11590);
nand U11620 (N_11620,N_11545,N_11409);
xor U11621 (N_11621,N_11543,N_11440);
or U11622 (N_11622,N_11464,N_11476);
and U11623 (N_11623,N_11445,N_11458);
or U11624 (N_11624,N_11402,N_11429);
xor U11625 (N_11625,N_11470,N_11467);
nor U11626 (N_11626,N_11495,N_11436);
xor U11627 (N_11627,N_11502,N_11569);
and U11628 (N_11628,N_11454,N_11463);
xor U11629 (N_11629,N_11488,N_11485);
nor U11630 (N_11630,N_11553,N_11526);
nor U11631 (N_11631,N_11483,N_11585);
nand U11632 (N_11632,N_11425,N_11420);
or U11633 (N_11633,N_11412,N_11418);
xnor U11634 (N_11634,N_11515,N_11587);
xnor U11635 (N_11635,N_11403,N_11562);
nand U11636 (N_11636,N_11477,N_11539);
nor U11637 (N_11637,N_11519,N_11447);
nand U11638 (N_11638,N_11405,N_11521);
nor U11639 (N_11639,N_11598,N_11555);
and U11640 (N_11640,N_11501,N_11580);
xor U11641 (N_11641,N_11509,N_11413);
nand U11642 (N_11642,N_11459,N_11536);
or U11643 (N_11643,N_11400,N_11441);
xnor U11644 (N_11644,N_11449,N_11577);
and U11645 (N_11645,N_11576,N_11434);
and U11646 (N_11646,N_11529,N_11535);
or U11647 (N_11647,N_11556,N_11490);
nor U11648 (N_11648,N_11524,N_11575);
xor U11649 (N_11649,N_11512,N_11408);
and U11650 (N_11650,N_11465,N_11560);
nor U11651 (N_11651,N_11438,N_11461);
or U11652 (N_11652,N_11544,N_11549);
nand U11653 (N_11653,N_11597,N_11583);
and U11654 (N_11654,N_11428,N_11530);
or U11655 (N_11655,N_11550,N_11468);
and U11656 (N_11656,N_11411,N_11586);
xnor U11657 (N_11657,N_11500,N_11491);
nor U11658 (N_11658,N_11533,N_11527);
nand U11659 (N_11659,N_11486,N_11599);
xnor U11660 (N_11660,N_11578,N_11554);
nand U11661 (N_11661,N_11516,N_11573);
xnor U11662 (N_11662,N_11456,N_11453);
and U11663 (N_11663,N_11571,N_11466);
or U11664 (N_11664,N_11564,N_11594);
and U11665 (N_11665,N_11432,N_11517);
xnor U11666 (N_11666,N_11538,N_11534);
xor U11667 (N_11667,N_11522,N_11518);
nor U11668 (N_11668,N_11531,N_11542);
xor U11669 (N_11669,N_11422,N_11508);
or U11670 (N_11670,N_11450,N_11478);
nor U11671 (N_11671,N_11506,N_11520);
nand U11672 (N_11672,N_11472,N_11574);
nor U11673 (N_11673,N_11591,N_11525);
nor U11674 (N_11674,N_11513,N_11589);
xor U11675 (N_11675,N_11593,N_11484);
nand U11676 (N_11676,N_11480,N_11595);
nor U11677 (N_11677,N_11437,N_11433);
or U11678 (N_11678,N_11559,N_11563);
xor U11679 (N_11679,N_11414,N_11444);
nor U11680 (N_11680,N_11532,N_11558);
nor U11681 (N_11681,N_11540,N_11421);
or U11682 (N_11682,N_11504,N_11462);
and U11683 (N_11683,N_11448,N_11546);
or U11684 (N_11684,N_11406,N_11514);
xor U11685 (N_11685,N_11567,N_11523);
xor U11686 (N_11686,N_11503,N_11510);
nor U11687 (N_11687,N_11499,N_11498);
nand U11688 (N_11688,N_11446,N_11415);
and U11689 (N_11689,N_11505,N_11473);
nor U11690 (N_11690,N_11507,N_11417);
nand U11691 (N_11691,N_11426,N_11557);
or U11692 (N_11692,N_11469,N_11581);
or U11693 (N_11693,N_11475,N_11561);
and U11694 (N_11694,N_11489,N_11592);
xnor U11695 (N_11695,N_11416,N_11451);
or U11696 (N_11696,N_11471,N_11439);
and U11697 (N_11697,N_11551,N_11452);
or U11698 (N_11698,N_11404,N_11457);
nor U11699 (N_11699,N_11579,N_11570);
and U11700 (N_11700,N_11574,N_11511);
or U11701 (N_11701,N_11512,N_11534);
nor U11702 (N_11702,N_11564,N_11590);
or U11703 (N_11703,N_11401,N_11588);
nand U11704 (N_11704,N_11496,N_11446);
nor U11705 (N_11705,N_11508,N_11536);
or U11706 (N_11706,N_11416,N_11491);
nor U11707 (N_11707,N_11468,N_11420);
and U11708 (N_11708,N_11406,N_11477);
nand U11709 (N_11709,N_11479,N_11474);
nor U11710 (N_11710,N_11505,N_11436);
nor U11711 (N_11711,N_11446,N_11510);
or U11712 (N_11712,N_11481,N_11537);
nor U11713 (N_11713,N_11509,N_11587);
and U11714 (N_11714,N_11591,N_11431);
or U11715 (N_11715,N_11435,N_11464);
nor U11716 (N_11716,N_11482,N_11461);
xor U11717 (N_11717,N_11449,N_11519);
and U11718 (N_11718,N_11445,N_11464);
nand U11719 (N_11719,N_11447,N_11577);
or U11720 (N_11720,N_11410,N_11442);
nor U11721 (N_11721,N_11482,N_11468);
nand U11722 (N_11722,N_11487,N_11440);
or U11723 (N_11723,N_11407,N_11538);
and U11724 (N_11724,N_11510,N_11566);
and U11725 (N_11725,N_11555,N_11495);
and U11726 (N_11726,N_11554,N_11505);
and U11727 (N_11727,N_11498,N_11418);
xor U11728 (N_11728,N_11504,N_11465);
nand U11729 (N_11729,N_11539,N_11599);
nor U11730 (N_11730,N_11554,N_11426);
or U11731 (N_11731,N_11516,N_11470);
xnor U11732 (N_11732,N_11462,N_11451);
and U11733 (N_11733,N_11481,N_11573);
nand U11734 (N_11734,N_11476,N_11538);
and U11735 (N_11735,N_11414,N_11400);
nor U11736 (N_11736,N_11547,N_11597);
and U11737 (N_11737,N_11528,N_11405);
nor U11738 (N_11738,N_11437,N_11487);
or U11739 (N_11739,N_11516,N_11494);
and U11740 (N_11740,N_11487,N_11453);
xnor U11741 (N_11741,N_11535,N_11553);
and U11742 (N_11742,N_11455,N_11568);
and U11743 (N_11743,N_11500,N_11559);
xnor U11744 (N_11744,N_11441,N_11452);
nand U11745 (N_11745,N_11463,N_11563);
nand U11746 (N_11746,N_11460,N_11486);
xnor U11747 (N_11747,N_11486,N_11508);
nor U11748 (N_11748,N_11475,N_11452);
nor U11749 (N_11749,N_11520,N_11531);
or U11750 (N_11750,N_11580,N_11409);
nor U11751 (N_11751,N_11596,N_11403);
xor U11752 (N_11752,N_11432,N_11425);
and U11753 (N_11753,N_11432,N_11532);
or U11754 (N_11754,N_11417,N_11577);
and U11755 (N_11755,N_11464,N_11494);
or U11756 (N_11756,N_11504,N_11555);
and U11757 (N_11757,N_11520,N_11428);
nand U11758 (N_11758,N_11562,N_11487);
nor U11759 (N_11759,N_11504,N_11558);
nand U11760 (N_11760,N_11486,N_11406);
xor U11761 (N_11761,N_11555,N_11511);
nand U11762 (N_11762,N_11596,N_11560);
xnor U11763 (N_11763,N_11488,N_11591);
xor U11764 (N_11764,N_11483,N_11514);
or U11765 (N_11765,N_11578,N_11424);
or U11766 (N_11766,N_11525,N_11482);
and U11767 (N_11767,N_11564,N_11418);
and U11768 (N_11768,N_11544,N_11496);
xnor U11769 (N_11769,N_11535,N_11593);
nor U11770 (N_11770,N_11568,N_11447);
or U11771 (N_11771,N_11433,N_11448);
nand U11772 (N_11772,N_11402,N_11415);
nor U11773 (N_11773,N_11425,N_11594);
nor U11774 (N_11774,N_11520,N_11416);
nor U11775 (N_11775,N_11436,N_11468);
xor U11776 (N_11776,N_11527,N_11420);
or U11777 (N_11777,N_11587,N_11495);
xor U11778 (N_11778,N_11480,N_11535);
nand U11779 (N_11779,N_11547,N_11478);
xor U11780 (N_11780,N_11429,N_11433);
or U11781 (N_11781,N_11542,N_11421);
xnor U11782 (N_11782,N_11529,N_11581);
xnor U11783 (N_11783,N_11478,N_11593);
and U11784 (N_11784,N_11448,N_11475);
and U11785 (N_11785,N_11551,N_11521);
nand U11786 (N_11786,N_11467,N_11403);
and U11787 (N_11787,N_11566,N_11427);
xor U11788 (N_11788,N_11516,N_11571);
nand U11789 (N_11789,N_11486,N_11487);
nor U11790 (N_11790,N_11562,N_11580);
nand U11791 (N_11791,N_11490,N_11583);
xnor U11792 (N_11792,N_11442,N_11448);
xor U11793 (N_11793,N_11569,N_11559);
or U11794 (N_11794,N_11519,N_11421);
nand U11795 (N_11795,N_11510,N_11499);
xor U11796 (N_11796,N_11486,N_11523);
or U11797 (N_11797,N_11493,N_11544);
and U11798 (N_11798,N_11445,N_11530);
nor U11799 (N_11799,N_11414,N_11565);
and U11800 (N_11800,N_11653,N_11731);
or U11801 (N_11801,N_11755,N_11756);
and U11802 (N_11802,N_11695,N_11689);
or U11803 (N_11803,N_11638,N_11719);
and U11804 (N_11804,N_11607,N_11778);
nand U11805 (N_11805,N_11779,N_11681);
and U11806 (N_11806,N_11616,N_11614);
or U11807 (N_11807,N_11669,N_11786);
nor U11808 (N_11808,N_11637,N_11691);
nand U11809 (N_11809,N_11643,N_11641);
nand U11810 (N_11810,N_11741,N_11792);
or U11811 (N_11811,N_11605,N_11795);
and U11812 (N_11812,N_11718,N_11721);
or U11813 (N_11813,N_11662,N_11749);
or U11814 (N_11814,N_11774,N_11712);
and U11815 (N_11815,N_11687,N_11720);
and U11816 (N_11816,N_11780,N_11738);
nor U11817 (N_11817,N_11652,N_11600);
xor U11818 (N_11818,N_11713,N_11690);
or U11819 (N_11819,N_11601,N_11745);
xor U11820 (N_11820,N_11644,N_11750);
and U11821 (N_11821,N_11751,N_11761);
and U11822 (N_11822,N_11760,N_11610);
xnor U11823 (N_11823,N_11602,N_11697);
nand U11824 (N_11824,N_11688,N_11724);
xor U11825 (N_11825,N_11753,N_11717);
nand U11826 (N_11826,N_11645,N_11722);
nor U11827 (N_11827,N_11618,N_11796);
and U11828 (N_11828,N_11651,N_11683);
and U11829 (N_11829,N_11708,N_11621);
xnor U11830 (N_11830,N_11673,N_11613);
and U11831 (N_11831,N_11622,N_11785);
or U11832 (N_11832,N_11677,N_11606);
and U11833 (N_11833,N_11740,N_11773);
nand U11834 (N_11834,N_11723,N_11647);
and U11835 (N_11835,N_11781,N_11646);
xnor U11836 (N_11836,N_11707,N_11709);
nor U11837 (N_11837,N_11725,N_11636);
and U11838 (N_11838,N_11770,N_11663);
nor U11839 (N_11839,N_11633,N_11629);
and U11840 (N_11840,N_11703,N_11776);
and U11841 (N_11841,N_11783,N_11706);
nor U11842 (N_11842,N_11676,N_11611);
nand U11843 (N_11843,N_11667,N_11728);
or U11844 (N_11844,N_11694,N_11692);
or U11845 (N_11845,N_11771,N_11682);
or U11846 (N_11846,N_11711,N_11767);
nor U11847 (N_11847,N_11631,N_11623);
xnor U11848 (N_11848,N_11639,N_11635);
nand U11849 (N_11849,N_11649,N_11699);
or U11850 (N_11850,N_11735,N_11769);
xnor U11851 (N_11851,N_11791,N_11793);
nor U11852 (N_11852,N_11757,N_11627);
or U11853 (N_11853,N_11619,N_11715);
nor U11854 (N_11854,N_11705,N_11626);
and U11855 (N_11855,N_11620,N_11668);
or U11856 (N_11856,N_11630,N_11609);
nor U11857 (N_11857,N_11799,N_11789);
and U11858 (N_11858,N_11762,N_11742);
xnor U11859 (N_11859,N_11768,N_11661);
or U11860 (N_11860,N_11678,N_11608);
nand U11861 (N_11861,N_11765,N_11790);
nand U11862 (N_11862,N_11714,N_11777);
or U11863 (N_11863,N_11612,N_11754);
nand U11864 (N_11864,N_11674,N_11732);
nand U11865 (N_11865,N_11746,N_11752);
nand U11866 (N_11866,N_11628,N_11734);
and U11867 (N_11867,N_11625,N_11710);
xor U11868 (N_11868,N_11666,N_11736);
xnor U11869 (N_11869,N_11798,N_11772);
or U11870 (N_11870,N_11675,N_11640);
xnor U11871 (N_11871,N_11648,N_11784);
and U11872 (N_11872,N_11684,N_11733);
or U11873 (N_11873,N_11671,N_11794);
nor U11874 (N_11874,N_11664,N_11726);
xnor U11875 (N_11875,N_11680,N_11716);
and U11876 (N_11876,N_11758,N_11782);
and U11877 (N_11877,N_11700,N_11696);
or U11878 (N_11878,N_11615,N_11693);
nand U11879 (N_11879,N_11658,N_11617);
nand U11880 (N_11880,N_11659,N_11727);
or U11881 (N_11881,N_11624,N_11698);
or U11882 (N_11882,N_11657,N_11730);
nand U11883 (N_11883,N_11747,N_11603);
nand U11884 (N_11884,N_11654,N_11670);
nor U11885 (N_11885,N_11763,N_11632);
xor U11886 (N_11886,N_11729,N_11788);
nor U11887 (N_11887,N_11642,N_11766);
xor U11888 (N_11888,N_11787,N_11797);
and U11889 (N_11889,N_11702,N_11739);
or U11890 (N_11890,N_11650,N_11744);
nor U11891 (N_11891,N_11701,N_11704);
nor U11892 (N_11892,N_11743,N_11737);
or U11893 (N_11893,N_11764,N_11686);
nand U11894 (N_11894,N_11759,N_11748);
nor U11895 (N_11895,N_11685,N_11679);
xor U11896 (N_11896,N_11604,N_11634);
xnor U11897 (N_11897,N_11656,N_11665);
or U11898 (N_11898,N_11672,N_11775);
nor U11899 (N_11899,N_11660,N_11655);
nand U11900 (N_11900,N_11610,N_11778);
or U11901 (N_11901,N_11696,N_11602);
xnor U11902 (N_11902,N_11731,N_11638);
nand U11903 (N_11903,N_11605,N_11727);
nand U11904 (N_11904,N_11761,N_11715);
nor U11905 (N_11905,N_11718,N_11739);
and U11906 (N_11906,N_11631,N_11743);
or U11907 (N_11907,N_11783,N_11631);
or U11908 (N_11908,N_11742,N_11761);
nand U11909 (N_11909,N_11655,N_11754);
nor U11910 (N_11910,N_11757,N_11727);
or U11911 (N_11911,N_11774,N_11627);
nand U11912 (N_11912,N_11648,N_11716);
and U11913 (N_11913,N_11706,N_11601);
nand U11914 (N_11914,N_11719,N_11739);
or U11915 (N_11915,N_11713,N_11789);
and U11916 (N_11916,N_11711,N_11726);
nand U11917 (N_11917,N_11627,N_11764);
and U11918 (N_11918,N_11712,N_11790);
and U11919 (N_11919,N_11694,N_11731);
and U11920 (N_11920,N_11636,N_11721);
and U11921 (N_11921,N_11791,N_11699);
or U11922 (N_11922,N_11665,N_11641);
nor U11923 (N_11923,N_11656,N_11788);
nor U11924 (N_11924,N_11726,N_11638);
nor U11925 (N_11925,N_11655,N_11622);
and U11926 (N_11926,N_11792,N_11662);
nor U11927 (N_11927,N_11627,N_11713);
or U11928 (N_11928,N_11718,N_11631);
nor U11929 (N_11929,N_11648,N_11638);
and U11930 (N_11930,N_11750,N_11743);
nand U11931 (N_11931,N_11736,N_11613);
or U11932 (N_11932,N_11666,N_11656);
and U11933 (N_11933,N_11726,N_11742);
nor U11934 (N_11934,N_11772,N_11762);
or U11935 (N_11935,N_11642,N_11633);
nor U11936 (N_11936,N_11787,N_11627);
and U11937 (N_11937,N_11750,N_11658);
nor U11938 (N_11938,N_11792,N_11791);
nand U11939 (N_11939,N_11785,N_11759);
and U11940 (N_11940,N_11686,N_11683);
or U11941 (N_11941,N_11634,N_11636);
or U11942 (N_11942,N_11782,N_11711);
xnor U11943 (N_11943,N_11783,N_11661);
xnor U11944 (N_11944,N_11744,N_11723);
or U11945 (N_11945,N_11687,N_11663);
and U11946 (N_11946,N_11706,N_11795);
or U11947 (N_11947,N_11673,N_11618);
xnor U11948 (N_11948,N_11613,N_11695);
and U11949 (N_11949,N_11683,N_11606);
and U11950 (N_11950,N_11622,N_11657);
nor U11951 (N_11951,N_11749,N_11629);
nor U11952 (N_11952,N_11643,N_11739);
nor U11953 (N_11953,N_11742,N_11704);
nor U11954 (N_11954,N_11663,N_11735);
nand U11955 (N_11955,N_11791,N_11780);
xnor U11956 (N_11956,N_11687,N_11721);
nand U11957 (N_11957,N_11619,N_11780);
nor U11958 (N_11958,N_11709,N_11772);
or U11959 (N_11959,N_11635,N_11655);
or U11960 (N_11960,N_11719,N_11629);
nand U11961 (N_11961,N_11630,N_11663);
nor U11962 (N_11962,N_11792,N_11715);
xor U11963 (N_11963,N_11611,N_11614);
nor U11964 (N_11964,N_11735,N_11738);
nor U11965 (N_11965,N_11609,N_11738);
nor U11966 (N_11966,N_11794,N_11796);
and U11967 (N_11967,N_11776,N_11736);
and U11968 (N_11968,N_11710,N_11789);
or U11969 (N_11969,N_11700,N_11643);
xor U11970 (N_11970,N_11655,N_11767);
xor U11971 (N_11971,N_11642,N_11661);
nor U11972 (N_11972,N_11617,N_11720);
or U11973 (N_11973,N_11682,N_11611);
and U11974 (N_11974,N_11773,N_11734);
or U11975 (N_11975,N_11722,N_11787);
and U11976 (N_11976,N_11730,N_11797);
nor U11977 (N_11977,N_11696,N_11761);
or U11978 (N_11978,N_11644,N_11766);
nand U11979 (N_11979,N_11774,N_11673);
and U11980 (N_11980,N_11648,N_11750);
xnor U11981 (N_11981,N_11795,N_11752);
nand U11982 (N_11982,N_11716,N_11674);
nand U11983 (N_11983,N_11642,N_11663);
xnor U11984 (N_11984,N_11797,N_11782);
nand U11985 (N_11985,N_11675,N_11612);
nand U11986 (N_11986,N_11731,N_11790);
nor U11987 (N_11987,N_11649,N_11616);
or U11988 (N_11988,N_11757,N_11625);
nand U11989 (N_11989,N_11671,N_11708);
xnor U11990 (N_11990,N_11652,N_11781);
xnor U11991 (N_11991,N_11611,N_11638);
nor U11992 (N_11992,N_11670,N_11647);
or U11993 (N_11993,N_11780,N_11754);
and U11994 (N_11994,N_11663,N_11743);
or U11995 (N_11995,N_11611,N_11770);
and U11996 (N_11996,N_11714,N_11681);
and U11997 (N_11997,N_11672,N_11663);
or U11998 (N_11998,N_11769,N_11632);
and U11999 (N_11999,N_11711,N_11688);
nand U12000 (N_12000,N_11996,N_11981);
xor U12001 (N_12001,N_11870,N_11963);
or U12002 (N_12002,N_11990,N_11975);
nor U12003 (N_12003,N_11946,N_11959);
xnor U12004 (N_12004,N_11833,N_11955);
or U12005 (N_12005,N_11889,N_11878);
nor U12006 (N_12006,N_11874,N_11911);
or U12007 (N_12007,N_11826,N_11979);
and U12008 (N_12008,N_11873,N_11988);
xnor U12009 (N_12009,N_11844,N_11853);
and U12010 (N_12010,N_11815,N_11830);
or U12011 (N_12011,N_11942,N_11887);
or U12012 (N_12012,N_11840,N_11993);
nor U12013 (N_12013,N_11822,N_11970);
and U12014 (N_12014,N_11901,N_11858);
nand U12015 (N_12015,N_11824,N_11848);
xnor U12016 (N_12016,N_11860,N_11890);
nor U12017 (N_12017,N_11888,N_11967);
nor U12018 (N_12018,N_11903,N_11954);
or U12019 (N_12019,N_11839,N_11987);
xor U12020 (N_12020,N_11929,N_11899);
nand U12021 (N_12021,N_11936,N_11968);
or U12022 (N_12022,N_11964,N_11800);
nor U12023 (N_12023,N_11875,N_11802);
nand U12024 (N_12024,N_11927,N_11881);
xnor U12025 (N_12025,N_11895,N_11953);
nand U12026 (N_12026,N_11947,N_11950);
and U12027 (N_12027,N_11882,N_11819);
nand U12028 (N_12028,N_11891,N_11814);
nor U12029 (N_12029,N_11969,N_11926);
nand U12030 (N_12030,N_11948,N_11810);
nor U12031 (N_12031,N_11921,N_11861);
nand U12032 (N_12032,N_11842,N_11821);
and U12033 (N_12033,N_11843,N_11999);
nand U12034 (N_12034,N_11896,N_11971);
or U12035 (N_12035,N_11806,N_11944);
nor U12036 (N_12036,N_11931,N_11864);
and U12037 (N_12037,N_11820,N_11908);
xnor U12038 (N_12038,N_11918,N_11836);
nor U12039 (N_12039,N_11912,N_11907);
xnor U12040 (N_12040,N_11977,N_11832);
nand U12041 (N_12041,N_11985,N_11933);
nand U12042 (N_12042,N_11976,N_11941);
nor U12043 (N_12043,N_11893,N_11823);
nand U12044 (N_12044,N_11919,N_11827);
xor U12045 (N_12045,N_11837,N_11872);
xnor U12046 (N_12046,N_11885,N_11894);
or U12047 (N_12047,N_11965,N_11851);
or U12048 (N_12048,N_11961,N_11940);
nor U12049 (N_12049,N_11974,N_11937);
nor U12050 (N_12050,N_11811,N_11852);
nor U12051 (N_12051,N_11915,N_11869);
nor U12052 (N_12052,N_11829,N_11904);
nand U12053 (N_12053,N_11897,N_11998);
or U12054 (N_12054,N_11883,N_11962);
xnor U12055 (N_12055,N_11935,N_11992);
or U12056 (N_12056,N_11978,N_11857);
nand U12057 (N_12057,N_11809,N_11973);
nand U12058 (N_12058,N_11945,N_11952);
nor U12059 (N_12059,N_11982,N_11960);
xor U12060 (N_12060,N_11983,N_11831);
nand U12061 (N_12061,N_11923,N_11867);
nor U12062 (N_12062,N_11924,N_11957);
nor U12063 (N_12063,N_11917,N_11855);
nand U12064 (N_12064,N_11939,N_11966);
nand U12065 (N_12065,N_11807,N_11808);
nand U12066 (N_12066,N_11943,N_11989);
or U12067 (N_12067,N_11812,N_11801);
nor U12068 (N_12068,N_11818,N_11835);
or U12069 (N_12069,N_11871,N_11856);
nand U12070 (N_12070,N_11910,N_11825);
xor U12071 (N_12071,N_11956,N_11991);
xnor U12072 (N_12072,N_11905,N_11909);
xor U12073 (N_12073,N_11816,N_11980);
xnor U12074 (N_12074,N_11850,N_11862);
and U12075 (N_12075,N_11834,N_11876);
and U12076 (N_12076,N_11949,N_11859);
nand U12077 (N_12077,N_11984,N_11884);
nand U12078 (N_12078,N_11817,N_11997);
nor U12079 (N_12079,N_11845,N_11877);
nand U12080 (N_12080,N_11986,N_11804);
nor U12081 (N_12081,N_11938,N_11868);
or U12082 (N_12082,N_11932,N_11920);
nand U12083 (N_12083,N_11900,N_11838);
and U12084 (N_12084,N_11879,N_11863);
nor U12085 (N_12085,N_11902,N_11828);
nor U12086 (N_12086,N_11930,N_11906);
nor U12087 (N_12087,N_11925,N_11916);
or U12088 (N_12088,N_11813,N_11898);
and U12089 (N_12089,N_11922,N_11805);
or U12090 (N_12090,N_11846,N_11994);
nand U12091 (N_12091,N_11951,N_11928);
nand U12092 (N_12092,N_11972,N_11866);
nand U12093 (N_12093,N_11914,N_11865);
nand U12094 (N_12094,N_11880,N_11854);
or U12095 (N_12095,N_11913,N_11841);
nand U12096 (N_12096,N_11892,N_11849);
or U12097 (N_12097,N_11886,N_11847);
and U12098 (N_12098,N_11958,N_11995);
xor U12099 (N_12099,N_11803,N_11934);
nand U12100 (N_12100,N_11917,N_11992);
xor U12101 (N_12101,N_11964,N_11955);
or U12102 (N_12102,N_11831,N_11891);
xor U12103 (N_12103,N_11897,N_11867);
or U12104 (N_12104,N_11808,N_11967);
xnor U12105 (N_12105,N_11807,N_11944);
or U12106 (N_12106,N_11923,N_11990);
and U12107 (N_12107,N_11936,N_11941);
nand U12108 (N_12108,N_11971,N_11910);
or U12109 (N_12109,N_11823,N_11924);
and U12110 (N_12110,N_11967,N_11836);
and U12111 (N_12111,N_11818,N_11871);
nor U12112 (N_12112,N_11964,N_11966);
and U12113 (N_12113,N_11902,N_11837);
nor U12114 (N_12114,N_11881,N_11896);
and U12115 (N_12115,N_11808,N_11863);
nor U12116 (N_12116,N_11816,N_11902);
and U12117 (N_12117,N_11992,N_11901);
or U12118 (N_12118,N_11830,N_11957);
and U12119 (N_12119,N_11919,N_11852);
nor U12120 (N_12120,N_11977,N_11903);
or U12121 (N_12121,N_11866,N_11834);
or U12122 (N_12122,N_11956,N_11966);
or U12123 (N_12123,N_11864,N_11905);
and U12124 (N_12124,N_11895,N_11872);
and U12125 (N_12125,N_11924,N_11953);
nor U12126 (N_12126,N_11817,N_11830);
xor U12127 (N_12127,N_11833,N_11871);
and U12128 (N_12128,N_11904,N_11885);
or U12129 (N_12129,N_11904,N_11942);
and U12130 (N_12130,N_11897,N_11841);
nor U12131 (N_12131,N_11913,N_11854);
nand U12132 (N_12132,N_11873,N_11877);
nand U12133 (N_12133,N_11900,N_11854);
and U12134 (N_12134,N_11980,N_11876);
and U12135 (N_12135,N_11993,N_11983);
and U12136 (N_12136,N_11915,N_11953);
or U12137 (N_12137,N_11864,N_11901);
nand U12138 (N_12138,N_11879,N_11824);
nor U12139 (N_12139,N_11879,N_11992);
or U12140 (N_12140,N_11990,N_11857);
xor U12141 (N_12141,N_11849,N_11981);
xnor U12142 (N_12142,N_11990,N_11818);
xor U12143 (N_12143,N_11906,N_11886);
xor U12144 (N_12144,N_11917,N_11933);
nand U12145 (N_12145,N_11926,N_11925);
nor U12146 (N_12146,N_11895,N_11808);
or U12147 (N_12147,N_11923,N_11807);
or U12148 (N_12148,N_11920,N_11938);
or U12149 (N_12149,N_11961,N_11823);
nor U12150 (N_12150,N_11820,N_11970);
and U12151 (N_12151,N_11818,N_11941);
xor U12152 (N_12152,N_11818,N_11984);
and U12153 (N_12153,N_11864,N_11805);
or U12154 (N_12154,N_11807,N_11851);
or U12155 (N_12155,N_11839,N_11994);
xnor U12156 (N_12156,N_11927,N_11843);
and U12157 (N_12157,N_11880,N_11850);
nand U12158 (N_12158,N_11876,N_11889);
and U12159 (N_12159,N_11895,N_11978);
nand U12160 (N_12160,N_11884,N_11954);
nor U12161 (N_12161,N_11913,N_11823);
or U12162 (N_12162,N_11943,N_11960);
nor U12163 (N_12163,N_11902,N_11956);
xnor U12164 (N_12164,N_11815,N_11909);
or U12165 (N_12165,N_11800,N_11835);
nor U12166 (N_12166,N_11999,N_11934);
xor U12167 (N_12167,N_11879,N_11925);
nor U12168 (N_12168,N_11922,N_11986);
or U12169 (N_12169,N_11945,N_11977);
or U12170 (N_12170,N_11966,N_11861);
and U12171 (N_12171,N_11943,N_11935);
and U12172 (N_12172,N_11853,N_11805);
xor U12173 (N_12173,N_11860,N_11978);
or U12174 (N_12174,N_11858,N_11982);
and U12175 (N_12175,N_11926,N_11880);
and U12176 (N_12176,N_11837,N_11813);
or U12177 (N_12177,N_11994,N_11837);
or U12178 (N_12178,N_11847,N_11865);
or U12179 (N_12179,N_11912,N_11862);
and U12180 (N_12180,N_11812,N_11877);
nor U12181 (N_12181,N_11800,N_11838);
xnor U12182 (N_12182,N_11961,N_11894);
nor U12183 (N_12183,N_11845,N_11981);
or U12184 (N_12184,N_11994,N_11955);
nor U12185 (N_12185,N_11805,N_11808);
or U12186 (N_12186,N_11820,N_11826);
or U12187 (N_12187,N_11908,N_11854);
nand U12188 (N_12188,N_11969,N_11863);
nor U12189 (N_12189,N_11892,N_11998);
and U12190 (N_12190,N_11915,N_11859);
nand U12191 (N_12191,N_11872,N_11890);
nor U12192 (N_12192,N_11996,N_11927);
nand U12193 (N_12193,N_11999,N_11828);
nand U12194 (N_12194,N_11879,N_11949);
xor U12195 (N_12195,N_11851,N_11854);
or U12196 (N_12196,N_11910,N_11909);
and U12197 (N_12197,N_11826,N_11866);
nor U12198 (N_12198,N_11965,N_11964);
xnor U12199 (N_12199,N_11827,N_11975);
or U12200 (N_12200,N_12133,N_12105);
or U12201 (N_12201,N_12199,N_12171);
nor U12202 (N_12202,N_12167,N_12029);
or U12203 (N_12203,N_12142,N_12150);
nor U12204 (N_12204,N_12129,N_12122);
or U12205 (N_12205,N_12135,N_12012);
xor U12206 (N_12206,N_12168,N_12076);
xnor U12207 (N_12207,N_12103,N_12050);
nand U12208 (N_12208,N_12104,N_12027);
nor U12209 (N_12209,N_12079,N_12075);
and U12210 (N_12210,N_12138,N_12155);
and U12211 (N_12211,N_12143,N_12198);
nor U12212 (N_12212,N_12173,N_12035);
and U12213 (N_12213,N_12019,N_12115);
or U12214 (N_12214,N_12088,N_12186);
or U12215 (N_12215,N_12040,N_12169);
or U12216 (N_12216,N_12023,N_12055);
xnor U12217 (N_12217,N_12126,N_12144);
and U12218 (N_12218,N_12125,N_12134);
or U12219 (N_12219,N_12187,N_12087);
nor U12220 (N_12220,N_12073,N_12082);
and U12221 (N_12221,N_12128,N_12059);
and U12222 (N_12222,N_12193,N_12149);
nor U12223 (N_12223,N_12045,N_12188);
nor U12224 (N_12224,N_12178,N_12097);
xor U12225 (N_12225,N_12030,N_12086);
nor U12226 (N_12226,N_12148,N_12051);
nand U12227 (N_12227,N_12197,N_12185);
nand U12228 (N_12228,N_12106,N_12114);
nand U12229 (N_12229,N_12170,N_12089);
xnor U12230 (N_12230,N_12189,N_12111);
and U12231 (N_12231,N_12101,N_12092);
and U12232 (N_12232,N_12110,N_12049);
and U12233 (N_12233,N_12192,N_12033);
and U12234 (N_12234,N_12151,N_12090);
nand U12235 (N_12235,N_12057,N_12043);
nor U12236 (N_12236,N_12118,N_12183);
and U12237 (N_12237,N_12081,N_12016);
and U12238 (N_12238,N_12176,N_12137);
or U12239 (N_12239,N_12174,N_12181);
xnor U12240 (N_12240,N_12044,N_12146);
nand U12241 (N_12241,N_12066,N_12136);
nand U12242 (N_12242,N_12147,N_12062);
nand U12243 (N_12243,N_12071,N_12085);
nand U12244 (N_12244,N_12037,N_12154);
nand U12245 (N_12245,N_12164,N_12119);
and U12246 (N_12246,N_12056,N_12011);
or U12247 (N_12247,N_12005,N_12007);
nor U12248 (N_12248,N_12179,N_12067);
and U12249 (N_12249,N_12026,N_12070);
or U12250 (N_12250,N_12161,N_12013);
and U12251 (N_12251,N_12194,N_12063);
nor U12252 (N_12252,N_12182,N_12031);
xor U12253 (N_12253,N_12131,N_12172);
nor U12254 (N_12254,N_12038,N_12163);
xnor U12255 (N_12255,N_12157,N_12020);
and U12256 (N_12256,N_12036,N_12107);
or U12257 (N_12257,N_12175,N_12121);
nand U12258 (N_12258,N_12021,N_12074);
nand U12259 (N_12259,N_12032,N_12080);
xnor U12260 (N_12260,N_12096,N_12091);
nor U12261 (N_12261,N_12078,N_12098);
and U12262 (N_12262,N_12004,N_12152);
or U12263 (N_12263,N_12054,N_12184);
xor U12264 (N_12264,N_12180,N_12060);
nand U12265 (N_12265,N_12022,N_12025);
or U12266 (N_12266,N_12018,N_12039);
or U12267 (N_12267,N_12156,N_12061);
and U12268 (N_12268,N_12064,N_12153);
and U12269 (N_12269,N_12117,N_12109);
nand U12270 (N_12270,N_12093,N_12014);
or U12271 (N_12271,N_12006,N_12165);
or U12272 (N_12272,N_12048,N_12001);
nand U12273 (N_12273,N_12046,N_12083);
and U12274 (N_12274,N_12102,N_12160);
xnor U12275 (N_12275,N_12113,N_12000);
or U12276 (N_12276,N_12177,N_12042);
xnor U12277 (N_12277,N_12017,N_12140);
xnor U12278 (N_12278,N_12162,N_12190);
and U12279 (N_12279,N_12116,N_12084);
xor U12280 (N_12280,N_12003,N_12065);
nand U12281 (N_12281,N_12094,N_12132);
and U12282 (N_12282,N_12130,N_12010);
and U12283 (N_12283,N_12095,N_12158);
xnor U12284 (N_12284,N_12024,N_12123);
xor U12285 (N_12285,N_12141,N_12112);
or U12286 (N_12286,N_12053,N_12008);
or U12287 (N_12287,N_12015,N_12196);
or U12288 (N_12288,N_12034,N_12100);
or U12289 (N_12289,N_12127,N_12120);
nor U12290 (N_12290,N_12058,N_12041);
nand U12291 (N_12291,N_12159,N_12145);
nor U12292 (N_12292,N_12052,N_12047);
and U12293 (N_12293,N_12139,N_12108);
or U12294 (N_12294,N_12009,N_12195);
or U12295 (N_12295,N_12077,N_12068);
or U12296 (N_12296,N_12191,N_12072);
or U12297 (N_12297,N_12028,N_12166);
and U12298 (N_12298,N_12099,N_12002);
nor U12299 (N_12299,N_12124,N_12069);
nand U12300 (N_12300,N_12077,N_12119);
nor U12301 (N_12301,N_12146,N_12135);
xnor U12302 (N_12302,N_12090,N_12042);
xnor U12303 (N_12303,N_12091,N_12196);
nor U12304 (N_12304,N_12057,N_12171);
and U12305 (N_12305,N_12094,N_12196);
or U12306 (N_12306,N_12141,N_12192);
or U12307 (N_12307,N_12120,N_12172);
xor U12308 (N_12308,N_12031,N_12040);
xnor U12309 (N_12309,N_12083,N_12100);
xor U12310 (N_12310,N_12184,N_12002);
and U12311 (N_12311,N_12122,N_12098);
nand U12312 (N_12312,N_12110,N_12154);
or U12313 (N_12313,N_12086,N_12043);
xor U12314 (N_12314,N_12188,N_12162);
or U12315 (N_12315,N_12096,N_12131);
xnor U12316 (N_12316,N_12072,N_12176);
or U12317 (N_12317,N_12000,N_12102);
xor U12318 (N_12318,N_12100,N_12096);
and U12319 (N_12319,N_12000,N_12052);
and U12320 (N_12320,N_12073,N_12195);
nand U12321 (N_12321,N_12087,N_12031);
nor U12322 (N_12322,N_12057,N_12021);
or U12323 (N_12323,N_12143,N_12165);
xor U12324 (N_12324,N_12132,N_12042);
nand U12325 (N_12325,N_12122,N_12022);
nor U12326 (N_12326,N_12086,N_12146);
or U12327 (N_12327,N_12183,N_12093);
nand U12328 (N_12328,N_12011,N_12129);
or U12329 (N_12329,N_12051,N_12062);
and U12330 (N_12330,N_12057,N_12017);
or U12331 (N_12331,N_12122,N_12111);
nand U12332 (N_12332,N_12160,N_12003);
xnor U12333 (N_12333,N_12128,N_12043);
nor U12334 (N_12334,N_12101,N_12156);
or U12335 (N_12335,N_12149,N_12131);
nand U12336 (N_12336,N_12170,N_12105);
xor U12337 (N_12337,N_12133,N_12066);
xor U12338 (N_12338,N_12049,N_12095);
nand U12339 (N_12339,N_12100,N_12143);
or U12340 (N_12340,N_12034,N_12039);
nand U12341 (N_12341,N_12123,N_12014);
and U12342 (N_12342,N_12125,N_12081);
nor U12343 (N_12343,N_12182,N_12029);
and U12344 (N_12344,N_12199,N_12150);
xnor U12345 (N_12345,N_12152,N_12128);
or U12346 (N_12346,N_12144,N_12041);
and U12347 (N_12347,N_12160,N_12044);
nor U12348 (N_12348,N_12093,N_12100);
xnor U12349 (N_12349,N_12174,N_12066);
and U12350 (N_12350,N_12036,N_12006);
xnor U12351 (N_12351,N_12189,N_12161);
and U12352 (N_12352,N_12189,N_12058);
nand U12353 (N_12353,N_12071,N_12030);
or U12354 (N_12354,N_12195,N_12113);
nand U12355 (N_12355,N_12171,N_12161);
xor U12356 (N_12356,N_12198,N_12135);
nor U12357 (N_12357,N_12039,N_12174);
nor U12358 (N_12358,N_12174,N_12142);
or U12359 (N_12359,N_12127,N_12186);
nand U12360 (N_12360,N_12073,N_12134);
and U12361 (N_12361,N_12124,N_12004);
nand U12362 (N_12362,N_12093,N_12173);
nor U12363 (N_12363,N_12091,N_12040);
or U12364 (N_12364,N_12078,N_12162);
xnor U12365 (N_12365,N_12094,N_12147);
xnor U12366 (N_12366,N_12002,N_12151);
nand U12367 (N_12367,N_12054,N_12012);
xnor U12368 (N_12368,N_12017,N_12142);
nor U12369 (N_12369,N_12136,N_12020);
and U12370 (N_12370,N_12091,N_12175);
and U12371 (N_12371,N_12185,N_12010);
xor U12372 (N_12372,N_12124,N_12061);
and U12373 (N_12373,N_12128,N_12166);
or U12374 (N_12374,N_12042,N_12158);
nand U12375 (N_12375,N_12060,N_12034);
nor U12376 (N_12376,N_12186,N_12042);
nor U12377 (N_12377,N_12124,N_12134);
nand U12378 (N_12378,N_12176,N_12108);
xnor U12379 (N_12379,N_12132,N_12168);
xor U12380 (N_12380,N_12013,N_12157);
nor U12381 (N_12381,N_12129,N_12171);
and U12382 (N_12382,N_12121,N_12146);
nand U12383 (N_12383,N_12095,N_12028);
nor U12384 (N_12384,N_12141,N_12136);
xnor U12385 (N_12385,N_12008,N_12189);
nor U12386 (N_12386,N_12140,N_12188);
nor U12387 (N_12387,N_12155,N_12118);
or U12388 (N_12388,N_12016,N_12113);
nand U12389 (N_12389,N_12155,N_12153);
or U12390 (N_12390,N_12119,N_12173);
xnor U12391 (N_12391,N_12141,N_12109);
nor U12392 (N_12392,N_12025,N_12124);
nor U12393 (N_12393,N_12193,N_12190);
nor U12394 (N_12394,N_12006,N_12060);
and U12395 (N_12395,N_12128,N_12033);
nand U12396 (N_12396,N_12180,N_12123);
and U12397 (N_12397,N_12031,N_12100);
nand U12398 (N_12398,N_12165,N_12081);
xnor U12399 (N_12399,N_12074,N_12100);
and U12400 (N_12400,N_12288,N_12365);
nor U12401 (N_12401,N_12389,N_12358);
and U12402 (N_12402,N_12260,N_12302);
nor U12403 (N_12403,N_12285,N_12239);
nor U12404 (N_12404,N_12298,N_12387);
nand U12405 (N_12405,N_12225,N_12265);
nand U12406 (N_12406,N_12290,N_12276);
and U12407 (N_12407,N_12201,N_12234);
nor U12408 (N_12408,N_12390,N_12224);
or U12409 (N_12409,N_12299,N_12381);
nor U12410 (N_12410,N_12316,N_12210);
or U12411 (N_12411,N_12277,N_12203);
xnor U12412 (N_12412,N_12398,N_12315);
or U12413 (N_12413,N_12331,N_12394);
nand U12414 (N_12414,N_12269,N_12388);
and U12415 (N_12415,N_12246,N_12371);
and U12416 (N_12416,N_12392,N_12206);
nor U12417 (N_12417,N_12374,N_12372);
and U12418 (N_12418,N_12244,N_12322);
nand U12419 (N_12419,N_12279,N_12295);
and U12420 (N_12420,N_12235,N_12230);
nand U12421 (N_12421,N_12251,N_12223);
xnor U12422 (N_12422,N_12350,N_12283);
nand U12423 (N_12423,N_12301,N_12297);
and U12424 (N_12424,N_12289,N_12249);
nor U12425 (N_12425,N_12382,N_12262);
and U12426 (N_12426,N_12347,N_12311);
xor U12427 (N_12427,N_12308,N_12329);
nor U12428 (N_12428,N_12378,N_12364);
nor U12429 (N_12429,N_12352,N_12384);
or U12430 (N_12430,N_12343,N_12214);
nor U12431 (N_12431,N_12280,N_12375);
and U12432 (N_12432,N_12231,N_12355);
or U12433 (N_12433,N_12304,N_12377);
or U12434 (N_12434,N_12253,N_12293);
nor U12435 (N_12435,N_12263,N_12273);
nor U12436 (N_12436,N_12266,N_12325);
and U12437 (N_12437,N_12391,N_12346);
nand U12438 (N_12438,N_12237,N_12335);
nand U12439 (N_12439,N_12305,N_12323);
xnor U12440 (N_12440,N_12267,N_12360);
nand U12441 (N_12441,N_12200,N_12205);
nor U12442 (N_12442,N_12354,N_12278);
nand U12443 (N_12443,N_12353,N_12281);
or U12444 (N_12444,N_12349,N_12261);
nor U12445 (N_12445,N_12208,N_12268);
xnor U12446 (N_12446,N_12257,N_12209);
xnor U12447 (N_12447,N_12217,N_12248);
nor U12448 (N_12448,N_12220,N_12212);
or U12449 (N_12449,N_12314,N_12337);
and U12450 (N_12450,N_12213,N_12336);
xor U12451 (N_12451,N_12227,N_12229);
nor U12452 (N_12452,N_12363,N_12321);
and U12453 (N_12453,N_12342,N_12271);
and U12454 (N_12454,N_12215,N_12370);
and U12455 (N_12455,N_12362,N_12380);
and U12456 (N_12456,N_12341,N_12287);
nor U12457 (N_12457,N_12236,N_12303);
nand U12458 (N_12458,N_12319,N_12238);
nor U12459 (N_12459,N_12356,N_12324);
nor U12460 (N_12460,N_12307,N_12256);
or U12461 (N_12461,N_12385,N_12284);
and U12462 (N_12462,N_12270,N_12241);
and U12463 (N_12463,N_12339,N_12361);
or U12464 (N_12464,N_12320,N_12300);
or U12465 (N_12465,N_12204,N_12291);
nor U12466 (N_12466,N_12313,N_12309);
xor U12467 (N_12467,N_12272,N_12226);
or U12468 (N_12468,N_12317,N_12373);
xor U12469 (N_12469,N_12219,N_12332);
nand U12470 (N_12470,N_12359,N_12328);
and U12471 (N_12471,N_12292,N_12211);
nor U12472 (N_12472,N_12233,N_12282);
or U12473 (N_12473,N_12326,N_12252);
xor U12474 (N_12474,N_12395,N_12275);
nand U12475 (N_12475,N_12232,N_12386);
nor U12476 (N_12476,N_12318,N_12344);
nor U12477 (N_12477,N_12393,N_12250);
and U12478 (N_12478,N_12366,N_12306);
and U12479 (N_12479,N_12368,N_12245);
nor U12480 (N_12480,N_12258,N_12242);
xnor U12481 (N_12481,N_12369,N_12357);
nand U12482 (N_12482,N_12243,N_12310);
nand U12483 (N_12483,N_12202,N_12330);
and U12484 (N_12484,N_12274,N_12338);
nand U12485 (N_12485,N_12379,N_12207);
nor U12486 (N_12486,N_12255,N_12399);
xnor U12487 (N_12487,N_12334,N_12383);
and U12488 (N_12488,N_12348,N_12240);
xor U12489 (N_12489,N_12345,N_12294);
or U12490 (N_12490,N_12247,N_12259);
nand U12491 (N_12491,N_12396,N_12376);
nand U12492 (N_12492,N_12216,N_12312);
nor U12493 (N_12493,N_12228,N_12264);
nor U12494 (N_12494,N_12222,N_12254);
or U12495 (N_12495,N_12397,N_12218);
nor U12496 (N_12496,N_12286,N_12221);
and U12497 (N_12497,N_12296,N_12367);
nand U12498 (N_12498,N_12327,N_12333);
nor U12499 (N_12499,N_12340,N_12351);
or U12500 (N_12500,N_12265,N_12202);
nand U12501 (N_12501,N_12347,N_12252);
nor U12502 (N_12502,N_12300,N_12378);
or U12503 (N_12503,N_12258,N_12385);
xnor U12504 (N_12504,N_12333,N_12235);
or U12505 (N_12505,N_12292,N_12228);
xor U12506 (N_12506,N_12364,N_12398);
nand U12507 (N_12507,N_12311,N_12385);
or U12508 (N_12508,N_12397,N_12209);
xnor U12509 (N_12509,N_12271,N_12211);
or U12510 (N_12510,N_12300,N_12227);
nand U12511 (N_12511,N_12217,N_12393);
nor U12512 (N_12512,N_12296,N_12381);
nor U12513 (N_12513,N_12284,N_12346);
nand U12514 (N_12514,N_12309,N_12335);
or U12515 (N_12515,N_12305,N_12383);
nand U12516 (N_12516,N_12338,N_12305);
nor U12517 (N_12517,N_12224,N_12360);
and U12518 (N_12518,N_12308,N_12221);
and U12519 (N_12519,N_12234,N_12242);
nor U12520 (N_12520,N_12350,N_12377);
and U12521 (N_12521,N_12240,N_12389);
nand U12522 (N_12522,N_12335,N_12234);
and U12523 (N_12523,N_12272,N_12339);
xor U12524 (N_12524,N_12352,N_12232);
xnor U12525 (N_12525,N_12221,N_12278);
and U12526 (N_12526,N_12352,N_12258);
nor U12527 (N_12527,N_12352,N_12247);
nor U12528 (N_12528,N_12333,N_12246);
or U12529 (N_12529,N_12363,N_12229);
nand U12530 (N_12530,N_12264,N_12311);
nor U12531 (N_12531,N_12223,N_12213);
nor U12532 (N_12532,N_12203,N_12337);
nor U12533 (N_12533,N_12216,N_12383);
or U12534 (N_12534,N_12381,N_12367);
nor U12535 (N_12535,N_12229,N_12388);
nor U12536 (N_12536,N_12332,N_12260);
and U12537 (N_12537,N_12249,N_12322);
and U12538 (N_12538,N_12206,N_12232);
or U12539 (N_12539,N_12296,N_12320);
nor U12540 (N_12540,N_12299,N_12341);
nand U12541 (N_12541,N_12214,N_12344);
or U12542 (N_12542,N_12227,N_12265);
xor U12543 (N_12543,N_12259,N_12261);
or U12544 (N_12544,N_12301,N_12245);
xor U12545 (N_12545,N_12309,N_12370);
or U12546 (N_12546,N_12399,N_12273);
nor U12547 (N_12547,N_12305,N_12378);
or U12548 (N_12548,N_12347,N_12209);
and U12549 (N_12549,N_12384,N_12272);
nand U12550 (N_12550,N_12296,N_12245);
and U12551 (N_12551,N_12301,N_12390);
nor U12552 (N_12552,N_12360,N_12361);
or U12553 (N_12553,N_12223,N_12376);
nor U12554 (N_12554,N_12262,N_12257);
nand U12555 (N_12555,N_12379,N_12229);
or U12556 (N_12556,N_12222,N_12211);
xnor U12557 (N_12557,N_12336,N_12327);
and U12558 (N_12558,N_12313,N_12389);
and U12559 (N_12559,N_12346,N_12217);
nor U12560 (N_12560,N_12212,N_12290);
or U12561 (N_12561,N_12389,N_12325);
and U12562 (N_12562,N_12355,N_12226);
or U12563 (N_12563,N_12368,N_12370);
nor U12564 (N_12564,N_12374,N_12228);
nand U12565 (N_12565,N_12394,N_12346);
nor U12566 (N_12566,N_12250,N_12316);
nor U12567 (N_12567,N_12216,N_12206);
or U12568 (N_12568,N_12396,N_12288);
xor U12569 (N_12569,N_12397,N_12276);
or U12570 (N_12570,N_12357,N_12230);
or U12571 (N_12571,N_12398,N_12328);
nand U12572 (N_12572,N_12399,N_12232);
nand U12573 (N_12573,N_12345,N_12285);
or U12574 (N_12574,N_12219,N_12385);
nor U12575 (N_12575,N_12327,N_12239);
xor U12576 (N_12576,N_12332,N_12375);
and U12577 (N_12577,N_12385,N_12207);
or U12578 (N_12578,N_12212,N_12268);
nor U12579 (N_12579,N_12201,N_12365);
xnor U12580 (N_12580,N_12298,N_12261);
xnor U12581 (N_12581,N_12316,N_12284);
nand U12582 (N_12582,N_12255,N_12354);
nor U12583 (N_12583,N_12279,N_12313);
xnor U12584 (N_12584,N_12386,N_12267);
and U12585 (N_12585,N_12308,N_12303);
nand U12586 (N_12586,N_12203,N_12205);
xnor U12587 (N_12587,N_12212,N_12231);
nor U12588 (N_12588,N_12338,N_12355);
nand U12589 (N_12589,N_12304,N_12246);
or U12590 (N_12590,N_12382,N_12325);
or U12591 (N_12591,N_12385,N_12294);
xor U12592 (N_12592,N_12320,N_12218);
xor U12593 (N_12593,N_12365,N_12251);
nor U12594 (N_12594,N_12257,N_12252);
xor U12595 (N_12595,N_12251,N_12253);
nand U12596 (N_12596,N_12260,N_12393);
nor U12597 (N_12597,N_12331,N_12374);
xor U12598 (N_12598,N_12267,N_12270);
or U12599 (N_12599,N_12224,N_12290);
and U12600 (N_12600,N_12482,N_12439);
nand U12601 (N_12601,N_12431,N_12518);
xor U12602 (N_12602,N_12566,N_12499);
nor U12603 (N_12603,N_12453,N_12575);
and U12604 (N_12604,N_12533,N_12494);
nand U12605 (N_12605,N_12591,N_12587);
nand U12606 (N_12606,N_12423,N_12551);
or U12607 (N_12607,N_12586,N_12595);
nand U12608 (N_12608,N_12483,N_12414);
nand U12609 (N_12609,N_12436,N_12465);
and U12610 (N_12610,N_12401,N_12599);
nand U12611 (N_12611,N_12590,N_12450);
or U12612 (N_12612,N_12412,N_12404);
xor U12613 (N_12613,N_12448,N_12527);
nand U12614 (N_12614,N_12493,N_12457);
nor U12615 (N_12615,N_12554,N_12567);
nand U12616 (N_12616,N_12492,N_12562);
or U12617 (N_12617,N_12564,N_12498);
or U12618 (N_12618,N_12413,N_12443);
nor U12619 (N_12619,N_12503,N_12532);
nor U12620 (N_12620,N_12410,N_12469);
nand U12621 (N_12621,N_12574,N_12539);
xor U12622 (N_12622,N_12466,N_12456);
nor U12623 (N_12623,N_12534,N_12481);
and U12624 (N_12624,N_12526,N_12407);
nor U12625 (N_12625,N_12542,N_12478);
or U12626 (N_12626,N_12415,N_12546);
xor U12627 (N_12627,N_12501,N_12454);
nor U12628 (N_12628,N_12577,N_12572);
nand U12629 (N_12629,N_12479,N_12578);
xor U12630 (N_12630,N_12496,N_12514);
or U12631 (N_12631,N_12583,N_12571);
nand U12632 (N_12632,N_12523,N_12459);
xor U12633 (N_12633,N_12584,N_12568);
xnor U12634 (N_12634,N_12455,N_12506);
nor U12635 (N_12635,N_12420,N_12530);
nor U12636 (N_12636,N_12426,N_12529);
nand U12637 (N_12637,N_12405,N_12576);
nand U12638 (N_12638,N_12507,N_12408);
and U12639 (N_12639,N_12422,N_12521);
xor U12640 (N_12640,N_12561,N_12515);
xnor U12641 (N_12641,N_12419,N_12573);
nand U12642 (N_12642,N_12438,N_12589);
nor U12643 (N_12643,N_12474,N_12458);
xor U12644 (N_12644,N_12559,N_12487);
nand U12645 (N_12645,N_12430,N_12588);
or U12646 (N_12646,N_12585,N_12495);
xor U12647 (N_12647,N_12464,N_12425);
or U12648 (N_12648,N_12504,N_12557);
xor U12649 (N_12649,N_12476,N_12556);
nor U12650 (N_12650,N_12593,N_12558);
nand U12651 (N_12651,N_12490,N_12462);
and U12652 (N_12652,N_12560,N_12549);
or U12653 (N_12653,N_12524,N_12500);
xor U12654 (N_12654,N_12520,N_12475);
or U12655 (N_12655,N_12451,N_12565);
nand U12656 (N_12656,N_12536,N_12452);
nand U12657 (N_12657,N_12472,N_12429);
or U12658 (N_12658,N_12528,N_12525);
and U12659 (N_12659,N_12416,N_12547);
and U12660 (N_12660,N_12444,N_12437);
nor U12661 (N_12661,N_12411,N_12402);
nor U12662 (N_12662,N_12540,N_12489);
nor U12663 (N_12663,N_12550,N_12424);
xnor U12664 (N_12664,N_12531,N_12505);
and U12665 (N_12665,N_12517,N_12512);
nand U12666 (N_12666,N_12597,N_12509);
nor U12667 (N_12667,N_12552,N_12488);
and U12668 (N_12668,N_12511,N_12417);
or U12669 (N_12669,N_12545,N_12480);
nor U12670 (N_12670,N_12519,N_12428);
nand U12671 (N_12671,N_12409,N_12598);
nand U12672 (N_12672,N_12468,N_12470);
nand U12673 (N_12673,N_12592,N_12563);
and U12674 (N_12674,N_12442,N_12467);
and U12675 (N_12675,N_12449,N_12535);
xor U12676 (N_12676,N_12445,N_12544);
nor U12677 (N_12677,N_12516,N_12461);
xnor U12678 (N_12678,N_12460,N_12522);
nand U12679 (N_12679,N_12441,N_12579);
nand U12680 (N_12680,N_12471,N_12508);
or U12681 (N_12681,N_12497,N_12580);
and U12682 (N_12682,N_12555,N_12484);
nor U12683 (N_12683,N_12502,N_12473);
xor U12684 (N_12684,N_12491,N_12421);
nor U12685 (N_12685,N_12485,N_12513);
and U12686 (N_12686,N_12406,N_12541);
xnor U12687 (N_12687,N_12553,N_12435);
or U12688 (N_12688,N_12400,N_12582);
or U12689 (N_12689,N_12548,N_12447);
xnor U12690 (N_12690,N_12581,N_12434);
and U12691 (N_12691,N_12569,N_12486);
xnor U12692 (N_12692,N_12477,N_12427);
nor U12693 (N_12693,N_12570,N_12446);
nor U12694 (N_12694,N_12403,N_12432);
and U12695 (N_12695,N_12510,N_12543);
or U12696 (N_12696,N_12537,N_12596);
or U12697 (N_12697,N_12418,N_12538);
nand U12698 (N_12698,N_12440,N_12463);
xor U12699 (N_12699,N_12594,N_12433);
xor U12700 (N_12700,N_12578,N_12475);
xor U12701 (N_12701,N_12490,N_12447);
nand U12702 (N_12702,N_12436,N_12459);
nand U12703 (N_12703,N_12513,N_12566);
or U12704 (N_12704,N_12443,N_12406);
nand U12705 (N_12705,N_12597,N_12463);
xor U12706 (N_12706,N_12544,N_12560);
xor U12707 (N_12707,N_12482,N_12514);
nand U12708 (N_12708,N_12525,N_12534);
or U12709 (N_12709,N_12582,N_12419);
and U12710 (N_12710,N_12583,N_12433);
nand U12711 (N_12711,N_12533,N_12544);
nor U12712 (N_12712,N_12506,N_12575);
or U12713 (N_12713,N_12478,N_12559);
nor U12714 (N_12714,N_12465,N_12511);
nand U12715 (N_12715,N_12502,N_12512);
nand U12716 (N_12716,N_12573,N_12413);
and U12717 (N_12717,N_12462,N_12549);
or U12718 (N_12718,N_12440,N_12465);
nand U12719 (N_12719,N_12589,N_12541);
or U12720 (N_12720,N_12462,N_12539);
nor U12721 (N_12721,N_12472,N_12528);
nand U12722 (N_12722,N_12522,N_12413);
xor U12723 (N_12723,N_12484,N_12435);
nor U12724 (N_12724,N_12514,N_12412);
xnor U12725 (N_12725,N_12488,N_12532);
xnor U12726 (N_12726,N_12526,N_12576);
and U12727 (N_12727,N_12503,N_12497);
xnor U12728 (N_12728,N_12489,N_12582);
xor U12729 (N_12729,N_12541,N_12599);
xor U12730 (N_12730,N_12442,N_12439);
and U12731 (N_12731,N_12495,N_12490);
xor U12732 (N_12732,N_12547,N_12462);
and U12733 (N_12733,N_12471,N_12554);
or U12734 (N_12734,N_12473,N_12586);
and U12735 (N_12735,N_12565,N_12400);
or U12736 (N_12736,N_12443,N_12577);
xnor U12737 (N_12737,N_12472,N_12554);
or U12738 (N_12738,N_12540,N_12596);
or U12739 (N_12739,N_12487,N_12453);
or U12740 (N_12740,N_12443,N_12486);
nand U12741 (N_12741,N_12546,N_12520);
and U12742 (N_12742,N_12561,N_12565);
and U12743 (N_12743,N_12409,N_12506);
and U12744 (N_12744,N_12473,N_12497);
or U12745 (N_12745,N_12529,N_12513);
nor U12746 (N_12746,N_12458,N_12568);
nor U12747 (N_12747,N_12471,N_12506);
xnor U12748 (N_12748,N_12447,N_12598);
and U12749 (N_12749,N_12501,N_12561);
nor U12750 (N_12750,N_12516,N_12586);
nor U12751 (N_12751,N_12586,N_12575);
or U12752 (N_12752,N_12593,N_12455);
nand U12753 (N_12753,N_12548,N_12595);
nor U12754 (N_12754,N_12518,N_12468);
and U12755 (N_12755,N_12546,N_12446);
nand U12756 (N_12756,N_12495,N_12503);
nand U12757 (N_12757,N_12404,N_12556);
and U12758 (N_12758,N_12498,N_12537);
or U12759 (N_12759,N_12480,N_12576);
or U12760 (N_12760,N_12413,N_12503);
nor U12761 (N_12761,N_12510,N_12514);
and U12762 (N_12762,N_12500,N_12504);
nand U12763 (N_12763,N_12527,N_12479);
nor U12764 (N_12764,N_12508,N_12406);
or U12765 (N_12765,N_12589,N_12478);
xnor U12766 (N_12766,N_12562,N_12404);
xnor U12767 (N_12767,N_12569,N_12512);
xnor U12768 (N_12768,N_12548,N_12568);
and U12769 (N_12769,N_12588,N_12490);
and U12770 (N_12770,N_12476,N_12558);
xnor U12771 (N_12771,N_12476,N_12512);
xnor U12772 (N_12772,N_12531,N_12471);
and U12773 (N_12773,N_12555,N_12526);
nand U12774 (N_12774,N_12501,N_12551);
or U12775 (N_12775,N_12531,N_12588);
and U12776 (N_12776,N_12551,N_12581);
or U12777 (N_12777,N_12521,N_12512);
xnor U12778 (N_12778,N_12458,N_12469);
xor U12779 (N_12779,N_12472,N_12500);
nor U12780 (N_12780,N_12559,N_12480);
nand U12781 (N_12781,N_12580,N_12529);
or U12782 (N_12782,N_12434,N_12445);
or U12783 (N_12783,N_12515,N_12500);
nand U12784 (N_12784,N_12455,N_12542);
and U12785 (N_12785,N_12407,N_12587);
nor U12786 (N_12786,N_12459,N_12450);
xnor U12787 (N_12787,N_12542,N_12540);
nor U12788 (N_12788,N_12490,N_12404);
xor U12789 (N_12789,N_12490,N_12464);
or U12790 (N_12790,N_12440,N_12447);
nor U12791 (N_12791,N_12486,N_12577);
or U12792 (N_12792,N_12448,N_12471);
xor U12793 (N_12793,N_12442,N_12496);
xor U12794 (N_12794,N_12452,N_12460);
nor U12795 (N_12795,N_12451,N_12545);
and U12796 (N_12796,N_12587,N_12548);
xor U12797 (N_12797,N_12440,N_12489);
xnor U12798 (N_12798,N_12582,N_12436);
nor U12799 (N_12799,N_12417,N_12405);
xor U12800 (N_12800,N_12740,N_12648);
and U12801 (N_12801,N_12680,N_12709);
and U12802 (N_12802,N_12640,N_12666);
nor U12803 (N_12803,N_12627,N_12730);
or U12804 (N_12804,N_12766,N_12658);
or U12805 (N_12805,N_12732,N_12737);
nor U12806 (N_12806,N_12610,N_12634);
and U12807 (N_12807,N_12619,N_12696);
nor U12808 (N_12808,N_12644,N_12786);
nor U12809 (N_12809,N_12753,N_12655);
nor U12810 (N_12810,N_12664,N_12768);
xor U12811 (N_12811,N_12757,N_12795);
and U12812 (N_12812,N_12657,N_12659);
nor U12813 (N_12813,N_12671,N_12739);
or U12814 (N_12814,N_12710,N_12733);
nor U12815 (N_12815,N_12751,N_12780);
xor U12816 (N_12816,N_12777,N_12678);
xor U12817 (N_12817,N_12603,N_12700);
and U12818 (N_12818,N_12693,N_12701);
xnor U12819 (N_12819,N_12735,N_12705);
xnor U12820 (N_12820,N_12647,N_12774);
and U12821 (N_12821,N_12745,N_12748);
nor U12822 (N_12822,N_12677,N_12797);
or U12823 (N_12823,N_12756,N_12719);
or U12824 (N_12824,N_12681,N_12772);
nand U12825 (N_12825,N_12635,N_12622);
nor U12826 (N_12826,N_12796,N_12661);
and U12827 (N_12827,N_12702,N_12760);
or U12828 (N_12828,N_12643,N_12776);
or U12829 (N_12829,N_12688,N_12604);
or U12830 (N_12830,N_12775,N_12625);
xnor U12831 (N_12831,N_12706,N_12653);
nor U12832 (N_12832,N_12749,N_12618);
and U12833 (N_12833,N_12689,N_12788);
nand U12834 (N_12834,N_12649,N_12674);
or U12835 (N_12835,N_12752,N_12793);
nand U12836 (N_12836,N_12720,N_12743);
nand U12837 (N_12837,N_12679,N_12632);
or U12838 (N_12838,N_12767,N_12669);
xor U12839 (N_12839,N_12773,N_12642);
nor U12840 (N_12840,N_12607,N_12602);
xor U12841 (N_12841,N_12697,N_12663);
nor U12842 (N_12842,N_12790,N_12638);
and U12843 (N_12843,N_12744,N_12781);
xor U12844 (N_12844,N_12676,N_12783);
or U12845 (N_12845,N_12727,N_12721);
nor U12846 (N_12846,N_12789,N_12631);
and U12847 (N_12847,N_12763,N_12782);
nand U12848 (N_12848,N_12685,N_12765);
xnor U12849 (N_12849,N_12734,N_12755);
nand U12850 (N_12850,N_12690,N_12794);
nand U12851 (N_12851,N_12656,N_12722);
nand U12852 (N_12852,N_12724,N_12615);
nor U12853 (N_12853,N_12718,N_12723);
nand U12854 (N_12854,N_12716,N_12764);
or U12855 (N_12855,N_12707,N_12667);
or U12856 (N_12856,N_12728,N_12633);
nand U12857 (N_12857,N_12601,N_12761);
nand U12858 (N_12858,N_12683,N_12750);
and U12859 (N_12859,N_12712,N_12742);
and U12860 (N_12860,N_12637,N_12792);
xnor U12861 (N_12861,N_12620,N_12673);
or U12862 (N_12862,N_12616,N_12646);
and U12863 (N_12863,N_12628,N_12645);
and U12864 (N_12864,N_12747,N_12798);
xor U12865 (N_12865,N_12762,N_12626);
nand U12866 (N_12866,N_12713,N_12746);
nand U12867 (N_12867,N_12699,N_12726);
or U12868 (N_12868,N_12729,N_12686);
and U12869 (N_12869,N_12731,N_12769);
and U12870 (N_12870,N_12652,N_12738);
or U12871 (N_12871,N_12695,N_12668);
nor U12872 (N_12872,N_12791,N_12670);
and U12873 (N_12873,N_12609,N_12708);
xnor U12874 (N_12874,N_12606,N_12660);
nand U12875 (N_12875,N_12629,N_12665);
nand U12876 (N_12876,N_12799,N_12758);
and U12877 (N_12877,N_12711,N_12600);
nand U12878 (N_12878,N_12613,N_12617);
or U12879 (N_12879,N_12698,N_12771);
nand U12880 (N_12880,N_12741,N_12694);
nor U12881 (N_12881,N_12641,N_12784);
or U12882 (N_12882,N_12630,N_12687);
and U12883 (N_12883,N_12611,N_12736);
and U12884 (N_12884,N_12787,N_12682);
xnor U12885 (N_12885,N_12650,N_12759);
nand U12886 (N_12886,N_12614,N_12624);
nor U12887 (N_12887,N_12639,N_12691);
nand U12888 (N_12888,N_12675,N_12651);
xor U12889 (N_12889,N_12779,N_12605);
or U12890 (N_12890,N_12754,N_12704);
or U12891 (N_12891,N_12612,N_12715);
or U12892 (N_12892,N_12717,N_12770);
or U12893 (N_12893,N_12672,N_12692);
or U12894 (N_12894,N_12636,N_12785);
and U12895 (N_12895,N_12778,N_12662);
and U12896 (N_12896,N_12714,N_12654);
nor U12897 (N_12897,N_12725,N_12684);
or U12898 (N_12898,N_12608,N_12621);
xor U12899 (N_12899,N_12703,N_12623);
and U12900 (N_12900,N_12663,N_12656);
nand U12901 (N_12901,N_12741,N_12663);
and U12902 (N_12902,N_12732,N_12727);
nand U12903 (N_12903,N_12716,N_12622);
xor U12904 (N_12904,N_12649,N_12764);
xnor U12905 (N_12905,N_12697,N_12690);
xnor U12906 (N_12906,N_12775,N_12607);
and U12907 (N_12907,N_12761,N_12727);
nor U12908 (N_12908,N_12692,N_12724);
or U12909 (N_12909,N_12740,N_12792);
and U12910 (N_12910,N_12638,N_12720);
xnor U12911 (N_12911,N_12699,N_12647);
xnor U12912 (N_12912,N_12611,N_12794);
and U12913 (N_12913,N_12726,N_12632);
xnor U12914 (N_12914,N_12608,N_12730);
nand U12915 (N_12915,N_12610,N_12609);
and U12916 (N_12916,N_12786,N_12682);
and U12917 (N_12917,N_12720,N_12681);
or U12918 (N_12918,N_12755,N_12692);
xnor U12919 (N_12919,N_12772,N_12784);
nand U12920 (N_12920,N_12745,N_12795);
nor U12921 (N_12921,N_12780,N_12722);
and U12922 (N_12922,N_12778,N_12681);
nand U12923 (N_12923,N_12769,N_12782);
nor U12924 (N_12924,N_12733,N_12633);
xnor U12925 (N_12925,N_12681,N_12714);
nor U12926 (N_12926,N_12672,N_12694);
and U12927 (N_12927,N_12727,N_12794);
or U12928 (N_12928,N_12682,N_12706);
nand U12929 (N_12929,N_12744,N_12684);
or U12930 (N_12930,N_12724,N_12610);
xnor U12931 (N_12931,N_12634,N_12779);
nand U12932 (N_12932,N_12715,N_12702);
and U12933 (N_12933,N_12792,N_12679);
xnor U12934 (N_12934,N_12618,N_12706);
nand U12935 (N_12935,N_12624,N_12647);
nor U12936 (N_12936,N_12667,N_12761);
nand U12937 (N_12937,N_12630,N_12625);
nand U12938 (N_12938,N_12717,N_12788);
and U12939 (N_12939,N_12792,N_12779);
and U12940 (N_12940,N_12666,N_12752);
xnor U12941 (N_12941,N_12725,N_12700);
nand U12942 (N_12942,N_12790,N_12688);
xor U12943 (N_12943,N_12634,N_12609);
nand U12944 (N_12944,N_12792,N_12647);
nand U12945 (N_12945,N_12657,N_12716);
nor U12946 (N_12946,N_12641,N_12675);
xor U12947 (N_12947,N_12603,N_12703);
nor U12948 (N_12948,N_12724,N_12634);
and U12949 (N_12949,N_12671,N_12696);
or U12950 (N_12950,N_12652,N_12762);
xor U12951 (N_12951,N_12676,N_12795);
nor U12952 (N_12952,N_12671,N_12689);
nand U12953 (N_12953,N_12712,N_12631);
or U12954 (N_12954,N_12733,N_12743);
nor U12955 (N_12955,N_12774,N_12784);
xnor U12956 (N_12956,N_12797,N_12625);
nand U12957 (N_12957,N_12606,N_12791);
or U12958 (N_12958,N_12739,N_12775);
and U12959 (N_12959,N_12681,N_12607);
xnor U12960 (N_12960,N_12710,N_12674);
and U12961 (N_12961,N_12676,N_12758);
nor U12962 (N_12962,N_12657,N_12655);
nand U12963 (N_12963,N_12604,N_12730);
xor U12964 (N_12964,N_12601,N_12787);
xor U12965 (N_12965,N_12756,N_12710);
nor U12966 (N_12966,N_12777,N_12634);
xnor U12967 (N_12967,N_12753,N_12632);
nand U12968 (N_12968,N_12704,N_12742);
xnor U12969 (N_12969,N_12731,N_12753);
nand U12970 (N_12970,N_12698,N_12678);
and U12971 (N_12971,N_12754,N_12779);
xor U12972 (N_12972,N_12602,N_12654);
and U12973 (N_12973,N_12695,N_12745);
xnor U12974 (N_12974,N_12778,N_12646);
nor U12975 (N_12975,N_12655,N_12728);
nand U12976 (N_12976,N_12660,N_12724);
xor U12977 (N_12977,N_12731,N_12618);
nand U12978 (N_12978,N_12693,N_12740);
nand U12979 (N_12979,N_12601,N_12686);
nor U12980 (N_12980,N_12791,N_12782);
or U12981 (N_12981,N_12661,N_12795);
nor U12982 (N_12982,N_12724,N_12686);
nand U12983 (N_12983,N_12759,N_12791);
and U12984 (N_12984,N_12616,N_12750);
or U12985 (N_12985,N_12678,N_12683);
or U12986 (N_12986,N_12655,N_12603);
nand U12987 (N_12987,N_12760,N_12643);
xnor U12988 (N_12988,N_12769,N_12642);
xnor U12989 (N_12989,N_12769,N_12724);
and U12990 (N_12990,N_12757,N_12777);
or U12991 (N_12991,N_12735,N_12701);
xnor U12992 (N_12992,N_12786,N_12788);
nand U12993 (N_12993,N_12718,N_12755);
and U12994 (N_12994,N_12781,N_12647);
nor U12995 (N_12995,N_12740,N_12602);
nor U12996 (N_12996,N_12605,N_12680);
and U12997 (N_12997,N_12687,N_12773);
xor U12998 (N_12998,N_12749,N_12681);
nand U12999 (N_12999,N_12717,N_12637);
nor U13000 (N_13000,N_12954,N_12843);
xnor U13001 (N_13001,N_12888,N_12913);
nand U13002 (N_13002,N_12946,N_12941);
or U13003 (N_13003,N_12898,N_12902);
or U13004 (N_13004,N_12829,N_12915);
or U13005 (N_13005,N_12921,N_12933);
xnor U13006 (N_13006,N_12849,N_12998);
nand U13007 (N_13007,N_12992,N_12995);
nor U13008 (N_13008,N_12863,N_12821);
and U13009 (N_13009,N_12800,N_12834);
or U13010 (N_13010,N_12872,N_12825);
and U13011 (N_13011,N_12994,N_12894);
or U13012 (N_13012,N_12895,N_12973);
and U13013 (N_13013,N_12847,N_12929);
xor U13014 (N_13014,N_12855,N_12832);
or U13015 (N_13015,N_12873,N_12835);
nand U13016 (N_13016,N_12807,N_12885);
nor U13017 (N_13017,N_12963,N_12896);
xor U13018 (N_13018,N_12818,N_12842);
or U13019 (N_13019,N_12904,N_12986);
nor U13020 (N_13020,N_12866,N_12816);
nor U13021 (N_13021,N_12813,N_12822);
nor U13022 (N_13022,N_12841,N_12903);
xnor U13023 (N_13023,N_12809,N_12999);
nor U13024 (N_13024,N_12907,N_12938);
nor U13025 (N_13025,N_12910,N_12922);
xor U13026 (N_13026,N_12893,N_12943);
xor U13027 (N_13027,N_12955,N_12857);
nand U13028 (N_13028,N_12883,N_12852);
nand U13029 (N_13029,N_12959,N_12856);
and U13030 (N_13030,N_12846,N_12936);
nor U13031 (N_13031,N_12909,N_12826);
and U13032 (N_13032,N_12869,N_12905);
or U13033 (N_13033,N_12802,N_12871);
and U13034 (N_13034,N_12882,N_12947);
nand U13035 (N_13035,N_12950,N_12874);
xor U13036 (N_13036,N_12880,N_12984);
and U13037 (N_13037,N_12952,N_12976);
or U13038 (N_13038,N_12981,N_12948);
nor U13039 (N_13039,N_12930,N_12931);
or U13040 (N_13040,N_12879,N_12912);
and U13041 (N_13041,N_12836,N_12853);
xnor U13042 (N_13042,N_12820,N_12977);
nor U13043 (N_13043,N_12899,N_12969);
nand U13044 (N_13044,N_12801,N_12953);
nand U13045 (N_13045,N_12886,N_12850);
nand U13046 (N_13046,N_12889,N_12861);
nor U13047 (N_13047,N_12840,N_12810);
nand U13048 (N_13048,N_12958,N_12854);
and U13049 (N_13049,N_12927,N_12827);
nand U13050 (N_13050,N_12925,N_12876);
xor U13051 (N_13051,N_12900,N_12877);
or U13052 (N_13052,N_12970,N_12972);
or U13053 (N_13053,N_12911,N_12919);
xor U13054 (N_13054,N_12917,N_12937);
nor U13055 (N_13055,N_12916,N_12993);
nand U13056 (N_13056,N_12858,N_12859);
or U13057 (N_13057,N_12860,N_12942);
nor U13058 (N_13058,N_12983,N_12920);
or U13059 (N_13059,N_12828,N_12837);
nand U13060 (N_13060,N_12965,N_12814);
nand U13061 (N_13061,N_12803,N_12817);
and U13062 (N_13062,N_12906,N_12957);
nand U13063 (N_13063,N_12908,N_12932);
or U13064 (N_13064,N_12940,N_12838);
and U13065 (N_13065,N_12926,N_12956);
or U13066 (N_13066,N_12812,N_12923);
and U13067 (N_13067,N_12968,N_12996);
xnor U13068 (N_13068,N_12960,N_12845);
nor U13069 (N_13069,N_12980,N_12951);
xor U13070 (N_13070,N_12833,N_12804);
or U13071 (N_13071,N_12862,N_12945);
or U13072 (N_13072,N_12979,N_12808);
nor U13073 (N_13073,N_12978,N_12966);
nand U13074 (N_13074,N_12875,N_12939);
xor U13075 (N_13075,N_12997,N_12867);
nand U13076 (N_13076,N_12897,N_12824);
or U13077 (N_13077,N_12971,N_12935);
nand U13078 (N_13078,N_12878,N_12844);
and U13079 (N_13079,N_12865,N_12988);
xor U13080 (N_13080,N_12918,N_12962);
nand U13081 (N_13081,N_12864,N_12839);
or U13082 (N_13082,N_12914,N_12901);
nor U13083 (N_13083,N_12848,N_12884);
or U13084 (N_13084,N_12815,N_12819);
or U13085 (N_13085,N_12891,N_12868);
or U13086 (N_13086,N_12989,N_12934);
nand U13087 (N_13087,N_12924,N_12928);
nand U13088 (N_13088,N_12991,N_12887);
xor U13089 (N_13089,N_12881,N_12967);
and U13090 (N_13090,N_12944,N_12982);
nand U13091 (N_13091,N_12974,N_12990);
nor U13092 (N_13092,N_12985,N_12830);
and U13093 (N_13093,N_12851,N_12961);
and U13094 (N_13094,N_12890,N_12949);
and U13095 (N_13095,N_12831,N_12892);
and U13096 (N_13096,N_12805,N_12811);
and U13097 (N_13097,N_12964,N_12975);
xnor U13098 (N_13098,N_12987,N_12806);
xor U13099 (N_13099,N_12870,N_12823);
xnor U13100 (N_13100,N_12899,N_12921);
nor U13101 (N_13101,N_12868,N_12853);
nor U13102 (N_13102,N_12989,N_12804);
nand U13103 (N_13103,N_12984,N_12849);
nand U13104 (N_13104,N_12925,N_12989);
xnor U13105 (N_13105,N_12832,N_12856);
xnor U13106 (N_13106,N_12922,N_12810);
xor U13107 (N_13107,N_12961,N_12981);
or U13108 (N_13108,N_12989,N_12943);
and U13109 (N_13109,N_12902,N_12958);
or U13110 (N_13110,N_12854,N_12997);
and U13111 (N_13111,N_12914,N_12852);
xnor U13112 (N_13112,N_12942,N_12890);
and U13113 (N_13113,N_12949,N_12933);
or U13114 (N_13114,N_12850,N_12820);
nor U13115 (N_13115,N_12966,N_12800);
or U13116 (N_13116,N_12837,N_12804);
nor U13117 (N_13117,N_12952,N_12914);
nand U13118 (N_13118,N_12936,N_12838);
nand U13119 (N_13119,N_12930,N_12991);
or U13120 (N_13120,N_12985,N_12954);
nor U13121 (N_13121,N_12939,N_12935);
nor U13122 (N_13122,N_12974,N_12972);
nand U13123 (N_13123,N_12969,N_12916);
and U13124 (N_13124,N_12919,N_12848);
xnor U13125 (N_13125,N_12966,N_12865);
xnor U13126 (N_13126,N_12919,N_12844);
nand U13127 (N_13127,N_12805,N_12907);
and U13128 (N_13128,N_12802,N_12944);
nor U13129 (N_13129,N_12990,N_12912);
xnor U13130 (N_13130,N_12933,N_12972);
xnor U13131 (N_13131,N_12801,N_12928);
or U13132 (N_13132,N_12950,N_12847);
nand U13133 (N_13133,N_12836,N_12924);
xor U13134 (N_13134,N_12868,N_12818);
or U13135 (N_13135,N_12992,N_12943);
or U13136 (N_13136,N_12932,N_12937);
and U13137 (N_13137,N_12976,N_12906);
and U13138 (N_13138,N_12959,N_12991);
or U13139 (N_13139,N_12804,N_12992);
nand U13140 (N_13140,N_12921,N_12823);
nor U13141 (N_13141,N_12993,N_12871);
nor U13142 (N_13142,N_12930,N_12901);
nand U13143 (N_13143,N_12885,N_12854);
nor U13144 (N_13144,N_12903,N_12896);
nor U13145 (N_13145,N_12936,N_12856);
and U13146 (N_13146,N_12951,N_12991);
nand U13147 (N_13147,N_12925,N_12961);
xnor U13148 (N_13148,N_12910,N_12833);
and U13149 (N_13149,N_12880,N_12858);
and U13150 (N_13150,N_12936,N_12908);
nor U13151 (N_13151,N_12829,N_12981);
nor U13152 (N_13152,N_12928,N_12998);
or U13153 (N_13153,N_12878,N_12997);
xnor U13154 (N_13154,N_12973,N_12845);
nand U13155 (N_13155,N_12819,N_12808);
nand U13156 (N_13156,N_12911,N_12941);
or U13157 (N_13157,N_12933,N_12968);
xnor U13158 (N_13158,N_12870,N_12878);
xor U13159 (N_13159,N_12921,N_12894);
nor U13160 (N_13160,N_12977,N_12933);
nand U13161 (N_13161,N_12930,N_12938);
nand U13162 (N_13162,N_12852,N_12953);
and U13163 (N_13163,N_12971,N_12870);
xor U13164 (N_13164,N_12930,N_12890);
nand U13165 (N_13165,N_12884,N_12978);
or U13166 (N_13166,N_12969,N_12835);
or U13167 (N_13167,N_12946,N_12990);
xor U13168 (N_13168,N_12967,N_12841);
or U13169 (N_13169,N_12812,N_12826);
and U13170 (N_13170,N_12995,N_12825);
nand U13171 (N_13171,N_12857,N_12915);
nand U13172 (N_13172,N_12825,N_12854);
nand U13173 (N_13173,N_12992,N_12882);
and U13174 (N_13174,N_12821,N_12997);
or U13175 (N_13175,N_12878,N_12854);
nor U13176 (N_13176,N_12979,N_12977);
xor U13177 (N_13177,N_12820,N_12880);
nor U13178 (N_13178,N_12863,N_12927);
nor U13179 (N_13179,N_12852,N_12867);
xor U13180 (N_13180,N_12962,N_12952);
nor U13181 (N_13181,N_12964,N_12984);
nand U13182 (N_13182,N_12921,N_12833);
nor U13183 (N_13183,N_12884,N_12968);
xnor U13184 (N_13184,N_12848,N_12880);
xor U13185 (N_13185,N_12867,N_12843);
and U13186 (N_13186,N_12938,N_12801);
and U13187 (N_13187,N_12922,N_12817);
and U13188 (N_13188,N_12907,N_12945);
or U13189 (N_13189,N_12801,N_12807);
nor U13190 (N_13190,N_12905,N_12884);
xor U13191 (N_13191,N_12901,N_12935);
xor U13192 (N_13192,N_12872,N_12837);
nand U13193 (N_13193,N_12846,N_12965);
xnor U13194 (N_13194,N_12891,N_12948);
nor U13195 (N_13195,N_12961,N_12977);
nand U13196 (N_13196,N_12988,N_12874);
xor U13197 (N_13197,N_12942,N_12846);
nor U13198 (N_13198,N_12961,N_12861);
or U13199 (N_13199,N_12851,N_12844);
xor U13200 (N_13200,N_13033,N_13065);
nor U13201 (N_13201,N_13183,N_13043);
nand U13202 (N_13202,N_13025,N_13071);
or U13203 (N_13203,N_13160,N_13187);
or U13204 (N_13204,N_13079,N_13013);
and U13205 (N_13205,N_13092,N_13045);
or U13206 (N_13206,N_13139,N_13036);
nor U13207 (N_13207,N_13007,N_13067);
and U13208 (N_13208,N_13099,N_13185);
xor U13209 (N_13209,N_13156,N_13031);
nand U13210 (N_13210,N_13129,N_13095);
or U13211 (N_13211,N_13080,N_13035);
nor U13212 (N_13212,N_13094,N_13073);
and U13213 (N_13213,N_13093,N_13141);
xnor U13214 (N_13214,N_13090,N_13006);
or U13215 (N_13215,N_13164,N_13062);
nor U13216 (N_13216,N_13127,N_13197);
or U13217 (N_13217,N_13102,N_13049);
nor U13218 (N_13218,N_13168,N_13017);
xnor U13219 (N_13219,N_13146,N_13148);
or U13220 (N_13220,N_13174,N_13053);
nor U13221 (N_13221,N_13177,N_13181);
and U13222 (N_13222,N_13042,N_13170);
and U13223 (N_13223,N_13110,N_13172);
nand U13224 (N_13224,N_13015,N_13107);
xor U13225 (N_13225,N_13122,N_13149);
nor U13226 (N_13226,N_13037,N_13081);
and U13227 (N_13227,N_13039,N_13186);
and U13228 (N_13228,N_13176,N_13109);
xor U13229 (N_13229,N_13084,N_13001);
and U13230 (N_13230,N_13135,N_13184);
nor U13231 (N_13231,N_13004,N_13194);
xor U13232 (N_13232,N_13152,N_13008);
nand U13233 (N_13233,N_13047,N_13024);
nor U13234 (N_13234,N_13096,N_13151);
nor U13235 (N_13235,N_13161,N_13076);
nor U13236 (N_13236,N_13121,N_13022);
nand U13237 (N_13237,N_13182,N_13021);
nor U13238 (N_13238,N_13190,N_13173);
nor U13239 (N_13239,N_13113,N_13027);
or U13240 (N_13240,N_13191,N_13188);
xor U13241 (N_13241,N_13050,N_13126);
or U13242 (N_13242,N_13055,N_13012);
xnor U13243 (N_13243,N_13124,N_13128);
and U13244 (N_13244,N_13167,N_13005);
nand U13245 (N_13245,N_13023,N_13058);
nand U13246 (N_13246,N_13030,N_13054);
nand U13247 (N_13247,N_13142,N_13180);
and U13248 (N_13248,N_13166,N_13154);
and U13249 (N_13249,N_13087,N_13145);
or U13250 (N_13250,N_13150,N_13046);
and U13251 (N_13251,N_13100,N_13175);
and U13252 (N_13252,N_13002,N_13134);
nand U13253 (N_13253,N_13153,N_13178);
nor U13254 (N_13254,N_13020,N_13018);
nor U13255 (N_13255,N_13119,N_13086);
nor U13256 (N_13256,N_13059,N_13069);
nand U13257 (N_13257,N_13196,N_13014);
nor U13258 (N_13258,N_13157,N_13130);
nand U13259 (N_13259,N_13143,N_13116);
and U13260 (N_13260,N_13057,N_13105);
or U13261 (N_13261,N_13044,N_13041);
nand U13262 (N_13262,N_13040,N_13104);
and U13263 (N_13263,N_13078,N_13179);
nand U13264 (N_13264,N_13155,N_13066);
xor U13265 (N_13265,N_13159,N_13101);
or U13266 (N_13266,N_13068,N_13098);
and U13267 (N_13267,N_13028,N_13077);
or U13268 (N_13268,N_13097,N_13140);
and U13269 (N_13269,N_13034,N_13112);
xnor U13270 (N_13270,N_13011,N_13199);
or U13271 (N_13271,N_13195,N_13082);
nand U13272 (N_13272,N_13048,N_13147);
xor U13273 (N_13273,N_13000,N_13009);
and U13274 (N_13274,N_13026,N_13131);
or U13275 (N_13275,N_13019,N_13192);
nand U13276 (N_13276,N_13123,N_13075);
nor U13277 (N_13277,N_13138,N_13029);
xnor U13278 (N_13278,N_13072,N_13118);
xnor U13279 (N_13279,N_13060,N_13106);
xor U13280 (N_13280,N_13074,N_13117);
and U13281 (N_13281,N_13137,N_13125);
nand U13282 (N_13282,N_13165,N_13056);
and U13283 (N_13283,N_13114,N_13169);
xor U13284 (N_13284,N_13193,N_13061);
nor U13285 (N_13285,N_13133,N_13120);
or U13286 (N_13286,N_13115,N_13162);
nand U13287 (N_13287,N_13198,N_13158);
nor U13288 (N_13288,N_13111,N_13083);
xor U13289 (N_13289,N_13070,N_13064);
nor U13290 (N_13290,N_13136,N_13171);
xnor U13291 (N_13291,N_13038,N_13010);
xnor U13292 (N_13292,N_13051,N_13063);
nand U13293 (N_13293,N_13052,N_13189);
nor U13294 (N_13294,N_13089,N_13088);
and U13295 (N_13295,N_13163,N_13091);
or U13296 (N_13296,N_13032,N_13016);
xnor U13297 (N_13297,N_13132,N_13003);
or U13298 (N_13298,N_13144,N_13103);
xor U13299 (N_13299,N_13108,N_13085);
nor U13300 (N_13300,N_13037,N_13000);
xor U13301 (N_13301,N_13128,N_13069);
xor U13302 (N_13302,N_13068,N_13130);
nor U13303 (N_13303,N_13018,N_13121);
xnor U13304 (N_13304,N_13037,N_13120);
nand U13305 (N_13305,N_13030,N_13145);
and U13306 (N_13306,N_13141,N_13021);
nor U13307 (N_13307,N_13186,N_13118);
nand U13308 (N_13308,N_13184,N_13048);
and U13309 (N_13309,N_13037,N_13119);
xnor U13310 (N_13310,N_13120,N_13188);
and U13311 (N_13311,N_13126,N_13080);
or U13312 (N_13312,N_13032,N_13010);
nand U13313 (N_13313,N_13062,N_13087);
and U13314 (N_13314,N_13110,N_13092);
or U13315 (N_13315,N_13092,N_13193);
nor U13316 (N_13316,N_13192,N_13056);
xor U13317 (N_13317,N_13070,N_13000);
nor U13318 (N_13318,N_13086,N_13017);
or U13319 (N_13319,N_13092,N_13156);
xnor U13320 (N_13320,N_13118,N_13176);
xor U13321 (N_13321,N_13190,N_13054);
and U13322 (N_13322,N_13130,N_13023);
xor U13323 (N_13323,N_13174,N_13035);
nor U13324 (N_13324,N_13061,N_13175);
nor U13325 (N_13325,N_13100,N_13051);
and U13326 (N_13326,N_13118,N_13101);
xnor U13327 (N_13327,N_13029,N_13133);
nand U13328 (N_13328,N_13084,N_13170);
or U13329 (N_13329,N_13056,N_13129);
or U13330 (N_13330,N_13183,N_13036);
nor U13331 (N_13331,N_13036,N_13144);
nand U13332 (N_13332,N_13196,N_13142);
nand U13333 (N_13333,N_13116,N_13031);
xnor U13334 (N_13334,N_13188,N_13057);
or U13335 (N_13335,N_13039,N_13022);
nand U13336 (N_13336,N_13171,N_13124);
nand U13337 (N_13337,N_13133,N_13041);
xnor U13338 (N_13338,N_13098,N_13008);
nand U13339 (N_13339,N_13119,N_13004);
nand U13340 (N_13340,N_13123,N_13138);
and U13341 (N_13341,N_13054,N_13095);
or U13342 (N_13342,N_13060,N_13081);
xor U13343 (N_13343,N_13185,N_13088);
and U13344 (N_13344,N_13002,N_13160);
nand U13345 (N_13345,N_13145,N_13157);
xnor U13346 (N_13346,N_13031,N_13068);
or U13347 (N_13347,N_13124,N_13182);
nand U13348 (N_13348,N_13129,N_13158);
and U13349 (N_13349,N_13042,N_13178);
xor U13350 (N_13350,N_13080,N_13002);
and U13351 (N_13351,N_13153,N_13048);
or U13352 (N_13352,N_13188,N_13076);
nand U13353 (N_13353,N_13147,N_13178);
or U13354 (N_13354,N_13164,N_13101);
xnor U13355 (N_13355,N_13072,N_13140);
and U13356 (N_13356,N_13097,N_13025);
xor U13357 (N_13357,N_13065,N_13168);
nor U13358 (N_13358,N_13104,N_13133);
or U13359 (N_13359,N_13007,N_13101);
xnor U13360 (N_13360,N_13133,N_13124);
and U13361 (N_13361,N_13142,N_13011);
and U13362 (N_13362,N_13171,N_13147);
or U13363 (N_13363,N_13124,N_13030);
nand U13364 (N_13364,N_13142,N_13169);
nand U13365 (N_13365,N_13031,N_13088);
nand U13366 (N_13366,N_13075,N_13192);
nand U13367 (N_13367,N_13080,N_13191);
xor U13368 (N_13368,N_13118,N_13150);
nand U13369 (N_13369,N_13088,N_13039);
nand U13370 (N_13370,N_13155,N_13077);
and U13371 (N_13371,N_13137,N_13144);
xor U13372 (N_13372,N_13130,N_13009);
xnor U13373 (N_13373,N_13024,N_13001);
nand U13374 (N_13374,N_13013,N_13167);
nand U13375 (N_13375,N_13157,N_13170);
nand U13376 (N_13376,N_13023,N_13119);
nand U13377 (N_13377,N_13014,N_13075);
and U13378 (N_13378,N_13173,N_13089);
nor U13379 (N_13379,N_13137,N_13196);
xor U13380 (N_13380,N_13074,N_13100);
nand U13381 (N_13381,N_13142,N_13106);
nand U13382 (N_13382,N_13185,N_13130);
or U13383 (N_13383,N_13166,N_13077);
or U13384 (N_13384,N_13180,N_13149);
xor U13385 (N_13385,N_13176,N_13062);
xnor U13386 (N_13386,N_13036,N_13008);
and U13387 (N_13387,N_13196,N_13167);
or U13388 (N_13388,N_13075,N_13040);
nor U13389 (N_13389,N_13051,N_13074);
nand U13390 (N_13390,N_13066,N_13187);
xnor U13391 (N_13391,N_13051,N_13028);
nand U13392 (N_13392,N_13057,N_13195);
xor U13393 (N_13393,N_13158,N_13042);
and U13394 (N_13394,N_13064,N_13102);
nor U13395 (N_13395,N_13133,N_13011);
xor U13396 (N_13396,N_13094,N_13000);
and U13397 (N_13397,N_13189,N_13108);
xor U13398 (N_13398,N_13026,N_13098);
and U13399 (N_13399,N_13075,N_13035);
and U13400 (N_13400,N_13277,N_13358);
or U13401 (N_13401,N_13205,N_13363);
and U13402 (N_13402,N_13333,N_13236);
nand U13403 (N_13403,N_13290,N_13383);
nor U13404 (N_13404,N_13304,N_13227);
xnor U13405 (N_13405,N_13356,N_13281);
and U13406 (N_13406,N_13334,N_13272);
nand U13407 (N_13407,N_13286,N_13246);
or U13408 (N_13408,N_13287,N_13251);
nand U13409 (N_13409,N_13395,N_13342);
xnor U13410 (N_13410,N_13374,N_13391);
and U13411 (N_13411,N_13359,N_13347);
xor U13412 (N_13412,N_13259,N_13309);
xor U13413 (N_13413,N_13206,N_13376);
nand U13414 (N_13414,N_13295,N_13280);
and U13415 (N_13415,N_13232,N_13297);
nor U13416 (N_13416,N_13241,N_13300);
xnor U13417 (N_13417,N_13312,N_13266);
xor U13418 (N_13418,N_13323,N_13217);
or U13419 (N_13419,N_13252,N_13273);
and U13420 (N_13420,N_13394,N_13382);
nor U13421 (N_13421,N_13220,N_13344);
or U13422 (N_13422,N_13293,N_13262);
nor U13423 (N_13423,N_13341,N_13263);
nor U13424 (N_13424,N_13257,N_13306);
xor U13425 (N_13425,N_13317,N_13237);
nand U13426 (N_13426,N_13310,N_13330);
and U13427 (N_13427,N_13329,N_13243);
nor U13428 (N_13428,N_13201,N_13324);
nand U13429 (N_13429,N_13238,N_13279);
xnor U13430 (N_13430,N_13360,N_13392);
nand U13431 (N_13431,N_13260,N_13299);
nand U13432 (N_13432,N_13223,N_13292);
nand U13433 (N_13433,N_13221,N_13276);
xor U13434 (N_13434,N_13255,N_13319);
and U13435 (N_13435,N_13332,N_13393);
nand U13436 (N_13436,N_13216,N_13240);
nor U13437 (N_13437,N_13322,N_13224);
xnor U13438 (N_13438,N_13225,N_13364);
nand U13439 (N_13439,N_13313,N_13242);
or U13440 (N_13440,N_13235,N_13307);
xor U13441 (N_13441,N_13267,N_13381);
xor U13442 (N_13442,N_13222,N_13377);
and U13443 (N_13443,N_13315,N_13369);
xnor U13444 (N_13444,N_13375,N_13254);
xnor U13445 (N_13445,N_13208,N_13202);
or U13446 (N_13446,N_13314,N_13250);
xnor U13447 (N_13447,N_13229,N_13239);
nor U13448 (N_13448,N_13284,N_13361);
nor U13449 (N_13449,N_13302,N_13389);
nor U13450 (N_13450,N_13219,N_13349);
and U13451 (N_13451,N_13270,N_13214);
and U13452 (N_13452,N_13207,N_13268);
nand U13453 (N_13453,N_13289,N_13283);
xor U13454 (N_13454,N_13303,N_13388);
nor U13455 (N_13455,N_13210,N_13366);
xor U13456 (N_13456,N_13230,N_13340);
nor U13457 (N_13457,N_13288,N_13275);
nand U13458 (N_13458,N_13212,N_13348);
nand U13459 (N_13459,N_13327,N_13269);
xnor U13460 (N_13460,N_13271,N_13218);
and U13461 (N_13461,N_13355,N_13367);
nor U13462 (N_13462,N_13245,N_13397);
nand U13463 (N_13463,N_13248,N_13370);
nand U13464 (N_13464,N_13265,N_13291);
xnor U13465 (N_13465,N_13211,N_13213);
and U13466 (N_13466,N_13357,N_13249);
nand U13467 (N_13467,N_13311,N_13371);
nand U13468 (N_13468,N_13261,N_13379);
and U13469 (N_13469,N_13244,N_13373);
or U13470 (N_13470,N_13350,N_13256);
or U13471 (N_13471,N_13346,N_13321);
xnor U13472 (N_13472,N_13386,N_13320);
xor U13473 (N_13473,N_13233,N_13234);
or U13474 (N_13474,N_13301,N_13226);
xnor U13475 (N_13475,N_13231,N_13296);
and U13476 (N_13476,N_13353,N_13343);
nand U13477 (N_13477,N_13345,N_13352);
and U13478 (N_13478,N_13305,N_13318);
and U13479 (N_13479,N_13247,N_13351);
nand U13480 (N_13480,N_13274,N_13316);
nor U13481 (N_13481,N_13325,N_13203);
and U13482 (N_13482,N_13282,N_13336);
and U13483 (N_13483,N_13278,N_13258);
nand U13484 (N_13484,N_13285,N_13384);
xnor U13485 (N_13485,N_13365,N_13339);
or U13486 (N_13486,N_13308,N_13387);
nor U13487 (N_13487,N_13380,N_13362);
or U13488 (N_13488,N_13204,N_13372);
or U13489 (N_13489,N_13354,N_13368);
nand U13490 (N_13490,N_13328,N_13399);
and U13491 (N_13491,N_13298,N_13200);
nor U13492 (N_13492,N_13378,N_13337);
nand U13493 (N_13493,N_13331,N_13335);
and U13494 (N_13494,N_13253,N_13228);
nand U13495 (N_13495,N_13209,N_13338);
and U13496 (N_13496,N_13390,N_13396);
and U13497 (N_13497,N_13264,N_13215);
and U13498 (N_13498,N_13326,N_13294);
or U13499 (N_13499,N_13398,N_13385);
and U13500 (N_13500,N_13214,N_13315);
nand U13501 (N_13501,N_13370,N_13268);
nor U13502 (N_13502,N_13257,N_13377);
nand U13503 (N_13503,N_13261,N_13224);
nand U13504 (N_13504,N_13303,N_13270);
xnor U13505 (N_13505,N_13377,N_13298);
and U13506 (N_13506,N_13281,N_13284);
nand U13507 (N_13507,N_13283,N_13397);
nor U13508 (N_13508,N_13364,N_13393);
xor U13509 (N_13509,N_13340,N_13359);
and U13510 (N_13510,N_13305,N_13313);
nand U13511 (N_13511,N_13240,N_13220);
nor U13512 (N_13512,N_13373,N_13237);
or U13513 (N_13513,N_13363,N_13269);
nand U13514 (N_13514,N_13299,N_13339);
and U13515 (N_13515,N_13212,N_13239);
nor U13516 (N_13516,N_13358,N_13359);
nor U13517 (N_13517,N_13373,N_13365);
nor U13518 (N_13518,N_13303,N_13344);
nor U13519 (N_13519,N_13216,N_13291);
and U13520 (N_13520,N_13251,N_13384);
and U13521 (N_13521,N_13289,N_13301);
or U13522 (N_13522,N_13339,N_13352);
nor U13523 (N_13523,N_13379,N_13222);
and U13524 (N_13524,N_13338,N_13202);
nor U13525 (N_13525,N_13350,N_13281);
nand U13526 (N_13526,N_13278,N_13326);
nand U13527 (N_13527,N_13276,N_13384);
xor U13528 (N_13528,N_13369,N_13358);
xnor U13529 (N_13529,N_13266,N_13307);
nand U13530 (N_13530,N_13287,N_13296);
nand U13531 (N_13531,N_13262,N_13239);
xor U13532 (N_13532,N_13271,N_13369);
xor U13533 (N_13533,N_13397,N_13356);
and U13534 (N_13534,N_13265,N_13382);
or U13535 (N_13535,N_13301,N_13308);
nand U13536 (N_13536,N_13374,N_13320);
or U13537 (N_13537,N_13269,N_13330);
xor U13538 (N_13538,N_13254,N_13226);
and U13539 (N_13539,N_13391,N_13228);
or U13540 (N_13540,N_13251,N_13361);
and U13541 (N_13541,N_13233,N_13267);
nand U13542 (N_13542,N_13311,N_13309);
and U13543 (N_13543,N_13362,N_13381);
and U13544 (N_13544,N_13317,N_13225);
or U13545 (N_13545,N_13246,N_13309);
xor U13546 (N_13546,N_13311,N_13306);
and U13547 (N_13547,N_13261,N_13227);
or U13548 (N_13548,N_13372,N_13352);
nor U13549 (N_13549,N_13357,N_13223);
xor U13550 (N_13550,N_13277,N_13235);
or U13551 (N_13551,N_13205,N_13348);
nand U13552 (N_13552,N_13208,N_13279);
or U13553 (N_13553,N_13248,N_13319);
nand U13554 (N_13554,N_13389,N_13371);
or U13555 (N_13555,N_13238,N_13347);
xnor U13556 (N_13556,N_13310,N_13363);
nand U13557 (N_13557,N_13240,N_13231);
or U13558 (N_13558,N_13354,N_13338);
or U13559 (N_13559,N_13316,N_13361);
nand U13560 (N_13560,N_13374,N_13274);
or U13561 (N_13561,N_13367,N_13360);
nor U13562 (N_13562,N_13205,N_13376);
nor U13563 (N_13563,N_13308,N_13320);
nand U13564 (N_13564,N_13301,N_13334);
and U13565 (N_13565,N_13230,N_13318);
xor U13566 (N_13566,N_13252,N_13302);
or U13567 (N_13567,N_13304,N_13279);
nor U13568 (N_13568,N_13246,N_13240);
or U13569 (N_13569,N_13381,N_13392);
and U13570 (N_13570,N_13270,N_13216);
nor U13571 (N_13571,N_13276,N_13358);
and U13572 (N_13572,N_13285,N_13361);
nand U13573 (N_13573,N_13335,N_13212);
and U13574 (N_13574,N_13324,N_13303);
or U13575 (N_13575,N_13236,N_13330);
or U13576 (N_13576,N_13390,N_13273);
xnor U13577 (N_13577,N_13260,N_13201);
xor U13578 (N_13578,N_13285,N_13258);
and U13579 (N_13579,N_13339,N_13274);
nor U13580 (N_13580,N_13255,N_13371);
xor U13581 (N_13581,N_13236,N_13343);
xnor U13582 (N_13582,N_13255,N_13262);
nor U13583 (N_13583,N_13276,N_13293);
xor U13584 (N_13584,N_13291,N_13325);
or U13585 (N_13585,N_13345,N_13354);
and U13586 (N_13586,N_13208,N_13224);
and U13587 (N_13587,N_13297,N_13238);
or U13588 (N_13588,N_13233,N_13213);
and U13589 (N_13589,N_13256,N_13226);
nand U13590 (N_13590,N_13334,N_13225);
nand U13591 (N_13591,N_13310,N_13289);
nor U13592 (N_13592,N_13364,N_13287);
xnor U13593 (N_13593,N_13204,N_13332);
and U13594 (N_13594,N_13303,N_13219);
nand U13595 (N_13595,N_13379,N_13275);
nand U13596 (N_13596,N_13349,N_13353);
or U13597 (N_13597,N_13387,N_13253);
xor U13598 (N_13598,N_13298,N_13296);
and U13599 (N_13599,N_13251,N_13226);
nand U13600 (N_13600,N_13538,N_13449);
and U13601 (N_13601,N_13590,N_13457);
xor U13602 (N_13602,N_13574,N_13584);
nand U13603 (N_13603,N_13581,N_13488);
nor U13604 (N_13604,N_13436,N_13463);
nand U13605 (N_13605,N_13508,N_13462);
xnor U13606 (N_13606,N_13517,N_13418);
or U13607 (N_13607,N_13546,N_13534);
or U13608 (N_13608,N_13568,N_13507);
or U13609 (N_13609,N_13555,N_13459);
and U13610 (N_13610,N_13441,N_13593);
nand U13611 (N_13611,N_13413,N_13419);
and U13612 (N_13612,N_13490,N_13594);
nor U13613 (N_13613,N_13473,N_13471);
nor U13614 (N_13614,N_13422,N_13482);
or U13615 (N_13615,N_13476,N_13589);
xnor U13616 (N_13616,N_13554,N_13526);
and U13617 (N_13617,N_13409,N_13578);
nand U13618 (N_13618,N_13530,N_13454);
nor U13619 (N_13619,N_13455,N_13465);
nand U13620 (N_13620,N_13469,N_13561);
nand U13621 (N_13621,N_13516,N_13424);
nand U13622 (N_13622,N_13575,N_13446);
nand U13623 (N_13623,N_13549,N_13520);
or U13624 (N_13624,N_13464,N_13518);
xor U13625 (N_13625,N_13514,N_13552);
xnor U13626 (N_13626,N_13501,N_13585);
nor U13627 (N_13627,N_13557,N_13591);
nand U13628 (N_13628,N_13492,N_13562);
xnor U13629 (N_13629,N_13503,N_13531);
nand U13630 (N_13630,N_13506,N_13499);
xor U13631 (N_13631,N_13540,N_13485);
or U13632 (N_13632,N_13525,N_13553);
or U13633 (N_13633,N_13401,N_13566);
or U13634 (N_13634,N_13411,N_13564);
and U13635 (N_13635,N_13505,N_13536);
xnor U13636 (N_13636,N_13543,N_13577);
and U13637 (N_13637,N_13431,N_13547);
nand U13638 (N_13638,N_13533,N_13541);
nor U13639 (N_13639,N_13524,N_13545);
nor U13640 (N_13640,N_13405,N_13597);
and U13641 (N_13641,N_13486,N_13513);
and U13642 (N_13642,N_13588,N_13480);
nand U13643 (N_13643,N_13556,N_13558);
or U13644 (N_13644,N_13544,N_13437);
nand U13645 (N_13645,N_13532,N_13448);
or U13646 (N_13646,N_13474,N_13410);
and U13647 (N_13647,N_13519,N_13407);
nor U13648 (N_13648,N_13414,N_13478);
nor U13649 (N_13649,N_13439,N_13559);
and U13650 (N_13650,N_13435,N_13595);
xnor U13651 (N_13651,N_13453,N_13512);
nand U13652 (N_13652,N_13452,N_13497);
and U13653 (N_13653,N_13494,N_13426);
xor U13654 (N_13654,N_13430,N_13515);
and U13655 (N_13655,N_13404,N_13444);
nor U13656 (N_13656,N_13472,N_13475);
nor U13657 (N_13657,N_13495,N_13458);
xor U13658 (N_13658,N_13598,N_13423);
nand U13659 (N_13659,N_13429,N_13402);
nand U13660 (N_13660,N_13567,N_13521);
or U13661 (N_13661,N_13550,N_13579);
and U13662 (N_13662,N_13522,N_13466);
xnor U13663 (N_13663,N_13504,N_13460);
nor U13664 (N_13664,N_13442,N_13481);
or U13665 (N_13665,N_13586,N_13582);
nor U13666 (N_13666,N_13461,N_13427);
nand U13667 (N_13667,N_13527,N_13509);
nand U13668 (N_13668,N_13491,N_13415);
xor U13669 (N_13669,N_13445,N_13416);
nor U13670 (N_13670,N_13451,N_13560);
and U13671 (N_13671,N_13583,N_13563);
and U13672 (N_13672,N_13523,N_13487);
or U13673 (N_13673,N_13498,N_13537);
nand U13674 (N_13674,N_13434,N_13599);
and U13675 (N_13675,N_13417,N_13510);
xnor U13676 (N_13676,N_13496,N_13428);
nor U13677 (N_13677,N_13470,N_13587);
or U13678 (N_13678,N_13400,N_13502);
and U13679 (N_13679,N_13479,N_13484);
and U13680 (N_13680,N_13596,N_13450);
nor U13681 (N_13681,N_13592,N_13565);
nand U13682 (N_13682,N_13572,N_13468);
xnor U13683 (N_13683,N_13535,N_13412);
and U13684 (N_13684,N_13528,N_13438);
nand U13685 (N_13685,N_13548,N_13489);
nand U13686 (N_13686,N_13573,N_13539);
or U13687 (N_13687,N_13551,N_13456);
and U13688 (N_13688,N_13440,N_13443);
and U13689 (N_13689,N_13447,N_13421);
xor U13690 (N_13690,N_13420,N_13483);
nand U13691 (N_13691,N_13576,N_13580);
nand U13692 (N_13692,N_13408,N_13511);
or U13693 (N_13693,N_13571,N_13467);
nor U13694 (N_13694,N_13570,N_13542);
xor U13695 (N_13695,N_13432,N_13500);
or U13696 (N_13696,N_13433,N_13493);
nor U13697 (N_13697,N_13569,N_13403);
and U13698 (N_13698,N_13477,N_13406);
and U13699 (N_13699,N_13529,N_13425);
and U13700 (N_13700,N_13586,N_13451);
and U13701 (N_13701,N_13502,N_13531);
nand U13702 (N_13702,N_13548,N_13451);
nand U13703 (N_13703,N_13492,N_13552);
xnor U13704 (N_13704,N_13426,N_13460);
xor U13705 (N_13705,N_13598,N_13441);
and U13706 (N_13706,N_13471,N_13535);
or U13707 (N_13707,N_13434,N_13470);
xor U13708 (N_13708,N_13486,N_13469);
or U13709 (N_13709,N_13578,N_13584);
and U13710 (N_13710,N_13435,N_13523);
and U13711 (N_13711,N_13414,N_13463);
and U13712 (N_13712,N_13489,N_13577);
or U13713 (N_13713,N_13515,N_13423);
or U13714 (N_13714,N_13538,N_13407);
nand U13715 (N_13715,N_13527,N_13459);
xnor U13716 (N_13716,N_13490,N_13441);
and U13717 (N_13717,N_13404,N_13555);
or U13718 (N_13718,N_13469,N_13507);
and U13719 (N_13719,N_13576,N_13455);
nor U13720 (N_13720,N_13542,N_13470);
xnor U13721 (N_13721,N_13416,N_13490);
and U13722 (N_13722,N_13416,N_13431);
nand U13723 (N_13723,N_13408,N_13547);
or U13724 (N_13724,N_13461,N_13450);
nor U13725 (N_13725,N_13432,N_13553);
or U13726 (N_13726,N_13468,N_13517);
xor U13727 (N_13727,N_13474,N_13512);
nor U13728 (N_13728,N_13597,N_13544);
or U13729 (N_13729,N_13512,N_13473);
nand U13730 (N_13730,N_13435,N_13445);
or U13731 (N_13731,N_13432,N_13523);
nor U13732 (N_13732,N_13457,N_13556);
nand U13733 (N_13733,N_13479,N_13453);
nand U13734 (N_13734,N_13538,N_13486);
and U13735 (N_13735,N_13498,N_13430);
nor U13736 (N_13736,N_13509,N_13496);
or U13737 (N_13737,N_13464,N_13550);
nor U13738 (N_13738,N_13593,N_13575);
or U13739 (N_13739,N_13469,N_13519);
xnor U13740 (N_13740,N_13450,N_13503);
nand U13741 (N_13741,N_13598,N_13573);
xor U13742 (N_13742,N_13432,N_13429);
nand U13743 (N_13743,N_13487,N_13400);
nor U13744 (N_13744,N_13582,N_13437);
or U13745 (N_13745,N_13404,N_13416);
xnor U13746 (N_13746,N_13400,N_13596);
nor U13747 (N_13747,N_13587,N_13597);
nand U13748 (N_13748,N_13571,N_13535);
or U13749 (N_13749,N_13410,N_13409);
and U13750 (N_13750,N_13556,N_13585);
nor U13751 (N_13751,N_13560,N_13453);
and U13752 (N_13752,N_13464,N_13421);
or U13753 (N_13753,N_13581,N_13574);
nand U13754 (N_13754,N_13525,N_13411);
nor U13755 (N_13755,N_13514,N_13404);
and U13756 (N_13756,N_13467,N_13560);
xnor U13757 (N_13757,N_13509,N_13570);
xnor U13758 (N_13758,N_13483,N_13425);
and U13759 (N_13759,N_13580,N_13495);
xor U13760 (N_13760,N_13488,N_13546);
nor U13761 (N_13761,N_13516,N_13532);
and U13762 (N_13762,N_13530,N_13465);
nand U13763 (N_13763,N_13475,N_13468);
and U13764 (N_13764,N_13439,N_13523);
and U13765 (N_13765,N_13490,N_13422);
nand U13766 (N_13766,N_13415,N_13410);
or U13767 (N_13767,N_13426,N_13567);
nand U13768 (N_13768,N_13430,N_13465);
and U13769 (N_13769,N_13558,N_13455);
nor U13770 (N_13770,N_13466,N_13439);
xnor U13771 (N_13771,N_13426,N_13422);
xor U13772 (N_13772,N_13475,N_13490);
nand U13773 (N_13773,N_13422,N_13512);
xnor U13774 (N_13774,N_13452,N_13544);
or U13775 (N_13775,N_13484,N_13420);
nor U13776 (N_13776,N_13490,N_13590);
xnor U13777 (N_13777,N_13419,N_13460);
nor U13778 (N_13778,N_13555,N_13597);
nand U13779 (N_13779,N_13480,N_13478);
or U13780 (N_13780,N_13404,N_13423);
nand U13781 (N_13781,N_13501,N_13444);
nor U13782 (N_13782,N_13440,N_13493);
or U13783 (N_13783,N_13513,N_13590);
nand U13784 (N_13784,N_13440,N_13456);
and U13785 (N_13785,N_13574,N_13488);
xor U13786 (N_13786,N_13589,N_13454);
nor U13787 (N_13787,N_13574,N_13449);
nor U13788 (N_13788,N_13408,N_13501);
or U13789 (N_13789,N_13411,N_13417);
or U13790 (N_13790,N_13513,N_13530);
nand U13791 (N_13791,N_13488,N_13540);
or U13792 (N_13792,N_13468,N_13547);
or U13793 (N_13793,N_13505,N_13525);
or U13794 (N_13794,N_13513,N_13403);
nand U13795 (N_13795,N_13498,N_13485);
and U13796 (N_13796,N_13478,N_13538);
nor U13797 (N_13797,N_13434,N_13401);
nand U13798 (N_13798,N_13593,N_13427);
and U13799 (N_13799,N_13537,N_13412);
xnor U13800 (N_13800,N_13663,N_13753);
nor U13801 (N_13801,N_13673,N_13649);
or U13802 (N_13802,N_13662,N_13766);
nand U13803 (N_13803,N_13729,N_13774);
xnor U13804 (N_13804,N_13623,N_13655);
and U13805 (N_13805,N_13606,N_13696);
nand U13806 (N_13806,N_13600,N_13769);
xor U13807 (N_13807,N_13653,N_13776);
nor U13808 (N_13808,N_13785,N_13795);
and U13809 (N_13809,N_13778,N_13726);
nor U13810 (N_13810,N_13618,N_13691);
or U13811 (N_13811,N_13683,N_13697);
and U13812 (N_13812,N_13602,N_13702);
nor U13813 (N_13813,N_13728,N_13615);
xor U13814 (N_13814,N_13799,N_13777);
xnor U13815 (N_13815,N_13742,N_13637);
nor U13816 (N_13816,N_13646,N_13724);
xor U13817 (N_13817,N_13695,N_13684);
nand U13818 (N_13818,N_13734,N_13666);
or U13819 (N_13819,N_13659,N_13676);
nand U13820 (N_13820,N_13711,N_13601);
xnor U13821 (N_13821,N_13796,N_13743);
nand U13822 (N_13822,N_13792,N_13678);
xnor U13823 (N_13823,N_13650,N_13668);
xor U13824 (N_13824,N_13715,N_13690);
and U13825 (N_13825,N_13750,N_13657);
xor U13826 (N_13826,N_13767,N_13698);
and U13827 (N_13827,N_13630,N_13773);
and U13828 (N_13828,N_13631,N_13675);
and U13829 (N_13829,N_13656,N_13620);
xnor U13830 (N_13830,N_13635,N_13755);
xnor U13831 (N_13831,N_13607,N_13626);
and U13832 (N_13832,N_13660,N_13692);
nor U13833 (N_13833,N_13701,N_13770);
xnor U13834 (N_13834,N_13710,N_13752);
and U13835 (N_13835,N_13794,N_13669);
xnor U13836 (N_13836,N_13786,N_13736);
and U13837 (N_13837,N_13705,N_13681);
nand U13838 (N_13838,N_13647,N_13643);
or U13839 (N_13839,N_13644,N_13761);
nor U13840 (N_13840,N_13689,N_13642);
and U13841 (N_13841,N_13745,N_13704);
or U13842 (N_13842,N_13735,N_13780);
or U13843 (N_13843,N_13763,N_13731);
xor U13844 (N_13844,N_13700,N_13699);
nor U13845 (N_13845,N_13665,N_13624);
nand U13846 (N_13846,N_13693,N_13740);
or U13847 (N_13847,N_13737,N_13640);
nor U13848 (N_13848,N_13775,N_13756);
or U13849 (N_13849,N_13732,N_13782);
xnor U13850 (N_13850,N_13664,N_13613);
and U13851 (N_13851,N_13757,N_13747);
or U13852 (N_13852,N_13648,N_13746);
and U13853 (N_13853,N_13614,N_13708);
nor U13854 (N_13854,N_13793,N_13687);
and U13855 (N_13855,N_13605,N_13719);
and U13856 (N_13856,N_13628,N_13765);
nor U13857 (N_13857,N_13720,N_13741);
xor U13858 (N_13858,N_13670,N_13603);
nand U13859 (N_13859,N_13682,N_13604);
or U13860 (N_13860,N_13622,N_13667);
nor U13861 (N_13861,N_13674,N_13771);
xor U13862 (N_13862,N_13654,N_13709);
nand U13863 (N_13863,N_13760,N_13749);
nor U13864 (N_13864,N_13787,N_13617);
or U13865 (N_13865,N_13712,N_13688);
xor U13866 (N_13866,N_13762,N_13636);
xnor U13867 (N_13867,N_13706,N_13797);
and U13868 (N_13868,N_13707,N_13629);
or U13869 (N_13869,N_13722,N_13661);
and U13870 (N_13870,N_13764,N_13612);
nand U13871 (N_13871,N_13625,N_13685);
or U13872 (N_13872,N_13759,N_13611);
nor U13873 (N_13873,N_13725,N_13677);
or U13874 (N_13874,N_13784,N_13694);
nor U13875 (N_13875,N_13672,N_13716);
nor U13876 (N_13876,N_13616,N_13790);
or U13877 (N_13877,N_13718,N_13723);
nor U13878 (N_13878,N_13730,N_13791);
nand U13879 (N_13879,N_13744,N_13751);
nand U13880 (N_13880,N_13714,N_13641);
nor U13881 (N_13881,N_13754,N_13634);
and U13882 (N_13882,N_13658,N_13610);
nand U13883 (N_13883,N_13633,N_13638);
nand U13884 (N_13884,N_13768,N_13627);
or U13885 (N_13885,N_13680,N_13645);
and U13886 (N_13886,N_13772,N_13621);
nor U13887 (N_13887,N_13758,N_13783);
nor U13888 (N_13888,N_13686,N_13703);
nor U13889 (N_13889,N_13713,N_13632);
or U13890 (N_13890,N_13789,N_13779);
nand U13891 (N_13891,N_13738,N_13651);
and U13892 (N_13892,N_13619,N_13798);
or U13893 (N_13893,N_13609,N_13748);
or U13894 (N_13894,N_13721,N_13733);
and U13895 (N_13895,N_13717,N_13727);
xor U13896 (N_13896,N_13679,N_13671);
and U13897 (N_13897,N_13788,N_13739);
and U13898 (N_13898,N_13639,N_13781);
and U13899 (N_13899,N_13652,N_13608);
xnor U13900 (N_13900,N_13624,N_13796);
nand U13901 (N_13901,N_13620,N_13660);
or U13902 (N_13902,N_13607,N_13658);
or U13903 (N_13903,N_13654,N_13655);
and U13904 (N_13904,N_13662,N_13777);
and U13905 (N_13905,N_13637,N_13796);
and U13906 (N_13906,N_13672,N_13641);
nand U13907 (N_13907,N_13645,N_13726);
or U13908 (N_13908,N_13658,N_13757);
or U13909 (N_13909,N_13630,N_13663);
and U13910 (N_13910,N_13679,N_13672);
nand U13911 (N_13911,N_13678,N_13614);
nand U13912 (N_13912,N_13712,N_13761);
nor U13913 (N_13913,N_13669,N_13613);
or U13914 (N_13914,N_13792,N_13740);
or U13915 (N_13915,N_13647,N_13751);
nand U13916 (N_13916,N_13649,N_13793);
or U13917 (N_13917,N_13754,N_13785);
nor U13918 (N_13918,N_13710,N_13723);
nand U13919 (N_13919,N_13714,N_13644);
xnor U13920 (N_13920,N_13720,N_13632);
and U13921 (N_13921,N_13755,N_13767);
or U13922 (N_13922,N_13656,N_13716);
nor U13923 (N_13923,N_13759,N_13713);
or U13924 (N_13924,N_13600,N_13720);
nand U13925 (N_13925,N_13710,N_13768);
nor U13926 (N_13926,N_13638,N_13733);
and U13927 (N_13927,N_13793,N_13704);
nand U13928 (N_13928,N_13693,N_13795);
xor U13929 (N_13929,N_13661,N_13689);
or U13930 (N_13930,N_13626,N_13632);
xnor U13931 (N_13931,N_13763,N_13603);
nand U13932 (N_13932,N_13793,N_13770);
and U13933 (N_13933,N_13738,N_13702);
xnor U13934 (N_13934,N_13752,N_13788);
xor U13935 (N_13935,N_13707,N_13764);
nand U13936 (N_13936,N_13623,N_13600);
or U13937 (N_13937,N_13604,N_13757);
or U13938 (N_13938,N_13615,N_13602);
nand U13939 (N_13939,N_13643,N_13722);
nor U13940 (N_13940,N_13757,N_13607);
and U13941 (N_13941,N_13693,N_13664);
nand U13942 (N_13942,N_13707,N_13711);
nor U13943 (N_13943,N_13723,N_13715);
and U13944 (N_13944,N_13702,N_13628);
xnor U13945 (N_13945,N_13643,N_13637);
or U13946 (N_13946,N_13612,N_13609);
and U13947 (N_13947,N_13756,N_13793);
xor U13948 (N_13948,N_13741,N_13752);
and U13949 (N_13949,N_13614,N_13689);
or U13950 (N_13950,N_13694,N_13699);
nor U13951 (N_13951,N_13745,N_13782);
and U13952 (N_13952,N_13799,N_13604);
or U13953 (N_13953,N_13601,N_13691);
nand U13954 (N_13954,N_13639,N_13741);
and U13955 (N_13955,N_13634,N_13796);
nor U13956 (N_13956,N_13618,N_13648);
xnor U13957 (N_13957,N_13722,N_13676);
nand U13958 (N_13958,N_13739,N_13643);
xor U13959 (N_13959,N_13723,N_13629);
or U13960 (N_13960,N_13653,N_13665);
and U13961 (N_13961,N_13625,N_13639);
and U13962 (N_13962,N_13645,N_13658);
nand U13963 (N_13963,N_13755,N_13628);
and U13964 (N_13964,N_13710,N_13640);
nor U13965 (N_13965,N_13649,N_13727);
and U13966 (N_13966,N_13618,N_13722);
xnor U13967 (N_13967,N_13721,N_13775);
xnor U13968 (N_13968,N_13792,N_13653);
nor U13969 (N_13969,N_13730,N_13634);
or U13970 (N_13970,N_13650,N_13687);
or U13971 (N_13971,N_13616,N_13744);
xor U13972 (N_13972,N_13646,N_13702);
or U13973 (N_13973,N_13798,N_13733);
or U13974 (N_13974,N_13725,N_13775);
and U13975 (N_13975,N_13733,N_13682);
xor U13976 (N_13976,N_13641,N_13720);
or U13977 (N_13977,N_13659,N_13642);
nor U13978 (N_13978,N_13678,N_13639);
xor U13979 (N_13979,N_13702,N_13749);
and U13980 (N_13980,N_13633,N_13639);
nor U13981 (N_13981,N_13719,N_13687);
or U13982 (N_13982,N_13655,N_13782);
nor U13983 (N_13983,N_13746,N_13792);
or U13984 (N_13984,N_13633,N_13772);
or U13985 (N_13985,N_13604,N_13623);
nand U13986 (N_13986,N_13782,N_13758);
nor U13987 (N_13987,N_13698,N_13628);
and U13988 (N_13988,N_13793,N_13733);
or U13989 (N_13989,N_13713,N_13662);
and U13990 (N_13990,N_13788,N_13782);
nor U13991 (N_13991,N_13621,N_13744);
nor U13992 (N_13992,N_13773,N_13674);
nor U13993 (N_13993,N_13734,N_13760);
xor U13994 (N_13994,N_13656,N_13706);
and U13995 (N_13995,N_13780,N_13649);
xor U13996 (N_13996,N_13625,N_13720);
nand U13997 (N_13997,N_13651,N_13709);
or U13998 (N_13998,N_13637,N_13712);
xor U13999 (N_13999,N_13634,N_13629);
xnor U14000 (N_14000,N_13880,N_13881);
and U14001 (N_14001,N_13828,N_13835);
xnor U14002 (N_14002,N_13874,N_13890);
xor U14003 (N_14003,N_13832,N_13856);
nor U14004 (N_14004,N_13816,N_13846);
xnor U14005 (N_14005,N_13903,N_13987);
or U14006 (N_14006,N_13933,N_13834);
or U14007 (N_14007,N_13859,N_13916);
or U14008 (N_14008,N_13914,N_13943);
xnor U14009 (N_14009,N_13857,N_13872);
or U14010 (N_14010,N_13968,N_13967);
nor U14011 (N_14011,N_13848,N_13887);
nor U14012 (N_14012,N_13882,N_13825);
nor U14013 (N_14013,N_13970,N_13869);
or U14014 (N_14014,N_13941,N_13830);
nor U14015 (N_14015,N_13958,N_13875);
xnor U14016 (N_14016,N_13862,N_13949);
xnor U14017 (N_14017,N_13801,N_13895);
and U14018 (N_14018,N_13854,N_13994);
nor U14019 (N_14019,N_13960,N_13999);
nand U14020 (N_14020,N_13946,N_13981);
and U14021 (N_14021,N_13847,N_13989);
and U14022 (N_14022,N_13991,N_13833);
or U14023 (N_14023,N_13986,N_13898);
or U14024 (N_14024,N_13858,N_13962);
and U14025 (N_14025,N_13923,N_13956);
nor U14026 (N_14026,N_13910,N_13924);
xnor U14027 (N_14027,N_13971,N_13906);
nor U14028 (N_14028,N_13879,N_13824);
and U14029 (N_14029,N_13827,N_13985);
or U14030 (N_14030,N_13809,N_13814);
and U14031 (N_14031,N_13915,N_13920);
xnor U14032 (N_14032,N_13839,N_13948);
or U14033 (N_14033,N_13978,N_13974);
or U14034 (N_14034,N_13852,N_13955);
xnor U14035 (N_14035,N_13865,N_13940);
xor U14036 (N_14036,N_13963,N_13947);
or U14037 (N_14037,N_13908,N_13892);
nand U14038 (N_14038,N_13953,N_13904);
and U14039 (N_14039,N_13817,N_13842);
or U14040 (N_14040,N_13819,N_13930);
xor U14041 (N_14041,N_13806,N_13829);
or U14042 (N_14042,N_13931,N_13871);
xor U14043 (N_14043,N_13850,N_13851);
nor U14044 (N_14044,N_13938,N_13804);
xnor U14045 (N_14045,N_13873,N_13934);
xor U14046 (N_14046,N_13861,N_13969);
and U14047 (N_14047,N_13918,N_13844);
nor U14048 (N_14048,N_13868,N_13870);
xor U14049 (N_14049,N_13821,N_13926);
or U14050 (N_14050,N_13928,N_13937);
nor U14051 (N_14051,N_13840,N_13936);
nor U14052 (N_14052,N_13973,N_13807);
nor U14053 (N_14053,N_13939,N_13883);
nor U14054 (N_14054,N_13925,N_13905);
and U14055 (N_14055,N_13866,N_13979);
nand U14056 (N_14056,N_13815,N_13876);
and U14057 (N_14057,N_13893,N_13803);
nand U14058 (N_14058,N_13823,N_13896);
nor U14059 (N_14059,N_13972,N_13957);
nor U14060 (N_14060,N_13959,N_13945);
and U14061 (N_14061,N_13867,N_13901);
nand U14062 (N_14062,N_13927,N_13849);
or U14063 (N_14063,N_13990,N_13808);
nand U14064 (N_14064,N_13884,N_13889);
or U14065 (N_14065,N_13950,N_13863);
and U14066 (N_14066,N_13894,N_13952);
and U14067 (N_14067,N_13961,N_13912);
or U14068 (N_14068,N_13984,N_13826);
nand U14069 (N_14069,N_13966,N_13855);
nand U14070 (N_14070,N_13951,N_13909);
xor U14071 (N_14071,N_13964,N_13836);
or U14072 (N_14072,N_13900,N_13998);
and U14073 (N_14073,N_13802,N_13954);
or U14074 (N_14074,N_13864,N_13878);
nand U14075 (N_14075,N_13992,N_13983);
and U14076 (N_14076,N_13935,N_13977);
or U14077 (N_14077,N_13902,N_13965);
and U14078 (N_14078,N_13919,N_13885);
xor U14079 (N_14079,N_13997,N_13843);
or U14080 (N_14080,N_13891,N_13888);
xor U14081 (N_14081,N_13993,N_13917);
nand U14082 (N_14082,N_13995,N_13899);
and U14083 (N_14083,N_13838,N_13805);
nand U14084 (N_14084,N_13897,N_13822);
or U14085 (N_14085,N_13877,N_13811);
or U14086 (N_14086,N_13886,N_13800);
nor U14087 (N_14087,N_13932,N_13944);
nand U14088 (N_14088,N_13812,N_13975);
nor U14089 (N_14089,N_13976,N_13988);
and U14090 (N_14090,N_13860,N_13845);
or U14091 (N_14091,N_13818,N_13837);
nand U14092 (N_14092,N_13982,N_13911);
or U14093 (N_14093,N_13907,N_13922);
xor U14094 (N_14094,N_13980,N_13853);
and U14095 (N_14095,N_13921,N_13841);
or U14096 (N_14096,N_13813,N_13929);
nand U14097 (N_14097,N_13820,N_13831);
nand U14098 (N_14098,N_13810,N_13996);
nor U14099 (N_14099,N_13913,N_13942);
nor U14100 (N_14100,N_13885,N_13887);
nand U14101 (N_14101,N_13938,N_13976);
or U14102 (N_14102,N_13963,N_13849);
nand U14103 (N_14103,N_13942,N_13818);
nor U14104 (N_14104,N_13962,N_13889);
xor U14105 (N_14105,N_13978,N_13925);
or U14106 (N_14106,N_13853,N_13876);
nor U14107 (N_14107,N_13933,N_13824);
and U14108 (N_14108,N_13839,N_13823);
or U14109 (N_14109,N_13808,N_13830);
and U14110 (N_14110,N_13875,N_13880);
nor U14111 (N_14111,N_13824,N_13863);
or U14112 (N_14112,N_13894,N_13842);
nor U14113 (N_14113,N_13866,N_13805);
nor U14114 (N_14114,N_13942,N_13884);
nor U14115 (N_14115,N_13911,N_13872);
nand U14116 (N_14116,N_13963,N_13995);
and U14117 (N_14117,N_13811,N_13905);
or U14118 (N_14118,N_13838,N_13947);
and U14119 (N_14119,N_13904,N_13869);
and U14120 (N_14120,N_13862,N_13866);
nor U14121 (N_14121,N_13946,N_13898);
or U14122 (N_14122,N_13894,N_13830);
and U14123 (N_14123,N_13986,N_13856);
nand U14124 (N_14124,N_13948,N_13951);
and U14125 (N_14125,N_13802,N_13947);
nand U14126 (N_14126,N_13925,N_13988);
xor U14127 (N_14127,N_13948,N_13909);
and U14128 (N_14128,N_13916,N_13963);
nand U14129 (N_14129,N_13874,N_13823);
xnor U14130 (N_14130,N_13979,N_13961);
nand U14131 (N_14131,N_13909,N_13875);
xnor U14132 (N_14132,N_13867,N_13951);
or U14133 (N_14133,N_13960,N_13886);
and U14134 (N_14134,N_13906,N_13809);
or U14135 (N_14135,N_13802,N_13882);
xor U14136 (N_14136,N_13802,N_13970);
xor U14137 (N_14137,N_13858,N_13802);
xor U14138 (N_14138,N_13823,N_13870);
nand U14139 (N_14139,N_13955,N_13999);
xnor U14140 (N_14140,N_13814,N_13804);
or U14141 (N_14141,N_13843,N_13856);
and U14142 (N_14142,N_13897,N_13930);
nand U14143 (N_14143,N_13843,N_13891);
nand U14144 (N_14144,N_13947,N_13845);
xnor U14145 (N_14145,N_13814,N_13853);
nand U14146 (N_14146,N_13922,N_13868);
xor U14147 (N_14147,N_13835,N_13832);
xnor U14148 (N_14148,N_13950,N_13844);
nand U14149 (N_14149,N_13834,N_13902);
nand U14150 (N_14150,N_13924,N_13850);
or U14151 (N_14151,N_13870,N_13853);
or U14152 (N_14152,N_13992,N_13920);
or U14153 (N_14153,N_13913,N_13948);
xor U14154 (N_14154,N_13993,N_13869);
nor U14155 (N_14155,N_13879,N_13905);
nand U14156 (N_14156,N_13855,N_13938);
and U14157 (N_14157,N_13930,N_13878);
nand U14158 (N_14158,N_13806,N_13970);
xnor U14159 (N_14159,N_13904,N_13863);
xor U14160 (N_14160,N_13935,N_13859);
nand U14161 (N_14161,N_13817,N_13925);
or U14162 (N_14162,N_13927,N_13817);
nor U14163 (N_14163,N_13934,N_13882);
and U14164 (N_14164,N_13805,N_13928);
or U14165 (N_14165,N_13909,N_13936);
nand U14166 (N_14166,N_13942,N_13844);
and U14167 (N_14167,N_13819,N_13973);
and U14168 (N_14168,N_13895,N_13832);
and U14169 (N_14169,N_13968,N_13896);
xnor U14170 (N_14170,N_13964,N_13886);
xor U14171 (N_14171,N_13966,N_13870);
nand U14172 (N_14172,N_13808,N_13982);
xor U14173 (N_14173,N_13981,N_13892);
xnor U14174 (N_14174,N_13870,N_13956);
or U14175 (N_14175,N_13859,N_13842);
or U14176 (N_14176,N_13932,N_13907);
nand U14177 (N_14177,N_13920,N_13911);
nand U14178 (N_14178,N_13819,N_13877);
and U14179 (N_14179,N_13843,N_13854);
or U14180 (N_14180,N_13967,N_13878);
nand U14181 (N_14181,N_13991,N_13923);
nor U14182 (N_14182,N_13924,N_13944);
nand U14183 (N_14183,N_13977,N_13998);
nand U14184 (N_14184,N_13851,N_13894);
nand U14185 (N_14185,N_13895,N_13955);
and U14186 (N_14186,N_13849,N_13907);
or U14187 (N_14187,N_13948,N_13815);
xnor U14188 (N_14188,N_13877,N_13867);
nor U14189 (N_14189,N_13997,N_13890);
xnor U14190 (N_14190,N_13943,N_13845);
nand U14191 (N_14191,N_13867,N_13853);
nand U14192 (N_14192,N_13809,N_13845);
nand U14193 (N_14193,N_13957,N_13868);
nor U14194 (N_14194,N_13913,N_13884);
and U14195 (N_14195,N_13920,N_13951);
xnor U14196 (N_14196,N_13876,N_13984);
and U14197 (N_14197,N_13846,N_13909);
xor U14198 (N_14198,N_13871,N_13832);
and U14199 (N_14199,N_13866,N_13909);
nand U14200 (N_14200,N_14128,N_14079);
nand U14201 (N_14201,N_14037,N_14002);
nand U14202 (N_14202,N_14036,N_14162);
xnor U14203 (N_14203,N_14053,N_14130);
or U14204 (N_14204,N_14015,N_14075);
nand U14205 (N_14205,N_14157,N_14050);
xnor U14206 (N_14206,N_14095,N_14011);
xnor U14207 (N_14207,N_14047,N_14061);
or U14208 (N_14208,N_14178,N_14042);
or U14209 (N_14209,N_14144,N_14136);
and U14210 (N_14210,N_14193,N_14152);
and U14211 (N_14211,N_14105,N_14124);
and U14212 (N_14212,N_14112,N_14173);
nor U14213 (N_14213,N_14141,N_14140);
xnor U14214 (N_14214,N_14022,N_14129);
or U14215 (N_14215,N_14096,N_14115);
nand U14216 (N_14216,N_14147,N_14143);
nor U14217 (N_14217,N_14060,N_14118);
and U14218 (N_14218,N_14001,N_14131);
nor U14219 (N_14219,N_14108,N_14039);
xnor U14220 (N_14220,N_14170,N_14066);
or U14221 (N_14221,N_14091,N_14122);
or U14222 (N_14222,N_14156,N_14146);
nor U14223 (N_14223,N_14084,N_14076);
nor U14224 (N_14224,N_14199,N_14114);
nand U14225 (N_14225,N_14113,N_14071);
xor U14226 (N_14226,N_14111,N_14164);
xnor U14227 (N_14227,N_14100,N_14010);
nor U14228 (N_14228,N_14139,N_14054);
nand U14229 (N_14229,N_14198,N_14080);
or U14230 (N_14230,N_14093,N_14025);
nor U14231 (N_14231,N_14196,N_14009);
and U14232 (N_14232,N_14000,N_14026);
and U14233 (N_14233,N_14135,N_14070);
xor U14234 (N_14234,N_14155,N_14192);
nand U14235 (N_14235,N_14167,N_14191);
nand U14236 (N_14236,N_14109,N_14003);
and U14237 (N_14237,N_14005,N_14094);
nand U14238 (N_14238,N_14125,N_14021);
xnor U14239 (N_14239,N_14177,N_14004);
nand U14240 (N_14240,N_14059,N_14158);
or U14241 (N_14241,N_14159,N_14045);
xnor U14242 (N_14242,N_14057,N_14064);
or U14243 (N_14243,N_14102,N_14018);
or U14244 (N_14244,N_14086,N_14148);
nor U14245 (N_14245,N_14194,N_14137);
nor U14246 (N_14246,N_14127,N_14073);
and U14247 (N_14247,N_14171,N_14081);
nor U14248 (N_14248,N_14013,N_14028);
and U14249 (N_14249,N_14068,N_14151);
nand U14250 (N_14250,N_14121,N_14163);
or U14251 (N_14251,N_14165,N_14085);
nor U14252 (N_14252,N_14008,N_14179);
xor U14253 (N_14253,N_14134,N_14174);
or U14254 (N_14254,N_14172,N_14123);
and U14255 (N_14255,N_14063,N_14078);
and U14256 (N_14256,N_14184,N_14023);
nor U14257 (N_14257,N_14024,N_14110);
or U14258 (N_14258,N_14154,N_14034);
and U14259 (N_14259,N_14012,N_14190);
and U14260 (N_14260,N_14195,N_14029);
xor U14261 (N_14261,N_14197,N_14187);
and U14262 (N_14262,N_14088,N_14117);
nor U14263 (N_14263,N_14067,N_14132);
and U14264 (N_14264,N_14186,N_14089);
xnor U14265 (N_14265,N_14126,N_14103);
xor U14266 (N_14266,N_14072,N_14056);
or U14267 (N_14267,N_14107,N_14176);
nand U14268 (N_14268,N_14188,N_14083);
nand U14269 (N_14269,N_14142,N_14104);
nand U14270 (N_14270,N_14160,N_14145);
or U14271 (N_14271,N_14106,N_14182);
nand U14272 (N_14272,N_14069,N_14120);
and U14273 (N_14273,N_14153,N_14058);
or U14274 (N_14274,N_14062,N_14065);
nor U14275 (N_14275,N_14051,N_14138);
xnor U14276 (N_14276,N_14181,N_14074);
or U14277 (N_14277,N_14116,N_14046);
or U14278 (N_14278,N_14092,N_14043);
nor U14279 (N_14279,N_14101,N_14168);
or U14280 (N_14280,N_14180,N_14035);
nand U14281 (N_14281,N_14133,N_14119);
or U14282 (N_14282,N_14055,N_14040);
xnor U14283 (N_14283,N_14020,N_14017);
nand U14284 (N_14284,N_14166,N_14049);
nor U14285 (N_14285,N_14082,N_14077);
xor U14286 (N_14286,N_14161,N_14183);
xnor U14287 (N_14287,N_14014,N_14048);
nand U14288 (N_14288,N_14052,N_14087);
nand U14289 (N_14289,N_14189,N_14019);
nand U14290 (N_14290,N_14007,N_14033);
and U14291 (N_14291,N_14030,N_14027);
nor U14292 (N_14292,N_14090,N_14016);
nor U14293 (N_14293,N_14038,N_14006);
or U14294 (N_14294,N_14097,N_14175);
nor U14295 (N_14295,N_14044,N_14169);
nor U14296 (N_14296,N_14041,N_14150);
nor U14297 (N_14297,N_14098,N_14149);
and U14298 (N_14298,N_14032,N_14099);
nand U14299 (N_14299,N_14185,N_14031);
and U14300 (N_14300,N_14113,N_14179);
nor U14301 (N_14301,N_14092,N_14057);
xor U14302 (N_14302,N_14029,N_14046);
xor U14303 (N_14303,N_14122,N_14099);
xor U14304 (N_14304,N_14044,N_14130);
or U14305 (N_14305,N_14063,N_14095);
nor U14306 (N_14306,N_14183,N_14126);
xnor U14307 (N_14307,N_14103,N_14195);
or U14308 (N_14308,N_14067,N_14037);
xor U14309 (N_14309,N_14053,N_14170);
nand U14310 (N_14310,N_14033,N_14036);
or U14311 (N_14311,N_14082,N_14076);
nand U14312 (N_14312,N_14035,N_14139);
or U14313 (N_14313,N_14076,N_14019);
nand U14314 (N_14314,N_14175,N_14164);
or U14315 (N_14315,N_14097,N_14176);
and U14316 (N_14316,N_14147,N_14102);
nor U14317 (N_14317,N_14115,N_14191);
or U14318 (N_14318,N_14100,N_14126);
nand U14319 (N_14319,N_14144,N_14150);
nor U14320 (N_14320,N_14139,N_14176);
or U14321 (N_14321,N_14105,N_14169);
and U14322 (N_14322,N_14079,N_14192);
and U14323 (N_14323,N_14072,N_14024);
nand U14324 (N_14324,N_14081,N_14123);
xor U14325 (N_14325,N_14065,N_14111);
xnor U14326 (N_14326,N_14151,N_14139);
xnor U14327 (N_14327,N_14079,N_14102);
or U14328 (N_14328,N_14164,N_14193);
or U14329 (N_14329,N_14047,N_14170);
or U14330 (N_14330,N_14031,N_14136);
and U14331 (N_14331,N_14152,N_14171);
and U14332 (N_14332,N_14160,N_14143);
or U14333 (N_14333,N_14060,N_14127);
and U14334 (N_14334,N_14177,N_14052);
and U14335 (N_14335,N_14002,N_14128);
xnor U14336 (N_14336,N_14190,N_14010);
xnor U14337 (N_14337,N_14096,N_14169);
nand U14338 (N_14338,N_14152,N_14190);
and U14339 (N_14339,N_14131,N_14097);
nor U14340 (N_14340,N_14039,N_14007);
and U14341 (N_14341,N_14171,N_14182);
nor U14342 (N_14342,N_14162,N_14133);
or U14343 (N_14343,N_14107,N_14046);
and U14344 (N_14344,N_14020,N_14139);
and U14345 (N_14345,N_14034,N_14146);
nor U14346 (N_14346,N_14032,N_14071);
nand U14347 (N_14347,N_14029,N_14138);
or U14348 (N_14348,N_14122,N_14165);
nor U14349 (N_14349,N_14109,N_14034);
nor U14350 (N_14350,N_14066,N_14009);
nor U14351 (N_14351,N_14198,N_14015);
and U14352 (N_14352,N_14118,N_14169);
and U14353 (N_14353,N_14063,N_14003);
nor U14354 (N_14354,N_14064,N_14085);
nor U14355 (N_14355,N_14072,N_14068);
nor U14356 (N_14356,N_14052,N_14089);
and U14357 (N_14357,N_14107,N_14055);
nand U14358 (N_14358,N_14136,N_14021);
xnor U14359 (N_14359,N_14085,N_14176);
or U14360 (N_14360,N_14075,N_14020);
nand U14361 (N_14361,N_14001,N_14015);
xnor U14362 (N_14362,N_14059,N_14011);
nand U14363 (N_14363,N_14125,N_14075);
or U14364 (N_14364,N_14022,N_14098);
xor U14365 (N_14365,N_14170,N_14182);
xnor U14366 (N_14366,N_14090,N_14047);
nand U14367 (N_14367,N_14120,N_14090);
and U14368 (N_14368,N_14104,N_14125);
nand U14369 (N_14369,N_14180,N_14077);
and U14370 (N_14370,N_14187,N_14098);
nor U14371 (N_14371,N_14047,N_14065);
nand U14372 (N_14372,N_14005,N_14162);
nand U14373 (N_14373,N_14085,N_14024);
and U14374 (N_14374,N_14092,N_14051);
and U14375 (N_14375,N_14170,N_14106);
or U14376 (N_14376,N_14143,N_14192);
nand U14377 (N_14377,N_14086,N_14140);
xor U14378 (N_14378,N_14071,N_14105);
xor U14379 (N_14379,N_14064,N_14132);
nor U14380 (N_14380,N_14153,N_14026);
nor U14381 (N_14381,N_14118,N_14136);
and U14382 (N_14382,N_14126,N_14195);
nor U14383 (N_14383,N_14025,N_14084);
or U14384 (N_14384,N_14032,N_14135);
nor U14385 (N_14385,N_14001,N_14130);
nor U14386 (N_14386,N_14108,N_14119);
nand U14387 (N_14387,N_14054,N_14173);
or U14388 (N_14388,N_14115,N_14085);
or U14389 (N_14389,N_14162,N_14179);
xor U14390 (N_14390,N_14157,N_14129);
nand U14391 (N_14391,N_14045,N_14174);
nor U14392 (N_14392,N_14169,N_14190);
xor U14393 (N_14393,N_14136,N_14142);
nor U14394 (N_14394,N_14105,N_14182);
xnor U14395 (N_14395,N_14110,N_14109);
and U14396 (N_14396,N_14186,N_14144);
or U14397 (N_14397,N_14024,N_14045);
xnor U14398 (N_14398,N_14105,N_14111);
or U14399 (N_14399,N_14155,N_14152);
xnor U14400 (N_14400,N_14224,N_14268);
and U14401 (N_14401,N_14361,N_14367);
and U14402 (N_14402,N_14347,N_14399);
or U14403 (N_14403,N_14333,N_14382);
or U14404 (N_14404,N_14337,N_14271);
or U14405 (N_14405,N_14247,N_14214);
and U14406 (N_14406,N_14205,N_14341);
and U14407 (N_14407,N_14216,N_14281);
nand U14408 (N_14408,N_14381,N_14338);
nand U14409 (N_14409,N_14204,N_14376);
and U14410 (N_14410,N_14379,N_14346);
xor U14411 (N_14411,N_14325,N_14237);
and U14412 (N_14412,N_14356,N_14295);
and U14413 (N_14413,N_14355,N_14318);
nor U14414 (N_14414,N_14296,N_14248);
nor U14415 (N_14415,N_14277,N_14293);
nor U14416 (N_14416,N_14349,N_14223);
and U14417 (N_14417,N_14396,N_14369);
nor U14418 (N_14418,N_14342,N_14315);
nand U14419 (N_14419,N_14284,N_14231);
nand U14420 (N_14420,N_14203,N_14253);
or U14421 (N_14421,N_14255,N_14229);
or U14422 (N_14422,N_14213,N_14371);
and U14423 (N_14423,N_14354,N_14220);
nand U14424 (N_14424,N_14285,N_14252);
nand U14425 (N_14425,N_14353,N_14336);
or U14426 (N_14426,N_14286,N_14388);
xnor U14427 (N_14427,N_14328,N_14215);
nor U14428 (N_14428,N_14391,N_14228);
and U14429 (N_14429,N_14352,N_14332);
or U14430 (N_14430,N_14266,N_14256);
and U14431 (N_14431,N_14257,N_14280);
nor U14432 (N_14432,N_14235,N_14313);
and U14433 (N_14433,N_14320,N_14201);
nand U14434 (N_14434,N_14304,N_14390);
nand U14435 (N_14435,N_14386,N_14339);
xor U14436 (N_14436,N_14294,N_14305);
and U14437 (N_14437,N_14289,N_14239);
nor U14438 (N_14438,N_14326,N_14331);
or U14439 (N_14439,N_14245,N_14207);
nor U14440 (N_14440,N_14316,N_14242);
and U14441 (N_14441,N_14350,N_14264);
nand U14442 (N_14442,N_14343,N_14241);
nor U14443 (N_14443,N_14322,N_14274);
or U14444 (N_14444,N_14238,N_14269);
or U14445 (N_14445,N_14323,N_14345);
nor U14446 (N_14446,N_14378,N_14377);
or U14447 (N_14447,N_14232,N_14324);
nor U14448 (N_14448,N_14221,N_14392);
or U14449 (N_14449,N_14344,N_14366);
nor U14450 (N_14450,N_14389,N_14329);
nor U14451 (N_14451,N_14373,N_14208);
and U14452 (N_14452,N_14312,N_14393);
nor U14453 (N_14453,N_14357,N_14210);
xor U14454 (N_14454,N_14383,N_14397);
and U14455 (N_14455,N_14360,N_14348);
xor U14456 (N_14456,N_14301,N_14374);
or U14457 (N_14457,N_14300,N_14298);
or U14458 (N_14458,N_14263,N_14363);
xnor U14459 (N_14459,N_14211,N_14327);
and U14460 (N_14460,N_14227,N_14306);
or U14461 (N_14461,N_14288,N_14311);
nor U14462 (N_14462,N_14275,N_14236);
or U14463 (N_14463,N_14335,N_14314);
xor U14464 (N_14464,N_14351,N_14270);
nor U14465 (N_14465,N_14375,N_14317);
nor U14466 (N_14466,N_14246,N_14278);
or U14467 (N_14467,N_14287,N_14398);
or U14468 (N_14468,N_14279,N_14359);
xnor U14469 (N_14469,N_14261,N_14262);
or U14470 (N_14470,N_14303,N_14385);
nand U14471 (N_14471,N_14291,N_14225);
nand U14472 (N_14472,N_14267,N_14309);
xor U14473 (N_14473,N_14260,N_14243);
and U14474 (N_14474,N_14387,N_14202);
or U14475 (N_14475,N_14330,N_14234);
or U14476 (N_14476,N_14250,N_14299);
xnor U14477 (N_14477,N_14368,N_14364);
xnor U14478 (N_14478,N_14290,N_14365);
xor U14479 (N_14479,N_14219,N_14370);
and U14480 (N_14480,N_14380,N_14230);
xor U14481 (N_14481,N_14321,N_14319);
nand U14482 (N_14482,N_14334,N_14358);
nand U14483 (N_14483,N_14302,N_14240);
nand U14484 (N_14484,N_14244,N_14394);
or U14485 (N_14485,N_14217,N_14307);
nor U14486 (N_14486,N_14226,N_14283);
xor U14487 (N_14487,N_14206,N_14272);
nand U14488 (N_14488,N_14372,N_14254);
nand U14489 (N_14489,N_14340,N_14259);
nor U14490 (N_14490,N_14209,N_14292);
nor U14491 (N_14491,N_14276,N_14222);
and U14492 (N_14492,N_14265,N_14200);
nand U14493 (N_14493,N_14308,N_14395);
or U14494 (N_14494,N_14310,N_14362);
or U14495 (N_14495,N_14384,N_14212);
nor U14496 (N_14496,N_14273,N_14297);
nor U14497 (N_14497,N_14218,N_14249);
nand U14498 (N_14498,N_14258,N_14251);
and U14499 (N_14499,N_14282,N_14233);
or U14500 (N_14500,N_14377,N_14360);
xor U14501 (N_14501,N_14291,N_14372);
and U14502 (N_14502,N_14289,N_14361);
and U14503 (N_14503,N_14204,N_14394);
nor U14504 (N_14504,N_14258,N_14230);
and U14505 (N_14505,N_14272,N_14247);
nand U14506 (N_14506,N_14231,N_14399);
nor U14507 (N_14507,N_14390,N_14379);
nand U14508 (N_14508,N_14243,N_14298);
nor U14509 (N_14509,N_14289,N_14382);
xnor U14510 (N_14510,N_14388,N_14285);
xnor U14511 (N_14511,N_14388,N_14229);
nand U14512 (N_14512,N_14376,N_14316);
nor U14513 (N_14513,N_14312,N_14304);
nor U14514 (N_14514,N_14315,N_14381);
nand U14515 (N_14515,N_14357,N_14212);
and U14516 (N_14516,N_14217,N_14378);
xnor U14517 (N_14517,N_14349,N_14374);
nand U14518 (N_14518,N_14207,N_14366);
or U14519 (N_14519,N_14289,N_14283);
xnor U14520 (N_14520,N_14380,N_14323);
or U14521 (N_14521,N_14369,N_14309);
and U14522 (N_14522,N_14396,N_14345);
nand U14523 (N_14523,N_14242,N_14236);
nor U14524 (N_14524,N_14329,N_14265);
xor U14525 (N_14525,N_14393,N_14341);
and U14526 (N_14526,N_14222,N_14230);
or U14527 (N_14527,N_14255,N_14233);
and U14528 (N_14528,N_14252,N_14276);
or U14529 (N_14529,N_14331,N_14396);
xnor U14530 (N_14530,N_14336,N_14354);
nand U14531 (N_14531,N_14366,N_14356);
nor U14532 (N_14532,N_14349,N_14279);
nor U14533 (N_14533,N_14399,N_14398);
and U14534 (N_14534,N_14221,N_14257);
nor U14535 (N_14535,N_14318,N_14225);
or U14536 (N_14536,N_14277,N_14279);
or U14537 (N_14537,N_14284,N_14267);
xnor U14538 (N_14538,N_14221,N_14315);
xnor U14539 (N_14539,N_14201,N_14297);
nand U14540 (N_14540,N_14243,N_14387);
nand U14541 (N_14541,N_14357,N_14311);
and U14542 (N_14542,N_14205,N_14250);
and U14543 (N_14543,N_14363,N_14297);
nor U14544 (N_14544,N_14349,N_14200);
nor U14545 (N_14545,N_14303,N_14332);
nand U14546 (N_14546,N_14283,N_14391);
or U14547 (N_14547,N_14278,N_14345);
and U14548 (N_14548,N_14384,N_14306);
nor U14549 (N_14549,N_14224,N_14329);
nor U14550 (N_14550,N_14353,N_14250);
xor U14551 (N_14551,N_14300,N_14270);
nand U14552 (N_14552,N_14367,N_14272);
or U14553 (N_14553,N_14296,N_14308);
nand U14554 (N_14554,N_14283,N_14210);
or U14555 (N_14555,N_14392,N_14325);
nor U14556 (N_14556,N_14390,N_14208);
and U14557 (N_14557,N_14300,N_14268);
and U14558 (N_14558,N_14259,N_14326);
or U14559 (N_14559,N_14310,N_14377);
and U14560 (N_14560,N_14333,N_14354);
nand U14561 (N_14561,N_14342,N_14329);
nand U14562 (N_14562,N_14393,N_14331);
and U14563 (N_14563,N_14273,N_14238);
nand U14564 (N_14564,N_14253,N_14316);
xnor U14565 (N_14565,N_14380,N_14337);
or U14566 (N_14566,N_14307,N_14335);
and U14567 (N_14567,N_14231,N_14346);
nor U14568 (N_14568,N_14238,N_14263);
xnor U14569 (N_14569,N_14313,N_14206);
xor U14570 (N_14570,N_14294,N_14325);
xnor U14571 (N_14571,N_14388,N_14242);
or U14572 (N_14572,N_14399,N_14261);
and U14573 (N_14573,N_14399,N_14244);
nor U14574 (N_14574,N_14285,N_14274);
and U14575 (N_14575,N_14318,N_14367);
xor U14576 (N_14576,N_14329,N_14385);
nor U14577 (N_14577,N_14366,N_14339);
nor U14578 (N_14578,N_14258,N_14273);
or U14579 (N_14579,N_14338,N_14255);
xnor U14580 (N_14580,N_14370,N_14390);
and U14581 (N_14581,N_14304,N_14230);
nand U14582 (N_14582,N_14202,N_14374);
xor U14583 (N_14583,N_14353,N_14266);
or U14584 (N_14584,N_14278,N_14249);
xor U14585 (N_14585,N_14299,N_14326);
and U14586 (N_14586,N_14363,N_14309);
and U14587 (N_14587,N_14251,N_14362);
and U14588 (N_14588,N_14287,N_14311);
and U14589 (N_14589,N_14342,N_14374);
nand U14590 (N_14590,N_14227,N_14368);
nand U14591 (N_14591,N_14323,N_14225);
nor U14592 (N_14592,N_14361,N_14283);
xor U14593 (N_14593,N_14370,N_14392);
xnor U14594 (N_14594,N_14317,N_14309);
xnor U14595 (N_14595,N_14220,N_14397);
xor U14596 (N_14596,N_14275,N_14267);
and U14597 (N_14597,N_14253,N_14208);
nor U14598 (N_14598,N_14372,N_14384);
nand U14599 (N_14599,N_14201,N_14362);
xnor U14600 (N_14600,N_14522,N_14528);
nand U14601 (N_14601,N_14524,N_14435);
or U14602 (N_14602,N_14513,N_14406);
nor U14603 (N_14603,N_14582,N_14558);
xor U14604 (N_14604,N_14447,N_14408);
nor U14605 (N_14605,N_14489,N_14465);
or U14606 (N_14606,N_14459,N_14490);
or U14607 (N_14607,N_14427,N_14595);
nand U14608 (N_14608,N_14552,N_14491);
xor U14609 (N_14609,N_14483,N_14419);
and U14610 (N_14610,N_14404,N_14423);
xor U14611 (N_14611,N_14461,N_14534);
and U14612 (N_14612,N_14498,N_14577);
nand U14613 (N_14613,N_14456,N_14551);
and U14614 (N_14614,N_14500,N_14583);
or U14615 (N_14615,N_14400,N_14514);
or U14616 (N_14616,N_14416,N_14542);
or U14617 (N_14617,N_14497,N_14414);
or U14618 (N_14618,N_14428,N_14563);
nand U14619 (N_14619,N_14469,N_14533);
and U14620 (N_14620,N_14562,N_14431);
nand U14621 (N_14621,N_14585,N_14474);
xor U14622 (N_14622,N_14550,N_14599);
or U14623 (N_14623,N_14467,N_14574);
or U14624 (N_14624,N_14426,N_14454);
and U14625 (N_14625,N_14412,N_14432);
nor U14626 (N_14626,N_14545,N_14557);
nor U14627 (N_14627,N_14564,N_14488);
xor U14628 (N_14628,N_14589,N_14567);
or U14629 (N_14629,N_14596,N_14548);
nor U14630 (N_14630,N_14455,N_14470);
nor U14631 (N_14631,N_14591,N_14410);
and U14632 (N_14632,N_14519,N_14578);
and U14633 (N_14633,N_14535,N_14573);
nor U14634 (N_14634,N_14468,N_14532);
nor U14635 (N_14635,N_14569,N_14521);
and U14636 (N_14636,N_14584,N_14531);
xnor U14637 (N_14637,N_14444,N_14553);
or U14638 (N_14638,N_14511,N_14429);
nand U14639 (N_14639,N_14415,N_14405);
or U14640 (N_14640,N_14523,N_14422);
nand U14641 (N_14641,N_14445,N_14592);
nor U14642 (N_14642,N_14438,N_14556);
xnor U14643 (N_14643,N_14440,N_14565);
nor U14644 (N_14644,N_14502,N_14443);
and U14645 (N_14645,N_14593,N_14417);
or U14646 (N_14646,N_14530,N_14418);
and U14647 (N_14647,N_14442,N_14499);
and U14648 (N_14648,N_14453,N_14590);
xor U14649 (N_14649,N_14463,N_14566);
and U14650 (N_14650,N_14407,N_14512);
or U14651 (N_14651,N_14402,N_14527);
nand U14652 (N_14652,N_14478,N_14568);
nor U14653 (N_14653,N_14559,N_14537);
xnor U14654 (N_14654,N_14579,N_14409);
nor U14655 (N_14655,N_14437,N_14554);
or U14656 (N_14656,N_14555,N_14525);
or U14657 (N_14657,N_14503,N_14448);
or U14658 (N_14658,N_14484,N_14581);
xor U14659 (N_14659,N_14520,N_14547);
nor U14660 (N_14660,N_14446,N_14403);
and U14661 (N_14661,N_14507,N_14411);
or U14662 (N_14662,N_14450,N_14439);
nor U14663 (N_14663,N_14496,N_14477);
and U14664 (N_14664,N_14560,N_14462);
nand U14665 (N_14665,N_14485,N_14549);
nor U14666 (N_14666,N_14433,N_14541);
nor U14667 (N_14667,N_14526,N_14480);
and U14668 (N_14668,N_14539,N_14586);
and U14669 (N_14669,N_14494,N_14505);
xnor U14670 (N_14670,N_14510,N_14451);
or U14671 (N_14671,N_14506,N_14464);
or U14672 (N_14672,N_14486,N_14504);
xnor U14673 (N_14673,N_14529,N_14436);
nand U14674 (N_14674,N_14473,N_14449);
nand U14675 (N_14675,N_14479,N_14430);
and U14676 (N_14676,N_14460,N_14466);
or U14677 (N_14677,N_14575,N_14472);
or U14678 (N_14678,N_14580,N_14594);
nor U14679 (N_14679,N_14536,N_14458);
nand U14680 (N_14680,N_14576,N_14561);
xor U14681 (N_14681,N_14475,N_14571);
or U14682 (N_14682,N_14441,N_14492);
and U14683 (N_14683,N_14413,N_14420);
nand U14684 (N_14684,N_14501,N_14597);
nor U14685 (N_14685,N_14495,N_14425);
or U14686 (N_14686,N_14570,N_14482);
or U14687 (N_14687,N_14515,N_14457);
xnor U14688 (N_14688,N_14509,N_14508);
nand U14689 (N_14689,N_14588,N_14572);
nor U14690 (N_14690,N_14517,N_14493);
xor U14691 (N_14691,N_14587,N_14476);
nand U14692 (N_14692,N_14424,N_14516);
or U14693 (N_14693,N_14421,N_14538);
or U14694 (N_14694,N_14543,N_14481);
nand U14695 (N_14695,N_14452,N_14518);
nor U14696 (N_14696,N_14434,N_14401);
and U14697 (N_14697,N_14471,N_14544);
and U14698 (N_14698,N_14540,N_14487);
nand U14699 (N_14699,N_14546,N_14598);
xor U14700 (N_14700,N_14556,N_14533);
nand U14701 (N_14701,N_14510,N_14549);
and U14702 (N_14702,N_14531,N_14445);
and U14703 (N_14703,N_14555,N_14421);
nor U14704 (N_14704,N_14487,N_14426);
and U14705 (N_14705,N_14472,N_14538);
nand U14706 (N_14706,N_14534,N_14507);
nor U14707 (N_14707,N_14439,N_14477);
and U14708 (N_14708,N_14475,N_14446);
and U14709 (N_14709,N_14410,N_14444);
nor U14710 (N_14710,N_14544,N_14494);
nor U14711 (N_14711,N_14432,N_14436);
nor U14712 (N_14712,N_14435,N_14505);
or U14713 (N_14713,N_14425,N_14491);
nor U14714 (N_14714,N_14448,N_14461);
nor U14715 (N_14715,N_14470,N_14583);
nor U14716 (N_14716,N_14434,N_14458);
nor U14717 (N_14717,N_14478,N_14411);
or U14718 (N_14718,N_14510,N_14588);
and U14719 (N_14719,N_14514,N_14430);
or U14720 (N_14720,N_14434,N_14496);
and U14721 (N_14721,N_14582,N_14456);
and U14722 (N_14722,N_14557,N_14504);
nand U14723 (N_14723,N_14417,N_14582);
and U14724 (N_14724,N_14469,N_14582);
nor U14725 (N_14725,N_14525,N_14577);
or U14726 (N_14726,N_14450,N_14567);
xnor U14727 (N_14727,N_14485,N_14538);
or U14728 (N_14728,N_14490,N_14584);
nor U14729 (N_14729,N_14518,N_14579);
nand U14730 (N_14730,N_14456,N_14486);
nor U14731 (N_14731,N_14570,N_14448);
xor U14732 (N_14732,N_14561,N_14430);
xnor U14733 (N_14733,N_14527,N_14557);
xor U14734 (N_14734,N_14411,N_14464);
and U14735 (N_14735,N_14537,N_14495);
nand U14736 (N_14736,N_14535,N_14507);
and U14737 (N_14737,N_14542,N_14565);
nand U14738 (N_14738,N_14459,N_14561);
and U14739 (N_14739,N_14444,N_14419);
or U14740 (N_14740,N_14471,N_14591);
and U14741 (N_14741,N_14458,N_14557);
nand U14742 (N_14742,N_14546,N_14437);
or U14743 (N_14743,N_14449,N_14499);
nand U14744 (N_14744,N_14504,N_14464);
and U14745 (N_14745,N_14571,N_14456);
nor U14746 (N_14746,N_14461,N_14445);
or U14747 (N_14747,N_14404,N_14525);
nor U14748 (N_14748,N_14584,N_14408);
nand U14749 (N_14749,N_14597,N_14419);
or U14750 (N_14750,N_14454,N_14449);
or U14751 (N_14751,N_14404,N_14471);
or U14752 (N_14752,N_14549,N_14558);
or U14753 (N_14753,N_14532,N_14566);
nand U14754 (N_14754,N_14492,N_14507);
nor U14755 (N_14755,N_14445,N_14454);
or U14756 (N_14756,N_14403,N_14546);
and U14757 (N_14757,N_14574,N_14543);
nor U14758 (N_14758,N_14457,N_14488);
nor U14759 (N_14759,N_14441,N_14402);
and U14760 (N_14760,N_14428,N_14550);
xor U14761 (N_14761,N_14414,N_14573);
xor U14762 (N_14762,N_14486,N_14535);
nor U14763 (N_14763,N_14503,N_14406);
nor U14764 (N_14764,N_14465,N_14522);
xnor U14765 (N_14765,N_14492,N_14593);
xnor U14766 (N_14766,N_14496,N_14419);
xnor U14767 (N_14767,N_14402,N_14545);
nor U14768 (N_14768,N_14587,N_14572);
or U14769 (N_14769,N_14412,N_14455);
xnor U14770 (N_14770,N_14557,N_14439);
nor U14771 (N_14771,N_14593,N_14596);
and U14772 (N_14772,N_14477,N_14513);
and U14773 (N_14773,N_14492,N_14400);
nand U14774 (N_14774,N_14420,N_14506);
nand U14775 (N_14775,N_14405,N_14596);
or U14776 (N_14776,N_14485,N_14405);
nand U14777 (N_14777,N_14581,N_14537);
and U14778 (N_14778,N_14597,N_14588);
xor U14779 (N_14779,N_14504,N_14521);
or U14780 (N_14780,N_14446,N_14552);
nor U14781 (N_14781,N_14427,N_14576);
or U14782 (N_14782,N_14511,N_14444);
nor U14783 (N_14783,N_14506,N_14554);
or U14784 (N_14784,N_14459,N_14592);
xor U14785 (N_14785,N_14415,N_14429);
and U14786 (N_14786,N_14567,N_14407);
nor U14787 (N_14787,N_14416,N_14469);
nand U14788 (N_14788,N_14563,N_14465);
nand U14789 (N_14789,N_14430,N_14429);
and U14790 (N_14790,N_14417,N_14543);
nand U14791 (N_14791,N_14471,N_14446);
nand U14792 (N_14792,N_14413,N_14523);
nor U14793 (N_14793,N_14542,N_14513);
nand U14794 (N_14794,N_14549,N_14530);
nand U14795 (N_14795,N_14509,N_14488);
nand U14796 (N_14796,N_14486,N_14437);
xnor U14797 (N_14797,N_14597,N_14506);
nor U14798 (N_14798,N_14447,N_14453);
nand U14799 (N_14799,N_14466,N_14533);
and U14800 (N_14800,N_14736,N_14757);
or U14801 (N_14801,N_14764,N_14679);
nor U14802 (N_14802,N_14718,N_14755);
and U14803 (N_14803,N_14789,N_14603);
nor U14804 (N_14804,N_14693,N_14681);
xnor U14805 (N_14805,N_14653,N_14624);
or U14806 (N_14806,N_14698,N_14713);
and U14807 (N_14807,N_14623,N_14708);
or U14808 (N_14808,N_14633,N_14619);
xor U14809 (N_14809,N_14786,N_14648);
nand U14810 (N_14810,N_14692,N_14672);
or U14811 (N_14811,N_14720,N_14735);
or U14812 (N_14812,N_14611,N_14750);
nand U14813 (N_14813,N_14643,N_14682);
nor U14814 (N_14814,N_14790,N_14635);
nand U14815 (N_14815,N_14730,N_14749);
xnor U14816 (N_14816,N_14765,N_14796);
nor U14817 (N_14817,N_14608,N_14724);
or U14818 (N_14818,N_14665,N_14660);
xnor U14819 (N_14819,N_14710,N_14671);
or U14820 (N_14820,N_14616,N_14719);
nor U14821 (N_14821,N_14763,N_14759);
or U14822 (N_14822,N_14678,N_14751);
nand U14823 (N_14823,N_14662,N_14631);
and U14824 (N_14824,N_14793,N_14715);
xnor U14825 (N_14825,N_14666,N_14744);
or U14826 (N_14826,N_14769,N_14747);
nor U14827 (N_14827,N_14761,N_14739);
or U14828 (N_14828,N_14798,N_14704);
nor U14829 (N_14829,N_14677,N_14687);
or U14830 (N_14830,N_14697,N_14756);
and U14831 (N_14831,N_14774,N_14647);
nor U14832 (N_14832,N_14770,N_14617);
and U14833 (N_14833,N_14725,N_14714);
nor U14834 (N_14834,N_14676,N_14620);
nor U14835 (N_14835,N_14614,N_14607);
nand U14836 (N_14836,N_14680,N_14783);
xnor U14837 (N_14837,N_14684,N_14663);
nand U14838 (N_14838,N_14615,N_14654);
nand U14839 (N_14839,N_14664,N_14667);
nand U14840 (N_14840,N_14705,N_14779);
nor U14841 (N_14841,N_14640,N_14722);
nor U14842 (N_14842,N_14748,N_14746);
and U14843 (N_14843,N_14696,N_14773);
xor U14844 (N_14844,N_14745,N_14772);
nor U14845 (N_14845,N_14702,N_14734);
nand U14846 (N_14846,N_14609,N_14797);
xnor U14847 (N_14847,N_14689,N_14784);
xnor U14848 (N_14848,N_14634,N_14733);
or U14849 (N_14849,N_14731,N_14629);
xnor U14850 (N_14850,N_14729,N_14781);
xnor U14851 (N_14851,N_14683,N_14659);
or U14852 (N_14852,N_14787,N_14741);
or U14853 (N_14853,N_14626,N_14701);
xor U14854 (N_14854,N_14602,N_14650);
or U14855 (N_14855,N_14776,N_14700);
or U14856 (N_14856,N_14768,N_14699);
nand U14857 (N_14857,N_14638,N_14632);
nand U14858 (N_14858,N_14760,N_14630);
nand U14859 (N_14859,N_14651,N_14613);
or U14860 (N_14860,N_14706,N_14782);
nor U14861 (N_14861,N_14743,N_14618);
nor U14862 (N_14862,N_14690,N_14775);
and U14863 (N_14863,N_14604,N_14753);
and U14864 (N_14864,N_14785,N_14726);
and U14865 (N_14865,N_14605,N_14661);
nand U14866 (N_14866,N_14621,N_14644);
xnor U14867 (N_14867,N_14754,N_14645);
nand U14868 (N_14868,N_14777,N_14709);
or U14869 (N_14869,N_14600,N_14766);
nor U14870 (N_14870,N_14762,N_14606);
nand U14871 (N_14871,N_14636,N_14742);
nand U14872 (N_14872,N_14794,N_14642);
or U14873 (N_14873,N_14688,N_14712);
nor U14874 (N_14874,N_14728,N_14727);
nor U14875 (N_14875,N_14788,N_14795);
nand U14876 (N_14876,N_14655,N_14691);
xor U14877 (N_14877,N_14639,N_14673);
xnor U14878 (N_14878,N_14695,N_14711);
and U14879 (N_14879,N_14658,N_14694);
xnor U14880 (N_14880,N_14792,N_14641);
xor U14881 (N_14881,N_14674,N_14601);
nor U14882 (N_14882,N_14652,N_14738);
and U14883 (N_14883,N_14737,N_14668);
xnor U14884 (N_14884,N_14675,N_14627);
and U14885 (N_14885,N_14740,N_14707);
nor U14886 (N_14886,N_14721,N_14732);
and U14887 (N_14887,N_14717,N_14685);
or U14888 (N_14888,N_14799,N_14622);
xor U14889 (N_14889,N_14752,N_14649);
nor U14890 (N_14890,N_14778,N_14771);
nor U14891 (N_14891,N_14791,N_14656);
nor U14892 (N_14892,N_14758,N_14612);
or U14893 (N_14893,N_14610,N_14686);
nand U14894 (N_14894,N_14767,N_14670);
nand U14895 (N_14895,N_14637,N_14723);
and U14896 (N_14896,N_14669,N_14703);
xor U14897 (N_14897,N_14646,N_14625);
or U14898 (N_14898,N_14716,N_14780);
or U14899 (N_14899,N_14628,N_14657);
xor U14900 (N_14900,N_14607,N_14611);
nand U14901 (N_14901,N_14740,N_14609);
nand U14902 (N_14902,N_14715,N_14697);
nand U14903 (N_14903,N_14726,N_14704);
nor U14904 (N_14904,N_14706,N_14615);
nand U14905 (N_14905,N_14775,N_14724);
nand U14906 (N_14906,N_14781,N_14683);
xor U14907 (N_14907,N_14729,N_14619);
nor U14908 (N_14908,N_14793,N_14620);
nand U14909 (N_14909,N_14748,N_14739);
nand U14910 (N_14910,N_14722,N_14724);
and U14911 (N_14911,N_14753,N_14736);
nand U14912 (N_14912,N_14732,N_14710);
nand U14913 (N_14913,N_14793,N_14744);
xnor U14914 (N_14914,N_14738,N_14773);
xnor U14915 (N_14915,N_14672,N_14682);
and U14916 (N_14916,N_14676,N_14765);
nor U14917 (N_14917,N_14765,N_14685);
or U14918 (N_14918,N_14683,N_14697);
nand U14919 (N_14919,N_14604,N_14623);
or U14920 (N_14920,N_14693,N_14649);
nand U14921 (N_14921,N_14612,N_14630);
nor U14922 (N_14922,N_14718,N_14633);
or U14923 (N_14923,N_14740,N_14616);
xnor U14924 (N_14924,N_14670,N_14642);
and U14925 (N_14925,N_14630,N_14795);
nor U14926 (N_14926,N_14712,N_14647);
or U14927 (N_14927,N_14699,N_14797);
and U14928 (N_14928,N_14619,N_14682);
nor U14929 (N_14929,N_14690,N_14722);
and U14930 (N_14930,N_14792,N_14684);
nor U14931 (N_14931,N_14639,N_14701);
xnor U14932 (N_14932,N_14784,N_14657);
and U14933 (N_14933,N_14717,N_14648);
and U14934 (N_14934,N_14653,N_14642);
xor U14935 (N_14935,N_14728,N_14785);
nand U14936 (N_14936,N_14732,N_14643);
xor U14937 (N_14937,N_14780,N_14753);
xnor U14938 (N_14938,N_14755,N_14642);
or U14939 (N_14939,N_14648,N_14791);
nand U14940 (N_14940,N_14781,N_14712);
nand U14941 (N_14941,N_14655,N_14750);
and U14942 (N_14942,N_14724,N_14755);
nand U14943 (N_14943,N_14653,N_14671);
and U14944 (N_14944,N_14605,N_14762);
and U14945 (N_14945,N_14682,N_14762);
xnor U14946 (N_14946,N_14613,N_14689);
and U14947 (N_14947,N_14714,N_14698);
and U14948 (N_14948,N_14750,N_14638);
nand U14949 (N_14949,N_14729,N_14761);
xor U14950 (N_14950,N_14769,N_14742);
nor U14951 (N_14951,N_14684,N_14642);
and U14952 (N_14952,N_14617,N_14790);
nand U14953 (N_14953,N_14682,N_14636);
nand U14954 (N_14954,N_14639,N_14742);
nor U14955 (N_14955,N_14704,N_14700);
nor U14956 (N_14956,N_14686,N_14659);
xor U14957 (N_14957,N_14737,N_14792);
nand U14958 (N_14958,N_14634,N_14729);
nand U14959 (N_14959,N_14777,N_14631);
nor U14960 (N_14960,N_14705,N_14656);
and U14961 (N_14961,N_14694,N_14786);
nor U14962 (N_14962,N_14687,N_14644);
or U14963 (N_14963,N_14677,N_14624);
or U14964 (N_14964,N_14649,N_14629);
nor U14965 (N_14965,N_14673,N_14640);
xor U14966 (N_14966,N_14781,N_14715);
and U14967 (N_14967,N_14701,N_14660);
or U14968 (N_14968,N_14798,N_14700);
and U14969 (N_14969,N_14663,N_14667);
or U14970 (N_14970,N_14660,N_14668);
and U14971 (N_14971,N_14780,N_14637);
nand U14972 (N_14972,N_14672,N_14656);
nand U14973 (N_14973,N_14676,N_14694);
or U14974 (N_14974,N_14608,N_14761);
nand U14975 (N_14975,N_14724,N_14679);
or U14976 (N_14976,N_14683,N_14731);
and U14977 (N_14977,N_14634,N_14645);
xnor U14978 (N_14978,N_14692,N_14696);
nand U14979 (N_14979,N_14777,N_14760);
nand U14980 (N_14980,N_14637,N_14763);
nand U14981 (N_14981,N_14694,N_14789);
nand U14982 (N_14982,N_14780,N_14713);
nand U14983 (N_14983,N_14680,N_14648);
nor U14984 (N_14984,N_14634,N_14714);
or U14985 (N_14985,N_14756,N_14641);
nor U14986 (N_14986,N_14763,N_14650);
nand U14987 (N_14987,N_14605,N_14741);
xnor U14988 (N_14988,N_14730,N_14607);
nand U14989 (N_14989,N_14767,N_14797);
nor U14990 (N_14990,N_14738,N_14799);
xor U14991 (N_14991,N_14727,N_14649);
nand U14992 (N_14992,N_14661,N_14658);
or U14993 (N_14993,N_14689,N_14619);
and U14994 (N_14994,N_14623,N_14701);
nor U14995 (N_14995,N_14781,N_14642);
xnor U14996 (N_14996,N_14743,N_14764);
or U14997 (N_14997,N_14700,N_14735);
nand U14998 (N_14998,N_14798,N_14614);
and U14999 (N_14999,N_14674,N_14680);
nand U15000 (N_15000,N_14986,N_14804);
nand U15001 (N_15001,N_14873,N_14963);
nor U15002 (N_15002,N_14938,N_14883);
and U15003 (N_15003,N_14815,N_14948);
or U15004 (N_15004,N_14824,N_14866);
or U15005 (N_15005,N_14863,N_14936);
nor U15006 (N_15006,N_14834,N_14969);
and U15007 (N_15007,N_14913,N_14980);
and U15008 (N_15008,N_14862,N_14809);
or U15009 (N_15009,N_14833,N_14868);
xnor U15010 (N_15010,N_14984,N_14922);
nand U15011 (N_15011,N_14907,N_14918);
nor U15012 (N_15012,N_14903,N_14819);
xnor U15013 (N_15013,N_14895,N_14844);
nor U15014 (N_15014,N_14972,N_14889);
nor U15015 (N_15015,N_14900,N_14941);
or U15016 (N_15016,N_14979,N_14995);
xnor U15017 (N_15017,N_14856,N_14961);
or U15018 (N_15018,N_14974,N_14964);
nor U15019 (N_15019,N_14908,N_14892);
nand U15020 (N_15020,N_14888,N_14827);
nand U15021 (N_15021,N_14914,N_14959);
and U15022 (N_15022,N_14848,N_14953);
xnor U15023 (N_15023,N_14939,N_14852);
xor U15024 (N_15024,N_14851,N_14929);
xnor U15025 (N_15025,N_14860,N_14812);
nand U15026 (N_15026,N_14949,N_14954);
and U15027 (N_15027,N_14957,N_14960);
xnor U15028 (N_15028,N_14881,N_14989);
or U15029 (N_15029,N_14885,N_14956);
or U15030 (N_15030,N_14991,N_14874);
and U15031 (N_15031,N_14917,N_14985);
nand U15032 (N_15032,N_14946,N_14968);
nor U15033 (N_15033,N_14909,N_14970);
nor U15034 (N_15034,N_14831,N_14951);
xor U15035 (N_15035,N_14867,N_14835);
xor U15036 (N_15036,N_14817,N_14988);
or U15037 (N_15037,N_14928,N_14864);
or U15038 (N_15038,N_14975,N_14923);
xnor U15039 (N_15039,N_14840,N_14807);
or U15040 (N_15040,N_14962,N_14933);
nor U15041 (N_15041,N_14816,N_14855);
nor U15042 (N_15042,N_14808,N_14967);
xnor U15043 (N_15043,N_14842,N_14832);
or U15044 (N_15044,N_14996,N_14841);
nor U15045 (N_15045,N_14976,N_14942);
nor U15046 (N_15046,N_14820,N_14994);
nor U15047 (N_15047,N_14981,N_14830);
xnor U15048 (N_15048,N_14891,N_14927);
nand U15049 (N_15049,N_14823,N_14875);
nand U15050 (N_15050,N_14910,N_14800);
and U15051 (N_15051,N_14806,N_14849);
xnor U15052 (N_15052,N_14897,N_14869);
nor U15053 (N_15053,N_14894,N_14836);
nand U15054 (N_15054,N_14999,N_14915);
or U15055 (N_15055,N_14876,N_14958);
xnor U15056 (N_15056,N_14886,N_14925);
nand U15057 (N_15057,N_14846,N_14983);
or U15058 (N_15058,N_14878,N_14802);
xor U15059 (N_15059,N_14921,N_14955);
xor U15060 (N_15060,N_14932,N_14977);
nand U15061 (N_15061,N_14896,N_14893);
nor U15062 (N_15062,N_14843,N_14839);
nor U15063 (N_15063,N_14899,N_14854);
and U15064 (N_15064,N_14850,N_14887);
nor U15065 (N_15065,N_14997,N_14898);
nor U15066 (N_15066,N_14947,N_14950);
nand U15067 (N_15067,N_14829,N_14879);
or U15068 (N_15068,N_14813,N_14814);
xnor U15069 (N_15069,N_14882,N_14890);
and U15070 (N_15070,N_14934,N_14987);
nor U15071 (N_15071,N_14911,N_14945);
or U15072 (N_15072,N_14861,N_14930);
or U15073 (N_15073,N_14828,N_14810);
nor U15074 (N_15074,N_14998,N_14912);
xnor U15075 (N_15075,N_14952,N_14931);
or U15076 (N_15076,N_14965,N_14811);
or U15077 (N_15077,N_14837,N_14880);
and U15078 (N_15078,N_14905,N_14982);
and U15079 (N_15079,N_14818,N_14966);
nand U15080 (N_15080,N_14884,N_14845);
xnor U15081 (N_15081,N_14902,N_14803);
and U15082 (N_15082,N_14920,N_14973);
nand U15083 (N_15083,N_14871,N_14877);
xnor U15084 (N_15084,N_14853,N_14857);
nand U15085 (N_15085,N_14978,N_14838);
or U15086 (N_15086,N_14971,N_14870);
nand U15087 (N_15087,N_14993,N_14865);
nor U15088 (N_15088,N_14935,N_14847);
xor U15089 (N_15089,N_14924,N_14992);
nor U15090 (N_15090,N_14826,N_14872);
nor U15091 (N_15091,N_14926,N_14916);
nand U15092 (N_15092,N_14919,N_14990);
xnor U15093 (N_15093,N_14822,N_14805);
nand U15094 (N_15094,N_14901,N_14937);
or U15095 (N_15095,N_14859,N_14904);
nor U15096 (N_15096,N_14825,N_14944);
nor U15097 (N_15097,N_14821,N_14858);
xor U15098 (N_15098,N_14940,N_14906);
xnor U15099 (N_15099,N_14943,N_14801);
and U15100 (N_15100,N_14812,N_14929);
xnor U15101 (N_15101,N_14913,N_14854);
nor U15102 (N_15102,N_14896,N_14984);
xnor U15103 (N_15103,N_14894,N_14921);
nand U15104 (N_15104,N_14892,N_14837);
or U15105 (N_15105,N_14849,N_14968);
or U15106 (N_15106,N_14840,N_14897);
nor U15107 (N_15107,N_14924,N_14953);
nand U15108 (N_15108,N_14917,N_14982);
nor U15109 (N_15109,N_14817,N_14839);
xor U15110 (N_15110,N_14907,N_14919);
and U15111 (N_15111,N_14982,N_14942);
nand U15112 (N_15112,N_14906,N_14856);
nand U15113 (N_15113,N_14811,N_14877);
nand U15114 (N_15114,N_14988,N_14979);
xnor U15115 (N_15115,N_14881,N_14923);
xnor U15116 (N_15116,N_14850,N_14873);
nor U15117 (N_15117,N_14947,N_14812);
nor U15118 (N_15118,N_14888,N_14971);
or U15119 (N_15119,N_14874,N_14857);
or U15120 (N_15120,N_14897,N_14973);
nand U15121 (N_15121,N_14900,N_14828);
or U15122 (N_15122,N_14924,N_14866);
or U15123 (N_15123,N_14845,N_14875);
or U15124 (N_15124,N_14867,N_14967);
or U15125 (N_15125,N_14870,N_14989);
nor U15126 (N_15126,N_14963,N_14962);
and U15127 (N_15127,N_14996,N_14845);
xnor U15128 (N_15128,N_14908,N_14931);
and U15129 (N_15129,N_14921,N_14918);
nor U15130 (N_15130,N_14879,N_14920);
and U15131 (N_15131,N_14902,N_14854);
nor U15132 (N_15132,N_14893,N_14954);
nand U15133 (N_15133,N_14836,N_14837);
xor U15134 (N_15134,N_14817,N_14813);
and U15135 (N_15135,N_14930,N_14969);
nor U15136 (N_15136,N_14985,N_14815);
nor U15137 (N_15137,N_14937,N_14859);
or U15138 (N_15138,N_14917,N_14829);
or U15139 (N_15139,N_14950,N_14849);
nor U15140 (N_15140,N_14848,N_14916);
nand U15141 (N_15141,N_14823,N_14877);
nand U15142 (N_15142,N_14931,N_14949);
or U15143 (N_15143,N_14985,N_14804);
nor U15144 (N_15144,N_14951,N_14927);
and U15145 (N_15145,N_14959,N_14800);
nor U15146 (N_15146,N_14848,N_14996);
nand U15147 (N_15147,N_14906,N_14827);
and U15148 (N_15148,N_14820,N_14868);
xnor U15149 (N_15149,N_14836,N_14847);
or U15150 (N_15150,N_14956,N_14981);
nor U15151 (N_15151,N_14916,N_14935);
nand U15152 (N_15152,N_14997,N_14860);
and U15153 (N_15153,N_14818,N_14821);
nor U15154 (N_15154,N_14871,N_14801);
xor U15155 (N_15155,N_14815,N_14859);
or U15156 (N_15156,N_14878,N_14908);
or U15157 (N_15157,N_14956,N_14882);
xnor U15158 (N_15158,N_14802,N_14865);
nand U15159 (N_15159,N_14893,N_14960);
or U15160 (N_15160,N_14982,N_14916);
and U15161 (N_15161,N_14828,N_14983);
nor U15162 (N_15162,N_14994,N_14936);
nor U15163 (N_15163,N_14811,N_14809);
nor U15164 (N_15164,N_14903,N_14954);
or U15165 (N_15165,N_14868,N_14858);
xor U15166 (N_15166,N_14888,N_14904);
xnor U15167 (N_15167,N_14826,N_14930);
nand U15168 (N_15168,N_14818,N_14907);
nand U15169 (N_15169,N_14807,N_14940);
nand U15170 (N_15170,N_14870,N_14939);
or U15171 (N_15171,N_14956,N_14922);
nor U15172 (N_15172,N_14806,N_14938);
nor U15173 (N_15173,N_14999,N_14861);
xor U15174 (N_15174,N_14955,N_14966);
and U15175 (N_15175,N_14930,N_14804);
nand U15176 (N_15176,N_14983,N_14894);
nor U15177 (N_15177,N_14903,N_14884);
nor U15178 (N_15178,N_14851,N_14994);
and U15179 (N_15179,N_14834,N_14870);
xnor U15180 (N_15180,N_14895,N_14938);
nand U15181 (N_15181,N_14872,N_14956);
xor U15182 (N_15182,N_14949,N_14942);
nor U15183 (N_15183,N_14984,N_14900);
nand U15184 (N_15184,N_14877,N_14980);
or U15185 (N_15185,N_14856,N_14912);
xor U15186 (N_15186,N_14833,N_14865);
nand U15187 (N_15187,N_14861,N_14913);
xor U15188 (N_15188,N_14913,N_14867);
nor U15189 (N_15189,N_14833,N_14843);
nor U15190 (N_15190,N_14837,N_14944);
nand U15191 (N_15191,N_14919,N_14880);
and U15192 (N_15192,N_14814,N_14924);
xnor U15193 (N_15193,N_14873,N_14836);
and U15194 (N_15194,N_14928,N_14952);
and U15195 (N_15195,N_14911,N_14981);
nand U15196 (N_15196,N_14802,N_14900);
nor U15197 (N_15197,N_14872,N_14937);
and U15198 (N_15198,N_14910,N_14801);
or U15199 (N_15199,N_14881,N_14876);
nor U15200 (N_15200,N_15092,N_15036);
nand U15201 (N_15201,N_15143,N_15152);
nor U15202 (N_15202,N_15177,N_15069);
xnor U15203 (N_15203,N_15073,N_15122);
or U15204 (N_15204,N_15068,N_15174);
nor U15205 (N_15205,N_15000,N_15017);
nand U15206 (N_15206,N_15136,N_15127);
nor U15207 (N_15207,N_15182,N_15134);
nor U15208 (N_15208,N_15018,N_15076);
and U15209 (N_15209,N_15031,N_15021);
nand U15210 (N_15210,N_15006,N_15121);
nand U15211 (N_15211,N_15113,N_15047);
xor U15212 (N_15212,N_15041,N_15198);
or U15213 (N_15213,N_15116,N_15057);
nor U15214 (N_15214,N_15070,N_15037);
or U15215 (N_15215,N_15150,N_15075);
and U15216 (N_15216,N_15154,N_15072);
nor U15217 (N_15217,N_15180,N_15137);
nand U15218 (N_15218,N_15146,N_15094);
and U15219 (N_15219,N_15188,N_15160);
and U15220 (N_15220,N_15176,N_15190);
or U15221 (N_15221,N_15118,N_15060);
or U15222 (N_15222,N_15003,N_15199);
nor U15223 (N_15223,N_15023,N_15084);
or U15224 (N_15224,N_15141,N_15131);
and U15225 (N_15225,N_15144,N_15055);
nand U15226 (N_15226,N_15033,N_15019);
and U15227 (N_15227,N_15042,N_15030);
nand U15228 (N_15228,N_15194,N_15135);
nor U15229 (N_15229,N_15096,N_15165);
and U15230 (N_15230,N_15081,N_15029);
nand U15231 (N_15231,N_15063,N_15022);
nand U15232 (N_15232,N_15120,N_15183);
xnor U15233 (N_15233,N_15139,N_15140);
xor U15234 (N_15234,N_15132,N_15123);
nand U15235 (N_15235,N_15151,N_15066);
or U15236 (N_15236,N_15192,N_15163);
xnor U15237 (N_15237,N_15179,N_15197);
or U15238 (N_15238,N_15125,N_15109);
or U15239 (N_15239,N_15166,N_15035);
and U15240 (N_15240,N_15161,N_15079);
or U15241 (N_15241,N_15027,N_15040);
xor U15242 (N_15242,N_15153,N_15115);
nand U15243 (N_15243,N_15148,N_15100);
nand U15244 (N_15244,N_15156,N_15046);
nor U15245 (N_15245,N_15053,N_15128);
and U15246 (N_15246,N_15196,N_15108);
xnor U15247 (N_15247,N_15187,N_15054);
and U15248 (N_15248,N_15039,N_15185);
xnor U15249 (N_15249,N_15082,N_15106);
nor U15250 (N_15250,N_15038,N_15062);
xor U15251 (N_15251,N_15104,N_15028);
or U15252 (N_15252,N_15168,N_15097);
nand U15253 (N_15253,N_15071,N_15091);
and U15254 (N_15254,N_15112,N_15184);
nand U15255 (N_15255,N_15189,N_15011);
xnor U15256 (N_15256,N_15049,N_15001);
and U15257 (N_15257,N_15181,N_15105);
or U15258 (N_15258,N_15119,N_15130);
or U15259 (N_15259,N_15157,N_15002);
nor U15260 (N_15260,N_15090,N_15102);
xor U15261 (N_15261,N_15064,N_15044);
nor U15262 (N_15262,N_15067,N_15024);
xor U15263 (N_15263,N_15186,N_15065);
and U15264 (N_15264,N_15142,N_15170);
xor U15265 (N_15265,N_15149,N_15074);
xnor U15266 (N_15266,N_15013,N_15010);
xor U15267 (N_15267,N_15095,N_15107);
and U15268 (N_15268,N_15009,N_15020);
nor U15269 (N_15269,N_15025,N_15159);
or U15270 (N_15270,N_15129,N_15083);
nand U15271 (N_15271,N_15193,N_15155);
nand U15272 (N_15272,N_15117,N_15147);
xor U15273 (N_15273,N_15012,N_15126);
or U15274 (N_15274,N_15026,N_15048);
nor U15275 (N_15275,N_15111,N_15171);
or U15276 (N_15276,N_15015,N_15110);
or U15277 (N_15277,N_15050,N_15089);
and U15278 (N_15278,N_15138,N_15167);
and U15279 (N_15279,N_15178,N_15034);
and U15280 (N_15280,N_15088,N_15043);
nand U15281 (N_15281,N_15191,N_15004);
nor U15282 (N_15282,N_15158,N_15169);
xnor U15283 (N_15283,N_15114,N_15059);
nor U15284 (N_15284,N_15016,N_15032);
nand U15285 (N_15285,N_15087,N_15078);
or U15286 (N_15286,N_15093,N_15051);
xnor U15287 (N_15287,N_15162,N_15103);
xor U15288 (N_15288,N_15085,N_15014);
or U15289 (N_15289,N_15145,N_15098);
nor U15290 (N_15290,N_15007,N_15175);
nor U15291 (N_15291,N_15172,N_15008);
nand U15292 (N_15292,N_15045,N_15124);
and U15293 (N_15293,N_15056,N_15133);
and U15294 (N_15294,N_15052,N_15080);
and U15295 (N_15295,N_15077,N_15005);
or U15296 (N_15296,N_15195,N_15061);
or U15297 (N_15297,N_15099,N_15101);
nand U15298 (N_15298,N_15164,N_15173);
nand U15299 (N_15299,N_15086,N_15058);
and U15300 (N_15300,N_15074,N_15195);
nor U15301 (N_15301,N_15010,N_15090);
nor U15302 (N_15302,N_15139,N_15080);
or U15303 (N_15303,N_15172,N_15127);
nand U15304 (N_15304,N_15112,N_15146);
nor U15305 (N_15305,N_15001,N_15114);
xor U15306 (N_15306,N_15037,N_15185);
xor U15307 (N_15307,N_15110,N_15088);
and U15308 (N_15308,N_15026,N_15072);
xor U15309 (N_15309,N_15062,N_15087);
nand U15310 (N_15310,N_15100,N_15133);
and U15311 (N_15311,N_15000,N_15191);
nand U15312 (N_15312,N_15032,N_15046);
or U15313 (N_15313,N_15072,N_15021);
and U15314 (N_15314,N_15019,N_15061);
nand U15315 (N_15315,N_15138,N_15028);
xnor U15316 (N_15316,N_15080,N_15006);
and U15317 (N_15317,N_15080,N_15128);
nor U15318 (N_15318,N_15095,N_15172);
nor U15319 (N_15319,N_15180,N_15170);
and U15320 (N_15320,N_15104,N_15065);
nand U15321 (N_15321,N_15140,N_15093);
xor U15322 (N_15322,N_15001,N_15075);
xnor U15323 (N_15323,N_15096,N_15098);
nand U15324 (N_15324,N_15128,N_15115);
nand U15325 (N_15325,N_15071,N_15151);
and U15326 (N_15326,N_15198,N_15067);
nor U15327 (N_15327,N_15169,N_15112);
and U15328 (N_15328,N_15057,N_15196);
xor U15329 (N_15329,N_15154,N_15138);
nand U15330 (N_15330,N_15001,N_15143);
and U15331 (N_15331,N_15078,N_15047);
and U15332 (N_15332,N_15069,N_15111);
and U15333 (N_15333,N_15120,N_15164);
nor U15334 (N_15334,N_15022,N_15036);
nor U15335 (N_15335,N_15101,N_15165);
or U15336 (N_15336,N_15049,N_15012);
xor U15337 (N_15337,N_15060,N_15144);
and U15338 (N_15338,N_15184,N_15194);
nand U15339 (N_15339,N_15165,N_15034);
and U15340 (N_15340,N_15118,N_15142);
xor U15341 (N_15341,N_15058,N_15043);
xor U15342 (N_15342,N_15043,N_15021);
or U15343 (N_15343,N_15159,N_15187);
xor U15344 (N_15344,N_15153,N_15114);
and U15345 (N_15345,N_15058,N_15047);
and U15346 (N_15346,N_15099,N_15035);
nor U15347 (N_15347,N_15128,N_15077);
nand U15348 (N_15348,N_15135,N_15034);
nor U15349 (N_15349,N_15067,N_15101);
xnor U15350 (N_15350,N_15106,N_15178);
or U15351 (N_15351,N_15195,N_15037);
nand U15352 (N_15352,N_15138,N_15184);
and U15353 (N_15353,N_15005,N_15035);
nor U15354 (N_15354,N_15067,N_15199);
nor U15355 (N_15355,N_15010,N_15091);
xnor U15356 (N_15356,N_15084,N_15130);
or U15357 (N_15357,N_15153,N_15127);
or U15358 (N_15358,N_15085,N_15096);
or U15359 (N_15359,N_15122,N_15026);
and U15360 (N_15360,N_15132,N_15087);
and U15361 (N_15361,N_15071,N_15125);
xor U15362 (N_15362,N_15103,N_15150);
xor U15363 (N_15363,N_15093,N_15180);
nor U15364 (N_15364,N_15034,N_15191);
or U15365 (N_15365,N_15110,N_15016);
and U15366 (N_15366,N_15034,N_15187);
nor U15367 (N_15367,N_15013,N_15081);
nor U15368 (N_15368,N_15125,N_15022);
nand U15369 (N_15369,N_15113,N_15196);
or U15370 (N_15370,N_15113,N_15170);
and U15371 (N_15371,N_15144,N_15104);
nand U15372 (N_15372,N_15085,N_15081);
and U15373 (N_15373,N_15153,N_15192);
or U15374 (N_15374,N_15078,N_15154);
xor U15375 (N_15375,N_15081,N_15108);
and U15376 (N_15376,N_15009,N_15097);
or U15377 (N_15377,N_15057,N_15081);
or U15378 (N_15378,N_15134,N_15114);
xor U15379 (N_15379,N_15003,N_15164);
nor U15380 (N_15380,N_15116,N_15078);
nor U15381 (N_15381,N_15080,N_15022);
and U15382 (N_15382,N_15088,N_15083);
xor U15383 (N_15383,N_15080,N_15196);
nor U15384 (N_15384,N_15122,N_15111);
nand U15385 (N_15385,N_15186,N_15039);
nor U15386 (N_15386,N_15191,N_15148);
nand U15387 (N_15387,N_15074,N_15042);
nor U15388 (N_15388,N_15076,N_15096);
or U15389 (N_15389,N_15125,N_15194);
and U15390 (N_15390,N_15144,N_15092);
nor U15391 (N_15391,N_15003,N_15080);
xor U15392 (N_15392,N_15048,N_15045);
and U15393 (N_15393,N_15100,N_15185);
and U15394 (N_15394,N_15195,N_15048);
and U15395 (N_15395,N_15044,N_15148);
and U15396 (N_15396,N_15181,N_15172);
nor U15397 (N_15397,N_15067,N_15044);
or U15398 (N_15398,N_15094,N_15143);
nor U15399 (N_15399,N_15191,N_15179);
nand U15400 (N_15400,N_15290,N_15367);
nor U15401 (N_15401,N_15259,N_15270);
xnor U15402 (N_15402,N_15256,N_15203);
nor U15403 (N_15403,N_15394,N_15271);
and U15404 (N_15404,N_15396,N_15248);
xor U15405 (N_15405,N_15235,N_15247);
and U15406 (N_15406,N_15294,N_15383);
or U15407 (N_15407,N_15331,N_15260);
and U15408 (N_15408,N_15308,N_15318);
nor U15409 (N_15409,N_15210,N_15324);
nor U15410 (N_15410,N_15232,N_15397);
or U15411 (N_15411,N_15365,N_15276);
xor U15412 (N_15412,N_15346,N_15336);
and U15413 (N_15413,N_15372,N_15305);
or U15414 (N_15414,N_15230,N_15373);
and U15415 (N_15415,N_15380,N_15381);
nand U15416 (N_15416,N_15240,N_15306);
nor U15417 (N_15417,N_15215,N_15309);
and U15418 (N_15418,N_15214,N_15272);
xnor U15419 (N_15419,N_15245,N_15342);
nand U15420 (N_15420,N_15241,N_15344);
xor U15421 (N_15421,N_15330,N_15275);
and U15422 (N_15422,N_15322,N_15281);
and U15423 (N_15423,N_15225,N_15224);
nor U15424 (N_15424,N_15303,N_15334);
xor U15425 (N_15425,N_15301,N_15356);
and U15426 (N_15426,N_15362,N_15253);
or U15427 (N_15427,N_15390,N_15277);
nand U15428 (N_15428,N_15384,N_15233);
nand U15429 (N_15429,N_15398,N_15350);
and U15430 (N_15430,N_15222,N_15218);
nand U15431 (N_15431,N_15378,N_15363);
nand U15432 (N_15432,N_15352,N_15343);
nand U15433 (N_15433,N_15300,N_15221);
xnor U15434 (N_15434,N_15286,N_15237);
nor U15435 (N_15435,N_15236,N_15246);
nor U15436 (N_15436,N_15377,N_15254);
xor U15437 (N_15437,N_15295,N_15202);
xnor U15438 (N_15438,N_15279,N_15333);
and U15439 (N_15439,N_15257,N_15291);
nor U15440 (N_15440,N_15302,N_15321);
and U15441 (N_15441,N_15311,N_15251);
xnor U15442 (N_15442,N_15340,N_15200);
nor U15443 (N_15443,N_15229,N_15348);
nand U15444 (N_15444,N_15347,N_15285);
nand U15445 (N_15445,N_15304,N_15369);
and U15446 (N_15446,N_15288,N_15274);
nand U15447 (N_15447,N_15354,N_15353);
and U15448 (N_15448,N_15283,N_15358);
or U15449 (N_15449,N_15375,N_15376);
and U15450 (N_15450,N_15234,N_15212);
nand U15451 (N_15451,N_15298,N_15357);
nor U15452 (N_15452,N_15307,N_15249);
and U15453 (N_15453,N_15223,N_15329);
nand U15454 (N_15454,N_15332,N_15255);
xor U15455 (N_15455,N_15266,N_15355);
or U15456 (N_15456,N_15287,N_15278);
or U15457 (N_15457,N_15268,N_15297);
nor U15458 (N_15458,N_15314,N_15361);
xnor U15459 (N_15459,N_15231,N_15315);
xnor U15460 (N_15460,N_15219,N_15360);
nor U15461 (N_15461,N_15280,N_15326);
nand U15462 (N_15462,N_15317,N_15393);
or U15463 (N_15463,N_15359,N_15216);
and U15464 (N_15464,N_15364,N_15328);
nor U15465 (N_15465,N_15220,N_15205);
nand U15466 (N_15466,N_15264,N_15292);
and U15467 (N_15467,N_15284,N_15258);
or U15468 (N_15468,N_15312,N_15267);
nor U15469 (N_15469,N_15389,N_15395);
nand U15470 (N_15470,N_15207,N_15316);
nand U15471 (N_15471,N_15265,N_15382);
nand U15472 (N_15472,N_15319,N_15368);
xnor U15473 (N_15473,N_15208,N_15327);
or U15474 (N_15474,N_15379,N_15226);
nand U15475 (N_15475,N_15320,N_15289);
or U15476 (N_15476,N_15388,N_15338);
or U15477 (N_15477,N_15341,N_15399);
and U15478 (N_15478,N_15228,N_15370);
xor U15479 (N_15479,N_15299,N_15293);
nor U15480 (N_15480,N_15325,N_15263);
nand U15481 (N_15481,N_15310,N_15201);
xor U15482 (N_15482,N_15204,N_15337);
or U15483 (N_15483,N_15313,N_15252);
xor U15484 (N_15484,N_15244,N_15261);
nand U15485 (N_15485,N_15211,N_15351);
or U15486 (N_15486,N_15349,N_15282);
xor U15487 (N_15487,N_15392,N_15243);
and U15488 (N_15488,N_15366,N_15262);
xor U15489 (N_15489,N_15385,N_15391);
or U15490 (N_15490,N_15335,N_15323);
or U15491 (N_15491,N_15227,N_15296);
or U15492 (N_15492,N_15213,N_15209);
xnor U15493 (N_15493,N_15371,N_15250);
nor U15494 (N_15494,N_15374,N_15206);
and U15495 (N_15495,N_15269,N_15217);
nor U15496 (N_15496,N_15387,N_15345);
and U15497 (N_15497,N_15238,N_15239);
xnor U15498 (N_15498,N_15273,N_15339);
nand U15499 (N_15499,N_15242,N_15386);
nand U15500 (N_15500,N_15367,N_15316);
nand U15501 (N_15501,N_15255,N_15267);
nand U15502 (N_15502,N_15374,N_15251);
and U15503 (N_15503,N_15208,N_15250);
or U15504 (N_15504,N_15295,N_15353);
or U15505 (N_15505,N_15267,N_15326);
nor U15506 (N_15506,N_15240,N_15245);
nand U15507 (N_15507,N_15392,N_15273);
or U15508 (N_15508,N_15342,N_15223);
and U15509 (N_15509,N_15256,N_15330);
nor U15510 (N_15510,N_15281,N_15328);
and U15511 (N_15511,N_15312,N_15284);
nor U15512 (N_15512,N_15325,N_15310);
xnor U15513 (N_15513,N_15335,N_15327);
nor U15514 (N_15514,N_15353,N_15381);
and U15515 (N_15515,N_15337,N_15314);
and U15516 (N_15516,N_15207,N_15210);
xnor U15517 (N_15517,N_15259,N_15252);
nand U15518 (N_15518,N_15292,N_15213);
nor U15519 (N_15519,N_15264,N_15315);
xor U15520 (N_15520,N_15211,N_15203);
nand U15521 (N_15521,N_15210,N_15384);
xnor U15522 (N_15522,N_15218,N_15316);
nand U15523 (N_15523,N_15239,N_15303);
xnor U15524 (N_15524,N_15338,N_15353);
xnor U15525 (N_15525,N_15304,N_15331);
nand U15526 (N_15526,N_15215,N_15297);
and U15527 (N_15527,N_15305,N_15223);
and U15528 (N_15528,N_15258,N_15253);
xor U15529 (N_15529,N_15218,N_15243);
xor U15530 (N_15530,N_15357,N_15355);
xnor U15531 (N_15531,N_15368,N_15366);
or U15532 (N_15532,N_15394,N_15379);
or U15533 (N_15533,N_15236,N_15216);
xor U15534 (N_15534,N_15286,N_15290);
xor U15535 (N_15535,N_15355,N_15367);
or U15536 (N_15536,N_15375,N_15216);
and U15537 (N_15537,N_15210,N_15385);
and U15538 (N_15538,N_15201,N_15336);
nor U15539 (N_15539,N_15355,N_15293);
nand U15540 (N_15540,N_15289,N_15287);
or U15541 (N_15541,N_15346,N_15364);
and U15542 (N_15542,N_15226,N_15316);
and U15543 (N_15543,N_15216,N_15237);
nor U15544 (N_15544,N_15308,N_15358);
or U15545 (N_15545,N_15369,N_15290);
xor U15546 (N_15546,N_15325,N_15220);
or U15547 (N_15547,N_15228,N_15234);
or U15548 (N_15548,N_15358,N_15381);
or U15549 (N_15549,N_15246,N_15397);
and U15550 (N_15550,N_15233,N_15211);
xor U15551 (N_15551,N_15240,N_15396);
and U15552 (N_15552,N_15248,N_15241);
nand U15553 (N_15553,N_15304,N_15367);
nand U15554 (N_15554,N_15329,N_15364);
nor U15555 (N_15555,N_15353,N_15341);
and U15556 (N_15556,N_15318,N_15244);
nand U15557 (N_15557,N_15237,N_15342);
and U15558 (N_15558,N_15220,N_15309);
nand U15559 (N_15559,N_15326,N_15324);
nand U15560 (N_15560,N_15394,N_15367);
nand U15561 (N_15561,N_15363,N_15349);
and U15562 (N_15562,N_15297,N_15219);
nand U15563 (N_15563,N_15246,N_15350);
and U15564 (N_15564,N_15293,N_15348);
or U15565 (N_15565,N_15329,N_15298);
xor U15566 (N_15566,N_15344,N_15272);
or U15567 (N_15567,N_15233,N_15203);
or U15568 (N_15568,N_15332,N_15324);
or U15569 (N_15569,N_15252,N_15341);
nand U15570 (N_15570,N_15382,N_15321);
and U15571 (N_15571,N_15364,N_15363);
and U15572 (N_15572,N_15365,N_15341);
xor U15573 (N_15573,N_15344,N_15260);
nand U15574 (N_15574,N_15342,N_15294);
xnor U15575 (N_15575,N_15217,N_15247);
nor U15576 (N_15576,N_15256,N_15214);
nand U15577 (N_15577,N_15375,N_15363);
nand U15578 (N_15578,N_15339,N_15395);
xor U15579 (N_15579,N_15266,N_15357);
nor U15580 (N_15580,N_15293,N_15345);
nor U15581 (N_15581,N_15325,N_15394);
or U15582 (N_15582,N_15220,N_15242);
nor U15583 (N_15583,N_15269,N_15353);
nor U15584 (N_15584,N_15388,N_15326);
and U15585 (N_15585,N_15223,N_15346);
xnor U15586 (N_15586,N_15204,N_15332);
or U15587 (N_15587,N_15396,N_15299);
nand U15588 (N_15588,N_15234,N_15237);
nor U15589 (N_15589,N_15210,N_15201);
nor U15590 (N_15590,N_15237,N_15259);
nor U15591 (N_15591,N_15374,N_15327);
and U15592 (N_15592,N_15280,N_15341);
nand U15593 (N_15593,N_15290,N_15291);
and U15594 (N_15594,N_15298,N_15211);
or U15595 (N_15595,N_15347,N_15379);
xnor U15596 (N_15596,N_15216,N_15353);
and U15597 (N_15597,N_15392,N_15250);
or U15598 (N_15598,N_15295,N_15214);
and U15599 (N_15599,N_15387,N_15257);
xor U15600 (N_15600,N_15572,N_15491);
nand U15601 (N_15601,N_15486,N_15476);
nor U15602 (N_15602,N_15426,N_15531);
nor U15603 (N_15603,N_15403,N_15550);
xnor U15604 (N_15604,N_15439,N_15582);
xnor U15605 (N_15605,N_15523,N_15433);
nand U15606 (N_15606,N_15505,N_15565);
nor U15607 (N_15607,N_15438,N_15463);
and U15608 (N_15608,N_15598,N_15448);
xnor U15609 (N_15609,N_15465,N_15497);
xor U15610 (N_15610,N_15455,N_15569);
and U15611 (N_15611,N_15578,N_15514);
or U15612 (N_15612,N_15493,N_15414);
xnor U15613 (N_15613,N_15545,N_15444);
xor U15614 (N_15614,N_15427,N_15561);
nand U15615 (N_15615,N_15404,N_15553);
xnor U15616 (N_15616,N_15466,N_15513);
nor U15617 (N_15617,N_15406,N_15434);
and U15618 (N_15618,N_15483,N_15554);
nor U15619 (N_15619,N_15504,N_15591);
and U15620 (N_15620,N_15415,N_15583);
nand U15621 (N_15621,N_15571,N_15492);
and U15622 (N_15622,N_15597,N_15515);
or U15623 (N_15623,N_15424,N_15484);
xor U15624 (N_15624,N_15435,N_15520);
nand U15625 (N_15625,N_15461,N_15447);
nor U15626 (N_15626,N_15499,N_15425);
or U15627 (N_15627,N_15446,N_15577);
and U15628 (N_15628,N_15579,N_15421);
and U15629 (N_15629,N_15451,N_15409);
nand U15630 (N_15630,N_15417,N_15580);
or U15631 (N_15631,N_15464,N_15459);
nand U15632 (N_15632,N_15538,N_15428);
xnor U15633 (N_15633,N_15477,N_15517);
and U15634 (N_15634,N_15462,N_15585);
or U15635 (N_15635,N_15423,N_15453);
and U15636 (N_15636,N_15599,N_15401);
nor U15637 (N_15637,N_15429,N_15593);
xor U15638 (N_15638,N_15402,N_15501);
and U15639 (N_15639,N_15551,N_15450);
or U15640 (N_15640,N_15460,N_15411);
xnor U15641 (N_15641,N_15524,N_15495);
and U15642 (N_15642,N_15546,N_15443);
and U15643 (N_15643,N_15519,N_15558);
nand U15644 (N_15644,N_15436,N_15416);
or U15645 (N_15645,N_15454,N_15563);
nand U15646 (N_15646,N_15407,N_15533);
and U15647 (N_15647,N_15543,N_15478);
and U15648 (N_15648,N_15473,N_15479);
nor U15649 (N_15649,N_15539,N_15573);
xor U15650 (N_15650,N_15430,N_15521);
xor U15651 (N_15651,N_15431,N_15456);
nor U15652 (N_15652,N_15555,N_15474);
nor U15653 (N_15653,N_15502,N_15516);
or U15654 (N_15654,N_15432,N_15467);
or U15655 (N_15655,N_15422,N_15472);
and U15656 (N_15656,N_15529,N_15544);
nand U15657 (N_15657,N_15511,N_15567);
nand U15658 (N_15658,N_15475,N_15530);
xor U15659 (N_15659,N_15413,N_15487);
and U15660 (N_15660,N_15595,N_15587);
nand U15661 (N_15661,N_15440,N_15457);
and U15662 (N_15662,N_15564,N_15522);
or U15663 (N_15663,N_15488,N_15468);
or U15664 (N_15664,N_15552,N_15542);
nor U15665 (N_15665,N_15452,N_15480);
nand U15666 (N_15666,N_15418,N_15449);
and U15667 (N_15667,N_15557,N_15586);
nand U15668 (N_15668,N_15471,N_15541);
and U15669 (N_15669,N_15581,N_15537);
xnor U15670 (N_15670,N_15548,N_15526);
and U15671 (N_15671,N_15534,N_15556);
or U15672 (N_15672,N_15496,N_15510);
and U15673 (N_15673,N_15420,N_15481);
and U15674 (N_15674,N_15584,N_15568);
nand U15675 (N_15675,N_15412,N_15528);
nand U15676 (N_15676,N_15527,N_15560);
nor U15677 (N_15677,N_15589,N_15574);
nand U15678 (N_15678,N_15503,N_15494);
nor U15679 (N_15679,N_15506,N_15470);
or U15680 (N_15680,N_15508,N_15535);
and U15681 (N_15681,N_15525,N_15559);
xor U15682 (N_15682,N_15490,N_15588);
nor U15683 (N_15683,N_15507,N_15498);
nand U15684 (N_15684,N_15445,N_15410);
nand U15685 (N_15685,N_15532,N_15576);
xor U15686 (N_15686,N_15518,N_15458);
or U15687 (N_15687,N_15592,N_15482);
or U15688 (N_15688,N_15419,N_15549);
xor U15689 (N_15689,N_15489,N_15400);
xor U15690 (N_15690,N_15566,N_15536);
or U15691 (N_15691,N_15469,N_15570);
nor U15692 (N_15692,N_15540,N_15562);
and U15693 (N_15693,N_15405,N_15485);
nand U15694 (N_15694,N_15437,N_15590);
nand U15695 (N_15695,N_15547,N_15575);
and U15696 (N_15696,N_15596,N_15441);
and U15697 (N_15697,N_15408,N_15500);
nand U15698 (N_15698,N_15442,N_15509);
nor U15699 (N_15699,N_15594,N_15512);
nand U15700 (N_15700,N_15414,N_15459);
xnor U15701 (N_15701,N_15562,N_15479);
or U15702 (N_15702,N_15554,N_15472);
or U15703 (N_15703,N_15503,N_15571);
nand U15704 (N_15704,N_15500,N_15554);
nor U15705 (N_15705,N_15591,N_15572);
xor U15706 (N_15706,N_15518,N_15558);
nor U15707 (N_15707,N_15491,N_15458);
or U15708 (N_15708,N_15504,N_15536);
and U15709 (N_15709,N_15432,N_15478);
nand U15710 (N_15710,N_15500,N_15414);
or U15711 (N_15711,N_15448,N_15501);
nor U15712 (N_15712,N_15415,N_15472);
and U15713 (N_15713,N_15448,N_15452);
nor U15714 (N_15714,N_15446,N_15505);
nor U15715 (N_15715,N_15554,N_15582);
or U15716 (N_15716,N_15543,N_15533);
nand U15717 (N_15717,N_15498,N_15459);
xor U15718 (N_15718,N_15489,N_15454);
nor U15719 (N_15719,N_15479,N_15583);
or U15720 (N_15720,N_15540,N_15439);
nor U15721 (N_15721,N_15477,N_15415);
nor U15722 (N_15722,N_15470,N_15404);
nand U15723 (N_15723,N_15563,N_15562);
xor U15724 (N_15724,N_15505,N_15400);
nor U15725 (N_15725,N_15575,N_15491);
nand U15726 (N_15726,N_15518,N_15500);
or U15727 (N_15727,N_15458,N_15463);
nand U15728 (N_15728,N_15506,N_15412);
nand U15729 (N_15729,N_15585,N_15599);
nand U15730 (N_15730,N_15585,N_15560);
or U15731 (N_15731,N_15530,N_15445);
xnor U15732 (N_15732,N_15516,N_15567);
nand U15733 (N_15733,N_15547,N_15442);
xnor U15734 (N_15734,N_15540,N_15538);
nor U15735 (N_15735,N_15516,N_15583);
xor U15736 (N_15736,N_15562,N_15448);
xnor U15737 (N_15737,N_15441,N_15590);
and U15738 (N_15738,N_15489,N_15455);
and U15739 (N_15739,N_15524,N_15585);
and U15740 (N_15740,N_15478,N_15505);
and U15741 (N_15741,N_15442,N_15531);
and U15742 (N_15742,N_15480,N_15507);
xnor U15743 (N_15743,N_15551,N_15481);
or U15744 (N_15744,N_15539,N_15557);
xor U15745 (N_15745,N_15542,N_15520);
or U15746 (N_15746,N_15592,N_15562);
or U15747 (N_15747,N_15480,N_15474);
nor U15748 (N_15748,N_15567,N_15584);
xnor U15749 (N_15749,N_15593,N_15484);
xnor U15750 (N_15750,N_15433,N_15563);
nand U15751 (N_15751,N_15521,N_15484);
nor U15752 (N_15752,N_15576,N_15421);
nor U15753 (N_15753,N_15526,N_15578);
and U15754 (N_15754,N_15495,N_15491);
and U15755 (N_15755,N_15463,N_15522);
nand U15756 (N_15756,N_15516,N_15507);
nand U15757 (N_15757,N_15479,N_15517);
xor U15758 (N_15758,N_15521,N_15453);
and U15759 (N_15759,N_15492,N_15406);
xnor U15760 (N_15760,N_15584,N_15534);
nand U15761 (N_15761,N_15568,N_15573);
or U15762 (N_15762,N_15415,N_15414);
nor U15763 (N_15763,N_15590,N_15583);
or U15764 (N_15764,N_15565,N_15576);
nor U15765 (N_15765,N_15400,N_15590);
and U15766 (N_15766,N_15436,N_15466);
xor U15767 (N_15767,N_15511,N_15490);
or U15768 (N_15768,N_15449,N_15456);
nand U15769 (N_15769,N_15545,N_15430);
nand U15770 (N_15770,N_15581,N_15597);
nor U15771 (N_15771,N_15507,N_15508);
nor U15772 (N_15772,N_15490,N_15465);
xnor U15773 (N_15773,N_15491,N_15597);
and U15774 (N_15774,N_15447,N_15542);
xnor U15775 (N_15775,N_15439,N_15404);
nand U15776 (N_15776,N_15497,N_15506);
or U15777 (N_15777,N_15552,N_15554);
and U15778 (N_15778,N_15425,N_15519);
nand U15779 (N_15779,N_15571,N_15535);
nor U15780 (N_15780,N_15440,N_15588);
and U15781 (N_15781,N_15415,N_15426);
or U15782 (N_15782,N_15465,N_15438);
nor U15783 (N_15783,N_15474,N_15473);
nand U15784 (N_15784,N_15457,N_15434);
nand U15785 (N_15785,N_15545,N_15539);
nand U15786 (N_15786,N_15517,N_15530);
nor U15787 (N_15787,N_15546,N_15577);
nor U15788 (N_15788,N_15463,N_15521);
and U15789 (N_15789,N_15529,N_15434);
and U15790 (N_15790,N_15576,N_15535);
nand U15791 (N_15791,N_15501,N_15405);
and U15792 (N_15792,N_15438,N_15468);
and U15793 (N_15793,N_15589,N_15573);
xor U15794 (N_15794,N_15514,N_15579);
or U15795 (N_15795,N_15555,N_15403);
nor U15796 (N_15796,N_15568,N_15462);
and U15797 (N_15797,N_15570,N_15410);
and U15798 (N_15798,N_15512,N_15499);
or U15799 (N_15799,N_15590,N_15472);
nor U15800 (N_15800,N_15705,N_15738);
xor U15801 (N_15801,N_15628,N_15683);
nand U15802 (N_15802,N_15758,N_15667);
nand U15803 (N_15803,N_15716,N_15782);
nor U15804 (N_15804,N_15687,N_15700);
nand U15805 (N_15805,N_15696,N_15650);
and U15806 (N_15806,N_15634,N_15702);
xnor U15807 (N_15807,N_15746,N_15659);
and U15808 (N_15808,N_15735,N_15772);
and U15809 (N_15809,N_15740,N_15610);
xor U15810 (N_15810,N_15651,N_15766);
and U15811 (N_15811,N_15707,N_15637);
and U15812 (N_15812,N_15642,N_15681);
nand U15813 (N_15813,N_15625,N_15655);
nor U15814 (N_15814,N_15682,N_15684);
and U15815 (N_15815,N_15711,N_15636);
xnor U15816 (N_15816,N_15670,N_15722);
and U15817 (N_15817,N_15741,N_15689);
xor U15818 (N_15818,N_15665,N_15754);
or U15819 (N_15819,N_15733,N_15720);
xor U15820 (N_15820,N_15619,N_15796);
nand U15821 (N_15821,N_15607,N_15676);
nor U15822 (N_15822,N_15747,N_15749);
and U15823 (N_15823,N_15729,N_15641);
nand U15824 (N_15824,N_15783,N_15752);
nor U15825 (N_15825,N_15627,N_15613);
nor U15826 (N_15826,N_15774,N_15620);
xor U15827 (N_15827,N_15664,N_15697);
nand U15828 (N_15828,N_15649,N_15715);
and U15829 (N_15829,N_15709,N_15694);
nor U15830 (N_15830,N_15653,N_15656);
or U15831 (N_15831,N_15616,N_15662);
and U15832 (N_15832,N_15635,N_15606);
nor U15833 (N_15833,N_15731,N_15660);
nor U15834 (N_15834,N_15788,N_15757);
nor U15835 (N_15835,N_15639,N_15703);
nand U15836 (N_15836,N_15767,N_15615);
or U15837 (N_15837,N_15668,N_15629);
nor U15838 (N_15838,N_15669,N_15604);
and U15839 (N_15839,N_15739,N_15602);
and U15840 (N_15840,N_15688,N_15623);
and U15841 (N_15841,N_15666,N_15730);
nand U15842 (N_15842,N_15727,N_15748);
xor U15843 (N_15843,N_15630,N_15769);
nand U15844 (N_15844,N_15719,N_15776);
nand U15845 (N_15845,N_15743,N_15793);
nand U15846 (N_15846,N_15777,N_15690);
and U15847 (N_15847,N_15771,N_15701);
xnor U15848 (N_15848,N_15675,N_15785);
nor U15849 (N_15849,N_15632,N_15732);
or U15850 (N_15850,N_15678,N_15768);
nor U15851 (N_15851,N_15618,N_15761);
or U15852 (N_15852,N_15611,N_15751);
xor U15853 (N_15853,N_15742,N_15648);
nor U15854 (N_15854,N_15646,N_15734);
nand U15855 (N_15855,N_15643,N_15764);
and U15856 (N_15856,N_15736,N_15704);
nand U15857 (N_15857,N_15721,N_15784);
nor U15858 (N_15858,N_15781,N_15633);
xnor U15859 (N_15859,N_15726,N_15755);
or U15860 (N_15860,N_15652,N_15760);
or U15861 (N_15861,N_15779,N_15685);
nand U15862 (N_15862,N_15798,N_15789);
xor U15863 (N_15863,N_15677,N_15797);
nand U15864 (N_15864,N_15601,N_15762);
nand U15865 (N_15865,N_15622,N_15644);
and U15866 (N_15866,N_15759,N_15647);
nor U15867 (N_15867,N_15708,N_15698);
xnor U15868 (N_15868,N_15718,N_15617);
or U15869 (N_15869,N_15737,N_15645);
and U15870 (N_15870,N_15671,N_15725);
or U15871 (N_15871,N_15672,N_15791);
or U15872 (N_15872,N_15706,N_15640);
nor U15873 (N_15873,N_15790,N_15614);
or U15874 (N_15874,N_15780,N_15608);
and U15875 (N_15875,N_15763,N_15673);
and U15876 (N_15876,N_15692,N_15654);
or U15877 (N_15877,N_15603,N_15714);
or U15878 (N_15878,N_15693,N_15723);
nand U15879 (N_15879,N_15679,N_15638);
or U15880 (N_15880,N_15699,N_15750);
or U15881 (N_15881,N_15728,N_15631);
or U15882 (N_15882,N_15663,N_15786);
nand U15883 (N_15883,N_15624,N_15756);
or U15884 (N_15884,N_15753,N_15745);
or U15885 (N_15885,N_15661,N_15600);
and U15886 (N_15886,N_15773,N_15657);
xnor U15887 (N_15887,N_15609,N_15724);
xnor U15888 (N_15888,N_15792,N_15710);
xnor U15889 (N_15889,N_15612,N_15775);
nand U15890 (N_15890,N_15778,N_15691);
or U15891 (N_15891,N_15695,N_15626);
nand U15892 (N_15892,N_15794,N_15713);
nor U15893 (N_15893,N_15686,N_15621);
or U15894 (N_15894,N_15717,N_15680);
nor U15895 (N_15895,N_15674,N_15744);
xor U15896 (N_15896,N_15795,N_15799);
xor U15897 (N_15897,N_15787,N_15765);
xor U15898 (N_15898,N_15712,N_15658);
or U15899 (N_15899,N_15605,N_15770);
xnor U15900 (N_15900,N_15614,N_15772);
nand U15901 (N_15901,N_15731,N_15728);
or U15902 (N_15902,N_15706,N_15780);
nor U15903 (N_15903,N_15676,N_15649);
nor U15904 (N_15904,N_15603,N_15693);
nand U15905 (N_15905,N_15764,N_15734);
nor U15906 (N_15906,N_15695,N_15741);
or U15907 (N_15907,N_15649,N_15678);
nor U15908 (N_15908,N_15735,N_15653);
and U15909 (N_15909,N_15687,N_15654);
xnor U15910 (N_15910,N_15632,N_15649);
and U15911 (N_15911,N_15786,N_15790);
or U15912 (N_15912,N_15784,N_15746);
nand U15913 (N_15913,N_15677,N_15695);
nor U15914 (N_15914,N_15794,N_15648);
or U15915 (N_15915,N_15737,N_15724);
and U15916 (N_15916,N_15792,N_15763);
nor U15917 (N_15917,N_15788,N_15716);
or U15918 (N_15918,N_15767,N_15750);
xor U15919 (N_15919,N_15664,N_15689);
and U15920 (N_15920,N_15629,N_15730);
nor U15921 (N_15921,N_15604,N_15751);
nand U15922 (N_15922,N_15717,N_15791);
nor U15923 (N_15923,N_15677,N_15673);
xnor U15924 (N_15924,N_15656,N_15684);
and U15925 (N_15925,N_15736,N_15790);
xor U15926 (N_15926,N_15667,N_15645);
xor U15927 (N_15927,N_15677,N_15765);
or U15928 (N_15928,N_15659,N_15764);
nor U15929 (N_15929,N_15702,N_15649);
nand U15930 (N_15930,N_15601,N_15661);
and U15931 (N_15931,N_15709,N_15655);
or U15932 (N_15932,N_15623,N_15612);
and U15933 (N_15933,N_15754,N_15758);
nor U15934 (N_15934,N_15635,N_15621);
nor U15935 (N_15935,N_15679,N_15630);
nand U15936 (N_15936,N_15667,N_15774);
xor U15937 (N_15937,N_15639,N_15610);
xor U15938 (N_15938,N_15631,N_15707);
nor U15939 (N_15939,N_15701,N_15662);
and U15940 (N_15940,N_15700,N_15690);
nand U15941 (N_15941,N_15642,N_15735);
or U15942 (N_15942,N_15763,N_15719);
nor U15943 (N_15943,N_15613,N_15705);
nand U15944 (N_15944,N_15795,N_15720);
xor U15945 (N_15945,N_15605,N_15750);
nand U15946 (N_15946,N_15646,N_15696);
nand U15947 (N_15947,N_15644,N_15666);
xnor U15948 (N_15948,N_15610,N_15702);
or U15949 (N_15949,N_15770,N_15702);
and U15950 (N_15950,N_15617,N_15664);
xor U15951 (N_15951,N_15619,N_15673);
nand U15952 (N_15952,N_15659,N_15675);
nor U15953 (N_15953,N_15771,N_15610);
nor U15954 (N_15954,N_15670,N_15693);
or U15955 (N_15955,N_15714,N_15743);
xnor U15956 (N_15956,N_15732,N_15675);
xor U15957 (N_15957,N_15720,N_15776);
nand U15958 (N_15958,N_15632,N_15678);
nor U15959 (N_15959,N_15626,N_15692);
and U15960 (N_15960,N_15732,N_15794);
or U15961 (N_15961,N_15696,N_15609);
xnor U15962 (N_15962,N_15742,N_15619);
or U15963 (N_15963,N_15787,N_15664);
or U15964 (N_15964,N_15612,N_15753);
xnor U15965 (N_15965,N_15625,N_15700);
nand U15966 (N_15966,N_15765,N_15663);
nor U15967 (N_15967,N_15641,N_15712);
nor U15968 (N_15968,N_15623,N_15776);
nand U15969 (N_15969,N_15644,N_15603);
nor U15970 (N_15970,N_15687,N_15716);
nor U15971 (N_15971,N_15744,N_15698);
xnor U15972 (N_15972,N_15647,N_15778);
xor U15973 (N_15973,N_15610,N_15665);
xnor U15974 (N_15974,N_15744,N_15782);
and U15975 (N_15975,N_15741,N_15633);
and U15976 (N_15976,N_15677,N_15766);
xor U15977 (N_15977,N_15613,N_15765);
xnor U15978 (N_15978,N_15665,N_15670);
and U15979 (N_15979,N_15601,N_15690);
nor U15980 (N_15980,N_15667,N_15764);
and U15981 (N_15981,N_15798,N_15757);
nor U15982 (N_15982,N_15799,N_15733);
nor U15983 (N_15983,N_15653,N_15651);
or U15984 (N_15984,N_15618,N_15711);
or U15985 (N_15985,N_15682,N_15775);
or U15986 (N_15986,N_15698,N_15751);
nor U15987 (N_15987,N_15731,N_15726);
or U15988 (N_15988,N_15797,N_15663);
and U15989 (N_15989,N_15772,N_15679);
nand U15990 (N_15990,N_15748,N_15777);
and U15991 (N_15991,N_15670,N_15765);
nor U15992 (N_15992,N_15623,N_15670);
nand U15993 (N_15993,N_15600,N_15680);
nor U15994 (N_15994,N_15640,N_15631);
nor U15995 (N_15995,N_15722,N_15770);
or U15996 (N_15996,N_15754,N_15685);
or U15997 (N_15997,N_15636,N_15786);
nand U15998 (N_15998,N_15644,N_15601);
or U15999 (N_15999,N_15617,N_15706);
nand U16000 (N_16000,N_15858,N_15974);
nand U16001 (N_16001,N_15920,N_15853);
xnor U16002 (N_16002,N_15895,N_15937);
and U16003 (N_16003,N_15868,N_15904);
or U16004 (N_16004,N_15813,N_15913);
nor U16005 (N_16005,N_15891,N_15875);
nor U16006 (N_16006,N_15983,N_15930);
nor U16007 (N_16007,N_15878,N_15941);
xnor U16008 (N_16008,N_15997,N_15899);
nand U16009 (N_16009,N_15900,N_15934);
nand U16010 (N_16010,N_15848,N_15940);
and U16011 (N_16011,N_15946,N_15885);
or U16012 (N_16012,N_15966,N_15821);
nand U16013 (N_16013,N_15811,N_15818);
and U16014 (N_16014,N_15842,N_15893);
or U16015 (N_16015,N_15881,N_15931);
nand U16016 (N_16016,N_15978,N_15854);
nor U16017 (N_16017,N_15929,N_15865);
nor U16018 (N_16018,N_15973,N_15877);
nand U16019 (N_16019,N_15950,N_15855);
or U16020 (N_16020,N_15820,N_15965);
and U16021 (N_16021,N_15844,N_15870);
or U16022 (N_16022,N_15898,N_15962);
and U16023 (N_16023,N_15902,N_15916);
nor U16024 (N_16024,N_15956,N_15847);
nor U16025 (N_16025,N_15939,N_15932);
nand U16026 (N_16026,N_15961,N_15824);
xnor U16027 (N_16027,N_15925,N_15955);
nand U16028 (N_16028,N_15918,N_15883);
and U16029 (N_16029,N_15839,N_15860);
xor U16030 (N_16030,N_15996,N_15981);
nand U16031 (N_16031,N_15863,N_15817);
nor U16032 (N_16032,N_15905,N_15910);
and U16033 (N_16033,N_15980,N_15917);
nor U16034 (N_16034,N_15985,N_15894);
nand U16035 (N_16035,N_15928,N_15835);
nor U16036 (N_16036,N_15810,N_15822);
nor U16037 (N_16037,N_15892,N_15846);
or U16038 (N_16038,N_15874,N_15942);
xor U16039 (N_16039,N_15889,N_15876);
nor U16040 (N_16040,N_15849,N_15919);
xnor U16041 (N_16041,N_15816,N_15888);
nand U16042 (N_16042,N_15924,N_15857);
nand U16043 (N_16043,N_15909,N_15958);
nand U16044 (N_16044,N_15825,N_15986);
or U16045 (N_16045,N_15836,N_15944);
and U16046 (N_16046,N_15989,N_15949);
nand U16047 (N_16047,N_15977,N_15993);
xnor U16048 (N_16048,N_15823,N_15968);
xor U16049 (N_16049,N_15851,N_15914);
nor U16050 (N_16050,N_15800,N_15880);
xor U16051 (N_16051,N_15864,N_15845);
or U16052 (N_16052,N_15871,N_15906);
nand U16053 (N_16053,N_15907,N_15819);
nor U16054 (N_16054,N_15938,N_15806);
and U16055 (N_16055,N_15945,N_15884);
nor U16056 (N_16056,N_15994,N_15867);
and U16057 (N_16057,N_15809,N_15984);
and U16058 (N_16058,N_15887,N_15943);
and U16059 (N_16059,N_15856,N_15999);
nand U16060 (N_16060,N_15990,N_15979);
nor U16061 (N_16061,N_15801,N_15843);
xor U16062 (N_16062,N_15890,N_15991);
nand U16063 (N_16063,N_15992,N_15897);
nand U16064 (N_16064,N_15953,N_15923);
nand U16065 (N_16065,N_15861,N_15969);
or U16066 (N_16066,N_15908,N_15982);
or U16067 (N_16067,N_15859,N_15911);
or U16068 (N_16068,N_15933,N_15957);
and U16069 (N_16069,N_15826,N_15869);
nand U16070 (N_16070,N_15840,N_15808);
and U16071 (N_16071,N_15954,N_15828);
xnor U16072 (N_16072,N_15952,N_15896);
xnor U16073 (N_16073,N_15995,N_15873);
nor U16074 (N_16074,N_15827,N_15951);
nand U16075 (N_16075,N_15832,N_15882);
nand U16076 (N_16076,N_15948,N_15830);
or U16077 (N_16077,N_15838,N_15936);
or U16078 (N_16078,N_15970,N_15975);
and U16079 (N_16079,N_15964,N_15915);
nor U16080 (N_16080,N_15972,N_15960);
xor U16081 (N_16081,N_15926,N_15862);
and U16082 (N_16082,N_15959,N_15922);
nand U16083 (N_16083,N_15852,N_15879);
and U16084 (N_16084,N_15805,N_15967);
nand U16085 (N_16085,N_15998,N_15837);
and U16086 (N_16086,N_15831,N_15872);
or U16087 (N_16087,N_15901,N_15834);
nor U16088 (N_16088,N_15815,N_15812);
xnor U16089 (N_16089,N_15976,N_15912);
or U16090 (N_16090,N_15921,N_15971);
nand U16091 (N_16091,N_15987,N_15903);
nor U16092 (N_16092,N_15850,N_15833);
xor U16093 (N_16093,N_15988,N_15841);
xnor U16094 (N_16094,N_15886,N_15866);
nand U16095 (N_16095,N_15802,N_15829);
or U16096 (N_16096,N_15935,N_15807);
xor U16097 (N_16097,N_15814,N_15803);
nor U16098 (N_16098,N_15947,N_15927);
and U16099 (N_16099,N_15963,N_15804);
nand U16100 (N_16100,N_15927,N_15939);
and U16101 (N_16101,N_15901,N_15884);
or U16102 (N_16102,N_15849,N_15938);
xnor U16103 (N_16103,N_15854,N_15990);
xor U16104 (N_16104,N_15953,N_15813);
nor U16105 (N_16105,N_15977,N_15985);
and U16106 (N_16106,N_15810,N_15832);
and U16107 (N_16107,N_15968,N_15812);
and U16108 (N_16108,N_15815,N_15962);
or U16109 (N_16109,N_15951,N_15995);
or U16110 (N_16110,N_15900,N_15935);
nor U16111 (N_16111,N_15974,N_15824);
nor U16112 (N_16112,N_15943,N_15987);
or U16113 (N_16113,N_15934,N_15941);
nor U16114 (N_16114,N_15986,N_15971);
nor U16115 (N_16115,N_15874,N_15983);
nand U16116 (N_16116,N_15977,N_15902);
nor U16117 (N_16117,N_15803,N_15996);
nand U16118 (N_16118,N_15930,N_15994);
nand U16119 (N_16119,N_15867,N_15856);
or U16120 (N_16120,N_15805,N_15974);
and U16121 (N_16121,N_15869,N_15898);
nor U16122 (N_16122,N_15825,N_15824);
nand U16123 (N_16123,N_15816,N_15978);
and U16124 (N_16124,N_15874,N_15902);
nand U16125 (N_16125,N_15866,N_15988);
xnor U16126 (N_16126,N_15866,N_15801);
nand U16127 (N_16127,N_15970,N_15802);
nor U16128 (N_16128,N_15848,N_15889);
and U16129 (N_16129,N_15906,N_15910);
and U16130 (N_16130,N_15933,N_15907);
nor U16131 (N_16131,N_15982,N_15999);
xor U16132 (N_16132,N_15890,N_15843);
nor U16133 (N_16133,N_15913,N_15987);
xor U16134 (N_16134,N_15809,N_15995);
nand U16135 (N_16135,N_15917,N_15889);
and U16136 (N_16136,N_15880,N_15986);
nand U16137 (N_16137,N_15968,N_15985);
and U16138 (N_16138,N_15942,N_15861);
nand U16139 (N_16139,N_15947,N_15814);
and U16140 (N_16140,N_15953,N_15935);
xor U16141 (N_16141,N_15991,N_15827);
nor U16142 (N_16142,N_15876,N_15826);
nand U16143 (N_16143,N_15808,N_15893);
nor U16144 (N_16144,N_15946,N_15836);
nor U16145 (N_16145,N_15914,N_15913);
nor U16146 (N_16146,N_15949,N_15995);
nand U16147 (N_16147,N_15935,N_15842);
nor U16148 (N_16148,N_15819,N_15897);
nor U16149 (N_16149,N_15838,N_15924);
and U16150 (N_16150,N_15867,N_15847);
and U16151 (N_16151,N_15924,N_15844);
or U16152 (N_16152,N_15837,N_15995);
xnor U16153 (N_16153,N_15942,N_15935);
or U16154 (N_16154,N_15928,N_15802);
nand U16155 (N_16155,N_15994,N_15964);
nor U16156 (N_16156,N_15821,N_15986);
nor U16157 (N_16157,N_15946,N_15802);
and U16158 (N_16158,N_15848,N_15927);
or U16159 (N_16159,N_15822,N_15917);
or U16160 (N_16160,N_15810,N_15872);
or U16161 (N_16161,N_15948,N_15825);
xor U16162 (N_16162,N_15891,N_15961);
or U16163 (N_16163,N_15874,N_15905);
or U16164 (N_16164,N_15873,N_15932);
nand U16165 (N_16165,N_15877,N_15969);
nor U16166 (N_16166,N_15995,N_15820);
nor U16167 (N_16167,N_15879,N_15883);
nand U16168 (N_16168,N_15903,N_15889);
or U16169 (N_16169,N_15858,N_15885);
xnor U16170 (N_16170,N_15881,N_15868);
nor U16171 (N_16171,N_15815,N_15916);
nand U16172 (N_16172,N_15997,N_15832);
xor U16173 (N_16173,N_15854,N_15931);
and U16174 (N_16174,N_15838,N_15912);
xor U16175 (N_16175,N_15849,N_15979);
or U16176 (N_16176,N_15916,N_15866);
nand U16177 (N_16177,N_15925,N_15850);
and U16178 (N_16178,N_15813,N_15925);
xor U16179 (N_16179,N_15870,N_15865);
or U16180 (N_16180,N_15970,N_15962);
xnor U16181 (N_16181,N_15943,N_15847);
or U16182 (N_16182,N_15922,N_15948);
nand U16183 (N_16183,N_15998,N_15980);
xor U16184 (N_16184,N_15935,N_15862);
nor U16185 (N_16185,N_15831,N_15916);
or U16186 (N_16186,N_15905,N_15952);
or U16187 (N_16187,N_15876,N_15801);
and U16188 (N_16188,N_15811,N_15822);
nand U16189 (N_16189,N_15840,N_15930);
or U16190 (N_16190,N_15902,N_15850);
and U16191 (N_16191,N_15880,N_15820);
xnor U16192 (N_16192,N_15817,N_15883);
nand U16193 (N_16193,N_15939,N_15854);
or U16194 (N_16194,N_15815,N_15952);
and U16195 (N_16195,N_15974,N_15925);
nor U16196 (N_16196,N_15812,N_15941);
nor U16197 (N_16197,N_15914,N_15992);
nor U16198 (N_16198,N_15801,N_15833);
xor U16199 (N_16199,N_15884,N_15876);
and U16200 (N_16200,N_16145,N_16160);
and U16201 (N_16201,N_16050,N_16091);
nand U16202 (N_16202,N_16189,N_16140);
nand U16203 (N_16203,N_16164,N_16194);
xnor U16204 (N_16204,N_16007,N_16128);
nor U16205 (N_16205,N_16174,N_16175);
or U16206 (N_16206,N_16073,N_16008);
and U16207 (N_16207,N_16019,N_16157);
or U16208 (N_16208,N_16125,N_16166);
xnor U16209 (N_16209,N_16100,N_16190);
and U16210 (N_16210,N_16184,N_16021);
xnor U16211 (N_16211,N_16047,N_16122);
xnor U16212 (N_16212,N_16120,N_16193);
nor U16213 (N_16213,N_16048,N_16144);
nand U16214 (N_16214,N_16037,N_16104);
or U16215 (N_16215,N_16153,N_16199);
or U16216 (N_16216,N_16110,N_16134);
nor U16217 (N_16217,N_16046,N_16126);
nand U16218 (N_16218,N_16023,N_16159);
or U16219 (N_16219,N_16163,N_16006);
xor U16220 (N_16220,N_16041,N_16105);
or U16221 (N_16221,N_16010,N_16026);
or U16222 (N_16222,N_16101,N_16152);
and U16223 (N_16223,N_16147,N_16085);
nor U16224 (N_16224,N_16186,N_16087);
nand U16225 (N_16225,N_16038,N_16177);
nor U16226 (N_16226,N_16055,N_16076);
xnor U16227 (N_16227,N_16098,N_16074);
xor U16228 (N_16228,N_16112,N_16197);
nor U16229 (N_16229,N_16158,N_16027);
and U16230 (N_16230,N_16011,N_16052);
and U16231 (N_16231,N_16078,N_16014);
nand U16232 (N_16232,N_16180,N_16179);
or U16233 (N_16233,N_16017,N_16141);
nor U16234 (N_16234,N_16151,N_16018);
xnor U16235 (N_16235,N_16167,N_16173);
nand U16236 (N_16236,N_16154,N_16040);
xor U16237 (N_16237,N_16088,N_16031);
or U16238 (N_16238,N_16139,N_16116);
nand U16239 (N_16239,N_16124,N_16161);
nor U16240 (N_16240,N_16070,N_16016);
nand U16241 (N_16241,N_16025,N_16115);
nand U16242 (N_16242,N_16036,N_16043);
nand U16243 (N_16243,N_16089,N_16168);
and U16244 (N_16244,N_16068,N_16042);
xnor U16245 (N_16245,N_16150,N_16107);
xnor U16246 (N_16246,N_16138,N_16015);
and U16247 (N_16247,N_16129,N_16072);
or U16248 (N_16248,N_16155,N_16066);
nand U16249 (N_16249,N_16001,N_16111);
xnor U16250 (N_16250,N_16137,N_16024);
nand U16251 (N_16251,N_16196,N_16080);
nand U16252 (N_16252,N_16192,N_16069);
and U16253 (N_16253,N_16053,N_16117);
nor U16254 (N_16254,N_16009,N_16132);
and U16255 (N_16255,N_16149,N_16049);
nand U16256 (N_16256,N_16058,N_16081);
nand U16257 (N_16257,N_16044,N_16012);
and U16258 (N_16258,N_16127,N_16004);
nand U16259 (N_16259,N_16002,N_16095);
nand U16260 (N_16260,N_16181,N_16035);
xnor U16261 (N_16261,N_16032,N_16030);
xor U16262 (N_16262,N_16109,N_16198);
and U16263 (N_16263,N_16057,N_16108);
nand U16264 (N_16264,N_16093,N_16013);
and U16265 (N_16265,N_16028,N_16133);
nor U16266 (N_16266,N_16079,N_16187);
xnor U16267 (N_16267,N_16106,N_16123);
and U16268 (N_16268,N_16195,N_16113);
xor U16269 (N_16269,N_16059,N_16082);
nor U16270 (N_16270,N_16130,N_16114);
xnor U16271 (N_16271,N_16103,N_16086);
nor U16272 (N_16272,N_16185,N_16062);
and U16273 (N_16273,N_16172,N_16063);
xor U16274 (N_16274,N_16099,N_16067);
or U16275 (N_16275,N_16084,N_16171);
xnor U16276 (N_16276,N_16170,N_16096);
xnor U16277 (N_16277,N_16065,N_16094);
nand U16278 (N_16278,N_16118,N_16136);
nand U16279 (N_16279,N_16119,N_16005);
and U16280 (N_16280,N_16188,N_16135);
nand U16281 (N_16281,N_16075,N_16156);
xor U16282 (N_16282,N_16003,N_16183);
nand U16283 (N_16283,N_16121,N_16022);
and U16284 (N_16284,N_16148,N_16131);
nor U16285 (N_16285,N_16029,N_16000);
nand U16286 (N_16286,N_16077,N_16165);
nand U16287 (N_16287,N_16039,N_16071);
xor U16288 (N_16288,N_16090,N_16020);
xor U16289 (N_16289,N_16143,N_16034);
xnor U16290 (N_16290,N_16083,N_16162);
nand U16291 (N_16291,N_16178,N_16142);
xor U16292 (N_16292,N_16191,N_16146);
xnor U16293 (N_16293,N_16051,N_16045);
xnor U16294 (N_16294,N_16102,N_16097);
nand U16295 (N_16295,N_16092,N_16061);
nand U16296 (N_16296,N_16176,N_16060);
nor U16297 (N_16297,N_16033,N_16056);
nand U16298 (N_16298,N_16182,N_16054);
nand U16299 (N_16299,N_16064,N_16169);
nand U16300 (N_16300,N_16151,N_16099);
nand U16301 (N_16301,N_16165,N_16153);
or U16302 (N_16302,N_16013,N_16047);
or U16303 (N_16303,N_16015,N_16037);
and U16304 (N_16304,N_16039,N_16023);
nor U16305 (N_16305,N_16099,N_16170);
nand U16306 (N_16306,N_16109,N_16017);
and U16307 (N_16307,N_16184,N_16044);
xor U16308 (N_16308,N_16163,N_16064);
nor U16309 (N_16309,N_16011,N_16020);
nor U16310 (N_16310,N_16038,N_16002);
nor U16311 (N_16311,N_16110,N_16059);
and U16312 (N_16312,N_16008,N_16163);
nor U16313 (N_16313,N_16193,N_16181);
nand U16314 (N_16314,N_16097,N_16052);
or U16315 (N_16315,N_16136,N_16122);
xnor U16316 (N_16316,N_16194,N_16110);
nand U16317 (N_16317,N_16181,N_16118);
nor U16318 (N_16318,N_16003,N_16098);
nand U16319 (N_16319,N_16042,N_16167);
or U16320 (N_16320,N_16130,N_16079);
nand U16321 (N_16321,N_16109,N_16179);
nor U16322 (N_16322,N_16079,N_16147);
nand U16323 (N_16323,N_16015,N_16183);
xor U16324 (N_16324,N_16064,N_16095);
nor U16325 (N_16325,N_16102,N_16131);
or U16326 (N_16326,N_16073,N_16045);
or U16327 (N_16327,N_16157,N_16188);
xnor U16328 (N_16328,N_16017,N_16020);
or U16329 (N_16329,N_16177,N_16006);
nand U16330 (N_16330,N_16094,N_16024);
nand U16331 (N_16331,N_16053,N_16122);
and U16332 (N_16332,N_16025,N_16015);
nand U16333 (N_16333,N_16046,N_16178);
nor U16334 (N_16334,N_16108,N_16154);
xnor U16335 (N_16335,N_16132,N_16074);
and U16336 (N_16336,N_16018,N_16191);
nor U16337 (N_16337,N_16006,N_16114);
nor U16338 (N_16338,N_16114,N_16064);
nor U16339 (N_16339,N_16171,N_16042);
xnor U16340 (N_16340,N_16017,N_16174);
and U16341 (N_16341,N_16162,N_16198);
xnor U16342 (N_16342,N_16001,N_16075);
nor U16343 (N_16343,N_16098,N_16195);
nand U16344 (N_16344,N_16155,N_16181);
and U16345 (N_16345,N_16069,N_16120);
xnor U16346 (N_16346,N_16117,N_16005);
xor U16347 (N_16347,N_16044,N_16174);
nor U16348 (N_16348,N_16167,N_16137);
nand U16349 (N_16349,N_16034,N_16004);
or U16350 (N_16350,N_16131,N_16147);
xnor U16351 (N_16351,N_16072,N_16097);
nand U16352 (N_16352,N_16184,N_16063);
or U16353 (N_16353,N_16110,N_16107);
and U16354 (N_16354,N_16004,N_16027);
nand U16355 (N_16355,N_16021,N_16060);
nor U16356 (N_16356,N_16051,N_16153);
nor U16357 (N_16357,N_16021,N_16120);
nor U16358 (N_16358,N_16106,N_16038);
and U16359 (N_16359,N_16105,N_16075);
xnor U16360 (N_16360,N_16185,N_16088);
nor U16361 (N_16361,N_16121,N_16124);
xnor U16362 (N_16362,N_16153,N_16132);
xnor U16363 (N_16363,N_16150,N_16175);
or U16364 (N_16364,N_16168,N_16059);
or U16365 (N_16365,N_16037,N_16177);
nor U16366 (N_16366,N_16016,N_16142);
nor U16367 (N_16367,N_16015,N_16161);
and U16368 (N_16368,N_16182,N_16044);
and U16369 (N_16369,N_16137,N_16103);
nand U16370 (N_16370,N_16175,N_16061);
nand U16371 (N_16371,N_16005,N_16120);
and U16372 (N_16372,N_16176,N_16011);
or U16373 (N_16373,N_16044,N_16180);
nor U16374 (N_16374,N_16053,N_16067);
nor U16375 (N_16375,N_16192,N_16047);
or U16376 (N_16376,N_16029,N_16004);
or U16377 (N_16377,N_16045,N_16106);
and U16378 (N_16378,N_16136,N_16051);
nand U16379 (N_16379,N_16192,N_16070);
or U16380 (N_16380,N_16026,N_16078);
nand U16381 (N_16381,N_16071,N_16046);
and U16382 (N_16382,N_16196,N_16130);
xnor U16383 (N_16383,N_16126,N_16052);
and U16384 (N_16384,N_16177,N_16016);
or U16385 (N_16385,N_16015,N_16171);
or U16386 (N_16386,N_16005,N_16004);
and U16387 (N_16387,N_16015,N_16097);
nand U16388 (N_16388,N_16129,N_16065);
or U16389 (N_16389,N_16195,N_16117);
and U16390 (N_16390,N_16105,N_16083);
or U16391 (N_16391,N_16091,N_16071);
and U16392 (N_16392,N_16089,N_16027);
nand U16393 (N_16393,N_16159,N_16075);
nand U16394 (N_16394,N_16037,N_16128);
nand U16395 (N_16395,N_16083,N_16121);
nand U16396 (N_16396,N_16128,N_16114);
nor U16397 (N_16397,N_16167,N_16144);
and U16398 (N_16398,N_16125,N_16191);
and U16399 (N_16399,N_16045,N_16178);
nand U16400 (N_16400,N_16388,N_16367);
nor U16401 (N_16401,N_16354,N_16283);
and U16402 (N_16402,N_16228,N_16278);
nand U16403 (N_16403,N_16356,N_16211);
and U16404 (N_16404,N_16339,N_16382);
nor U16405 (N_16405,N_16243,N_16311);
nor U16406 (N_16406,N_16365,N_16391);
nor U16407 (N_16407,N_16234,N_16351);
xor U16408 (N_16408,N_16308,N_16309);
xnor U16409 (N_16409,N_16397,N_16380);
xnor U16410 (N_16410,N_16205,N_16390);
or U16411 (N_16411,N_16206,N_16305);
xor U16412 (N_16412,N_16338,N_16257);
nor U16413 (N_16413,N_16302,N_16252);
xor U16414 (N_16414,N_16202,N_16284);
xnor U16415 (N_16415,N_16248,N_16345);
nand U16416 (N_16416,N_16393,N_16240);
or U16417 (N_16417,N_16220,N_16370);
and U16418 (N_16418,N_16296,N_16207);
or U16419 (N_16419,N_16265,N_16259);
and U16420 (N_16420,N_16256,N_16232);
nand U16421 (N_16421,N_16327,N_16251);
xnor U16422 (N_16422,N_16363,N_16294);
nor U16423 (N_16423,N_16225,N_16318);
and U16424 (N_16424,N_16263,N_16316);
nand U16425 (N_16425,N_16266,N_16239);
or U16426 (N_16426,N_16314,N_16340);
nor U16427 (N_16427,N_16379,N_16281);
nor U16428 (N_16428,N_16262,N_16387);
xor U16429 (N_16429,N_16398,N_16396);
or U16430 (N_16430,N_16261,N_16291);
xor U16431 (N_16431,N_16204,N_16324);
xor U16432 (N_16432,N_16213,N_16233);
nand U16433 (N_16433,N_16229,N_16353);
nor U16434 (N_16434,N_16306,N_16389);
and U16435 (N_16435,N_16369,N_16272);
and U16436 (N_16436,N_16254,N_16292);
and U16437 (N_16437,N_16235,N_16384);
xor U16438 (N_16438,N_16315,N_16226);
and U16439 (N_16439,N_16361,N_16275);
or U16440 (N_16440,N_16344,N_16212);
or U16441 (N_16441,N_16303,N_16236);
xnor U16442 (N_16442,N_16210,N_16383);
nor U16443 (N_16443,N_16376,N_16289);
and U16444 (N_16444,N_16279,N_16224);
nand U16445 (N_16445,N_16247,N_16322);
and U16446 (N_16446,N_16216,N_16313);
xor U16447 (N_16447,N_16374,N_16246);
nand U16448 (N_16448,N_16310,N_16218);
nor U16449 (N_16449,N_16343,N_16319);
and U16450 (N_16450,N_16372,N_16375);
or U16451 (N_16451,N_16268,N_16307);
or U16452 (N_16452,N_16200,N_16287);
or U16453 (N_16453,N_16300,N_16337);
or U16454 (N_16454,N_16295,N_16329);
xor U16455 (N_16455,N_16215,N_16352);
nor U16456 (N_16456,N_16342,N_16255);
nor U16457 (N_16457,N_16341,N_16323);
or U16458 (N_16458,N_16333,N_16286);
nor U16459 (N_16459,N_16317,N_16273);
or U16460 (N_16460,N_16325,N_16260);
and U16461 (N_16461,N_16399,N_16222);
and U16462 (N_16462,N_16395,N_16368);
nand U16463 (N_16463,N_16297,N_16330);
or U16464 (N_16464,N_16230,N_16270);
or U16465 (N_16465,N_16385,N_16238);
or U16466 (N_16466,N_16277,N_16299);
nor U16467 (N_16467,N_16364,N_16274);
and U16468 (N_16468,N_16269,N_16386);
xor U16469 (N_16469,N_16201,N_16332);
or U16470 (N_16470,N_16366,N_16392);
and U16471 (N_16471,N_16231,N_16326);
nand U16472 (N_16472,N_16328,N_16250);
or U16473 (N_16473,N_16267,N_16336);
nor U16474 (N_16474,N_16355,N_16357);
xnor U16475 (N_16475,N_16237,N_16264);
nand U16476 (N_16476,N_16242,N_16362);
nand U16477 (N_16477,N_16301,N_16358);
nand U16478 (N_16478,N_16290,N_16217);
nand U16479 (N_16479,N_16394,N_16282);
nor U16480 (N_16480,N_16304,N_16223);
xor U16481 (N_16481,N_16249,N_16335);
or U16482 (N_16482,N_16298,N_16214);
nand U16483 (N_16483,N_16293,N_16244);
xnor U16484 (N_16484,N_16377,N_16258);
or U16485 (N_16485,N_16373,N_16203);
xnor U16486 (N_16486,N_16360,N_16285);
or U16487 (N_16487,N_16271,N_16221);
nand U16488 (N_16488,N_16227,N_16334);
nor U16489 (N_16489,N_16371,N_16349);
nand U16490 (N_16490,N_16321,N_16381);
or U16491 (N_16491,N_16378,N_16346);
nand U16492 (N_16492,N_16320,N_16245);
nor U16493 (N_16493,N_16241,N_16209);
nor U16494 (N_16494,N_16288,N_16348);
and U16495 (N_16495,N_16359,N_16350);
xor U16496 (N_16496,N_16253,N_16219);
xor U16497 (N_16497,N_16208,N_16331);
and U16498 (N_16498,N_16347,N_16312);
xor U16499 (N_16499,N_16276,N_16280);
or U16500 (N_16500,N_16336,N_16264);
nand U16501 (N_16501,N_16385,N_16220);
and U16502 (N_16502,N_16230,N_16351);
nand U16503 (N_16503,N_16278,N_16358);
xor U16504 (N_16504,N_16348,N_16200);
nand U16505 (N_16505,N_16252,N_16207);
xnor U16506 (N_16506,N_16297,N_16218);
and U16507 (N_16507,N_16352,N_16369);
or U16508 (N_16508,N_16310,N_16278);
xnor U16509 (N_16509,N_16294,N_16329);
or U16510 (N_16510,N_16338,N_16371);
and U16511 (N_16511,N_16277,N_16369);
nand U16512 (N_16512,N_16274,N_16243);
or U16513 (N_16513,N_16359,N_16254);
or U16514 (N_16514,N_16323,N_16234);
xnor U16515 (N_16515,N_16263,N_16372);
nand U16516 (N_16516,N_16231,N_16291);
nand U16517 (N_16517,N_16363,N_16236);
nand U16518 (N_16518,N_16247,N_16214);
nand U16519 (N_16519,N_16366,N_16231);
xor U16520 (N_16520,N_16280,N_16348);
or U16521 (N_16521,N_16316,N_16341);
nor U16522 (N_16522,N_16379,N_16243);
nor U16523 (N_16523,N_16232,N_16211);
xnor U16524 (N_16524,N_16380,N_16396);
or U16525 (N_16525,N_16211,N_16398);
and U16526 (N_16526,N_16357,N_16312);
nand U16527 (N_16527,N_16310,N_16281);
and U16528 (N_16528,N_16269,N_16224);
or U16529 (N_16529,N_16307,N_16281);
nand U16530 (N_16530,N_16372,N_16350);
nor U16531 (N_16531,N_16256,N_16238);
nand U16532 (N_16532,N_16200,N_16333);
nor U16533 (N_16533,N_16228,N_16279);
nor U16534 (N_16534,N_16319,N_16302);
nor U16535 (N_16535,N_16245,N_16363);
nor U16536 (N_16536,N_16247,N_16346);
xor U16537 (N_16537,N_16281,N_16360);
nor U16538 (N_16538,N_16355,N_16231);
and U16539 (N_16539,N_16376,N_16372);
xnor U16540 (N_16540,N_16284,N_16317);
or U16541 (N_16541,N_16375,N_16308);
nand U16542 (N_16542,N_16330,N_16220);
xor U16543 (N_16543,N_16319,N_16321);
or U16544 (N_16544,N_16283,N_16288);
and U16545 (N_16545,N_16376,N_16229);
nor U16546 (N_16546,N_16348,N_16246);
xor U16547 (N_16547,N_16251,N_16259);
or U16548 (N_16548,N_16380,N_16258);
and U16549 (N_16549,N_16329,N_16278);
or U16550 (N_16550,N_16278,N_16347);
xnor U16551 (N_16551,N_16300,N_16247);
nand U16552 (N_16552,N_16397,N_16224);
nand U16553 (N_16553,N_16351,N_16307);
or U16554 (N_16554,N_16349,N_16270);
or U16555 (N_16555,N_16214,N_16258);
xnor U16556 (N_16556,N_16319,N_16285);
and U16557 (N_16557,N_16241,N_16311);
nand U16558 (N_16558,N_16328,N_16238);
xor U16559 (N_16559,N_16248,N_16243);
nor U16560 (N_16560,N_16315,N_16230);
and U16561 (N_16561,N_16282,N_16299);
nor U16562 (N_16562,N_16383,N_16305);
and U16563 (N_16563,N_16280,N_16309);
xor U16564 (N_16564,N_16263,N_16225);
nor U16565 (N_16565,N_16274,N_16215);
and U16566 (N_16566,N_16323,N_16325);
and U16567 (N_16567,N_16284,N_16362);
nor U16568 (N_16568,N_16330,N_16212);
or U16569 (N_16569,N_16262,N_16351);
or U16570 (N_16570,N_16202,N_16382);
or U16571 (N_16571,N_16311,N_16396);
xnor U16572 (N_16572,N_16210,N_16294);
or U16573 (N_16573,N_16377,N_16314);
xor U16574 (N_16574,N_16330,N_16262);
or U16575 (N_16575,N_16298,N_16274);
nor U16576 (N_16576,N_16368,N_16293);
and U16577 (N_16577,N_16393,N_16293);
or U16578 (N_16578,N_16271,N_16320);
nand U16579 (N_16579,N_16390,N_16228);
or U16580 (N_16580,N_16245,N_16307);
xor U16581 (N_16581,N_16209,N_16381);
and U16582 (N_16582,N_16300,N_16353);
nor U16583 (N_16583,N_16388,N_16331);
nor U16584 (N_16584,N_16269,N_16382);
nor U16585 (N_16585,N_16377,N_16283);
xor U16586 (N_16586,N_16209,N_16389);
and U16587 (N_16587,N_16387,N_16371);
nor U16588 (N_16588,N_16319,N_16204);
xor U16589 (N_16589,N_16390,N_16344);
nand U16590 (N_16590,N_16243,N_16384);
nand U16591 (N_16591,N_16227,N_16215);
xor U16592 (N_16592,N_16310,N_16394);
nor U16593 (N_16593,N_16326,N_16258);
and U16594 (N_16594,N_16240,N_16395);
or U16595 (N_16595,N_16359,N_16319);
and U16596 (N_16596,N_16260,N_16206);
nor U16597 (N_16597,N_16319,N_16211);
nor U16598 (N_16598,N_16279,N_16324);
or U16599 (N_16599,N_16348,N_16388);
nand U16600 (N_16600,N_16483,N_16428);
nand U16601 (N_16601,N_16499,N_16575);
nand U16602 (N_16602,N_16524,N_16487);
nand U16603 (N_16603,N_16564,N_16450);
and U16604 (N_16604,N_16508,N_16597);
nor U16605 (N_16605,N_16584,N_16580);
and U16606 (N_16606,N_16406,N_16594);
xnor U16607 (N_16607,N_16542,N_16573);
and U16608 (N_16608,N_16417,N_16460);
xnor U16609 (N_16609,N_16457,N_16449);
nand U16610 (N_16610,N_16528,N_16545);
or U16611 (N_16611,N_16434,N_16492);
and U16612 (N_16612,N_16431,N_16405);
and U16613 (N_16613,N_16489,N_16536);
and U16614 (N_16614,N_16500,N_16469);
and U16615 (N_16615,N_16415,N_16538);
or U16616 (N_16616,N_16433,N_16541);
nor U16617 (N_16617,N_16470,N_16485);
xnor U16618 (N_16618,N_16570,N_16518);
nor U16619 (N_16619,N_16586,N_16446);
nand U16620 (N_16620,N_16421,N_16409);
xnor U16621 (N_16621,N_16475,N_16474);
xnor U16622 (N_16622,N_16582,N_16526);
nor U16623 (N_16623,N_16407,N_16402);
xnor U16624 (N_16624,N_16412,N_16523);
nor U16625 (N_16625,N_16496,N_16583);
or U16626 (N_16626,N_16529,N_16441);
nor U16627 (N_16627,N_16546,N_16550);
and U16628 (N_16628,N_16426,N_16553);
and U16629 (N_16629,N_16501,N_16557);
nor U16630 (N_16630,N_16543,N_16444);
and U16631 (N_16631,N_16569,N_16559);
nand U16632 (N_16632,N_16462,N_16439);
xor U16633 (N_16633,N_16522,N_16576);
nor U16634 (N_16634,N_16561,N_16532);
and U16635 (N_16635,N_16587,N_16525);
and U16636 (N_16636,N_16438,N_16497);
xnor U16637 (N_16637,N_16411,N_16507);
and U16638 (N_16638,N_16481,N_16521);
or U16639 (N_16639,N_16555,N_16494);
nand U16640 (N_16640,N_16520,N_16568);
xor U16641 (N_16641,N_16579,N_16552);
and U16642 (N_16642,N_16596,N_16595);
or U16643 (N_16643,N_16516,N_16551);
or U16644 (N_16644,N_16514,N_16539);
or U16645 (N_16645,N_16425,N_16598);
nand U16646 (N_16646,N_16537,N_16506);
nor U16647 (N_16647,N_16478,N_16427);
or U16648 (N_16648,N_16566,N_16477);
or U16649 (N_16649,N_16563,N_16548);
nor U16650 (N_16650,N_16577,N_16533);
xnor U16651 (N_16651,N_16484,N_16414);
and U16652 (N_16652,N_16540,N_16401);
nor U16653 (N_16653,N_16509,N_16410);
nor U16654 (N_16654,N_16488,N_16556);
nand U16655 (N_16655,N_16544,N_16589);
or U16656 (N_16656,N_16472,N_16403);
nor U16657 (N_16657,N_16513,N_16422);
xor U16658 (N_16658,N_16430,N_16585);
or U16659 (N_16659,N_16416,N_16599);
nor U16660 (N_16660,N_16581,N_16510);
nor U16661 (N_16661,N_16429,N_16571);
or U16662 (N_16662,N_16454,N_16404);
and U16663 (N_16663,N_16447,N_16503);
nor U16664 (N_16664,N_16572,N_16466);
nor U16665 (N_16665,N_16519,N_16459);
nor U16666 (N_16666,N_16432,N_16531);
xor U16667 (N_16667,N_16480,N_16505);
xnor U16668 (N_16668,N_16562,N_16471);
or U16669 (N_16669,N_16420,N_16408);
nor U16670 (N_16670,N_16527,N_16588);
nand U16671 (N_16671,N_16502,N_16451);
nor U16672 (N_16672,N_16419,N_16413);
and U16673 (N_16673,N_16534,N_16486);
or U16674 (N_16674,N_16440,N_16465);
or U16675 (N_16675,N_16445,N_16593);
nand U16676 (N_16676,N_16479,N_16442);
or U16677 (N_16677,N_16464,N_16591);
and U16678 (N_16678,N_16467,N_16453);
or U16679 (N_16679,N_16535,N_16590);
or U16680 (N_16680,N_16549,N_16482);
and U16681 (N_16681,N_16565,N_16530);
nand U16682 (N_16682,N_16463,N_16424);
nor U16683 (N_16683,N_16458,N_16468);
or U16684 (N_16684,N_16491,N_16435);
and U16685 (N_16685,N_16504,N_16423);
xnor U16686 (N_16686,N_16574,N_16512);
xnor U16687 (N_16687,N_16400,N_16455);
and U16688 (N_16688,N_16560,N_16452);
nor U16689 (N_16689,N_16461,N_16517);
xor U16690 (N_16690,N_16448,N_16578);
and U16691 (N_16691,N_16515,N_16592);
nor U16692 (N_16692,N_16554,N_16567);
or U16693 (N_16693,N_16436,N_16498);
nor U16694 (N_16694,N_16456,N_16437);
or U16695 (N_16695,N_16443,N_16547);
or U16696 (N_16696,N_16495,N_16418);
nor U16697 (N_16697,N_16473,N_16490);
nand U16698 (N_16698,N_16511,N_16558);
or U16699 (N_16699,N_16476,N_16493);
nor U16700 (N_16700,N_16583,N_16403);
nand U16701 (N_16701,N_16569,N_16476);
nor U16702 (N_16702,N_16478,N_16529);
and U16703 (N_16703,N_16410,N_16578);
xor U16704 (N_16704,N_16551,N_16458);
xor U16705 (N_16705,N_16522,N_16514);
or U16706 (N_16706,N_16528,N_16504);
or U16707 (N_16707,N_16451,N_16503);
nand U16708 (N_16708,N_16408,N_16495);
nor U16709 (N_16709,N_16506,N_16523);
or U16710 (N_16710,N_16556,N_16408);
nand U16711 (N_16711,N_16414,N_16594);
or U16712 (N_16712,N_16549,N_16411);
nand U16713 (N_16713,N_16487,N_16447);
xor U16714 (N_16714,N_16518,N_16429);
or U16715 (N_16715,N_16485,N_16444);
xor U16716 (N_16716,N_16404,N_16553);
xnor U16717 (N_16717,N_16445,N_16420);
xor U16718 (N_16718,N_16587,N_16548);
xor U16719 (N_16719,N_16453,N_16512);
nand U16720 (N_16720,N_16586,N_16418);
nor U16721 (N_16721,N_16443,N_16593);
nand U16722 (N_16722,N_16481,N_16459);
nor U16723 (N_16723,N_16572,N_16548);
or U16724 (N_16724,N_16597,N_16510);
nor U16725 (N_16725,N_16456,N_16521);
or U16726 (N_16726,N_16463,N_16559);
nor U16727 (N_16727,N_16568,N_16577);
or U16728 (N_16728,N_16405,N_16485);
or U16729 (N_16729,N_16474,N_16571);
nor U16730 (N_16730,N_16522,N_16460);
nand U16731 (N_16731,N_16557,N_16462);
nor U16732 (N_16732,N_16558,N_16449);
and U16733 (N_16733,N_16579,N_16584);
or U16734 (N_16734,N_16537,N_16437);
nor U16735 (N_16735,N_16543,N_16587);
or U16736 (N_16736,N_16578,N_16479);
nor U16737 (N_16737,N_16482,N_16404);
nand U16738 (N_16738,N_16408,N_16539);
or U16739 (N_16739,N_16435,N_16504);
nor U16740 (N_16740,N_16516,N_16463);
nor U16741 (N_16741,N_16546,N_16599);
xor U16742 (N_16742,N_16591,N_16477);
and U16743 (N_16743,N_16581,N_16500);
xnor U16744 (N_16744,N_16528,N_16440);
and U16745 (N_16745,N_16582,N_16568);
nand U16746 (N_16746,N_16450,N_16520);
nand U16747 (N_16747,N_16565,N_16538);
nand U16748 (N_16748,N_16585,N_16597);
or U16749 (N_16749,N_16408,N_16452);
xor U16750 (N_16750,N_16511,N_16440);
and U16751 (N_16751,N_16562,N_16407);
nand U16752 (N_16752,N_16531,N_16459);
xnor U16753 (N_16753,N_16441,N_16416);
and U16754 (N_16754,N_16417,N_16436);
and U16755 (N_16755,N_16568,N_16534);
and U16756 (N_16756,N_16431,N_16446);
xor U16757 (N_16757,N_16418,N_16512);
nor U16758 (N_16758,N_16421,N_16422);
or U16759 (N_16759,N_16523,N_16595);
or U16760 (N_16760,N_16473,N_16407);
or U16761 (N_16761,N_16529,N_16509);
xor U16762 (N_16762,N_16516,N_16405);
nand U16763 (N_16763,N_16465,N_16586);
nor U16764 (N_16764,N_16444,N_16590);
and U16765 (N_16765,N_16445,N_16590);
nor U16766 (N_16766,N_16534,N_16591);
or U16767 (N_16767,N_16554,N_16598);
and U16768 (N_16768,N_16425,N_16427);
nor U16769 (N_16769,N_16416,N_16420);
and U16770 (N_16770,N_16459,N_16522);
and U16771 (N_16771,N_16408,N_16417);
and U16772 (N_16772,N_16453,N_16412);
xnor U16773 (N_16773,N_16560,N_16455);
or U16774 (N_16774,N_16562,N_16466);
nor U16775 (N_16775,N_16487,N_16523);
and U16776 (N_16776,N_16590,N_16586);
or U16777 (N_16777,N_16485,N_16466);
xnor U16778 (N_16778,N_16565,N_16553);
and U16779 (N_16779,N_16523,N_16413);
xnor U16780 (N_16780,N_16449,N_16468);
nand U16781 (N_16781,N_16488,N_16585);
xnor U16782 (N_16782,N_16488,N_16558);
xnor U16783 (N_16783,N_16557,N_16479);
and U16784 (N_16784,N_16520,N_16426);
and U16785 (N_16785,N_16470,N_16459);
nand U16786 (N_16786,N_16500,N_16549);
nand U16787 (N_16787,N_16436,N_16471);
and U16788 (N_16788,N_16580,N_16555);
and U16789 (N_16789,N_16537,N_16426);
nor U16790 (N_16790,N_16558,N_16422);
or U16791 (N_16791,N_16413,N_16482);
xnor U16792 (N_16792,N_16541,N_16592);
or U16793 (N_16793,N_16570,N_16463);
and U16794 (N_16794,N_16409,N_16541);
or U16795 (N_16795,N_16475,N_16444);
nor U16796 (N_16796,N_16522,N_16506);
or U16797 (N_16797,N_16458,N_16555);
nor U16798 (N_16798,N_16509,N_16523);
xor U16799 (N_16799,N_16404,N_16468);
xor U16800 (N_16800,N_16762,N_16775);
or U16801 (N_16801,N_16613,N_16768);
nor U16802 (N_16802,N_16627,N_16730);
nand U16803 (N_16803,N_16674,N_16788);
nand U16804 (N_16804,N_16625,N_16628);
and U16805 (N_16805,N_16622,N_16740);
nor U16806 (N_16806,N_16701,N_16731);
xor U16807 (N_16807,N_16721,N_16758);
nor U16808 (N_16808,N_16666,N_16634);
xnor U16809 (N_16809,N_16669,N_16741);
and U16810 (N_16810,N_16771,N_16635);
xor U16811 (N_16811,N_16732,N_16682);
or U16812 (N_16812,N_16645,N_16636);
xnor U16813 (N_16813,N_16705,N_16699);
nand U16814 (N_16814,N_16601,N_16757);
nand U16815 (N_16815,N_16617,N_16734);
nor U16816 (N_16816,N_16772,N_16716);
nand U16817 (N_16817,N_16702,N_16664);
xnor U16818 (N_16818,N_16733,N_16720);
nor U16819 (N_16819,N_16602,N_16773);
xnor U16820 (N_16820,N_16719,N_16651);
nand U16821 (N_16821,N_16735,N_16646);
nor U16822 (N_16822,N_16605,N_16755);
xor U16823 (N_16823,N_16667,N_16630);
nor U16824 (N_16824,N_16609,N_16763);
nand U16825 (N_16825,N_16767,N_16652);
and U16826 (N_16826,N_16658,N_16656);
and U16827 (N_16827,N_16789,N_16706);
and U16828 (N_16828,N_16684,N_16714);
nand U16829 (N_16829,N_16633,N_16754);
nor U16830 (N_16830,N_16765,N_16791);
nor U16831 (N_16831,N_16726,N_16737);
and U16832 (N_16832,N_16774,N_16671);
nor U16833 (N_16833,N_16744,N_16695);
or U16834 (N_16834,N_16778,N_16614);
and U16835 (N_16835,N_16603,N_16647);
or U16836 (N_16836,N_16661,N_16686);
and U16837 (N_16837,N_16712,N_16707);
and U16838 (N_16838,N_16689,N_16709);
nor U16839 (N_16839,N_16786,N_16787);
or U16840 (N_16840,N_16655,N_16711);
nand U16841 (N_16841,N_16692,N_16640);
and U16842 (N_16842,N_16698,N_16766);
and U16843 (N_16843,N_16697,N_16792);
and U16844 (N_16844,N_16660,N_16696);
nor U16845 (N_16845,N_16797,N_16639);
xor U16846 (N_16846,N_16675,N_16673);
xnor U16847 (N_16847,N_16690,N_16668);
nand U16848 (N_16848,N_16703,N_16672);
or U16849 (N_16849,N_16648,N_16747);
and U16850 (N_16850,N_16727,N_16704);
xor U16851 (N_16851,N_16677,N_16691);
nand U16852 (N_16852,N_16615,N_16620);
and U16853 (N_16853,N_16795,N_16718);
xnor U16854 (N_16854,N_16626,N_16750);
or U16855 (N_16855,N_16724,N_16618);
xor U16856 (N_16856,N_16752,N_16748);
nand U16857 (N_16857,N_16738,N_16723);
and U16858 (N_16858,N_16756,N_16659);
or U16859 (N_16859,N_16623,N_16612);
nand U16860 (N_16860,N_16610,N_16687);
or U16861 (N_16861,N_16681,N_16759);
nor U16862 (N_16862,N_16779,N_16653);
xor U16863 (N_16863,N_16708,N_16796);
nor U16864 (N_16864,N_16638,N_16688);
and U16865 (N_16865,N_16642,N_16781);
nor U16866 (N_16866,N_16693,N_16751);
and U16867 (N_16867,N_16761,N_16745);
or U16868 (N_16868,N_16629,N_16604);
nor U16869 (N_16869,N_16725,N_16785);
xnor U16870 (N_16870,N_16742,N_16619);
xnor U16871 (N_16871,N_16713,N_16784);
nand U16872 (N_16872,N_16715,N_16662);
or U16873 (N_16873,N_16600,N_16743);
or U16874 (N_16874,N_16694,N_16798);
nand U16875 (N_16875,N_16760,N_16799);
and U16876 (N_16876,N_16783,N_16670);
xor U16877 (N_16877,N_16770,N_16606);
or U16878 (N_16878,N_16632,N_16616);
or U16879 (N_16879,N_16764,N_16680);
xnor U16880 (N_16880,N_16676,N_16739);
xnor U16881 (N_16881,N_16607,N_16608);
and U16882 (N_16882,N_16722,N_16644);
xor U16883 (N_16883,N_16621,N_16685);
and U16884 (N_16884,N_16683,N_16710);
and U16885 (N_16885,N_16793,N_16657);
nand U16886 (N_16886,N_16665,N_16753);
or U16887 (N_16887,N_16631,N_16777);
nor U16888 (N_16888,N_16624,N_16679);
xor U16889 (N_16889,N_16717,N_16769);
xnor U16890 (N_16890,N_16641,N_16780);
xnor U16891 (N_16891,N_16790,N_16663);
nor U16892 (N_16892,N_16782,N_16637);
and U16893 (N_16893,N_16776,N_16700);
or U16894 (N_16894,N_16611,N_16649);
and U16895 (N_16895,N_16736,N_16650);
nor U16896 (N_16896,N_16749,N_16746);
and U16897 (N_16897,N_16729,N_16654);
xnor U16898 (N_16898,N_16728,N_16678);
and U16899 (N_16899,N_16643,N_16794);
and U16900 (N_16900,N_16696,N_16631);
xnor U16901 (N_16901,N_16650,N_16722);
or U16902 (N_16902,N_16744,N_16685);
nand U16903 (N_16903,N_16772,N_16690);
nand U16904 (N_16904,N_16635,N_16727);
and U16905 (N_16905,N_16731,N_16619);
and U16906 (N_16906,N_16629,N_16658);
xnor U16907 (N_16907,N_16797,N_16604);
or U16908 (N_16908,N_16627,N_16646);
xor U16909 (N_16909,N_16619,N_16790);
nand U16910 (N_16910,N_16720,N_16756);
nand U16911 (N_16911,N_16721,N_16657);
and U16912 (N_16912,N_16707,N_16774);
and U16913 (N_16913,N_16610,N_16674);
and U16914 (N_16914,N_16618,N_16628);
and U16915 (N_16915,N_16737,N_16700);
nor U16916 (N_16916,N_16770,N_16696);
and U16917 (N_16917,N_16787,N_16756);
or U16918 (N_16918,N_16707,N_16745);
nor U16919 (N_16919,N_16757,N_16620);
nand U16920 (N_16920,N_16684,N_16769);
xor U16921 (N_16921,N_16626,N_16621);
nor U16922 (N_16922,N_16634,N_16777);
xnor U16923 (N_16923,N_16785,N_16724);
xor U16924 (N_16924,N_16611,N_16733);
nand U16925 (N_16925,N_16751,N_16763);
and U16926 (N_16926,N_16708,N_16710);
and U16927 (N_16927,N_16663,N_16623);
nor U16928 (N_16928,N_16661,N_16605);
nand U16929 (N_16929,N_16653,N_16659);
or U16930 (N_16930,N_16675,N_16703);
nor U16931 (N_16931,N_16736,N_16653);
xnor U16932 (N_16932,N_16615,N_16679);
nand U16933 (N_16933,N_16672,N_16676);
nand U16934 (N_16934,N_16631,N_16707);
nand U16935 (N_16935,N_16609,N_16639);
nor U16936 (N_16936,N_16749,N_16701);
nand U16937 (N_16937,N_16619,N_16754);
and U16938 (N_16938,N_16602,N_16770);
and U16939 (N_16939,N_16792,N_16759);
nand U16940 (N_16940,N_16690,N_16716);
or U16941 (N_16941,N_16610,N_16702);
and U16942 (N_16942,N_16750,N_16759);
or U16943 (N_16943,N_16763,N_16685);
xor U16944 (N_16944,N_16689,N_16711);
nor U16945 (N_16945,N_16733,N_16624);
and U16946 (N_16946,N_16738,N_16774);
nor U16947 (N_16947,N_16610,N_16696);
nor U16948 (N_16948,N_16655,N_16780);
nor U16949 (N_16949,N_16759,N_16672);
nor U16950 (N_16950,N_16647,N_16626);
nor U16951 (N_16951,N_16798,N_16749);
and U16952 (N_16952,N_16605,N_16692);
nand U16953 (N_16953,N_16627,N_16615);
and U16954 (N_16954,N_16636,N_16788);
or U16955 (N_16955,N_16794,N_16696);
nand U16956 (N_16956,N_16605,N_16609);
nand U16957 (N_16957,N_16670,N_16664);
or U16958 (N_16958,N_16603,N_16684);
nor U16959 (N_16959,N_16751,N_16616);
xor U16960 (N_16960,N_16665,N_16718);
nand U16961 (N_16961,N_16786,N_16644);
nor U16962 (N_16962,N_16661,N_16647);
and U16963 (N_16963,N_16785,N_16637);
nor U16964 (N_16964,N_16743,N_16720);
nor U16965 (N_16965,N_16700,N_16690);
nand U16966 (N_16966,N_16730,N_16619);
xor U16967 (N_16967,N_16694,N_16642);
nor U16968 (N_16968,N_16735,N_16702);
nor U16969 (N_16969,N_16659,N_16610);
xor U16970 (N_16970,N_16798,N_16667);
nand U16971 (N_16971,N_16744,N_16757);
xnor U16972 (N_16972,N_16727,N_16639);
nor U16973 (N_16973,N_16768,N_16779);
nor U16974 (N_16974,N_16760,N_16622);
xor U16975 (N_16975,N_16613,N_16746);
nor U16976 (N_16976,N_16731,N_16602);
or U16977 (N_16977,N_16641,N_16684);
or U16978 (N_16978,N_16625,N_16694);
or U16979 (N_16979,N_16688,N_16643);
nand U16980 (N_16980,N_16754,N_16734);
and U16981 (N_16981,N_16781,N_16762);
nor U16982 (N_16982,N_16721,N_16735);
xnor U16983 (N_16983,N_16731,N_16605);
or U16984 (N_16984,N_16687,N_16704);
xor U16985 (N_16985,N_16635,N_16742);
xor U16986 (N_16986,N_16689,N_16698);
and U16987 (N_16987,N_16778,N_16621);
nor U16988 (N_16988,N_16677,N_16786);
or U16989 (N_16989,N_16713,N_16793);
nor U16990 (N_16990,N_16759,N_16703);
and U16991 (N_16991,N_16686,N_16651);
or U16992 (N_16992,N_16791,N_16666);
and U16993 (N_16993,N_16639,N_16776);
nor U16994 (N_16994,N_16671,N_16654);
nand U16995 (N_16995,N_16689,N_16744);
xnor U16996 (N_16996,N_16703,N_16763);
and U16997 (N_16997,N_16753,N_16685);
and U16998 (N_16998,N_16772,N_16698);
nand U16999 (N_16999,N_16662,N_16757);
nor U17000 (N_17000,N_16850,N_16859);
nand U17001 (N_17001,N_16843,N_16935);
and U17002 (N_17002,N_16846,N_16807);
and U17003 (N_17003,N_16908,N_16986);
or U17004 (N_17004,N_16802,N_16883);
and U17005 (N_17005,N_16996,N_16887);
nor U17006 (N_17006,N_16889,N_16911);
or U17007 (N_17007,N_16939,N_16963);
and U17008 (N_17008,N_16819,N_16916);
or U17009 (N_17009,N_16849,N_16810);
xnor U17010 (N_17010,N_16860,N_16993);
nand U17011 (N_17011,N_16985,N_16878);
nor U17012 (N_17012,N_16989,N_16924);
nor U17013 (N_17013,N_16998,N_16968);
or U17014 (N_17014,N_16928,N_16994);
or U17015 (N_17015,N_16904,N_16899);
nor U17016 (N_17016,N_16814,N_16995);
nor U17017 (N_17017,N_16932,N_16881);
and U17018 (N_17018,N_16971,N_16902);
nand U17019 (N_17019,N_16840,N_16870);
nand U17020 (N_17020,N_16955,N_16925);
and U17021 (N_17021,N_16943,N_16954);
or U17022 (N_17022,N_16893,N_16969);
xor U17023 (N_17023,N_16871,N_16847);
nand U17024 (N_17024,N_16833,N_16826);
nand U17025 (N_17025,N_16944,N_16997);
xor U17026 (N_17026,N_16875,N_16901);
nor U17027 (N_17027,N_16880,N_16811);
and U17028 (N_17028,N_16922,N_16805);
or U17029 (N_17029,N_16817,N_16966);
nand U17030 (N_17030,N_16895,N_16981);
and U17031 (N_17031,N_16837,N_16832);
or U17032 (N_17032,N_16909,N_16951);
xnor U17033 (N_17033,N_16841,N_16931);
nand U17034 (N_17034,N_16930,N_16947);
or U17035 (N_17035,N_16813,N_16890);
or U17036 (N_17036,N_16938,N_16824);
xor U17037 (N_17037,N_16978,N_16907);
and U17038 (N_17038,N_16949,N_16831);
xnor U17039 (N_17039,N_16933,N_16877);
nor U17040 (N_17040,N_16953,N_16958);
nand U17041 (N_17041,N_16914,N_16867);
nor U17042 (N_17042,N_16919,N_16835);
or U17043 (N_17043,N_16865,N_16823);
xor U17044 (N_17044,N_16855,N_16973);
nand U17045 (N_17045,N_16917,N_16941);
xnor U17046 (N_17046,N_16836,N_16929);
nand U17047 (N_17047,N_16977,N_16838);
nand U17048 (N_17048,N_16903,N_16915);
nand U17049 (N_17049,N_16976,N_16983);
or U17050 (N_17050,N_16913,N_16853);
or U17051 (N_17051,N_16905,N_16808);
xnor U17052 (N_17052,N_16897,N_16921);
nor U17053 (N_17053,N_16804,N_16987);
or U17054 (N_17054,N_16945,N_16991);
nor U17055 (N_17055,N_16964,N_16854);
nand U17056 (N_17056,N_16975,N_16872);
or U17057 (N_17057,N_16866,N_16864);
and U17058 (N_17058,N_16942,N_16815);
nor U17059 (N_17059,N_16959,N_16830);
xnor U17060 (N_17060,N_16923,N_16999);
nand U17061 (N_17061,N_16851,N_16876);
nor U17062 (N_17062,N_16821,N_16957);
nand U17063 (N_17063,N_16948,N_16972);
nor U17064 (N_17064,N_16898,N_16825);
nand U17065 (N_17065,N_16856,N_16884);
xnor U17066 (N_17066,N_16910,N_16937);
nand U17067 (N_17067,N_16822,N_16839);
and U17068 (N_17068,N_16888,N_16803);
or U17069 (N_17069,N_16848,N_16806);
or U17070 (N_17070,N_16800,N_16906);
xnor U17071 (N_17071,N_16979,N_16962);
nor U17072 (N_17072,N_16950,N_16845);
xor U17073 (N_17073,N_16874,N_16984);
and U17074 (N_17074,N_16974,N_16992);
or U17075 (N_17075,N_16961,N_16801);
and U17076 (N_17076,N_16862,N_16892);
and U17077 (N_17077,N_16827,N_16812);
or U17078 (N_17078,N_16828,N_16934);
nor U17079 (N_17079,N_16967,N_16912);
or U17080 (N_17080,N_16869,N_16894);
nand U17081 (N_17081,N_16927,N_16844);
or U17082 (N_17082,N_16965,N_16936);
and U17083 (N_17083,N_16858,N_16816);
or U17084 (N_17084,N_16956,N_16873);
and U17085 (N_17085,N_16863,N_16926);
xnor U17086 (N_17086,N_16852,N_16842);
or U17087 (N_17087,N_16896,N_16891);
and U17088 (N_17088,N_16868,N_16900);
or U17089 (N_17089,N_16818,N_16861);
nor U17090 (N_17090,N_16820,N_16982);
nand U17091 (N_17091,N_16879,N_16920);
nor U17092 (N_17092,N_16980,N_16809);
or U17093 (N_17093,N_16990,N_16834);
and U17094 (N_17094,N_16960,N_16946);
nor U17095 (N_17095,N_16886,N_16988);
or U17096 (N_17096,N_16857,N_16940);
nor U17097 (N_17097,N_16952,N_16885);
or U17098 (N_17098,N_16882,N_16970);
nor U17099 (N_17099,N_16918,N_16829);
nand U17100 (N_17100,N_16931,N_16811);
or U17101 (N_17101,N_16920,N_16876);
nor U17102 (N_17102,N_16994,N_16993);
nand U17103 (N_17103,N_16925,N_16967);
xnor U17104 (N_17104,N_16873,N_16983);
xnor U17105 (N_17105,N_16827,N_16962);
xnor U17106 (N_17106,N_16809,N_16945);
nand U17107 (N_17107,N_16806,N_16937);
nand U17108 (N_17108,N_16821,N_16831);
or U17109 (N_17109,N_16914,N_16964);
xor U17110 (N_17110,N_16882,N_16851);
nor U17111 (N_17111,N_16825,N_16951);
nor U17112 (N_17112,N_16825,N_16900);
or U17113 (N_17113,N_16874,N_16914);
nand U17114 (N_17114,N_16970,N_16931);
and U17115 (N_17115,N_16908,N_16948);
and U17116 (N_17116,N_16887,N_16930);
nor U17117 (N_17117,N_16885,N_16968);
xor U17118 (N_17118,N_16831,N_16902);
or U17119 (N_17119,N_16932,N_16927);
or U17120 (N_17120,N_16935,N_16873);
nand U17121 (N_17121,N_16933,N_16952);
and U17122 (N_17122,N_16991,N_16935);
and U17123 (N_17123,N_16893,N_16927);
xor U17124 (N_17124,N_16915,N_16892);
or U17125 (N_17125,N_16851,N_16814);
nand U17126 (N_17126,N_16893,N_16860);
nand U17127 (N_17127,N_16830,N_16891);
xor U17128 (N_17128,N_16928,N_16931);
nor U17129 (N_17129,N_16926,N_16909);
xor U17130 (N_17130,N_16846,N_16872);
xnor U17131 (N_17131,N_16968,N_16811);
nor U17132 (N_17132,N_16969,N_16915);
nor U17133 (N_17133,N_16972,N_16857);
nor U17134 (N_17134,N_16872,N_16980);
nand U17135 (N_17135,N_16967,N_16985);
and U17136 (N_17136,N_16852,N_16883);
nand U17137 (N_17137,N_16968,N_16881);
and U17138 (N_17138,N_16894,N_16933);
nor U17139 (N_17139,N_16845,N_16941);
and U17140 (N_17140,N_16979,N_16951);
nor U17141 (N_17141,N_16969,N_16979);
nand U17142 (N_17142,N_16811,N_16903);
or U17143 (N_17143,N_16816,N_16897);
xor U17144 (N_17144,N_16867,N_16988);
xnor U17145 (N_17145,N_16995,N_16957);
and U17146 (N_17146,N_16880,N_16928);
and U17147 (N_17147,N_16978,N_16888);
xnor U17148 (N_17148,N_16874,N_16960);
and U17149 (N_17149,N_16810,N_16830);
nor U17150 (N_17150,N_16972,N_16894);
xor U17151 (N_17151,N_16831,N_16964);
nor U17152 (N_17152,N_16837,N_16895);
and U17153 (N_17153,N_16868,N_16978);
or U17154 (N_17154,N_16851,N_16917);
nand U17155 (N_17155,N_16963,N_16946);
nor U17156 (N_17156,N_16943,N_16846);
nand U17157 (N_17157,N_16863,N_16873);
or U17158 (N_17158,N_16945,N_16994);
xnor U17159 (N_17159,N_16867,N_16816);
nor U17160 (N_17160,N_16932,N_16896);
and U17161 (N_17161,N_16953,N_16851);
nand U17162 (N_17162,N_16996,N_16878);
and U17163 (N_17163,N_16982,N_16882);
nor U17164 (N_17164,N_16801,N_16898);
xor U17165 (N_17165,N_16880,N_16904);
xor U17166 (N_17166,N_16881,N_16991);
nor U17167 (N_17167,N_16849,N_16920);
nand U17168 (N_17168,N_16922,N_16919);
or U17169 (N_17169,N_16968,N_16908);
and U17170 (N_17170,N_16897,N_16859);
and U17171 (N_17171,N_16995,N_16952);
nand U17172 (N_17172,N_16853,N_16928);
or U17173 (N_17173,N_16942,N_16810);
xor U17174 (N_17174,N_16988,N_16924);
nand U17175 (N_17175,N_16850,N_16822);
and U17176 (N_17176,N_16848,N_16978);
nand U17177 (N_17177,N_16806,N_16952);
nand U17178 (N_17178,N_16978,N_16972);
nand U17179 (N_17179,N_16927,N_16981);
or U17180 (N_17180,N_16966,N_16997);
or U17181 (N_17181,N_16845,N_16898);
nor U17182 (N_17182,N_16919,N_16904);
nand U17183 (N_17183,N_16823,N_16807);
and U17184 (N_17184,N_16958,N_16835);
nor U17185 (N_17185,N_16848,N_16856);
xor U17186 (N_17186,N_16809,N_16958);
and U17187 (N_17187,N_16945,N_16839);
and U17188 (N_17188,N_16966,N_16869);
or U17189 (N_17189,N_16871,N_16980);
nand U17190 (N_17190,N_16989,N_16800);
nand U17191 (N_17191,N_16811,N_16836);
or U17192 (N_17192,N_16888,N_16872);
and U17193 (N_17193,N_16964,N_16878);
nand U17194 (N_17194,N_16809,N_16814);
nand U17195 (N_17195,N_16918,N_16991);
nor U17196 (N_17196,N_16829,N_16878);
xnor U17197 (N_17197,N_16854,N_16956);
and U17198 (N_17198,N_16871,N_16948);
nor U17199 (N_17199,N_16928,N_16989);
nor U17200 (N_17200,N_17129,N_17168);
nand U17201 (N_17201,N_17199,N_17066);
nor U17202 (N_17202,N_17015,N_17026);
xnor U17203 (N_17203,N_17115,N_17173);
xnor U17204 (N_17204,N_17031,N_17106);
and U17205 (N_17205,N_17036,N_17161);
nor U17206 (N_17206,N_17060,N_17035);
nand U17207 (N_17207,N_17050,N_17042);
or U17208 (N_17208,N_17192,N_17084);
and U17209 (N_17209,N_17113,N_17059);
and U17210 (N_17210,N_17073,N_17108);
xor U17211 (N_17211,N_17017,N_17072);
or U17212 (N_17212,N_17146,N_17148);
nand U17213 (N_17213,N_17170,N_17166);
nand U17214 (N_17214,N_17003,N_17088);
or U17215 (N_17215,N_17077,N_17016);
nand U17216 (N_17216,N_17132,N_17184);
and U17217 (N_17217,N_17189,N_17163);
and U17218 (N_17218,N_17012,N_17071);
nor U17219 (N_17219,N_17019,N_17171);
or U17220 (N_17220,N_17116,N_17196);
xor U17221 (N_17221,N_17020,N_17049);
and U17222 (N_17222,N_17011,N_17058);
xor U17223 (N_17223,N_17118,N_17028);
nor U17224 (N_17224,N_17109,N_17096);
xor U17225 (N_17225,N_17025,N_17154);
nor U17226 (N_17226,N_17069,N_17091);
xnor U17227 (N_17227,N_17177,N_17053);
xnor U17228 (N_17228,N_17052,N_17085);
or U17229 (N_17229,N_17006,N_17158);
xor U17230 (N_17230,N_17137,N_17029);
and U17231 (N_17231,N_17014,N_17070);
xor U17232 (N_17232,N_17141,N_17005);
nor U17233 (N_17233,N_17187,N_17023);
and U17234 (N_17234,N_17067,N_17044);
or U17235 (N_17235,N_17027,N_17061);
nand U17236 (N_17236,N_17092,N_17099);
nor U17237 (N_17237,N_17120,N_17155);
or U17238 (N_17238,N_17140,N_17034);
nand U17239 (N_17239,N_17068,N_17082);
xor U17240 (N_17240,N_17039,N_17138);
or U17241 (N_17241,N_17119,N_17183);
xnor U17242 (N_17242,N_17062,N_17030);
nor U17243 (N_17243,N_17051,N_17133);
xor U17244 (N_17244,N_17008,N_17101);
and U17245 (N_17245,N_17000,N_17122);
nor U17246 (N_17246,N_17024,N_17167);
nor U17247 (N_17247,N_17086,N_17046);
or U17248 (N_17248,N_17124,N_17157);
or U17249 (N_17249,N_17093,N_17047);
xor U17250 (N_17250,N_17130,N_17131);
nor U17251 (N_17251,N_17064,N_17078);
nand U17252 (N_17252,N_17004,N_17107);
or U17253 (N_17253,N_17089,N_17010);
nand U17254 (N_17254,N_17013,N_17112);
nor U17255 (N_17255,N_17079,N_17048);
or U17256 (N_17256,N_17094,N_17156);
nand U17257 (N_17257,N_17123,N_17063);
and U17258 (N_17258,N_17038,N_17074);
and U17259 (N_17259,N_17145,N_17181);
or U17260 (N_17260,N_17143,N_17095);
nand U17261 (N_17261,N_17134,N_17054);
and U17262 (N_17262,N_17194,N_17190);
or U17263 (N_17263,N_17188,N_17022);
nand U17264 (N_17264,N_17105,N_17041);
nand U17265 (N_17265,N_17114,N_17126);
nor U17266 (N_17266,N_17197,N_17033);
and U17267 (N_17267,N_17135,N_17102);
nand U17268 (N_17268,N_17136,N_17178);
nand U17269 (N_17269,N_17037,N_17198);
and U17270 (N_17270,N_17065,N_17144);
or U17271 (N_17271,N_17193,N_17172);
or U17272 (N_17272,N_17175,N_17056);
nor U17273 (N_17273,N_17075,N_17174);
nor U17274 (N_17274,N_17152,N_17142);
and U17275 (N_17275,N_17043,N_17100);
nand U17276 (N_17276,N_17040,N_17195);
nand U17277 (N_17277,N_17180,N_17128);
and U17278 (N_17278,N_17147,N_17164);
or U17279 (N_17279,N_17057,N_17179);
or U17280 (N_17280,N_17018,N_17159);
or U17281 (N_17281,N_17001,N_17186);
xnor U17282 (N_17282,N_17007,N_17176);
and U17283 (N_17283,N_17150,N_17160);
and U17284 (N_17284,N_17090,N_17104);
or U17285 (N_17285,N_17045,N_17165);
xor U17286 (N_17286,N_17103,N_17087);
xnor U17287 (N_17287,N_17185,N_17153);
nand U17288 (N_17288,N_17162,N_17009);
nor U17289 (N_17289,N_17169,N_17125);
or U17290 (N_17290,N_17139,N_17083);
or U17291 (N_17291,N_17117,N_17080);
nand U17292 (N_17292,N_17127,N_17121);
xnor U17293 (N_17293,N_17002,N_17021);
nor U17294 (N_17294,N_17098,N_17110);
nand U17295 (N_17295,N_17182,N_17076);
xor U17296 (N_17296,N_17097,N_17081);
and U17297 (N_17297,N_17149,N_17111);
xor U17298 (N_17298,N_17151,N_17191);
or U17299 (N_17299,N_17032,N_17055);
nand U17300 (N_17300,N_17131,N_17141);
nand U17301 (N_17301,N_17100,N_17179);
nand U17302 (N_17302,N_17144,N_17083);
nand U17303 (N_17303,N_17142,N_17008);
xor U17304 (N_17304,N_17087,N_17134);
and U17305 (N_17305,N_17015,N_17159);
nand U17306 (N_17306,N_17041,N_17054);
xnor U17307 (N_17307,N_17012,N_17151);
and U17308 (N_17308,N_17043,N_17120);
or U17309 (N_17309,N_17117,N_17010);
nand U17310 (N_17310,N_17140,N_17152);
nor U17311 (N_17311,N_17031,N_17078);
xor U17312 (N_17312,N_17168,N_17053);
nand U17313 (N_17313,N_17016,N_17177);
or U17314 (N_17314,N_17127,N_17187);
nor U17315 (N_17315,N_17199,N_17064);
or U17316 (N_17316,N_17073,N_17043);
nor U17317 (N_17317,N_17175,N_17159);
and U17318 (N_17318,N_17006,N_17033);
and U17319 (N_17319,N_17069,N_17011);
xor U17320 (N_17320,N_17098,N_17136);
nand U17321 (N_17321,N_17132,N_17180);
nor U17322 (N_17322,N_17120,N_17111);
xor U17323 (N_17323,N_17005,N_17178);
xnor U17324 (N_17324,N_17103,N_17162);
nand U17325 (N_17325,N_17178,N_17184);
and U17326 (N_17326,N_17014,N_17111);
and U17327 (N_17327,N_17006,N_17114);
or U17328 (N_17328,N_17177,N_17045);
xor U17329 (N_17329,N_17073,N_17175);
xor U17330 (N_17330,N_17074,N_17109);
or U17331 (N_17331,N_17112,N_17071);
nand U17332 (N_17332,N_17045,N_17159);
and U17333 (N_17333,N_17074,N_17062);
nor U17334 (N_17334,N_17118,N_17058);
or U17335 (N_17335,N_17193,N_17079);
and U17336 (N_17336,N_17088,N_17014);
and U17337 (N_17337,N_17175,N_17082);
and U17338 (N_17338,N_17091,N_17074);
and U17339 (N_17339,N_17182,N_17153);
xnor U17340 (N_17340,N_17108,N_17155);
nor U17341 (N_17341,N_17178,N_17098);
and U17342 (N_17342,N_17134,N_17121);
nor U17343 (N_17343,N_17157,N_17012);
nor U17344 (N_17344,N_17104,N_17071);
nor U17345 (N_17345,N_17171,N_17070);
or U17346 (N_17346,N_17041,N_17023);
nor U17347 (N_17347,N_17097,N_17126);
nand U17348 (N_17348,N_17137,N_17044);
nor U17349 (N_17349,N_17009,N_17108);
nor U17350 (N_17350,N_17039,N_17052);
xnor U17351 (N_17351,N_17155,N_17119);
nand U17352 (N_17352,N_17036,N_17060);
nor U17353 (N_17353,N_17183,N_17012);
xor U17354 (N_17354,N_17186,N_17109);
nand U17355 (N_17355,N_17188,N_17025);
nand U17356 (N_17356,N_17147,N_17155);
xnor U17357 (N_17357,N_17074,N_17067);
or U17358 (N_17358,N_17199,N_17164);
or U17359 (N_17359,N_17148,N_17162);
xor U17360 (N_17360,N_17165,N_17025);
or U17361 (N_17361,N_17031,N_17153);
and U17362 (N_17362,N_17092,N_17189);
and U17363 (N_17363,N_17183,N_17095);
and U17364 (N_17364,N_17016,N_17009);
and U17365 (N_17365,N_17025,N_17183);
nor U17366 (N_17366,N_17187,N_17008);
nor U17367 (N_17367,N_17151,N_17179);
or U17368 (N_17368,N_17130,N_17010);
xor U17369 (N_17369,N_17163,N_17092);
or U17370 (N_17370,N_17165,N_17162);
nand U17371 (N_17371,N_17151,N_17125);
nor U17372 (N_17372,N_17008,N_17136);
nand U17373 (N_17373,N_17036,N_17054);
nor U17374 (N_17374,N_17067,N_17057);
xor U17375 (N_17375,N_17004,N_17125);
xor U17376 (N_17376,N_17103,N_17128);
or U17377 (N_17377,N_17006,N_17062);
xnor U17378 (N_17378,N_17144,N_17120);
and U17379 (N_17379,N_17079,N_17138);
nor U17380 (N_17380,N_17153,N_17137);
or U17381 (N_17381,N_17149,N_17070);
and U17382 (N_17382,N_17174,N_17000);
or U17383 (N_17383,N_17185,N_17031);
nor U17384 (N_17384,N_17103,N_17176);
or U17385 (N_17385,N_17043,N_17055);
xor U17386 (N_17386,N_17176,N_17080);
xnor U17387 (N_17387,N_17182,N_17197);
xor U17388 (N_17388,N_17161,N_17085);
nor U17389 (N_17389,N_17043,N_17149);
or U17390 (N_17390,N_17002,N_17058);
nand U17391 (N_17391,N_17059,N_17094);
and U17392 (N_17392,N_17080,N_17002);
nand U17393 (N_17393,N_17153,N_17134);
or U17394 (N_17394,N_17031,N_17032);
or U17395 (N_17395,N_17181,N_17194);
nor U17396 (N_17396,N_17108,N_17046);
nand U17397 (N_17397,N_17167,N_17175);
and U17398 (N_17398,N_17064,N_17138);
xnor U17399 (N_17399,N_17109,N_17108);
and U17400 (N_17400,N_17232,N_17315);
xor U17401 (N_17401,N_17359,N_17291);
xor U17402 (N_17402,N_17231,N_17348);
or U17403 (N_17403,N_17225,N_17327);
xor U17404 (N_17404,N_17385,N_17204);
or U17405 (N_17405,N_17271,N_17278);
nand U17406 (N_17406,N_17210,N_17398);
or U17407 (N_17407,N_17281,N_17230);
and U17408 (N_17408,N_17279,N_17286);
or U17409 (N_17409,N_17370,N_17219);
or U17410 (N_17410,N_17202,N_17255);
nand U17411 (N_17411,N_17346,N_17357);
xnor U17412 (N_17412,N_17273,N_17206);
and U17413 (N_17413,N_17361,N_17350);
nor U17414 (N_17414,N_17274,N_17209);
or U17415 (N_17415,N_17257,N_17395);
and U17416 (N_17416,N_17383,N_17250);
nand U17417 (N_17417,N_17310,N_17277);
and U17418 (N_17418,N_17246,N_17358);
nor U17419 (N_17419,N_17259,N_17311);
nand U17420 (N_17420,N_17308,N_17290);
and U17421 (N_17421,N_17388,N_17347);
or U17422 (N_17422,N_17365,N_17295);
nand U17423 (N_17423,N_17276,N_17377);
nand U17424 (N_17424,N_17317,N_17294);
and U17425 (N_17425,N_17356,N_17390);
nand U17426 (N_17426,N_17318,N_17305);
nor U17427 (N_17427,N_17260,N_17287);
nand U17428 (N_17428,N_17392,N_17234);
xor U17429 (N_17429,N_17387,N_17298);
nand U17430 (N_17430,N_17341,N_17328);
nor U17431 (N_17431,N_17284,N_17227);
xnor U17432 (N_17432,N_17268,N_17380);
and U17433 (N_17433,N_17244,N_17337);
or U17434 (N_17434,N_17282,N_17252);
nand U17435 (N_17435,N_17253,N_17334);
nand U17436 (N_17436,N_17243,N_17391);
and U17437 (N_17437,N_17366,N_17293);
or U17438 (N_17438,N_17256,N_17314);
nor U17439 (N_17439,N_17263,N_17235);
nor U17440 (N_17440,N_17303,N_17323);
xor U17441 (N_17441,N_17301,N_17381);
and U17442 (N_17442,N_17296,N_17267);
nand U17443 (N_17443,N_17242,N_17349);
nor U17444 (N_17444,N_17247,N_17221);
or U17445 (N_17445,N_17211,N_17362);
and U17446 (N_17446,N_17322,N_17332);
nor U17447 (N_17447,N_17228,N_17382);
or U17448 (N_17448,N_17236,N_17354);
nor U17449 (N_17449,N_17223,N_17352);
xnor U17450 (N_17450,N_17212,N_17321);
nor U17451 (N_17451,N_17229,N_17275);
nor U17452 (N_17452,N_17272,N_17369);
or U17453 (N_17453,N_17238,N_17222);
nand U17454 (N_17454,N_17262,N_17335);
xor U17455 (N_17455,N_17344,N_17304);
nand U17456 (N_17456,N_17205,N_17351);
and U17457 (N_17457,N_17367,N_17285);
nand U17458 (N_17458,N_17331,N_17336);
or U17459 (N_17459,N_17389,N_17313);
and U17460 (N_17460,N_17378,N_17340);
and U17461 (N_17461,N_17316,N_17309);
xnor U17462 (N_17462,N_17394,N_17326);
nand U17463 (N_17463,N_17375,N_17333);
nor U17464 (N_17464,N_17224,N_17374);
nor U17465 (N_17465,N_17249,N_17306);
nand U17466 (N_17466,N_17266,N_17208);
xnor U17467 (N_17467,N_17393,N_17218);
and U17468 (N_17468,N_17292,N_17363);
xor U17469 (N_17469,N_17338,N_17345);
or U17470 (N_17470,N_17289,N_17207);
and U17471 (N_17471,N_17233,N_17280);
or U17472 (N_17472,N_17376,N_17270);
nand U17473 (N_17473,N_17353,N_17254);
nor U17474 (N_17474,N_17258,N_17386);
or U17475 (N_17475,N_17217,N_17241);
or U17476 (N_17476,N_17300,N_17342);
and U17477 (N_17477,N_17261,N_17302);
xor U17478 (N_17478,N_17215,N_17372);
or U17479 (N_17479,N_17203,N_17355);
nand U17480 (N_17480,N_17319,N_17297);
xor U17481 (N_17481,N_17283,N_17245);
nor U17482 (N_17482,N_17373,N_17397);
nor U17483 (N_17483,N_17360,N_17320);
nor U17484 (N_17484,N_17213,N_17329);
xor U17485 (N_17485,N_17307,N_17201);
and U17486 (N_17486,N_17214,N_17339);
nor U17487 (N_17487,N_17216,N_17237);
xor U17488 (N_17488,N_17240,N_17399);
or U17489 (N_17489,N_17269,N_17368);
nor U17490 (N_17490,N_17396,N_17379);
nor U17491 (N_17491,N_17288,N_17371);
xor U17492 (N_17492,N_17248,N_17239);
or U17493 (N_17493,N_17265,N_17251);
or U17494 (N_17494,N_17312,N_17226);
and U17495 (N_17495,N_17264,N_17220);
or U17496 (N_17496,N_17299,N_17330);
nand U17497 (N_17497,N_17343,N_17384);
nor U17498 (N_17498,N_17200,N_17325);
nor U17499 (N_17499,N_17324,N_17364);
nor U17500 (N_17500,N_17250,N_17268);
xnor U17501 (N_17501,N_17378,N_17244);
or U17502 (N_17502,N_17389,N_17363);
or U17503 (N_17503,N_17397,N_17398);
and U17504 (N_17504,N_17305,N_17366);
or U17505 (N_17505,N_17290,N_17280);
xor U17506 (N_17506,N_17389,N_17255);
nor U17507 (N_17507,N_17331,N_17382);
nor U17508 (N_17508,N_17257,N_17272);
or U17509 (N_17509,N_17347,N_17248);
nor U17510 (N_17510,N_17333,N_17221);
nand U17511 (N_17511,N_17348,N_17331);
or U17512 (N_17512,N_17231,N_17221);
nand U17513 (N_17513,N_17220,N_17393);
or U17514 (N_17514,N_17376,N_17304);
xnor U17515 (N_17515,N_17227,N_17307);
nand U17516 (N_17516,N_17336,N_17373);
nor U17517 (N_17517,N_17367,N_17236);
and U17518 (N_17518,N_17278,N_17222);
nor U17519 (N_17519,N_17237,N_17368);
and U17520 (N_17520,N_17394,N_17312);
and U17521 (N_17521,N_17267,N_17355);
nor U17522 (N_17522,N_17371,N_17246);
nand U17523 (N_17523,N_17287,N_17264);
xor U17524 (N_17524,N_17284,N_17251);
and U17525 (N_17525,N_17328,N_17205);
xnor U17526 (N_17526,N_17244,N_17267);
and U17527 (N_17527,N_17323,N_17202);
or U17528 (N_17528,N_17273,N_17241);
xor U17529 (N_17529,N_17228,N_17230);
and U17530 (N_17530,N_17366,N_17303);
and U17531 (N_17531,N_17226,N_17272);
or U17532 (N_17532,N_17387,N_17299);
and U17533 (N_17533,N_17315,N_17276);
nor U17534 (N_17534,N_17289,N_17249);
xor U17535 (N_17535,N_17316,N_17273);
nor U17536 (N_17536,N_17291,N_17312);
and U17537 (N_17537,N_17318,N_17395);
nand U17538 (N_17538,N_17383,N_17240);
and U17539 (N_17539,N_17235,N_17244);
nand U17540 (N_17540,N_17317,N_17214);
xnor U17541 (N_17541,N_17333,N_17289);
xor U17542 (N_17542,N_17259,N_17312);
xnor U17543 (N_17543,N_17306,N_17341);
or U17544 (N_17544,N_17261,N_17288);
or U17545 (N_17545,N_17347,N_17344);
xnor U17546 (N_17546,N_17215,N_17294);
and U17547 (N_17547,N_17261,N_17294);
or U17548 (N_17548,N_17314,N_17253);
or U17549 (N_17549,N_17368,N_17242);
and U17550 (N_17550,N_17391,N_17255);
nand U17551 (N_17551,N_17276,N_17386);
or U17552 (N_17552,N_17355,N_17279);
xnor U17553 (N_17553,N_17353,N_17264);
nand U17554 (N_17554,N_17216,N_17202);
nor U17555 (N_17555,N_17236,N_17366);
or U17556 (N_17556,N_17357,N_17340);
and U17557 (N_17557,N_17331,N_17380);
xnor U17558 (N_17558,N_17298,N_17222);
nor U17559 (N_17559,N_17285,N_17222);
xnor U17560 (N_17560,N_17368,N_17224);
nand U17561 (N_17561,N_17285,N_17246);
and U17562 (N_17562,N_17334,N_17369);
and U17563 (N_17563,N_17382,N_17348);
or U17564 (N_17564,N_17245,N_17214);
xnor U17565 (N_17565,N_17231,N_17351);
xnor U17566 (N_17566,N_17263,N_17392);
xnor U17567 (N_17567,N_17202,N_17389);
nand U17568 (N_17568,N_17280,N_17326);
xnor U17569 (N_17569,N_17324,N_17331);
and U17570 (N_17570,N_17203,N_17383);
nand U17571 (N_17571,N_17346,N_17265);
or U17572 (N_17572,N_17396,N_17200);
nor U17573 (N_17573,N_17335,N_17350);
nand U17574 (N_17574,N_17383,N_17362);
xor U17575 (N_17575,N_17250,N_17210);
xnor U17576 (N_17576,N_17391,N_17315);
nand U17577 (N_17577,N_17286,N_17397);
nor U17578 (N_17578,N_17386,N_17266);
nand U17579 (N_17579,N_17339,N_17259);
nand U17580 (N_17580,N_17309,N_17210);
xor U17581 (N_17581,N_17378,N_17341);
nor U17582 (N_17582,N_17205,N_17235);
xor U17583 (N_17583,N_17292,N_17215);
or U17584 (N_17584,N_17282,N_17205);
or U17585 (N_17585,N_17201,N_17315);
nor U17586 (N_17586,N_17272,N_17388);
nand U17587 (N_17587,N_17394,N_17357);
xor U17588 (N_17588,N_17384,N_17322);
xnor U17589 (N_17589,N_17338,N_17253);
and U17590 (N_17590,N_17367,N_17214);
nand U17591 (N_17591,N_17246,N_17303);
or U17592 (N_17592,N_17391,N_17378);
and U17593 (N_17593,N_17229,N_17321);
or U17594 (N_17594,N_17211,N_17240);
and U17595 (N_17595,N_17245,N_17345);
xnor U17596 (N_17596,N_17334,N_17345);
and U17597 (N_17597,N_17370,N_17354);
nor U17598 (N_17598,N_17266,N_17290);
or U17599 (N_17599,N_17253,N_17374);
xnor U17600 (N_17600,N_17432,N_17564);
nand U17601 (N_17601,N_17510,N_17473);
nor U17602 (N_17602,N_17552,N_17595);
and U17603 (N_17603,N_17433,N_17486);
nand U17604 (N_17604,N_17539,N_17435);
nand U17605 (N_17605,N_17573,N_17576);
and U17606 (N_17606,N_17481,N_17519);
nor U17607 (N_17607,N_17494,N_17518);
nand U17608 (N_17608,N_17590,N_17580);
and U17609 (N_17609,N_17463,N_17467);
nand U17610 (N_17610,N_17440,N_17599);
nand U17611 (N_17611,N_17410,N_17415);
or U17612 (N_17612,N_17511,N_17500);
or U17613 (N_17613,N_17563,N_17548);
nand U17614 (N_17614,N_17516,N_17547);
nor U17615 (N_17615,N_17584,N_17478);
nor U17616 (N_17616,N_17567,N_17487);
xor U17617 (N_17617,N_17549,N_17420);
and U17618 (N_17618,N_17565,N_17581);
and U17619 (N_17619,N_17587,N_17468);
nor U17620 (N_17620,N_17483,N_17508);
or U17621 (N_17621,N_17528,N_17401);
xnor U17622 (N_17622,N_17459,N_17489);
nor U17623 (N_17623,N_17436,N_17570);
and U17624 (N_17624,N_17534,N_17502);
and U17625 (N_17625,N_17521,N_17480);
xnor U17626 (N_17626,N_17556,N_17588);
nor U17627 (N_17627,N_17495,N_17560);
or U17628 (N_17628,N_17562,N_17477);
xnor U17629 (N_17629,N_17566,N_17474);
nand U17630 (N_17630,N_17558,N_17479);
nand U17631 (N_17631,N_17499,N_17428);
nand U17632 (N_17632,N_17520,N_17491);
or U17633 (N_17633,N_17464,N_17461);
nand U17634 (N_17634,N_17405,N_17404);
xor U17635 (N_17635,N_17542,N_17422);
or U17636 (N_17636,N_17561,N_17450);
or U17637 (N_17637,N_17575,N_17466);
or U17638 (N_17638,N_17523,N_17598);
nand U17639 (N_17639,N_17439,N_17460);
xnor U17640 (N_17640,N_17557,N_17417);
nand U17641 (N_17641,N_17543,N_17579);
nand U17642 (N_17642,N_17476,N_17462);
xnor U17643 (N_17643,N_17513,N_17569);
nand U17644 (N_17644,N_17424,N_17515);
or U17645 (N_17645,N_17475,N_17472);
nor U17646 (N_17646,N_17501,N_17445);
xnor U17647 (N_17647,N_17470,N_17414);
nand U17648 (N_17648,N_17426,N_17506);
and U17649 (N_17649,N_17592,N_17488);
and U17650 (N_17650,N_17525,N_17536);
nand U17651 (N_17651,N_17541,N_17507);
and U17652 (N_17652,N_17555,N_17532);
and U17653 (N_17653,N_17568,N_17582);
or U17654 (N_17654,N_17514,N_17545);
nor U17655 (N_17655,N_17448,N_17456);
xor U17656 (N_17656,N_17431,N_17438);
and U17657 (N_17657,N_17484,N_17416);
and U17658 (N_17658,N_17411,N_17526);
nand U17659 (N_17659,N_17441,N_17423);
nor U17660 (N_17660,N_17497,N_17589);
xnor U17661 (N_17661,N_17453,N_17504);
nand U17662 (N_17662,N_17442,N_17402);
and U17663 (N_17663,N_17454,N_17452);
nand U17664 (N_17664,N_17427,N_17577);
nor U17665 (N_17665,N_17586,N_17457);
and U17666 (N_17666,N_17498,N_17493);
nor U17667 (N_17667,N_17597,N_17583);
nor U17668 (N_17668,N_17403,N_17413);
nand U17669 (N_17669,N_17572,N_17585);
xnor U17670 (N_17670,N_17443,N_17496);
xnor U17671 (N_17671,N_17553,N_17544);
nand U17672 (N_17672,N_17429,N_17458);
and U17673 (N_17673,N_17409,N_17425);
xnor U17674 (N_17674,N_17451,N_17512);
or U17675 (N_17675,N_17527,N_17482);
and U17676 (N_17676,N_17593,N_17400);
and U17677 (N_17677,N_17522,N_17537);
xor U17678 (N_17678,N_17492,N_17591);
or U17679 (N_17679,N_17419,N_17550);
or U17680 (N_17680,N_17469,N_17449);
xnor U17681 (N_17681,N_17533,N_17418);
xor U17682 (N_17682,N_17406,N_17465);
or U17683 (N_17683,N_17434,N_17531);
nor U17684 (N_17684,N_17509,N_17596);
or U17685 (N_17685,N_17407,N_17578);
or U17686 (N_17686,N_17412,N_17490);
and U17687 (N_17687,N_17455,N_17571);
and U17688 (N_17688,N_17444,N_17485);
nand U17689 (N_17689,N_17530,N_17503);
and U17690 (N_17690,N_17430,N_17554);
nor U17691 (N_17691,N_17551,N_17437);
or U17692 (N_17692,N_17446,N_17574);
nand U17693 (N_17693,N_17505,N_17529);
nand U17694 (N_17694,N_17524,N_17594);
nor U17695 (N_17695,N_17447,N_17421);
and U17696 (N_17696,N_17471,N_17540);
nand U17697 (N_17697,N_17546,N_17538);
xnor U17698 (N_17698,N_17559,N_17517);
nand U17699 (N_17699,N_17535,N_17408);
nor U17700 (N_17700,N_17577,N_17523);
and U17701 (N_17701,N_17420,N_17482);
nor U17702 (N_17702,N_17548,N_17585);
xor U17703 (N_17703,N_17452,N_17536);
nor U17704 (N_17704,N_17510,N_17420);
nand U17705 (N_17705,N_17447,N_17516);
and U17706 (N_17706,N_17502,N_17587);
and U17707 (N_17707,N_17463,N_17435);
nor U17708 (N_17708,N_17507,N_17447);
nand U17709 (N_17709,N_17507,N_17448);
and U17710 (N_17710,N_17456,N_17452);
and U17711 (N_17711,N_17507,N_17410);
nand U17712 (N_17712,N_17582,N_17579);
and U17713 (N_17713,N_17585,N_17463);
xor U17714 (N_17714,N_17569,N_17576);
nor U17715 (N_17715,N_17567,N_17587);
nor U17716 (N_17716,N_17531,N_17574);
or U17717 (N_17717,N_17583,N_17425);
xnor U17718 (N_17718,N_17530,N_17558);
or U17719 (N_17719,N_17492,N_17539);
nor U17720 (N_17720,N_17567,N_17446);
or U17721 (N_17721,N_17501,N_17584);
nand U17722 (N_17722,N_17517,N_17589);
nor U17723 (N_17723,N_17522,N_17441);
or U17724 (N_17724,N_17587,N_17431);
and U17725 (N_17725,N_17437,N_17524);
or U17726 (N_17726,N_17582,N_17445);
nand U17727 (N_17727,N_17576,N_17501);
and U17728 (N_17728,N_17438,N_17527);
xnor U17729 (N_17729,N_17460,N_17501);
nand U17730 (N_17730,N_17547,N_17529);
nor U17731 (N_17731,N_17566,N_17406);
nand U17732 (N_17732,N_17463,N_17419);
and U17733 (N_17733,N_17489,N_17431);
nor U17734 (N_17734,N_17478,N_17443);
xor U17735 (N_17735,N_17508,N_17493);
and U17736 (N_17736,N_17401,N_17456);
and U17737 (N_17737,N_17516,N_17591);
nor U17738 (N_17738,N_17505,N_17517);
or U17739 (N_17739,N_17402,N_17589);
nor U17740 (N_17740,N_17598,N_17552);
nor U17741 (N_17741,N_17461,N_17518);
and U17742 (N_17742,N_17504,N_17480);
and U17743 (N_17743,N_17402,N_17445);
nor U17744 (N_17744,N_17439,N_17569);
nand U17745 (N_17745,N_17502,N_17514);
and U17746 (N_17746,N_17409,N_17416);
nor U17747 (N_17747,N_17441,N_17420);
nor U17748 (N_17748,N_17595,N_17525);
nor U17749 (N_17749,N_17407,N_17445);
or U17750 (N_17750,N_17440,N_17575);
and U17751 (N_17751,N_17480,N_17401);
and U17752 (N_17752,N_17475,N_17422);
or U17753 (N_17753,N_17563,N_17473);
and U17754 (N_17754,N_17413,N_17471);
nand U17755 (N_17755,N_17565,N_17443);
or U17756 (N_17756,N_17441,N_17551);
and U17757 (N_17757,N_17570,N_17534);
or U17758 (N_17758,N_17581,N_17458);
nor U17759 (N_17759,N_17438,N_17547);
or U17760 (N_17760,N_17478,N_17507);
nor U17761 (N_17761,N_17563,N_17419);
and U17762 (N_17762,N_17539,N_17574);
nor U17763 (N_17763,N_17504,N_17582);
nand U17764 (N_17764,N_17490,N_17445);
or U17765 (N_17765,N_17487,N_17437);
xnor U17766 (N_17766,N_17470,N_17531);
or U17767 (N_17767,N_17421,N_17598);
xnor U17768 (N_17768,N_17538,N_17593);
nand U17769 (N_17769,N_17512,N_17563);
xor U17770 (N_17770,N_17588,N_17413);
or U17771 (N_17771,N_17440,N_17592);
or U17772 (N_17772,N_17493,N_17574);
or U17773 (N_17773,N_17579,N_17469);
or U17774 (N_17774,N_17425,N_17438);
and U17775 (N_17775,N_17416,N_17458);
or U17776 (N_17776,N_17504,N_17403);
or U17777 (N_17777,N_17513,N_17577);
xor U17778 (N_17778,N_17443,N_17429);
and U17779 (N_17779,N_17421,N_17452);
or U17780 (N_17780,N_17518,N_17568);
nor U17781 (N_17781,N_17553,N_17518);
xor U17782 (N_17782,N_17552,N_17524);
nand U17783 (N_17783,N_17479,N_17575);
and U17784 (N_17784,N_17494,N_17483);
nand U17785 (N_17785,N_17449,N_17569);
or U17786 (N_17786,N_17471,N_17581);
nor U17787 (N_17787,N_17510,N_17554);
nand U17788 (N_17788,N_17547,N_17501);
nand U17789 (N_17789,N_17454,N_17576);
xor U17790 (N_17790,N_17523,N_17532);
or U17791 (N_17791,N_17560,N_17511);
nand U17792 (N_17792,N_17450,N_17580);
and U17793 (N_17793,N_17400,N_17455);
nor U17794 (N_17794,N_17424,N_17563);
nand U17795 (N_17795,N_17515,N_17511);
and U17796 (N_17796,N_17443,N_17468);
nor U17797 (N_17797,N_17449,N_17464);
nand U17798 (N_17798,N_17573,N_17425);
nand U17799 (N_17799,N_17427,N_17465);
or U17800 (N_17800,N_17674,N_17663);
or U17801 (N_17801,N_17621,N_17729);
nor U17802 (N_17802,N_17619,N_17794);
nor U17803 (N_17803,N_17625,N_17661);
or U17804 (N_17804,N_17638,N_17787);
and U17805 (N_17805,N_17693,N_17760);
nor U17806 (N_17806,N_17700,N_17730);
and U17807 (N_17807,N_17649,N_17716);
or U17808 (N_17808,N_17659,N_17669);
nand U17809 (N_17809,N_17768,N_17713);
nor U17810 (N_17810,N_17746,N_17632);
or U17811 (N_17811,N_17622,N_17680);
nand U17812 (N_17812,N_17782,N_17670);
nor U17813 (N_17813,N_17792,N_17747);
and U17814 (N_17814,N_17645,N_17714);
and U17815 (N_17815,N_17718,N_17676);
nor U17816 (N_17816,N_17725,N_17634);
xor U17817 (N_17817,N_17648,N_17675);
nor U17818 (N_17818,N_17607,N_17699);
xnor U17819 (N_17819,N_17751,N_17686);
nand U17820 (N_17820,N_17604,N_17743);
xor U17821 (N_17821,N_17709,N_17600);
nand U17822 (N_17822,N_17650,N_17641);
nand U17823 (N_17823,N_17658,N_17797);
nand U17824 (N_17824,N_17754,N_17708);
nand U17825 (N_17825,N_17673,N_17613);
nor U17826 (N_17826,N_17762,N_17770);
xnor U17827 (N_17827,N_17707,N_17652);
nor U17828 (N_17828,N_17742,N_17627);
or U17829 (N_17829,N_17734,N_17732);
xnor U17830 (N_17830,N_17609,N_17712);
and U17831 (N_17831,N_17655,N_17636);
or U17832 (N_17832,N_17735,N_17776);
and U17833 (N_17833,N_17785,N_17720);
nor U17834 (N_17834,N_17642,N_17705);
or U17835 (N_17835,N_17733,N_17710);
nand U17836 (N_17836,N_17647,N_17790);
nand U17837 (N_17837,N_17653,N_17767);
nand U17838 (N_17838,N_17623,N_17701);
nand U17839 (N_17839,N_17715,N_17774);
nor U17840 (N_17840,N_17692,N_17799);
nor U17841 (N_17841,N_17689,N_17711);
xor U17842 (N_17842,N_17786,N_17656);
and U17843 (N_17843,N_17706,N_17603);
nand U17844 (N_17844,N_17761,N_17796);
nor U17845 (N_17845,N_17795,N_17740);
nor U17846 (N_17846,N_17660,N_17775);
or U17847 (N_17847,N_17688,N_17657);
xnor U17848 (N_17848,N_17777,N_17752);
xnor U17849 (N_17849,N_17757,N_17783);
nand U17850 (N_17850,N_17608,N_17618);
xor U17851 (N_17851,N_17788,N_17697);
xnor U17852 (N_17852,N_17672,N_17764);
and U17853 (N_17853,N_17694,N_17704);
and U17854 (N_17854,N_17643,N_17690);
xnor U17855 (N_17855,N_17696,N_17611);
nand U17856 (N_17856,N_17681,N_17624);
or U17857 (N_17857,N_17798,N_17756);
or U17858 (N_17858,N_17620,N_17639);
or U17859 (N_17859,N_17668,N_17703);
and U17860 (N_17860,N_17749,N_17606);
and U17861 (N_17861,N_17671,N_17773);
xnor U17862 (N_17862,N_17630,N_17772);
and U17863 (N_17863,N_17605,N_17781);
nand U17864 (N_17864,N_17695,N_17698);
or U17865 (N_17865,N_17646,N_17679);
or U17866 (N_17866,N_17666,N_17612);
or U17867 (N_17867,N_17739,N_17737);
nor U17868 (N_17868,N_17702,N_17662);
xnor U17869 (N_17869,N_17723,N_17766);
xnor U17870 (N_17870,N_17722,N_17687);
xor U17871 (N_17871,N_17779,N_17684);
nand U17872 (N_17872,N_17741,N_17721);
and U17873 (N_17873,N_17717,N_17629);
or U17874 (N_17874,N_17626,N_17665);
nand U17875 (N_17875,N_17726,N_17683);
nand U17876 (N_17876,N_17748,N_17614);
and U17877 (N_17877,N_17789,N_17780);
nor U17878 (N_17878,N_17778,N_17719);
xnor U17879 (N_17879,N_17755,N_17602);
or U17880 (N_17880,N_17654,N_17750);
xor U17881 (N_17881,N_17724,N_17784);
xor U17882 (N_17882,N_17617,N_17637);
xnor U17883 (N_17883,N_17744,N_17745);
xnor U17884 (N_17884,N_17664,N_17736);
nor U17885 (N_17885,N_17738,N_17758);
nand U17886 (N_17886,N_17763,N_17667);
or U17887 (N_17887,N_17677,N_17753);
nand U17888 (N_17888,N_17685,N_17678);
xor U17889 (N_17889,N_17610,N_17644);
and U17890 (N_17890,N_17759,N_17633);
nand U17891 (N_17891,N_17615,N_17628);
nand U17892 (N_17892,N_17731,N_17635);
or U17893 (N_17893,N_17682,N_17727);
nand U17894 (N_17894,N_17771,N_17728);
nor U17895 (N_17895,N_17691,N_17651);
xor U17896 (N_17896,N_17793,N_17791);
or U17897 (N_17897,N_17769,N_17616);
and U17898 (N_17898,N_17631,N_17640);
nor U17899 (N_17899,N_17765,N_17601);
and U17900 (N_17900,N_17794,N_17746);
nand U17901 (N_17901,N_17620,N_17734);
nor U17902 (N_17902,N_17614,N_17784);
nand U17903 (N_17903,N_17722,N_17701);
xnor U17904 (N_17904,N_17667,N_17735);
xnor U17905 (N_17905,N_17746,N_17639);
or U17906 (N_17906,N_17601,N_17623);
and U17907 (N_17907,N_17617,N_17795);
and U17908 (N_17908,N_17767,N_17700);
nor U17909 (N_17909,N_17644,N_17637);
or U17910 (N_17910,N_17764,N_17688);
or U17911 (N_17911,N_17744,N_17633);
and U17912 (N_17912,N_17627,N_17658);
nand U17913 (N_17913,N_17787,N_17763);
nor U17914 (N_17914,N_17659,N_17670);
nor U17915 (N_17915,N_17788,N_17665);
xnor U17916 (N_17916,N_17689,N_17668);
nor U17917 (N_17917,N_17635,N_17750);
nor U17918 (N_17918,N_17691,N_17703);
nand U17919 (N_17919,N_17690,N_17621);
nand U17920 (N_17920,N_17642,N_17785);
xnor U17921 (N_17921,N_17639,N_17618);
and U17922 (N_17922,N_17698,N_17611);
and U17923 (N_17923,N_17616,N_17743);
nand U17924 (N_17924,N_17733,N_17645);
or U17925 (N_17925,N_17643,N_17608);
and U17926 (N_17926,N_17631,N_17744);
and U17927 (N_17927,N_17707,N_17620);
xor U17928 (N_17928,N_17717,N_17784);
nand U17929 (N_17929,N_17632,N_17637);
xnor U17930 (N_17930,N_17646,N_17763);
or U17931 (N_17931,N_17646,N_17715);
and U17932 (N_17932,N_17733,N_17689);
xor U17933 (N_17933,N_17763,N_17731);
nor U17934 (N_17934,N_17748,N_17740);
nand U17935 (N_17935,N_17735,N_17731);
nand U17936 (N_17936,N_17703,N_17750);
xnor U17937 (N_17937,N_17620,N_17785);
nor U17938 (N_17938,N_17615,N_17635);
nor U17939 (N_17939,N_17724,N_17628);
nor U17940 (N_17940,N_17783,N_17706);
or U17941 (N_17941,N_17689,N_17706);
and U17942 (N_17942,N_17772,N_17747);
nand U17943 (N_17943,N_17624,N_17709);
or U17944 (N_17944,N_17761,N_17798);
nand U17945 (N_17945,N_17608,N_17769);
and U17946 (N_17946,N_17713,N_17657);
nor U17947 (N_17947,N_17616,N_17633);
nand U17948 (N_17948,N_17644,N_17707);
xor U17949 (N_17949,N_17726,N_17737);
xor U17950 (N_17950,N_17758,N_17798);
nand U17951 (N_17951,N_17687,N_17638);
xor U17952 (N_17952,N_17756,N_17631);
and U17953 (N_17953,N_17711,N_17655);
or U17954 (N_17954,N_17751,N_17760);
or U17955 (N_17955,N_17620,N_17611);
or U17956 (N_17956,N_17680,N_17615);
nor U17957 (N_17957,N_17797,N_17710);
nor U17958 (N_17958,N_17726,N_17796);
or U17959 (N_17959,N_17680,N_17734);
nand U17960 (N_17960,N_17743,N_17639);
and U17961 (N_17961,N_17686,N_17696);
nor U17962 (N_17962,N_17644,N_17744);
or U17963 (N_17963,N_17745,N_17759);
xor U17964 (N_17964,N_17756,N_17788);
nor U17965 (N_17965,N_17657,N_17788);
or U17966 (N_17966,N_17777,N_17667);
nand U17967 (N_17967,N_17660,N_17796);
xor U17968 (N_17968,N_17610,N_17750);
and U17969 (N_17969,N_17646,N_17628);
and U17970 (N_17970,N_17754,N_17600);
nand U17971 (N_17971,N_17711,N_17632);
and U17972 (N_17972,N_17708,N_17710);
xor U17973 (N_17973,N_17746,N_17652);
or U17974 (N_17974,N_17728,N_17798);
or U17975 (N_17975,N_17695,N_17748);
or U17976 (N_17976,N_17693,N_17644);
nor U17977 (N_17977,N_17744,N_17715);
and U17978 (N_17978,N_17634,N_17648);
or U17979 (N_17979,N_17734,N_17648);
or U17980 (N_17980,N_17741,N_17656);
nand U17981 (N_17981,N_17790,N_17665);
nor U17982 (N_17982,N_17728,N_17622);
xnor U17983 (N_17983,N_17651,N_17799);
xnor U17984 (N_17984,N_17720,N_17732);
nor U17985 (N_17985,N_17778,N_17605);
nand U17986 (N_17986,N_17729,N_17744);
and U17987 (N_17987,N_17699,N_17665);
or U17988 (N_17988,N_17671,N_17719);
nand U17989 (N_17989,N_17742,N_17623);
nand U17990 (N_17990,N_17620,N_17691);
or U17991 (N_17991,N_17786,N_17762);
xnor U17992 (N_17992,N_17694,N_17791);
xor U17993 (N_17993,N_17793,N_17688);
nand U17994 (N_17994,N_17756,N_17644);
and U17995 (N_17995,N_17625,N_17655);
or U17996 (N_17996,N_17677,N_17674);
or U17997 (N_17997,N_17770,N_17763);
xnor U17998 (N_17998,N_17759,N_17787);
nand U17999 (N_17999,N_17700,N_17749);
and U18000 (N_18000,N_17872,N_17895);
nor U18001 (N_18001,N_17838,N_17892);
and U18002 (N_18002,N_17949,N_17999);
nand U18003 (N_18003,N_17985,N_17964);
nor U18004 (N_18004,N_17906,N_17902);
and U18005 (N_18005,N_17973,N_17947);
or U18006 (N_18006,N_17917,N_17825);
nand U18007 (N_18007,N_17846,N_17827);
and U18008 (N_18008,N_17831,N_17970);
or U18009 (N_18009,N_17922,N_17866);
or U18010 (N_18010,N_17974,N_17855);
or U18011 (N_18011,N_17994,N_17891);
nand U18012 (N_18012,N_17993,N_17839);
or U18013 (N_18013,N_17890,N_17988);
xor U18014 (N_18014,N_17908,N_17863);
or U18015 (N_18015,N_17894,N_17904);
or U18016 (N_18016,N_17942,N_17929);
or U18017 (N_18017,N_17806,N_17998);
nand U18018 (N_18018,N_17923,N_17856);
or U18019 (N_18019,N_17840,N_17927);
or U18020 (N_18020,N_17953,N_17980);
or U18021 (N_18021,N_17842,N_17885);
and U18022 (N_18022,N_17975,N_17990);
nand U18023 (N_18023,N_17939,N_17926);
nor U18024 (N_18024,N_17830,N_17898);
or U18025 (N_18025,N_17971,N_17861);
nor U18026 (N_18026,N_17919,N_17886);
xnor U18027 (N_18027,N_17905,N_17805);
and U18028 (N_18028,N_17811,N_17996);
nor U18029 (N_18029,N_17884,N_17835);
nand U18030 (N_18030,N_17916,N_17967);
or U18031 (N_18031,N_17948,N_17984);
nand U18032 (N_18032,N_17911,N_17935);
xor U18033 (N_18033,N_17937,N_17944);
nand U18034 (N_18034,N_17918,N_17818);
or U18035 (N_18035,N_17871,N_17897);
nand U18036 (N_18036,N_17828,N_17879);
nand U18037 (N_18037,N_17834,N_17819);
and U18038 (N_18038,N_17938,N_17857);
xor U18039 (N_18039,N_17934,N_17941);
and U18040 (N_18040,N_17849,N_17848);
or U18041 (N_18041,N_17976,N_17946);
nor U18042 (N_18042,N_17957,N_17921);
nand U18043 (N_18043,N_17931,N_17820);
and U18044 (N_18044,N_17950,N_17854);
nor U18045 (N_18045,N_17968,N_17829);
and U18046 (N_18046,N_17837,N_17865);
nand U18047 (N_18047,N_17961,N_17997);
and U18048 (N_18048,N_17809,N_17982);
nor U18049 (N_18049,N_17862,N_17932);
xor U18050 (N_18050,N_17876,N_17903);
and U18051 (N_18051,N_17943,N_17992);
xor U18052 (N_18052,N_17928,N_17966);
nor U18053 (N_18053,N_17845,N_17877);
nor U18054 (N_18054,N_17962,N_17989);
xor U18055 (N_18055,N_17882,N_17987);
and U18056 (N_18056,N_17815,N_17878);
xor U18057 (N_18057,N_17914,N_17844);
xor U18058 (N_18058,N_17813,N_17870);
nand U18059 (N_18059,N_17873,N_17958);
nor U18060 (N_18060,N_17801,N_17956);
nor U18061 (N_18061,N_17913,N_17858);
and U18062 (N_18062,N_17812,N_17960);
or U18063 (N_18063,N_17954,N_17802);
nand U18064 (N_18064,N_17851,N_17883);
or U18065 (N_18065,N_17940,N_17816);
xnor U18066 (N_18066,N_17853,N_17807);
nand U18067 (N_18067,N_17945,N_17821);
xor U18068 (N_18068,N_17983,N_17907);
or U18069 (N_18069,N_17869,N_17981);
or U18070 (N_18070,N_17887,N_17823);
xnor U18071 (N_18071,N_17965,N_17868);
nor U18072 (N_18072,N_17836,N_17955);
and U18073 (N_18073,N_17874,N_17850);
or U18074 (N_18074,N_17817,N_17893);
xnor U18075 (N_18075,N_17889,N_17930);
xor U18076 (N_18076,N_17952,N_17824);
or U18077 (N_18077,N_17909,N_17822);
xnor U18078 (N_18078,N_17832,N_17852);
xor U18079 (N_18079,N_17978,N_17833);
nand U18080 (N_18080,N_17826,N_17875);
nand U18081 (N_18081,N_17900,N_17963);
or U18082 (N_18082,N_17979,N_17888);
nor U18083 (N_18083,N_17860,N_17925);
nand U18084 (N_18084,N_17843,N_17814);
xnor U18085 (N_18085,N_17808,N_17951);
nand U18086 (N_18086,N_17804,N_17867);
or U18087 (N_18087,N_17991,N_17920);
or U18088 (N_18088,N_17896,N_17880);
or U18089 (N_18089,N_17847,N_17936);
or U18090 (N_18090,N_17803,N_17995);
xor U18091 (N_18091,N_17800,N_17841);
xor U18092 (N_18092,N_17810,N_17910);
and U18093 (N_18093,N_17859,N_17986);
nor U18094 (N_18094,N_17924,N_17881);
nand U18095 (N_18095,N_17901,N_17969);
and U18096 (N_18096,N_17912,N_17915);
nor U18097 (N_18097,N_17977,N_17959);
nor U18098 (N_18098,N_17972,N_17933);
nand U18099 (N_18099,N_17864,N_17899);
xnor U18100 (N_18100,N_17859,N_17832);
nor U18101 (N_18101,N_17935,N_17883);
xnor U18102 (N_18102,N_17917,N_17895);
nand U18103 (N_18103,N_17881,N_17903);
nor U18104 (N_18104,N_17903,N_17967);
nor U18105 (N_18105,N_17998,N_17919);
and U18106 (N_18106,N_17937,N_17886);
nand U18107 (N_18107,N_17949,N_17973);
nand U18108 (N_18108,N_17987,N_17989);
nand U18109 (N_18109,N_17879,N_17935);
nand U18110 (N_18110,N_17962,N_17835);
and U18111 (N_18111,N_17902,N_17907);
and U18112 (N_18112,N_17834,N_17916);
nand U18113 (N_18113,N_17923,N_17948);
nand U18114 (N_18114,N_17959,N_17932);
and U18115 (N_18115,N_17924,N_17986);
or U18116 (N_18116,N_17809,N_17876);
xor U18117 (N_18117,N_17959,N_17929);
or U18118 (N_18118,N_17894,N_17986);
and U18119 (N_18119,N_17876,N_17977);
or U18120 (N_18120,N_17932,N_17863);
nor U18121 (N_18121,N_17866,N_17835);
xnor U18122 (N_18122,N_17966,N_17957);
xor U18123 (N_18123,N_17959,N_17884);
nor U18124 (N_18124,N_17860,N_17832);
xnor U18125 (N_18125,N_17906,N_17961);
and U18126 (N_18126,N_17989,N_17985);
nor U18127 (N_18127,N_17943,N_17999);
xnor U18128 (N_18128,N_17854,N_17892);
nand U18129 (N_18129,N_17843,N_17826);
nand U18130 (N_18130,N_17836,N_17986);
nand U18131 (N_18131,N_17944,N_17851);
xor U18132 (N_18132,N_17917,N_17922);
and U18133 (N_18133,N_17951,N_17874);
nor U18134 (N_18134,N_17914,N_17931);
or U18135 (N_18135,N_17999,N_17817);
nor U18136 (N_18136,N_17905,N_17943);
nand U18137 (N_18137,N_17953,N_17806);
nand U18138 (N_18138,N_17820,N_17824);
nor U18139 (N_18139,N_17876,N_17842);
nor U18140 (N_18140,N_17895,N_17972);
or U18141 (N_18141,N_17909,N_17941);
xnor U18142 (N_18142,N_17991,N_17959);
nor U18143 (N_18143,N_17961,N_17994);
nand U18144 (N_18144,N_17994,N_17858);
nor U18145 (N_18145,N_17893,N_17981);
or U18146 (N_18146,N_17935,N_17932);
nand U18147 (N_18147,N_17974,N_17867);
xnor U18148 (N_18148,N_17872,N_17960);
nand U18149 (N_18149,N_17942,N_17904);
and U18150 (N_18150,N_17841,N_17819);
nor U18151 (N_18151,N_17861,N_17879);
or U18152 (N_18152,N_17830,N_17835);
and U18153 (N_18153,N_17882,N_17912);
or U18154 (N_18154,N_17969,N_17861);
nor U18155 (N_18155,N_17903,N_17819);
and U18156 (N_18156,N_17917,N_17970);
and U18157 (N_18157,N_17802,N_17928);
and U18158 (N_18158,N_17925,N_17812);
and U18159 (N_18159,N_17826,N_17937);
or U18160 (N_18160,N_17951,N_17996);
and U18161 (N_18161,N_17851,N_17863);
nand U18162 (N_18162,N_17852,N_17880);
nor U18163 (N_18163,N_17963,N_17823);
nor U18164 (N_18164,N_17804,N_17869);
and U18165 (N_18165,N_17993,N_17845);
nor U18166 (N_18166,N_17943,N_17869);
xnor U18167 (N_18167,N_17954,N_17816);
nand U18168 (N_18168,N_17858,N_17969);
or U18169 (N_18169,N_17961,N_17918);
xor U18170 (N_18170,N_17979,N_17916);
xor U18171 (N_18171,N_17994,N_17905);
or U18172 (N_18172,N_17845,N_17889);
xnor U18173 (N_18173,N_17844,N_17918);
nor U18174 (N_18174,N_17969,N_17804);
and U18175 (N_18175,N_17866,N_17820);
nor U18176 (N_18176,N_17866,N_17885);
nand U18177 (N_18177,N_17904,N_17992);
and U18178 (N_18178,N_17875,N_17801);
or U18179 (N_18179,N_17819,N_17963);
or U18180 (N_18180,N_17913,N_17845);
nand U18181 (N_18181,N_17931,N_17940);
and U18182 (N_18182,N_17909,N_17859);
nor U18183 (N_18183,N_17860,N_17899);
or U18184 (N_18184,N_17979,N_17910);
xnor U18185 (N_18185,N_17828,N_17893);
or U18186 (N_18186,N_17839,N_17898);
or U18187 (N_18187,N_17997,N_17927);
or U18188 (N_18188,N_17929,N_17996);
or U18189 (N_18189,N_17992,N_17989);
xor U18190 (N_18190,N_17907,N_17875);
nand U18191 (N_18191,N_17894,N_17993);
xor U18192 (N_18192,N_17858,N_17907);
nand U18193 (N_18193,N_17903,N_17850);
nor U18194 (N_18194,N_17818,N_17810);
and U18195 (N_18195,N_17908,N_17802);
and U18196 (N_18196,N_17942,N_17952);
and U18197 (N_18197,N_17826,N_17829);
xnor U18198 (N_18198,N_17829,N_17924);
xor U18199 (N_18199,N_17921,N_17938);
nor U18200 (N_18200,N_18146,N_18085);
or U18201 (N_18201,N_18124,N_18129);
nor U18202 (N_18202,N_18041,N_18040);
xnor U18203 (N_18203,N_18172,N_18127);
xnor U18204 (N_18204,N_18029,N_18187);
and U18205 (N_18205,N_18070,N_18120);
and U18206 (N_18206,N_18123,N_18084);
and U18207 (N_18207,N_18034,N_18073);
nor U18208 (N_18208,N_18173,N_18000);
or U18209 (N_18209,N_18079,N_18076);
nand U18210 (N_18210,N_18038,N_18068);
or U18211 (N_18211,N_18052,N_18153);
xor U18212 (N_18212,N_18134,N_18167);
nand U18213 (N_18213,N_18077,N_18180);
xor U18214 (N_18214,N_18069,N_18031);
and U18215 (N_18215,N_18022,N_18020);
and U18216 (N_18216,N_18138,N_18116);
nor U18217 (N_18217,N_18025,N_18036);
nor U18218 (N_18218,N_18039,N_18092);
or U18219 (N_18219,N_18062,N_18166);
nor U18220 (N_18220,N_18192,N_18179);
nor U18221 (N_18221,N_18051,N_18198);
and U18222 (N_18222,N_18049,N_18004);
nor U18223 (N_18223,N_18033,N_18016);
or U18224 (N_18224,N_18121,N_18067);
nand U18225 (N_18225,N_18193,N_18074);
and U18226 (N_18226,N_18024,N_18154);
or U18227 (N_18227,N_18135,N_18071);
nor U18228 (N_18228,N_18018,N_18139);
xnor U18229 (N_18229,N_18042,N_18053);
nand U18230 (N_18230,N_18065,N_18059);
and U18231 (N_18231,N_18086,N_18001);
nand U18232 (N_18232,N_18005,N_18132);
nand U18233 (N_18233,N_18112,N_18155);
or U18234 (N_18234,N_18054,N_18117);
xnor U18235 (N_18235,N_18027,N_18147);
or U18236 (N_18236,N_18111,N_18044);
and U18237 (N_18237,N_18082,N_18103);
nand U18238 (N_18238,N_18028,N_18133);
nand U18239 (N_18239,N_18099,N_18056);
and U18240 (N_18240,N_18108,N_18094);
or U18241 (N_18241,N_18162,N_18128);
and U18242 (N_18242,N_18100,N_18197);
nand U18243 (N_18243,N_18095,N_18021);
nand U18244 (N_18244,N_18131,N_18159);
nand U18245 (N_18245,N_18168,N_18194);
nand U18246 (N_18246,N_18157,N_18115);
and U18247 (N_18247,N_18126,N_18150);
xor U18248 (N_18248,N_18149,N_18188);
nand U18249 (N_18249,N_18089,N_18081);
xnor U18250 (N_18250,N_18106,N_18195);
nand U18251 (N_18251,N_18019,N_18156);
nor U18252 (N_18252,N_18017,N_18143);
nor U18253 (N_18253,N_18110,N_18118);
nor U18254 (N_18254,N_18045,N_18190);
nor U18255 (N_18255,N_18169,N_18043);
or U18256 (N_18256,N_18015,N_18060);
nor U18257 (N_18257,N_18098,N_18144);
or U18258 (N_18258,N_18023,N_18160);
or U18259 (N_18259,N_18032,N_18148);
xor U18260 (N_18260,N_18184,N_18058);
and U18261 (N_18261,N_18072,N_18008);
nand U18262 (N_18262,N_18189,N_18191);
nor U18263 (N_18263,N_18006,N_18090);
or U18264 (N_18264,N_18122,N_18141);
or U18265 (N_18265,N_18183,N_18105);
xnor U18266 (N_18266,N_18152,N_18174);
or U18267 (N_18267,N_18030,N_18151);
nor U18268 (N_18268,N_18002,N_18171);
nand U18269 (N_18269,N_18145,N_18158);
nor U18270 (N_18270,N_18064,N_18012);
or U18271 (N_18271,N_18137,N_18080);
nand U18272 (N_18272,N_18182,N_18164);
nand U18273 (N_18273,N_18011,N_18007);
xnor U18274 (N_18274,N_18199,N_18136);
and U18275 (N_18275,N_18101,N_18009);
or U18276 (N_18276,N_18075,N_18026);
and U18277 (N_18277,N_18104,N_18175);
and U18278 (N_18278,N_18050,N_18013);
and U18279 (N_18279,N_18097,N_18055);
and U18280 (N_18280,N_18078,N_18063);
nand U18281 (N_18281,N_18125,N_18186);
xnor U18282 (N_18282,N_18178,N_18014);
nor U18283 (N_18283,N_18142,N_18003);
xnor U18284 (N_18284,N_18140,N_18181);
and U18285 (N_18285,N_18102,N_18185);
and U18286 (N_18286,N_18176,N_18161);
or U18287 (N_18287,N_18083,N_18165);
nand U18288 (N_18288,N_18114,N_18177);
or U18289 (N_18289,N_18109,N_18093);
xnor U18290 (N_18290,N_18066,N_18096);
xnor U18291 (N_18291,N_18119,N_18046);
xor U18292 (N_18292,N_18037,N_18107);
or U18293 (N_18293,N_18061,N_18113);
and U18294 (N_18294,N_18010,N_18057);
or U18295 (N_18295,N_18087,N_18163);
nor U18296 (N_18296,N_18196,N_18088);
and U18297 (N_18297,N_18048,N_18130);
or U18298 (N_18298,N_18035,N_18091);
nand U18299 (N_18299,N_18047,N_18170);
or U18300 (N_18300,N_18176,N_18000);
xnor U18301 (N_18301,N_18159,N_18057);
nor U18302 (N_18302,N_18012,N_18006);
nand U18303 (N_18303,N_18086,N_18087);
nand U18304 (N_18304,N_18178,N_18055);
xor U18305 (N_18305,N_18026,N_18092);
or U18306 (N_18306,N_18057,N_18064);
and U18307 (N_18307,N_18027,N_18120);
or U18308 (N_18308,N_18188,N_18110);
and U18309 (N_18309,N_18155,N_18061);
or U18310 (N_18310,N_18185,N_18124);
xnor U18311 (N_18311,N_18151,N_18027);
xnor U18312 (N_18312,N_18086,N_18006);
nor U18313 (N_18313,N_18070,N_18041);
nor U18314 (N_18314,N_18182,N_18051);
nand U18315 (N_18315,N_18109,N_18148);
or U18316 (N_18316,N_18068,N_18017);
or U18317 (N_18317,N_18136,N_18173);
nor U18318 (N_18318,N_18089,N_18085);
and U18319 (N_18319,N_18055,N_18024);
nand U18320 (N_18320,N_18110,N_18070);
and U18321 (N_18321,N_18196,N_18153);
and U18322 (N_18322,N_18148,N_18085);
nand U18323 (N_18323,N_18147,N_18024);
or U18324 (N_18324,N_18035,N_18178);
nand U18325 (N_18325,N_18086,N_18023);
nand U18326 (N_18326,N_18077,N_18131);
and U18327 (N_18327,N_18190,N_18170);
nor U18328 (N_18328,N_18145,N_18081);
xnor U18329 (N_18329,N_18038,N_18050);
and U18330 (N_18330,N_18181,N_18101);
or U18331 (N_18331,N_18034,N_18047);
and U18332 (N_18332,N_18063,N_18009);
nor U18333 (N_18333,N_18059,N_18024);
xnor U18334 (N_18334,N_18072,N_18085);
nand U18335 (N_18335,N_18179,N_18093);
xnor U18336 (N_18336,N_18194,N_18077);
and U18337 (N_18337,N_18105,N_18065);
nand U18338 (N_18338,N_18071,N_18040);
and U18339 (N_18339,N_18129,N_18162);
or U18340 (N_18340,N_18174,N_18176);
xor U18341 (N_18341,N_18182,N_18106);
nand U18342 (N_18342,N_18106,N_18101);
nor U18343 (N_18343,N_18072,N_18026);
nor U18344 (N_18344,N_18051,N_18032);
and U18345 (N_18345,N_18159,N_18011);
xnor U18346 (N_18346,N_18149,N_18113);
nor U18347 (N_18347,N_18094,N_18008);
or U18348 (N_18348,N_18137,N_18172);
xnor U18349 (N_18349,N_18069,N_18177);
or U18350 (N_18350,N_18083,N_18010);
or U18351 (N_18351,N_18033,N_18030);
xnor U18352 (N_18352,N_18066,N_18091);
or U18353 (N_18353,N_18120,N_18157);
nor U18354 (N_18354,N_18103,N_18198);
or U18355 (N_18355,N_18164,N_18035);
xor U18356 (N_18356,N_18018,N_18156);
or U18357 (N_18357,N_18061,N_18015);
xnor U18358 (N_18358,N_18181,N_18178);
nand U18359 (N_18359,N_18070,N_18165);
nor U18360 (N_18360,N_18094,N_18092);
and U18361 (N_18361,N_18091,N_18165);
nor U18362 (N_18362,N_18107,N_18088);
nor U18363 (N_18363,N_18133,N_18114);
nor U18364 (N_18364,N_18119,N_18128);
xnor U18365 (N_18365,N_18050,N_18157);
nand U18366 (N_18366,N_18057,N_18122);
nand U18367 (N_18367,N_18028,N_18042);
nand U18368 (N_18368,N_18029,N_18185);
nand U18369 (N_18369,N_18169,N_18011);
nor U18370 (N_18370,N_18051,N_18121);
nand U18371 (N_18371,N_18008,N_18101);
or U18372 (N_18372,N_18161,N_18042);
xor U18373 (N_18373,N_18003,N_18114);
nor U18374 (N_18374,N_18163,N_18188);
nor U18375 (N_18375,N_18160,N_18121);
and U18376 (N_18376,N_18184,N_18113);
nand U18377 (N_18377,N_18082,N_18026);
xor U18378 (N_18378,N_18085,N_18079);
xor U18379 (N_18379,N_18082,N_18024);
and U18380 (N_18380,N_18189,N_18133);
xnor U18381 (N_18381,N_18137,N_18074);
nor U18382 (N_18382,N_18073,N_18184);
or U18383 (N_18383,N_18185,N_18024);
and U18384 (N_18384,N_18055,N_18113);
xnor U18385 (N_18385,N_18087,N_18003);
nand U18386 (N_18386,N_18169,N_18174);
nand U18387 (N_18387,N_18143,N_18086);
nand U18388 (N_18388,N_18019,N_18060);
nor U18389 (N_18389,N_18114,N_18126);
or U18390 (N_18390,N_18019,N_18155);
or U18391 (N_18391,N_18175,N_18174);
or U18392 (N_18392,N_18056,N_18187);
nor U18393 (N_18393,N_18055,N_18198);
xor U18394 (N_18394,N_18017,N_18174);
xnor U18395 (N_18395,N_18164,N_18043);
nand U18396 (N_18396,N_18123,N_18021);
or U18397 (N_18397,N_18007,N_18119);
or U18398 (N_18398,N_18147,N_18122);
nand U18399 (N_18399,N_18071,N_18038);
or U18400 (N_18400,N_18258,N_18294);
or U18401 (N_18401,N_18340,N_18377);
nand U18402 (N_18402,N_18396,N_18283);
nand U18403 (N_18403,N_18398,N_18260);
nor U18404 (N_18404,N_18221,N_18382);
or U18405 (N_18405,N_18239,N_18323);
nand U18406 (N_18406,N_18364,N_18250);
xor U18407 (N_18407,N_18228,N_18225);
xor U18408 (N_18408,N_18261,N_18298);
and U18409 (N_18409,N_18305,N_18238);
or U18410 (N_18410,N_18244,N_18234);
and U18411 (N_18411,N_18203,N_18275);
or U18412 (N_18412,N_18263,N_18278);
nand U18413 (N_18413,N_18277,N_18303);
nor U18414 (N_18414,N_18350,N_18297);
or U18415 (N_18415,N_18265,N_18246);
xor U18416 (N_18416,N_18249,N_18227);
nor U18417 (N_18417,N_18206,N_18339);
nand U18418 (N_18418,N_18213,N_18372);
nor U18419 (N_18419,N_18326,N_18317);
nand U18420 (N_18420,N_18272,N_18200);
xnor U18421 (N_18421,N_18355,N_18360);
nor U18422 (N_18422,N_18208,N_18229);
or U18423 (N_18423,N_18352,N_18368);
or U18424 (N_18424,N_18286,N_18300);
and U18425 (N_18425,N_18365,N_18346);
xor U18426 (N_18426,N_18344,N_18395);
xor U18427 (N_18427,N_18212,N_18321);
and U18428 (N_18428,N_18222,N_18388);
nor U18429 (N_18429,N_18356,N_18308);
nand U18430 (N_18430,N_18370,N_18271);
nand U18431 (N_18431,N_18391,N_18288);
nor U18432 (N_18432,N_18373,N_18330);
xor U18433 (N_18433,N_18349,N_18306);
and U18434 (N_18434,N_18361,N_18386);
nand U18435 (N_18435,N_18320,N_18209);
xor U18436 (N_18436,N_18245,N_18367);
and U18437 (N_18437,N_18231,N_18270);
xor U18438 (N_18438,N_18290,N_18287);
xor U18439 (N_18439,N_18313,N_18211);
and U18440 (N_18440,N_18215,N_18338);
nand U18441 (N_18441,N_18279,N_18237);
xor U18442 (N_18442,N_18289,N_18241);
or U18443 (N_18443,N_18273,N_18334);
or U18444 (N_18444,N_18274,N_18374);
xor U18445 (N_18445,N_18375,N_18337);
nor U18446 (N_18446,N_18366,N_18207);
nor U18447 (N_18447,N_18210,N_18235);
and U18448 (N_18448,N_18315,N_18316);
or U18449 (N_18449,N_18304,N_18332);
xor U18450 (N_18450,N_18387,N_18399);
nand U18451 (N_18451,N_18363,N_18259);
nand U18452 (N_18452,N_18312,N_18240);
and U18453 (N_18453,N_18379,N_18351);
xor U18454 (N_18454,N_18353,N_18291);
nor U18455 (N_18455,N_18264,N_18299);
nand U18456 (N_18456,N_18295,N_18281);
nor U18457 (N_18457,N_18219,N_18383);
and U18458 (N_18458,N_18226,N_18285);
and U18459 (N_18459,N_18310,N_18218);
xnor U18460 (N_18460,N_18301,N_18384);
and U18461 (N_18461,N_18394,N_18343);
xnor U18462 (N_18462,N_18393,N_18202);
and U18463 (N_18463,N_18223,N_18341);
xor U18464 (N_18464,N_18284,N_18268);
and U18465 (N_18465,N_18381,N_18276);
xor U18466 (N_18466,N_18233,N_18314);
nand U18467 (N_18467,N_18369,N_18307);
and U18468 (N_18468,N_18224,N_18201);
nor U18469 (N_18469,N_18214,N_18335);
xnor U18470 (N_18470,N_18309,N_18266);
nand U18471 (N_18471,N_18280,N_18282);
nor U18472 (N_18472,N_18236,N_18357);
nor U18473 (N_18473,N_18232,N_18253);
and U18474 (N_18474,N_18358,N_18230);
or U18475 (N_18475,N_18354,N_18220);
xnor U18476 (N_18476,N_18324,N_18342);
xor U18477 (N_18477,N_18302,N_18251);
and U18478 (N_18478,N_18347,N_18242);
and U18479 (N_18479,N_18359,N_18322);
nor U18480 (N_18480,N_18257,N_18378);
nand U18481 (N_18481,N_18267,N_18397);
and U18482 (N_18482,N_18255,N_18345);
nand U18483 (N_18483,N_18389,N_18325);
and U18484 (N_18484,N_18385,N_18319);
nand U18485 (N_18485,N_18204,N_18256);
xor U18486 (N_18486,N_18243,N_18390);
and U18487 (N_18487,N_18336,N_18327);
nand U18488 (N_18488,N_18362,N_18254);
or U18489 (N_18489,N_18376,N_18217);
nand U18490 (N_18490,N_18216,N_18348);
or U18491 (N_18491,N_18380,N_18252);
or U18492 (N_18492,N_18329,N_18292);
nor U18493 (N_18493,N_18328,N_18311);
xor U18494 (N_18494,N_18205,N_18331);
xnor U18495 (N_18495,N_18262,N_18371);
nor U18496 (N_18496,N_18248,N_18296);
nor U18497 (N_18497,N_18392,N_18247);
and U18498 (N_18498,N_18293,N_18318);
or U18499 (N_18499,N_18333,N_18269);
or U18500 (N_18500,N_18297,N_18360);
or U18501 (N_18501,N_18261,N_18320);
xor U18502 (N_18502,N_18300,N_18341);
nand U18503 (N_18503,N_18340,N_18342);
and U18504 (N_18504,N_18202,N_18396);
and U18505 (N_18505,N_18398,N_18282);
xor U18506 (N_18506,N_18273,N_18215);
nand U18507 (N_18507,N_18201,N_18236);
nand U18508 (N_18508,N_18385,N_18315);
nor U18509 (N_18509,N_18274,N_18291);
and U18510 (N_18510,N_18277,N_18213);
nor U18511 (N_18511,N_18280,N_18298);
xnor U18512 (N_18512,N_18262,N_18319);
and U18513 (N_18513,N_18288,N_18291);
xor U18514 (N_18514,N_18343,N_18346);
xor U18515 (N_18515,N_18380,N_18293);
and U18516 (N_18516,N_18366,N_18209);
and U18517 (N_18517,N_18357,N_18201);
nor U18518 (N_18518,N_18315,N_18323);
or U18519 (N_18519,N_18213,N_18304);
nor U18520 (N_18520,N_18268,N_18351);
nand U18521 (N_18521,N_18257,N_18284);
xor U18522 (N_18522,N_18320,N_18233);
xor U18523 (N_18523,N_18221,N_18364);
or U18524 (N_18524,N_18301,N_18241);
and U18525 (N_18525,N_18365,N_18211);
or U18526 (N_18526,N_18370,N_18200);
or U18527 (N_18527,N_18381,N_18228);
nand U18528 (N_18528,N_18201,N_18228);
nor U18529 (N_18529,N_18302,N_18241);
and U18530 (N_18530,N_18260,N_18337);
nor U18531 (N_18531,N_18317,N_18380);
or U18532 (N_18532,N_18356,N_18239);
or U18533 (N_18533,N_18331,N_18254);
or U18534 (N_18534,N_18259,N_18257);
and U18535 (N_18535,N_18398,N_18242);
and U18536 (N_18536,N_18202,N_18227);
or U18537 (N_18537,N_18287,N_18276);
and U18538 (N_18538,N_18202,N_18300);
and U18539 (N_18539,N_18274,N_18309);
xnor U18540 (N_18540,N_18363,N_18251);
xnor U18541 (N_18541,N_18287,N_18254);
and U18542 (N_18542,N_18256,N_18392);
and U18543 (N_18543,N_18285,N_18312);
nand U18544 (N_18544,N_18333,N_18382);
nor U18545 (N_18545,N_18282,N_18389);
xnor U18546 (N_18546,N_18294,N_18312);
nand U18547 (N_18547,N_18290,N_18303);
nand U18548 (N_18548,N_18365,N_18283);
and U18549 (N_18549,N_18344,N_18343);
or U18550 (N_18550,N_18385,N_18200);
nand U18551 (N_18551,N_18397,N_18293);
and U18552 (N_18552,N_18388,N_18215);
xnor U18553 (N_18553,N_18228,N_18278);
nor U18554 (N_18554,N_18365,N_18302);
and U18555 (N_18555,N_18301,N_18299);
or U18556 (N_18556,N_18217,N_18312);
nand U18557 (N_18557,N_18291,N_18237);
and U18558 (N_18558,N_18391,N_18376);
xnor U18559 (N_18559,N_18380,N_18331);
nand U18560 (N_18560,N_18387,N_18219);
or U18561 (N_18561,N_18288,N_18385);
nor U18562 (N_18562,N_18343,N_18257);
or U18563 (N_18563,N_18241,N_18244);
nand U18564 (N_18564,N_18296,N_18312);
nand U18565 (N_18565,N_18274,N_18368);
and U18566 (N_18566,N_18224,N_18387);
nor U18567 (N_18567,N_18257,N_18287);
or U18568 (N_18568,N_18282,N_18374);
or U18569 (N_18569,N_18312,N_18320);
nor U18570 (N_18570,N_18291,N_18392);
and U18571 (N_18571,N_18317,N_18353);
nand U18572 (N_18572,N_18263,N_18376);
and U18573 (N_18573,N_18261,N_18230);
and U18574 (N_18574,N_18326,N_18276);
nor U18575 (N_18575,N_18306,N_18238);
and U18576 (N_18576,N_18322,N_18375);
nor U18577 (N_18577,N_18275,N_18318);
xor U18578 (N_18578,N_18330,N_18319);
nand U18579 (N_18579,N_18285,N_18372);
nand U18580 (N_18580,N_18242,N_18325);
nand U18581 (N_18581,N_18261,N_18233);
nand U18582 (N_18582,N_18388,N_18253);
or U18583 (N_18583,N_18386,N_18305);
xor U18584 (N_18584,N_18241,N_18243);
or U18585 (N_18585,N_18370,N_18260);
and U18586 (N_18586,N_18215,N_18351);
or U18587 (N_18587,N_18366,N_18211);
xnor U18588 (N_18588,N_18318,N_18356);
and U18589 (N_18589,N_18309,N_18379);
nor U18590 (N_18590,N_18381,N_18205);
and U18591 (N_18591,N_18234,N_18366);
nand U18592 (N_18592,N_18256,N_18355);
or U18593 (N_18593,N_18238,N_18278);
nor U18594 (N_18594,N_18334,N_18282);
nor U18595 (N_18595,N_18335,N_18207);
or U18596 (N_18596,N_18208,N_18270);
nor U18597 (N_18597,N_18347,N_18368);
nand U18598 (N_18598,N_18386,N_18258);
nand U18599 (N_18599,N_18308,N_18209);
or U18600 (N_18600,N_18493,N_18593);
nand U18601 (N_18601,N_18478,N_18468);
nor U18602 (N_18602,N_18489,N_18544);
xor U18603 (N_18603,N_18559,N_18416);
xor U18604 (N_18604,N_18558,N_18466);
nor U18605 (N_18605,N_18449,N_18402);
or U18606 (N_18606,N_18508,N_18506);
nand U18607 (N_18607,N_18497,N_18500);
and U18608 (N_18608,N_18487,N_18457);
or U18609 (N_18609,N_18503,N_18565);
and U18610 (N_18610,N_18407,N_18527);
xor U18611 (N_18611,N_18513,N_18479);
or U18612 (N_18612,N_18461,N_18456);
and U18613 (N_18613,N_18471,N_18514);
nor U18614 (N_18614,N_18473,N_18566);
nand U18615 (N_18615,N_18425,N_18539);
and U18616 (N_18616,N_18502,N_18597);
and U18617 (N_18617,N_18531,N_18447);
or U18618 (N_18618,N_18554,N_18572);
nand U18619 (N_18619,N_18547,N_18525);
nor U18620 (N_18620,N_18437,N_18589);
nand U18621 (N_18621,N_18580,N_18486);
and U18622 (N_18622,N_18534,N_18577);
or U18623 (N_18623,N_18451,N_18418);
xnor U18624 (N_18624,N_18442,N_18480);
or U18625 (N_18625,N_18518,N_18515);
xnor U18626 (N_18626,N_18519,N_18408);
and U18627 (N_18627,N_18439,N_18469);
xnor U18628 (N_18628,N_18549,N_18595);
nand U18629 (N_18629,N_18538,N_18536);
or U18630 (N_18630,N_18511,N_18452);
and U18631 (N_18631,N_18507,N_18555);
nor U18632 (N_18632,N_18415,N_18522);
nand U18633 (N_18633,N_18550,N_18448);
nand U18634 (N_18634,N_18584,N_18533);
or U18635 (N_18635,N_18564,N_18464);
nor U18636 (N_18636,N_18477,N_18470);
or U18637 (N_18637,N_18495,N_18474);
or U18638 (N_18638,N_18516,N_18412);
xor U18639 (N_18639,N_18510,N_18585);
and U18640 (N_18640,N_18557,N_18587);
and U18641 (N_18641,N_18501,N_18560);
nor U18642 (N_18642,N_18460,N_18496);
and U18643 (N_18643,N_18575,N_18440);
nand U18644 (N_18644,N_18484,N_18405);
xor U18645 (N_18645,N_18552,N_18462);
and U18646 (N_18646,N_18488,N_18530);
and U18647 (N_18647,N_18443,N_18433);
and U18648 (N_18648,N_18521,N_18472);
nor U18649 (N_18649,N_18411,N_18517);
and U18650 (N_18650,N_18588,N_18561);
nor U18651 (N_18651,N_18582,N_18567);
xor U18652 (N_18652,N_18563,N_18524);
nor U18653 (N_18653,N_18435,N_18494);
or U18654 (N_18654,N_18401,N_18568);
xnor U18655 (N_18655,N_18546,N_18453);
and U18656 (N_18656,N_18436,N_18537);
nor U18657 (N_18657,N_18512,N_18482);
or U18658 (N_18658,N_18463,N_18490);
nor U18659 (N_18659,N_18543,N_18410);
nor U18660 (N_18660,N_18432,N_18576);
and U18661 (N_18661,N_18545,N_18476);
nand U18662 (N_18662,N_18520,N_18505);
nor U18663 (N_18663,N_18592,N_18417);
and U18664 (N_18664,N_18483,N_18562);
xnor U18665 (N_18665,N_18509,N_18553);
nor U18666 (N_18666,N_18404,N_18498);
xnor U18667 (N_18667,N_18598,N_18570);
and U18668 (N_18668,N_18481,N_18591);
xnor U18669 (N_18669,N_18428,N_18403);
nand U18670 (N_18670,N_18526,N_18419);
nand U18671 (N_18671,N_18581,N_18571);
or U18672 (N_18672,N_18467,N_18504);
nand U18673 (N_18673,N_18523,N_18422);
nor U18674 (N_18674,N_18583,N_18424);
or U18675 (N_18675,N_18413,N_18421);
and U18676 (N_18676,N_18475,N_18450);
nor U18677 (N_18677,N_18455,N_18429);
nor U18678 (N_18678,N_18599,N_18541);
or U18679 (N_18679,N_18431,N_18556);
nor U18680 (N_18680,N_18573,N_18548);
nor U18681 (N_18681,N_18578,N_18438);
or U18682 (N_18682,N_18459,N_18542);
xnor U18683 (N_18683,N_18400,N_18590);
or U18684 (N_18684,N_18529,N_18444);
nand U18685 (N_18685,N_18454,N_18532);
nor U18686 (N_18686,N_18492,N_18579);
xnor U18687 (N_18687,N_18569,N_18406);
or U18688 (N_18688,N_18540,N_18596);
and U18689 (N_18689,N_18465,N_18434);
and U18690 (N_18690,N_18430,N_18423);
xnor U18691 (N_18691,N_18441,N_18458);
and U18692 (N_18692,N_18414,N_18528);
nand U18693 (N_18693,N_18551,N_18446);
nand U18694 (N_18694,N_18426,N_18409);
nand U18695 (N_18695,N_18574,N_18485);
xor U18696 (N_18696,N_18586,N_18420);
xor U18697 (N_18697,N_18594,N_18491);
and U18698 (N_18698,N_18445,N_18427);
and U18699 (N_18699,N_18499,N_18535);
or U18700 (N_18700,N_18517,N_18451);
and U18701 (N_18701,N_18572,N_18589);
and U18702 (N_18702,N_18564,N_18543);
nand U18703 (N_18703,N_18499,N_18467);
or U18704 (N_18704,N_18591,N_18580);
nand U18705 (N_18705,N_18527,N_18416);
and U18706 (N_18706,N_18536,N_18540);
xor U18707 (N_18707,N_18539,N_18548);
xnor U18708 (N_18708,N_18575,N_18420);
nand U18709 (N_18709,N_18430,N_18594);
xor U18710 (N_18710,N_18545,N_18541);
or U18711 (N_18711,N_18506,N_18556);
and U18712 (N_18712,N_18541,N_18400);
nand U18713 (N_18713,N_18438,N_18489);
and U18714 (N_18714,N_18534,N_18406);
xnor U18715 (N_18715,N_18554,N_18567);
nor U18716 (N_18716,N_18577,N_18587);
and U18717 (N_18717,N_18429,N_18562);
or U18718 (N_18718,N_18464,N_18503);
or U18719 (N_18719,N_18584,N_18482);
nand U18720 (N_18720,N_18513,N_18561);
or U18721 (N_18721,N_18439,N_18483);
or U18722 (N_18722,N_18499,N_18599);
nand U18723 (N_18723,N_18541,N_18489);
or U18724 (N_18724,N_18486,N_18480);
nand U18725 (N_18725,N_18466,N_18411);
nand U18726 (N_18726,N_18487,N_18403);
nand U18727 (N_18727,N_18598,N_18545);
xnor U18728 (N_18728,N_18454,N_18447);
and U18729 (N_18729,N_18455,N_18448);
xnor U18730 (N_18730,N_18464,N_18508);
nand U18731 (N_18731,N_18451,N_18565);
nand U18732 (N_18732,N_18555,N_18448);
nand U18733 (N_18733,N_18578,N_18530);
nor U18734 (N_18734,N_18565,N_18447);
nor U18735 (N_18735,N_18438,N_18409);
and U18736 (N_18736,N_18491,N_18407);
nand U18737 (N_18737,N_18590,N_18500);
xnor U18738 (N_18738,N_18517,N_18420);
nand U18739 (N_18739,N_18579,N_18526);
xnor U18740 (N_18740,N_18533,N_18567);
nand U18741 (N_18741,N_18544,N_18554);
nor U18742 (N_18742,N_18533,N_18418);
nor U18743 (N_18743,N_18519,N_18543);
and U18744 (N_18744,N_18567,N_18460);
or U18745 (N_18745,N_18585,N_18590);
nor U18746 (N_18746,N_18578,N_18441);
nand U18747 (N_18747,N_18508,N_18468);
and U18748 (N_18748,N_18447,N_18575);
or U18749 (N_18749,N_18470,N_18493);
nand U18750 (N_18750,N_18441,N_18498);
xor U18751 (N_18751,N_18469,N_18418);
or U18752 (N_18752,N_18535,N_18560);
nor U18753 (N_18753,N_18507,N_18534);
or U18754 (N_18754,N_18467,N_18523);
nor U18755 (N_18755,N_18554,N_18518);
nand U18756 (N_18756,N_18587,N_18529);
nand U18757 (N_18757,N_18406,N_18520);
nand U18758 (N_18758,N_18556,N_18488);
xnor U18759 (N_18759,N_18454,N_18569);
or U18760 (N_18760,N_18561,N_18520);
nand U18761 (N_18761,N_18503,N_18491);
nand U18762 (N_18762,N_18487,N_18530);
or U18763 (N_18763,N_18569,N_18440);
xor U18764 (N_18764,N_18545,N_18564);
xnor U18765 (N_18765,N_18432,N_18408);
nor U18766 (N_18766,N_18581,N_18548);
and U18767 (N_18767,N_18585,N_18516);
xnor U18768 (N_18768,N_18439,N_18515);
nor U18769 (N_18769,N_18478,N_18540);
xor U18770 (N_18770,N_18421,N_18464);
and U18771 (N_18771,N_18468,N_18549);
nor U18772 (N_18772,N_18494,N_18566);
nand U18773 (N_18773,N_18493,N_18572);
and U18774 (N_18774,N_18537,N_18497);
xor U18775 (N_18775,N_18574,N_18519);
and U18776 (N_18776,N_18511,N_18443);
xnor U18777 (N_18777,N_18557,N_18518);
and U18778 (N_18778,N_18502,N_18589);
nand U18779 (N_18779,N_18563,N_18558);
xnor U18780 (N_18780,N_18539,N_18483);
nand U18781 (N_18781,N_18497,N_18423);
nor U18782 (N_18782,N_18556,N_18425);
nor U18783 (N_18783,N_18470,N_18462);
nand U18784 (N_18784,N_18432,N_18471);
xor U18785 (N_18785,N_18598,N_18471);
xor U18786 (N_18786,N_18551,N_18458);
or U18787 (N_18787,N_18406,N_18478);
nor U18788 (N_18788,N_18421,N_18537);
nor U18789 (N_18789,N_18526,N_18434);
nor U18790 (N_18790,N_18521,N_18520);
and U18791 (N_18791,N_18580,N_18415);
nor U18792 (N_18792,N_18402,N_18510);
xor U18793 (N_18793,N_18492,N_18420);
or U18794 (N_18794,N_18506,N_18590);
xnor U18795 (N_18795,N_18441,N_18592);
and U18796 (N_18796,N_18472,N_18545);
or U18797 (N_18797,N_18518,N_18584);
nand U18798 (N_18798,N_18524,N_18536);
nor U18799 (N_18799,N_18430,N_18598);
xor U18800 (N_18800,N_18600,N_18746);
xnor U18801 (N_18801,N_18692,N_18650);
or U18802 (N_18802,N_18694,N_18748);
nand U18803 (N_18803,N_18760,N_18763);
nor U18804 (N_18804,N_18625,N_18645);
nor U18805 (N_18805,N_18767,N_18668);
xor U18806 (N_18806,N_18734,N_18718);
nand U18807 (N_18807,N_18751,N_18784);
and U18808 (N_18808,N_18674,N_18644);
xor U18809 (N_18809,N_18612,N_18745);
and U18810 (N_18810,N_18611,N_18621);
nand U18811 (N_18811,N_18619,N_18770);
and U18812 (N_18812,N_18682,N_18780);
xor U18813 (N_18813,N_18620,N_18779);
nor U18814 (N_18814,N_18605,N_18678);
and U18815 (N_18815,N_18696,N_18688);
nand U18816 (N_18816,N_18783,N_18638);
and U18817 (N_18817,N_18691,N_18624);
xor U18818 (N_18818,N_18643,N_18686);
nor U18819 (N_18819,N_18733,N_18609);
nor U18820 (N_18820,N_18680,N_18735);
and U18821 (N_18821,N_18613,N_18663);
and U18822 (N_18822,N_18657,N_18737);
nand U18823 (N_18823,N_18704,N_18654);
or U18824 (N_18824,N_18789,N_18772);
xnor U18825 (N_18825,N_18679,N_18701);
xor U18826 (N_18826,N_18653,N_18790);
or U18827 (N_18827,N_18673,N_18604);
nand U18828 (N_18828,N_18787,N_18699);
nor U18829 (N_18829,N_18689,N_18753);
xor U18830 (N_18830,N_18670,N_18723);
nand U18831 (N_18831,N_18736,N_18616);
or U18832 (N_18832,N_18658,N_18750);
and U18833 (N_18833,N_18744,N_18759);
or U18834 (N_18834,N_18747,N_18785);
nand U18835 (N_18835,N_18626,N_18719);
and U18836 (N_18836,N_18683,N_18708);
nand U18837 (N_18837,N_18738,N_18607);
nand U18838 (N_18838,N_18603,N_18788);
and U18839 (N_18839,N_18659,N_18703);
and U18840 (N_18840,N_18637,N_18608);
xor U18841 (N_18841,N_18667,N_18728);
nand U18842 (N_18842,N_18687,N_18797);
nor U18843 (N_18843,N_18634,N_18642);
or U18844 (N_18844,N_18752,N_18690);
nor U18845 (N_18845,N_18755,N_18766);
xnor U18846 (N_18846,N_18671,N_18754);
or U18847 (N_18847,N_18666,N_18649);
nor U18848 (N_18848,N_18631,N_18618);
xnor U18849 (N_18849,N_18794,N_18676);
nor U18850 (N_18850,N_18757,N_18606);
and U18851 (N_18851,N_18622,N_18617);
nor U18852 (N_18852,N_18726,N_18672);
xnor U18853 (N_18853,N_18720,N_18707);
and U18854 (N_18854,N_18739,N_18727);
and U18855 (N_18855,N_18721,N_18773);
and U18856 (N_18856,N_18702,N_18732);
nand U18857 (N_18857,N_18652,N_18795);
nor U18858 (N_18858,N_18610,N_18695);
nor U18859 (N_18859,N_18651,N_18661);
nand U18860 (N_18860,N_18782,N_18615);
and U18861 (N_18861,N_18771,N_18633);
xnor U18862 (N_18862,N_18697,N_18778);
and U18863 (N_18863,N_18628,N_18706);
or U18864 (N_18864,N_18722,N_18709);
xnor U18865 (N_18865,N_18715,N_18640);
and U18866 (N_18866,N_18776,N_18705);
nor U18867 (N_18867,N_18698,N_18614);
and U18868 (N_18868,N_18665,N_18677);
and U18869 (N_18869,N_18742,N_18664);
xnor U18870 (N_18870,N_18791,N_18655);
nand U18871 (N_18871,N_18700,N_18675);
nor U18872 (N_18872,N_18714,N_18717);
xor U18873 (N_18873,N_18756,N_18749);
nand U18874 (N_18874,N_18775,N_18796);
xnor U18875 (N_18875,N_18710,N_18725);
nand U18876 (N_18876,N_18761,N_18636);
or U18877 (N_18877,N_18765,N_18758);
and U18878 (N_18878,N_18711,N_18669);
or U18879 (N_18879,N_18648,N_18769);
or U18880 (N_18880,N_18743,N_18635);
or U18881 (N_18881,N_18660,N_18762);
and U18882 (N_18882,N_18777,N_18740);
nor U18883 (N_18883,N_18685,N_18639);
and U18884 (N_18884,N_18729,N_18713);
nor U18885 (N_18885,N_18630,N_18793);
xor U18886 (N_18886,N_18693,N_18656);
and U18887 (N_18887,N_18641,N_18798);
nor U18888 (N_18888,N_18792,N_18774);
and U18889 (N_18889,N_18684,N_18781);
nor U18890 (N_18890,N_18768,N_18716);
nor U18891 (N_18891,N_18764,N_18712);
xor U18892 (N_18892,N_18724,N_18799);
and U18893 (N_18893,N_18601,N_18741);
nand U18894 (N_18894,N_18629,N_18647);
or U18895 (N_18895,N_18602,N_18662);
nand U18896 (N_18896,N_18646,N_18627);
nand U18897 (N_18897,N_18730,N_18632);
xor U18898 (N_18898,N_18786,N_18731);
or U18899 (N_18899,N_18623,N_18681);
or U18900 (N_18900,N_18686,N_18647);
or U18901 (N_18901,N_18617,N_18715);
xor U18902 (N_18902,N_18618,N_18637);
or U18903 (N_18903,N_18784,N_18708);
xor U18904 (N_18904,N_18785,N_18733);
nand U18905 (N_18905,N_18756,N_18794);
nand U18906 (N_18906,N_18656,N_18794);
or U18907 (N_18907,N_18732,N_18642);
nor U18908 (N_18908,N_18730,N_18654);
xnor U18909 (N_18909,N_18779,N_18718);
xnor U18910 (N_18910,N_18609,N_18792);
xnor U18911 (N_18911,N_18755,N_18784);
and U18912 (N_18912,N_18752,N_18677);
nand U18913 (N_18913,N_18637,N_18741);
or U18914 (N_18914,N_18645,N_18714);
nor U18915 (N_18915,N_18640,N_18688);
or U18916 (N_18916,N_18713,N_18768);
xnor U18917 (N_18917,N_18633,N_18630);
nand U18918 (N_18918,N_18641,N_18784);
xnor U18919 (N_18919,N_18682,N_18692);
and U18920 (N_18920,N_18606,N_18628);
and U18921 (N_18921,N_18603,N_18773);
nor U18922 (N_18922,N_18714,N_18633);
and U18923 (N_18923,N_18754,N_18635);
nand U18924 (N_18924,N_18618,N_18765);
or U18925 (N_18925,N_18786,N_18770);
nor U18926 (N_18926,N_18736,N_18653);
or U18927 (N_18927,N_18653,N_18695);
or U18928 (N_18928,N_18740,N_18737);
nor U18929 (N_18929,N_18742,N_18782);
xor U18930 (N_18930,N_18721,N_18684);
or U18931 (N_18931,N_18708,N_18627);
nor U18932 (N_18932,N_18694,N_18607);
and U18933 (N_18933,N_18630,N_18785);
xnor U18934 (N_18934,N_18794,N_18735);
or U18935 (N_18935,N_18725,N_18625);
nor U18936 (N_18936,N_18653,N_18716);
or U18937 (N_18937,N_18610,N_18740);
nor U18938 (N_18938,N_18755,N_18686);
xor U18939 (N_18939,N_18665,N_18658);
nand U18940 (N_18940,N_18660,N_18638);
nor U18941 (N_18941,N_18768,N_18682);
or U18942 (N_18942,N_18643,N_18608);
and U18943 (N_18943,N_18682,N_18743);
xor U18944 (N_18944,N_18644,N_18613);
or U18945 (N_18945,N_18741,N_18704);
nor U18946 (N_18946,N_18725,N_18708);
nor U18947 (N_18947,N_18676,N_18772);
and U18948 (N_18948,N_18628,N_18654);
nand U18949 (N_18949,N_18773,N_18665);
nor U18950 (N_18950,N_18664,N_18653);
and U18951 (N_18951,N_18794,N_18632);
xor U18952 (N_18952,N_18623,N_18767);
and U18953 (N_18953,N_18753,N_18640);
and U18954 (N_18954,N_18605,N_18776);
or U18955 (N_18955,N_18667,N_18787);
or U18956 (N_18956,N_18708,N_18621);
and U18957 (N_18957,N_18617,N_18790);
xnor U18958 (N_18958,N_18681,N_18635);
nand U18959 (N_18959,N_18716,N_18656);
nor U18960 (N_18960,N_18675,N_18713);
xor U18961 (N_18961,N_18619,N_18704);
or U18962 (N_18962,N_18670,N_18775);
nand U18963 (N_18963,N_18747,N_18616);
xor U18964 (N_18964,N_18639,N_18650);
or U18965 (N_18965,N_18691,N_18695);
xor U18966 (N_18966,N_18741,N_18609);
and U18967 (N_18967,N_18741,N_18711);
nand U18968 (N_18968,N_18779,N_18686);
or U18969 (N_18969,N_18642,N_18720);
nand U18970 (N_18970,N_18774,N_18665);
or U18971 (N_18971,N_18650,N_18756);
xnor U18972 (N_18972,N_18796,N_18718);
xor U18973 (N_18973,N_18714,N_18635);
xnor U18974 (N_18974,N_18690,N_18686);
or U18975 (N_18975,N_18787,N_18732);
nor U18976 (N_18976,N_18634,N_18622);
nor U18977 (N_18977,N_18720,N_18644);
xnor U18978 (N_18978,N_18677,N_18607);
nand U18979 (N_18979,N_18721,N_18652);
or U18980 (N_18980,N_18741,N_18761);
nor U18981 (N_18981,N_18724,N_18781);
nor U18982 (N_18982,N_18648,N_18752);
nor U18983 (N_18983,N_18695,N_18742);
xor U18984 (N_18984,N_18742,N_18610);
nand U18985 (N_18985,N_18604,N_18776);
xor U18986 (N_18986,N_18774,N_18636);
xnor U18987 (N_18987,N_18736,N_18669);
xor U18988 (N_18988,N_18790,N_18760);
or U18989 (N_18989,N_18680,N_18764);
and U18990 (N_18990,N_18660,N_18634);
nand U18991 (N_18991,N_18603,N_18655);
or U18992 (N_18992,N_18647,N_18668);
nor U18993 (N_18993,N_18799,N_18627);
nor U18994 (N_18994,N_18787,N_18778);
or U18995 (N_18995,N_18663,N_18636);
nor U18996 (N_18996,N_18787,N_18600);
xnor U18997 (N_18997,N_18624,N_18755);
and U18998 (N_18998,N_18723,N_18711);
nand U18999 (N_18999,N_18620,N_18667);
or U19000 (N_19000,N_18878,N_18984);
or U19001 (N_19001,N_18889,N_18829);
or U19002 (N_19002,N_18876,N_18817);
nor U19003 (N_19003,N_18820,N_18886);
nor U19004 (N_19004,N_18899,N_18806);
and U19005 (N_19005,N_18906,N_18840);
and U19006 (N_19006,N_18975,N_18846);
nand U19007 (N_19007,N_18935,N_18967);
or U19008 (N_19008,N_18986,N_18887);
nor U19009 (N_19009,N_18849,N_18873);
and U19010 (N_19010,N_18892,N_18924);
nand U19011 (N_19011,N_18801,N_18996);
nand U19012 (N_19012,N_18859,N_18913);
and U19013 (N_19013,N_18896,N_18860);
xor U19014 (N_19014,N_18912,N_18917);
xor U19015 (N_19015,N_18958,N_18841);
nor U19016 (N_19016,N_18865,N_18895);
and U19017 (N_19017,N_18925,N_18898);
nand U19018 (N_19018,N_18989,N_18845);
or U19019 (N_19019,N_18811,N_18982);
xnor U19020 (N_19020,N_18883,N_18914);
nor U19021 (N_19021,N_18930,N_18812);
nand U19022 (N_19022,N_18833,N_18993);
and U19023 (N_19023,N_18947,N_18923);
nand U19024 (N_19024,N_18819,N_18940);
nand U19025 (N_19025,N_18861,N_18905);
xnor U19026 (N_19026,N_18891,N_18863);
and U19027 (N_19027,N_18884,N_18866);
nor U19028 (N_19028,N_18858,N_18988);
nand U19029 (N_19029,N_18952,N_18921);
or U19030 (N_19030,N_18971,N_18918);
and U19031 (N_19031,N_18908,N_18965);
or U19032 (N_19032,N_18992,N_18962);
xor U19033 (N_19033,N_18943,N_18959);
xor U19034 (N_19034,N_18997,N_18950);
nand U19035 (N_19035,N_18948,N_18870);
xor U19036 (N_19036,N_18915,N_18844);
or U19037 (N_19037,N_18855,N_18904);
and U19038 (N_19038,N_18972,N_18832);
xnor U19039 (N_19039,N_18910,N_18807);
xor U19040 (N_19040,N_18902,N_18909);
or U19041 (N_19041,N_18871,N_18907);
xor U19042 (N_19042,N_18964,N_18903);
or U19043 (N_19043,N_18804,N_18825);
or U19044 (N_19044,N_18955,N_18837);
xor U19045 (N_19045,N_18998,N_18800);
nand U19046 (N_19046,N_18879,N_18961);
or U19047 (N_19047,N_18848,N_18979);
xnor U19048 (N_19048,N_18926,N_18803);
or U19049 (N_19049,N_18938,N_18839);
nand U19050 (N_19050,N_18953,N_18805);
and U19051 (N_19051,N_18809,N_18853);
or U19052 (N_19052,N_18927,N_18893);
xnor U19053 (N_19053,N_18963,N_18956);
or U19054 (N_19054,N_18821,N_18872);
xor U19055 (N_19055,N_18808,N_18838);
nor U19056 (N_19056,N_18995,N_18864);
nand U19057 (N_19057,N_18862,N_18868);
xnor U19058 (N_19058,N_18929,N_18932);
or U19059 (N_19059,N_18936,N_18919);
nand U19060 (N_19060,N_18968,N_18920);
xnor U19061 (N_19061,N_18810,N_18957);
nand U19062 (N_19062,N_18885,N_18877);
nand U19063 (N_19063,N_18922,N_18897);
nor U19064 (N_19064,N_18830,N_18928);
xor U19065 (N_19065,N_18983,N_18880);
nor U19066 (N_19066,N_18831,N_18847);
or U19067 (N_19067,N_18882,N_18843);
xnor U19068 (N_19068,N_18852,N_18869);
nor U19069 (N_19069,N_18974,N_18990);
or U19070 (N_19070,N_18981,N_18842);
nand U19071 (N_19071,N_18802,N_18954);
or U19072 (N_19072,N_18894,N_18857);
nor U19073 (N_19073,N_18850,N_18969);
nand U19074 (N_19074,N_18931,N_18978);
xnor U19075 (N_19075,N_18828,N_18874);
nor U19076 (N_19076,N_18881,N_18890);
nor U19077 (N_19077,N_18941,N_18966);
and U19078 (N_19078,N_18818,N_18970);
xnor U19079 (N_19079,N_18951,N_18942);
xnor U19080 (N_19080,N_18944,N_18867);
or U19081 (N_19081,N_18888,N_18822);
xnor U19082 (N_19082,N_18985,N_18939);
or U19083 (N_19083,N_18987,N_18834);
and U19084 (N_19084,N_18815,N_18916);
and U19085 (N_19085,N_18875,N_18973);
xnor U19086 (N_19086,N_18980,N_18946);
and U19087 (N_19087,N_18994,N_18824);
nand U19088 (N_19088,N_18827,N_18816);
and U19089 (N_19089,N_18851,N_18949);
nand U19090 (N_19090,N_18960,N_18854);
or U19091 (N_19091,N_18826,N_18856);
or U19092 (N_19092,N_18934,N_18945);
xnor U19093 (N_19093,N_18991,N_18977);
nand U19094 (N_19094,N_18901,N_18900);
nand U19095 (N_19095,N_18813,N_18835);
and U19096 (N_19096,N_18999,N_18911);
and U19097 (N_19097,N_18814,N_18933);
nor U19098 (N_19098,N_18976,N_18937);
nor U19099 (N_19099,N_18823,N_18836);
nand U19100 (N_19100,N_18839,N_18866);
nand U19101 (N_19101,N_18908,N_18934);
and U19102 (N_19102,N_18956,N_18873);
nor U19103 (N_19103,N_18833,N_18972);
or U19104 (N_19104,N_18971,N_18968);
xor U19105 (N_19105,N_18853,N_18931);
or U19106 (N_19106,N_18860,N_18814);
xnor U19107 (N_19107,N_18860,N_18972);
xnor U19108 (N_19108,N_18951,N_18827);
nor U19109 (N_19109,N_18844,N_18963);
nor U19110 (N_19110,N_18801,N_18991);
and U19111 (N_19111,N_18912,N_18880);
nand U19112 (N_19112,N_18895,N_18890);
nor U19113 (N_19113,N_18819,N_18973);
or U19114 (N_19114,N_18973,N_18920);
or U19115 (N_19115,N_18911,N_18847);
xnor U19116 (N_19116,N_18963,N_18988);
and U19117 (N_19117,N_18863,N_18856);
nor U19118 (N_19118,N_18855,N_18957);
or U19119 (N_19119,N_18918,N_18840);
xor U19120 (N_19120,N_18870,N_18995);
or U19121 (N_19121,N_18851,N_18968);
nor U19122 (N_19122,N_18885,N_18947);
xnor U19123 (N_19123,N_18801,N_18975);
and U19124 (N_19124,N_18876,N_18989);
nand U19125 (N_19125,N_18966,N_18820);
xnor U19126 (N_19126,N_18822,N_18840);
xnor U19127 (N_19127,N_18815,N_18898);
xnor U19128 (N_19128,N_18842,N_18888);
nand U19129 (N_19129,N_18916,N_18926);
and U19130 (N_19130,N_18854,N_18963);
nor U19131 (N_19131,N_18893,N_18967);
or U19132 (N_19132,N_18916,N_18803);
nor U19133 (N_19133,N_18884,N_18861);
or U19134 (N_19134,N_18809,N_18932);
or U19135 (N_19135,N_18936,N_18865);
xor U19136 (N_19136,N_18920,N_18998);
xor U19137 (N_19137,N_18843,N_18946);
nor U19138 (N_19138,N_18808,N_18813);
and U19139 (N_19139,N_18837,N_18942);
and U19140 (N_19140,N_18957,N_18811);
nor U19141 (N_19141,N_18831,N_18825);
nor U19142 (N_19142,N_18919,N_18859);
nor U19143 (N_19143,N_18843,N_18981);
and U19144 (N_19144,N_18951,N_18868);
xnor U19145 (N_19145,N_18802,N_18864);
xor U19146 (N_19146,N_18954,N_18811);
nor U19147 (N_19147,N_18910,N_18893);
nor U19148 (N_19148,N_18975,N_18941);
nor U19149 (N_19149,N_18992,N_18989);
or U19150 (N_19150,N_18961,N_18828);
nor U19151 (N_19151,N_18801,N_18874);
nand U19152 (N_19152,N_18804,N_18968);
xor U19153 (N_19153,N_18940,N_18965);
and U19154 (N_19154,N_18885,N_18931);
nor U19155 (N_19155,N_18997,N_18996);
xor U19156 (N_19156,N_18869,N_18862);
and U19157 (N_19157,N_18843,N_18962);
nand U19158 (N_19158,N_18893,N_18869);
nand U19159 (N_19159,N_18962,N_18997);
xor U19160 (N_19160,N_18987,N_18968);
and U19161 (N_19161,N_18804,N_18983);
xor U19162 (N_19162,N_18932,N_18801);
and U19163 (N_19163,N_18841,N_18936);
and U19164 (N_19164,N_18893,N_18848);
nand U19165 (N_19165,N_18812,N_18857);
nor U19166 (N_19166,N_18863,N_18841);
or U19167 (N_19167,N_18839,N_18990);
and U19168 (N_19168,N_18958,N_18971);
and U19169 (N_19169,N_18843,N_18951);
and U19170 (N_19170,N_18865,N_18843);
xnor U19171 (N_19171,N_18874,N_18863);
nand U19172 (N_19172,N_18926,N_18998);
nand U19173 (N_19173,N_18895,N_18835);
or U19174 (N_19174,N_18929,N_18915);
nand U19175 (N_19175,N_18894,N_18970);
xnor U19176 (N_19176,N_18844,N_18996);
and U19177 (N_19177,N_18880,N_18853);
and U19178 (N_19178,N_18937,N_18814);
xor U19179 (N_19179,N_18888,N_18801);
nor U19180 (N_19180,N_18997,N_18988);
nand U19181 (N_19181,N_18854,N_18953);
xor U19182 (N_19182,N_18952,N_18995);
or U19183 (N_19183,N_18909,N_18943);
and U19184 (N_19184,N_18821,N_18851);
and U19185 (N_19185,N_18887,N_18954);
nor U19186 (N_19186,N_18925,N_18965);
or U19187 (N_19187,N_18914,N_18819);
or U19188 (N_19188,N_18981,N_18913);
nand U19189 (N_19189,N_18820,N_18892);
nor U19190 (N_19190,N_18965,N_18849);
and U19191 (N_19191,N_18884,N_18988);
or U19192 (N_19192,N_18899,N_18837);
or U19193 (N_19193,N_18897,N_18830);
nand U19194 (N_19194,N_18977,N_18939);
xor U19195 (N_19195,N_18926,N_18855);
or U19196 (N_19196,N_18914,N_18880);
nor U19197 (N_19197,N_18954,N_18977);
nor U19198 (N_19198,N_18985,N_18802);
or U19199 (N_19199,N_18864,N_18958);
xor U19200 (N_19200,N_19070,N_19078);
xor U19201 (N_19201,N_19173,N_19042);
xnor U19202 (N_19202,N_19037,N_19016);
nand U19203 (N_19203,N_19030,N_19004);
and U19204 (N_19204,N_19179,N_19147);
nand U19205 (N_19205,N_19154,N_19089);
nor U19206 (N_19206,N_19056,N_19075);
and U19207 (N_19207,N_19000,N_19140);
and U19208 (N_19208,N_19033,N_19093);
or U19209 (N_19209,N_19097,N_19192);
or U19210 (N_19210,N_19131,N_19189);
xor U19211 (N_19211,N_19003,N_19157);
or U19212 (N_19212,N_19086,N_19048);
nor U19213 (N_19213,N_19074,N_19105);
nand U19214 (N_19214,N_19170,N_19072);
and U19215 (N_19215,N_19191,N_19190);
and U19216 (N_19216,N_19178,N_19138);
nand U19217 (N_19217,N_19002,N_19038);
nand U19218 (N_19218,N_19025,N_19186);
and U19219 (N_19219,N_19009,N_19064);
and U19220 (N_19220,N_19013,N_19020);
and U19221 (N_19221,N_19068,N_19132);
nand U19222 (N_19222,N_19195,N_19171);
or U19223 (N_19223,N_19159,N_19017);
nand U19224 (N_19224,N_19098,N_19183);
nand U19225 (N_19225,N_19092,N_19036);
and U19226 (N_19226,N_19001,N_19032);
xnor U19227 (N_19227,N_19120,N_19180);
or U19228 (N_19228,N_19166,N_19160);
xor U19229 (N_19229,N_19175,N_19015);
nor U19230 (N_19230,N_19126,N_19109);
and U19231 (N_19231,N_19145,N_19077);
and U19232 (N_19232,N_19134,N_19148);
and U19233 (N_19233,N_19144,N_19123);
nand U19234 (N_19234,N_19185,N_19081);
nand U19235 (N_19235,N_19018,N_19057);
or U19236 (N_19236,N_19193,N_19102);
or U19237 (N_19237,N_19150,N_19096);
xnor U19238 (N_19238,N_19167,N_19153);
and U19239 (N_19239,N_19127,N_19165);
or U19240 (N_19240,N_19113,N_19034);
nor U19241 (N_19241,N_19080,N_19114);
nand U19242 (N_19242,N_19043,N_19040);
nand U19243 (N_19243,N_19100,N_19168);
xor U19244 (N_19244,N_19091,N_19039);
or U19245 (N_19245,N_19006,N_19106);
or U19246 (N_19246,N_19061,N_19054);
xor U19247 (N_19247,N_19047,N_19196);
xnor U19248 (N_19248,N_19095,N_19158);
or U19249 (N_19249,N_19076,N_19130);
and U19250 (N_19250,N_19176,N_19103);
xor U19251 (N_19251,N_19059,N_19125);
xor U19252 (N_19252,N_19062,N_19199);
xor U19253 (N_19253,N_19162,N_19188);
or U19254 (N_19254,N_19021,N_19084);
xnor U19255 (N_19255,N_19045,N_19065);
nor U19256 (N_19256,N_19137,N_19060);
nor U19257 (N_19257,N_19029,N_19161);
xor U19258 (N_19258,N_19046,N_19022);
nand U19259 (N_19259,N_19151,N_19141);
or U19260 (N_19260,N_19149,N_19010);
and U19261 (N_19261,N_19012,N_19142);
and U19262 (N_19262,N_19146,N_19110);
nand U19263 (N_19263,N_19182,N_19049);
or U19264 (N_19264,N_19116,N_19101);
nor U19265 (N_19265,N_19027,N_19128);
and U19266 (N_19266,N_19079,N_19031);
xor U19267 (N_19267,N_19108,N_19051);
nor U19268 (N_19268,N_19023,N_19088);
xnor U19269 (N_19269,N_19169,N_19053);
nand U19270 (N_19270,N_19014,N_19111);
xnor U19271 (N_19271,N_19024,N_19044);
nand U19272 (N_19272,N_19198,N_19194);
or U19273 (N_19273,N_19099,N_19115);
or U19274 (N_19274,N_19026,N_19163);
nor U19275 (N_19275,N_19011,N_19124);
nand U19276 (N_19276,N_19041,N_19087);
nand U19277 (N_19277,N_19143,N_19155);
nand U19278 (N_19278,N_19139,N_19117);
and U19279 (N_19279,N_19058,N_19063);
and U19280 (N_19280,N_19181,N_19107);
or U19281 (N_19281,N_19067,N_19119);
nand U19282 (N_19282,N_19028,N_19094);
or U19283 (N_19283,N_19069,N_19055);
nor U19284 (N_19284,N_19112,N_19066);
nand U19285 (N_19285,N_19085,N_19083);
or U19286 (N_19286,N_19007,N_19122);
nand U19287 (N_19287,N_19118,N_19050);
xnor U19288 (N_19288,N_19035,N_19156);
and U19289 (N_19289,N_19052,N_19129);
nand U19290 (N_19290,N_19152,N_19136);
and U19291 (N_19291,N_19071,N_19174);
nor U19292 (N_19292,N_19135,N_19184);
nand U19293 (N_19293,N_19104,N_19187);
xnor U19294 (N_19294,N_19197,N_19073);
nand U19295 (N_19295,N_19121,N_19133);
or U19296 (N_19296,N_19172,N_19177);
nand U19297 (N_19297,N_19090,N_19082);
and U19298 (N_19298,N_19019,N_19008);
xnor U19299 (N_19299,N_19164,N_19005);
xor U19300 (N_19300,N_19100,N_19009);
or U19301 (N_19301,N_19131,N_19075);
and U19302 (N_19302,N_19137,N_19158);
xor U19303 (N_19303,N_19042,N_19192);
or U19304 (N_19304,N_19136,N_19133);
xor U19305 (N_19305,N_19004,N_19079);
or U19306 (N_19306,N_19092,N_19014);
nand U19307 (N_19307,N_19072,N_19050);
nor U19308 (N_19308,N_19126,N_19162);
and U19309 (N_19309,N_19061,N_19166);
and U19310 (N_19310,N_19082,N_19135);
xnor U19311 (N_19311,N_19176,N_19057);
nor U19312 (N_19312,N_19191,N_19123);
or U19313 (N_19313,N_19054,N_19052);
and U19314 (N_19314,N_19098,N_19177);
xnor U19315 (N_19315,N_19046,N_19115);
nor U19316 (N_19316,N_19101,N_19066);
or U19317 (N_19317,N_19120,N_19065);
xnor U19318 (N_19318,N_19167,N_19020);
nand U19319 (N_19319,N_19028,N_19035);
or U19320 (N_19320,N_19188,N_19046);
or U19321 (N_19321,N_19087,N_19106);
xnor U19322 (N_19322,N_19179,N_19046);
or U19323 (N_19323,N_19014,N_19139);
and U19324 (N_19324,N_19003,N_19014);
and U19325 (N_19325,N_19171,N_19091);
nor U19326 (N_19326,N_19119,N_19193);
xor U19327 (N_19327,N_19184,N_19041);
or U19328 (N_19328,N_19160,N_19079);
xnor U19329 (N_19329,N_19052,N_19114);
and U19330 (N_19330,N_19032,N_19023);
and U19331 (N_19331,N_19115,N_19132);
xor U19332 (N_19332,N_19087,N_19057);
and U19333 (N_19333,N_19167,N_19189);
nor U19334 (N_19334,N_19055,N_19071);
and U19335 (N_19335,N_19014,N_19084);
nand U19336 (N_19336,N_19130,N_19165);
or U19337 (N_19337,N_19081,N_19173);
and U19338 (N_19338,N_19142,N_19091);
nor U19339 (N_19339,N_19167,N_19152);
nor U19340 (N_19340,N_19023,N_19093);
and U19341 (N_19341,N_19112,N_19157);
and U19342 (N_19342,N_19031,N_19066);
and U19343 (N_19343,N_19033,N_19021);
nand U19344 (N_19344,N_19038,N_19145);
or U19345 (N_19345,N_19035,N_19072);
xor U19346 (N_19346,N_19151,N_19191);
nor U19347 (N_19347,N_19132,N_19050);
nor U19348 (N_19348,N_19019,N_19043);
nor U19349 (N_19349,N_19009,N_19030);
xnor U19350 (N_19350,N_19085,N_19023);
and U19351 (N_19351,N_19067,N_19009);
and U19352 (N_19352,N_19013,N_19087);
xor U19353 (N_19353,N_19124,N_19182);
xnor U19354 (N_19354,N_19054,N_19149);
or U19355 (N_19355,N_19047,N_19189);
xnor U19356 (N_19356,N_19159,N_19108);
and U19357 (N_19357,N_19078,N_19107);
xor U19358 (N_19358,N_19019,N_19121);
xor U19359 (N_19359,N_19112,N_19063);
nor U19360 (N_19360,N_19034,N_19089);
nand U19361 (N_19361,N_19042,N_19097);
nor U19362 (N_19362,N_19026,N_19158);
nand U19363 (N_19363,N_19125,N_19001);
or U19364 (N_19364,N_19031,N_19043);
nor U19365 (N_19365,N_19024,N_19074);
nor U19366 (N_19366,N_19123,N_19035);
or U19367 (N_19367,N_19090,N_19043);
xor U19368 (N_19368,N_19100,N_19092);
and U19369 (N_19369,N_19146,N_19095);
and U19370 (N_19370,N_19129,N_19002);
or U19371 (N_19371,N_19184,N_19192);
nand U19372 (N_19372,N_19146,N_19178);
nor U19373 (N_19373,N_19194,N_19129);
xor U19374 (N_19374,N_19121,N_19111);
and U19375 (N_19375,N_19165,N_19066);
nand U19376 (N_19376,N_19083,N_19187);
and U19377 (N_19377,N_19183,N_19168);
or U19378 (N_19378,N_19001,N_19184);
xnor U19379 (N_19379,N_19174,N_19170);
nand U19380 (N_19380,N_19020,N_19030);
or U19381 (N_19381,N_19077,N_19175);
or U19382 (N_19382,N_19115,N_19035);
or U19383 (N_19383,N_19068,N_19085);
xnor U19384 (N_19384,N_19111,N_19163);
and U19385 (N_19385,N_19093,N_19178);
xor U19386 (N_19386,N_19182,N_19183);
nand U19387 (N_19387,N_19129,N_19010);
or U19388 (N_19388,N_19105,N_19153);
and U19389 (N_19389,N_19047,N_19192);
xor U19390 (N_19390,N_19120,N_19010);
nand U19391 (N_19391,N_19082,N_19145);
or U19392 (N_19392,N_19018,N_19023);
or U19393 (N_19393,N_19138,N_19129);
nand U19394 (N_19394,N_19038,N_19129);
and U19395 (N_19395,N_19091,N_19092);
or U19396 (N_19396,N_19129,N_19088);
xnor U19397 (N_19397,N_19068,N_19106);
and U19398 (N_19398,N_19187,N_19088);
nand U19399 (N_19399,N_19014,N_19048);
and U19400 (N_19400,N_19356,N_19374);
nand U19401 (N_19401,N_19379,N_19278);
and U19402 (N_19402,N_19389,N_19248);
xnor U19403 (N_19403,N_19375,N_19265);
nand U19404 (N_19404,N_19376,N_19299);
xor U19405 (N_19405,N_19233,N_19357);
nand U19406 (N_19406,N_19235,N_19322);
xnor U19407 (N_19407,N_19334,N_19259);
or U19408 (N_19408,N_19347,N_19254);
and U19409 (N_19409,N_19345,N_19384);
and U19410 (N_19410,N_19243,N_19213);
nand U19411 (N_19411,N_19367,N_19263);
and U19412 (N_19412,N_19242,N_19330);
nand U19413 (N_19413,N_19383,N_19274);
nor U19414 (N_19414,N_19360,N_19369);
or U19415 (N_19415,N_19268,N_19361);
and U19416 (N_19416,N_19364,N_19277);
nand U19417 (N_19417,N_19349,N_19294);
or U19418 (N_19418,N_19339,N_19210);
nor U19419 (N_19419,N_19332,N_19276);
and U19420 (N_19420,N_19288,N_19314);
nand U19421 (N_19421,N_19396,N_19269);
nor U19422 (N_19422,N_19208,N_19273);
xor U19423 (N_19423,N_19366,N_19318);
xnor U19424 (N_19424,N_19282,N_19222);
and U19425 (N_19425,N_19267,N_19342);
and U19426 (N_19426,N_19386,N_19310);
xor U19427 (N_19427,N_19202,N_19230);
xnor U19428 (N_19428,N_19315,N_19225);
nor U19429 (N_19429,N_19355,N_19283);
xnor U19430 (N_19430,N_19304,N_19371);
nand U19431 (N_19431,N_19341,N_19284);
nand U19432 (N_19432,N_19394,N_19296);
xor U19433 (N_19433,N_19214,N_19290);
and U19434 (N_19434,N_19239,N_19316);
and U19435 (N_19435,N_19253,N_19348);
xnor U19436 (N_19436,N_19237,N_19390);
nand U19437 (N_19437,N_19399,N_19325);
nor U19438 (N_19438,N_19302,N_19264);
or U19439 (N_19439,N_19311,N_19324);
nand U19440 (N_19440,N_19397,N_19216);
or U19441 (N_19441,N_19350,N_19319);
nand U19442 (N_19442,N_19368,N_19280);
nand U19443 (N_19443,N_19321,N_19295);
nor U19444 (N_19444,N_19209,N_19380);
xnor U19445 (N_19445,N_19307,N_19305);
xor U19446 (N_19446,N_19309,N_19228);
nor U19447 (N_19447,N_19272,N_19312);
and U19448 (N_19448,N_19336,N_19218);
and U19449 (N_19449,N_19281,N_19252);
or U19450 (N_19450,N_19303,N_19234);
nor U19451 (N_19451,N_19232,N_19338);
nand U19452 (N_19452,N_19240,N_19344);
and U19453 (N_19453,N_19354,N_19378);
nand U19454 (N_19454,N_19352,N_19212);
nand U19455 (N_19455,N_19298,N_19219);
xnor U19456 (N_19456,N_19293,N_19246);
nor U19457 (N_19457,N_19377,N_19285);
or U19458 (N_19458,N_19247,N_19392);
nand U19459 (N_19459,N_19211,N_19365);
and U19460 (N_19460,N_19382,N_19335);
nor U19461 (N_19461,N_19223,N_19203);
and U19462 (N_19462,N_19244,N_19358);
nor U19463 (N_19463,N_19286,N_19224);
or U19464 (N_19464,N_19217,N_19275);
and U19465 (N_19465,N_19245,N_19226);
xor U19466 (N_19466,N_19291,N_19370);
nand U19467 (N_19467,N_19231,N_19262);
or U19468 (N_19468,N_19340,N_19255);
and U19469 (N_19469,N_19346,N_19221);
nor U19470 (N_19470,N_19270,N_19317);
or U19471 (N_19471,N_19258,N_19393);
nand U19472 (N_19472,N_19292,N_19205);
or U19473 (N_19473,N_19359,N_19289);
nor U19474 (N_19474,N_19200,N_19353);
or U19475 (N_19475,N_19328,N_19320);
nor U19476 (N_19476,N_19398,N_19388);
and U19477 (N_19477,N_19207,N_19206);
nor U19478 (N_19478,N_19363,N_19251);
nor U19479 (N_19479,N_19327,N_19215);
nand U19480 (N_19480,N_19227,N_19229);
nor U19481 (N_19481,N_19313,N_19204);
xnor U19482 (N_19482,N_19381,N_19297);
or U19483 (N_19483,N_19257,N_19266);
and U19484 (N_19484,N_19261,N_19271);
and U19485 (N_19485,N_19351,N_19238);
or U19486 (N_19486,N_19337,N_19331);
nor U19487 (N_19487,N_19250,N_19326);
nand U19488 (N_19488,N_19329,N_19260);
or U19489 (N_19489,N_19241,N_19333);
or U19490 (N_19490,N_19395,N_19201);
xnor U19491 (N_19491,N_19343,N_19256);
nor U19492 (N_19492,N_19387,N_19373);
nor U19493 (N_19493,N_19300,N_19287);
and U19494 (N_19494,N_19391,N_19308);
nand U19495 (N_19495,N_19279,N_19236);
and U19496 (N_19496,N_19372,N_19301);
or U19497 (N_19497,N_19385,N_19306);
nand U19498 (N_19498,N_19249,N_19362);
xnor U19499 (N_19499,N_19323,N_19220);
xnor U19500 (N_19500,N_19260,N_19299);
xor U19501 (N_19501,N_19346,N_19353);
xor U19502 (N_19502,N_19390,N_19224);
nor U19503 (N_19503,N_19214,N_19267);
xnor U19504 (N_19504,N_19361,N_19284);
or U19505 (N_19505,N_19230,N_19357);
or U19506 (N_19506,N_19290,N_19329);
and U19507 (N_19507,N_19217,N_19220);
xnor U19508 (N_19508,N_19395,N_19247);
nor U19509 (N_19509,N_19239,N_19254);
nor U19510 (N_19510,N_19388,N_19307);
xnor U19511 (N_19511,N_19379,N_19213);
or U19512 (N_19512,N_19381,N_19369);
nor U19513 (N_19513,N_19271,N_19217);
nand U19514 (N_19514,N_19253,N_19269);
nand U19515 (N_19515,N_19288,N_19296);
xor U19516 (N_19516,N_19292,N_19320);
or U19517 (N_19517,N_19292,N_19291);
and U19518 (N_19518,N_19345,N_19360);
nor U19519 (N_19519,N_19268,N_19369);
or U19520 (N_19520,N_19251,N_19220);
nor U19521 (N_19521,N_19337,N_19213);
nor U19522 (N_19522,N_19206,N_19264);
nor U19523 (N_19523,N_19376,N_19303);
xor U19524 (N_19524,N_19388,N_19369);
nand U19525 (N_19525,N_19394,N_19206);
and U19526 (N_19526,N_19205,N_19250);
and U19527 (N_19527,N_19250,N_19261);
or U19528 (N_19528,N_19295,N_19344);
nor U19529 (N_19529,N_19334,N_19389);
nand U19530 (N_19530,N_19393,N_19371);
xor U19531 (N_19531,N_19378,N_19363);
or U19532 (N_19532,N_19248,N_19289);
or U19533 (N_19533,N_19257,N_19224);
and U19534 (N_19534,N_19290,N_19211);
xor U19535 (N_19535,N_19396,N_19227);
nor U19536 (N_19536,N_19220,N_19212);
nor U19537 (N_19537,N_19261,N_19282);
and U19538 (N_19538,N_19261,N_19332);
and U19539 (N_19539,N_19299,N_19347);
xor U19540 (N_19540,N_19322,N_19275);
nand U19541 (N_19541,N_19354,N_19247);
xnor U19542 (N_19542,N_19296,N_19270);
and U19543 (N_19543,N_19244,N_19213);
and U19544 (N_19544,N_19237,N_19394);
and U19545 (N_19545,N_19324,N_19221);
xnor U19546 (N_19546,N_19214,N_19255);
xnor U19547 (N_19547,N_19235,N_19284);
nand U19548 (N_19548,N_19373,N_19222);
nor U19549 (N_19549,N_19299,N_19385);
and U19550 (N_19550,N_19231,N_19344);
nand U19551 (N_19551,N_19248,N_19303);
nand U19552 (N_19552,N_19286,N_19230);
nand U19553 (N_19553,N_19308,N_19333);
and U19554 (N_19554,N_19274,N_19237);
and U19555 (N_19555,N_19309,N_19301);
xnor U19556 (N_19556,N_19318,N_19273);
xor U19557 (N_19557,N_19230,N_19211);
nor U19558 (N_19558,N_19358,N_19383);
or U19559 (N_19559,N_19253,N_19212);
xnor U19560 (N_19560,N_19361,N_19350);
or U19561 (N_19561,N_19329,N_19279);
and U19562 (N_19562,N_19322,N_19261);
nand U19563 (N_19563,N_19341,N_19229);
xnor U19564 (N_19564,N_19372,N_19338);
and U19565 (N_19565,N_19260,N_19376);
or U19566 (N_19566,N_19296,N_19385);
nand U19567 (N_19567,N_19337,N_19382);
nand U19568 (N_19568,N_19349,N_19299);
nand U19569 (N_19569,N_19280,N_19373);
nand U19570 (N_19570,N_19373,N_19377);
xor U19571 (N_19571,N_19277,N_19229);
or U19572 (N_19572,N_19219,N_19317);
and U19573 (N_19573,N_19305,N_19266);
nand U19574 (N_19574,N_19332,N_19262);
or U19575 (N_19575,N_19368,N_19215);
nor U19576 (N_19576,N_19201,N_19397);
and U19577 (N_19577,N_19233,N_19211);
and U19578 (N_19578,N_19314,N_19323);
nor U19579 (N_19579,N_19334,N_19344);
nor U19580 (N_19580,N_19301,N_19202);
and U19581 (N_19581,N_19324,N_19265);
nor U19582 (N_19582,N_19269,N_19259);
nand U19583 (N_19583,N_19289,N_19277);
nand U19584 (N_19584,N_19360,N_19269);
nor U19585 (N_19585,N_19370,N_19279);
and U19586 (N_19586,N_19256,N_19302);
nand U19587 (N_19587,N_19208,N_19337);
and U19588 (N_19588,N_19277,N_19290);
nand U19589 (N_19589,N_19359,N_19203);
or U19590 (N_19590,N_19237,N_19245);
nor U19591 (N_19591,N_19224,N_19328);
nor U19592 (N_19592,N_19262,N_19275);
or U19593 (N_19593,N_19329,N_19314);
or U19594 (N_19594,N_19201,N_19304);
nand U19595 (N_19595,N_19361,N_19349);
xnor U19596 (N_19596,N_19312,N_19313);
nor U19597 (N_19597,N_19375,N_19293);
nand U19598 (N_19598,N_19251,N_19267);
or U19599 (N_19599,N_19251,N_19223);
or U19600 (N_19600,N_19498,N_19415);
or U19601 (N_19601,N_19469,N_19508);
and U19602 (N_19602,N_19449,N_19569);
nand U19603 (N_19603,N_19473,N_19542);
nor U19604 (N_19604,N_19475,N_19464);
and U19605 (N_19605,N_19533,N_19543);
nand U19606 (N_19606,N_19593,N_19400);
nand U19607 (N_19607,N_19575,N_19579);
xor U19608 (N_19608,N_19513,N_19439);
nor U19609 (N_19609,N_19490,N_19483);
or U19610 (N_19610,N_19560,N_19445);
and U19611 (N_19611,N_19417,N_19590);
and U19612 (N_19612,N_19516,N_19520);
and U19613 (N_19613,N_19489,N_19450);
nand U19614 (N_19614,N_19536,N_19587);
or U19615 (N_19615,N_19567,N_19467);
or U19616 (N_19616,N_19535,N_19563);
xor U19617 (N_19617,N_19544,N_19444);
nor U19618 (N_19618,N_19554,N_19411);
or U19619 (N_19619,N_19452,N_19486);
and U19620 (N_19620,N_19453,N_19438);
nor U19621 (N_19621,N_19568,N_19495);
nand U19622 (N_19622,N_19426,N_19523);
nand U19623 (N_19623,N_19423,N_19455);
and U19624 (N_19624,N_19401,N_19451);
nand U19625 (N_19625,N_19592,N_19532);
nor U19626 (N_19626,N_19539,N_19570);
and U19627 (N_19627,N_19443,N_19447);
nand U19628 (N_19628,N_19463,N_19441);
and U19629 (N_19629,N_19431,N_19515);
nand U19630 (N_19630,N_19484,N_19429);
nand U19631 (N_19631,N_19472,N_19573);
and U19632 (N_19632,N_19476,N_19459);
nor U19633 (N_19633,N_19514,N_19446);
nor U19634 (N_19634,N_19525,N_19481);
nor U19635 (N_19635,N_19500,N_19497);
or U19636 (N_19636,N_19440,N_19499);
xnor U19637 (N_19637,N_19419,N_19565);
xor U19638 (N_19638,N_19437,N_19583);
nand U19639 (N_19639,N_19502,N_19482);
and U19640 (N_19640,N_19537,N_19588);
nand U19641 (N_19641,N_19404,N_19549);
nand U19642 (N_19642,N_19466,N_19433);
nor U19643 (N_19643,N_19510,N_19557);
nor U19644 (N_19644,N_19435,N_19501);
nor U19645 (N_19645,N_19561,N_19555);
xor U19646 (N_19646,N_19477,N_19442);
and U19647 (N_19647,N_19492,N_19408);
or U19648 (N_19648,N_19558,N_19491);
nand U19649 (N_19649,N_19518,N_19522);
and U19650 (N_19650,N_19405,N_19530);
xor U19651 (N_19651,N_19553,N_19572);
or U19652 (N_19652,N_19428,N_19454);
xnor U19653 (N_19653,N_19578,N_19504);
and U19654 (N_19654,N_19599,N_19434);
xnor U19655 (N_19655,N_19521,N_19527);
xor U19656 (N_19656,N_19550,N_19503);
nor U19657 (N_19657,N_19571,N_19487);
or U19658 (N_19658,N_19585,N_19529);
or U19659 (N_19659,N_19511,N_19595);
and U19660 (N_19660,N_19406,N_19403);
or U19661 (N_19661,N_19574,N_19540);
and U19662 (N_19662,N_19551,N_19448);
and U19663 (N_19663,N_19432,N_19460);
and U19664 (N_19664,N_19556,N_19421);
nor U19665 (N_19665,N_19598,N_19509);
xnor U19666 (N_19666,N_19422,N_19581);
or U19667 (N_19667,N_19418,N_19468);
nand U19668 (N_19668,N_19416,N_19409);
xnor U19669 (N_19669,N_19538,N_19505);
nand U19670 (N_19670,N_19480,N_19412);
xnor U19671 (N_19671,N_19506,N_19414);
nand U19672 (N_19672,N_19494,N_19496);
and U19673 (N_19673,N_19479,N_19596);
or U19674 (N_19674,N_19456,N_19564);
or U19675 (N_19675,N_19512,N_19470);
xor U19676 (N_19676,N_19559,N_19430);
nor U19677 (N_19677,N_19471,N_19407);
nand U19678 (N_19678,N_19425,N_19474);
nand U19679 (N_19679,N_19548,N_19526);
xnor U19680 (N_19680,N_19517,N_19584);
nand U19681 (N_19681,N_19534,N_19589);
nor U19682 (N_19682,N_19586,N_19528);
and U19683 (N_19683,N_19420,N_19580);
xnor U19684 (N_19684,N_19410,N_19597);
nand U19685 (N_19685,N_19582,N_19546);
xnor U19686 (N_19686,N_19465,N_19576);
xnor U19687 (N_19687,N_19594,N_19402);
nand U19688 (N_19688,N_19488,N_19562);
and U19689 (N_19689,N_19552,N_19424);
nand U19690 (N_19690,N_19577,N_19493);
xor U19691 (N_19691,N_19545,N_19413);
xor U19692 (N_19692,N_19478,N_19531);
nor U19693 (N_19693,N_19507,N_19457);
and U19694 (N_19694,N_19524,N_19436);
xor U19695 (N_19695,N_19519,N_19566);
and U19696 (N_19696,N_19458,N_19462);
xor U19697 (N_19697,N_19591,N_19461);
nand U19698 (N_19698,N_19547,N_19541);
and U19699 (N_19699,N_19427,N_19485);
or U19700 (N_19700,N_19494,N_19547);
nand U19701 (N_19701,N_19401,N_19509);
xor U19702 (N_19702,N_19597,N_19598);
or U19703 (N_19703,N_19435,N_19452);
and U19704 (N_19704,N_19553,N_19581);
xnor U19705 (N_19705,N_19466,N_19452);
or U19706 (N_19706,N_19429,N_19461);
xnor U19707 (N_19707,N_19577,N_19428);
and U19708 (N_19708,N_19553,N_19506);
nor U19709 (N_19709,N_19524,N_19552);
and U19710 (N_19710,N_19547,N_19596);
and U19711 (N_19711,N_19546,N_19586);
or U19712 (N_19712,N_19459,N_19575);
xor U19713 (N_19713,N_19556,N_19580);
nand U19714 (N_19714,N_19444,N_19439);
and U19715 (N_19715,N_19428,N_19557);
xor U19716 (N_19716,N_19519,N_19573);
nand U19717 (N_19717,N_19586,N_19490);
nor U19718 (N_19718,N_19448,N_19463);
and U19719 (N_19719,N_19470,N_19484);
and U19720 (N_19720,N_19534,N_19469);
and U19721 (N_19721,N_19507,N_19523);
nand U19722 (N_19722,N_19527,N_19590);
xnor U19723 (N_19723,N_19406,N_19480);
nand U19724 (N_19724,N_19560,N_19557);
xnor U19725 (N_19725,N_19403,N_19474);
nor U19726 (N_19726,N_19403,N_19581);
nand U19727 (N_19727,N_19428,N_19596);
and U19728 (N_19728,N_19415,N_19584);
nand U19729 (N_19729,N_19483,N_19449);
nor U19730 (N_19730,N_19533,N_19513);
nor U19731 (N_19731,N_19554,N_19497);
and U19732 (N_19732,N_19565,N_19543);
xor U19733 (N_19733,N_19413,N_19505);
and U19734 (N_19734,N_19429,N_19590);
nand U19735 (N_19735,N_19576,N_19478);
nand U19736 (N_19736,N_19546,N_19555);
or U19737 (N_19737,N_19501,N_19553);
and U19738 (N_19738,N_19401,N_19498);
and U19739 (N_19739,N_19573,N_19442);
nor U19740 (N_19740,N_19440,N_19515);
xnor U19741 (N_19741,N_19457,N_19532);
xor U19742 (N_19742,N_19520,N_19554);
xnor U19743 (N_19743,N_19445,N_19495);
nand U19744 (N_19744,N_19588,N_19565);
nand U19745 (N_19745,N_19564,N_19560);
and U19746 (N_19746,N_19510,N_19582);
nor U19747 (N_19747,N_19598,N_19584);
nand U19748 (N_19748,N_19492,N_19546);
nand U19749 (N_19749,N_19465,N_19584);
xnor U19750 (N_19750,N_19497,N_19528);
nand U19751 (N_19751,N_19509,N_19499);
or U19752 (N_19752,N_19501,N_19434);
and U19753 (N_19753,N_19520,N_19413);
xnor U19754 (N_19754,N_19558,N_19506);
nor U19755 (N_19755,N_19417,N_19478);
and U19756 (N_19756,N_19490,N_19466);
or U19757 (N_19757,N_19488,N_19416);
nor U19758 (N_19758,N_19516,N_19513);
nand U19759 (N_19759,N_19591,N_19450);
xnor U19760 (N_19760,N_19570,N_19401);
nor U19761 (N_19761,N_19444,N_19407);
or U19762 (N_19762,N_19416,N_19510);
and U19763 (N_19763,N_19569,N_19495);
and U19764 (N_19764,N_19523,N_19441);
nor U19765 (N_19765,N_19589,N_19488);
nor U19766 (N_19766,N_19401,N_19454);
and U19767 (N_19767,N_19490,N_19599);
and U19768 (N_19768,N_19413,N_19578);
nand U19769 (N_19769,N_19437,N_19573);
or U19770 (N_19770,N_19453,N_19467);
nand U19771 (N_19771,N_19468,N_19476);
or U19772 (N_19772,N_19482,N_19407);
and U19773 (N_19773,N_19517,N_19554);
xor U19774 (N_19774,N_19487,N_19588);
nor U19775 (N_19775,N_19476,N_19588);
and U19776 (N_19776,N_19461,N_19438);
and U19777 (N_19777,N_19593,N_19452);
or U19778 (N_19778,N_19548,N_19591);
or U19779 (N_19779,N_19418,N_19462);
and U19780 (N_19780,N_19581,N_19419);
or U19781 (N_19781,N_19581,N_19599);
nand U19782 (N_19782,N_19421,N_19460);
and U19783 (N_19783,N_19411,N_19454);
xnor U19784 (N_19784,N_19497,N_19571);
nor U19785 (N_19785,N_19450,N_19530);
and U19786 (N_19786,N_19417,N_19486);
or U19787 (N_19787,N_19472,N_19445);
nor U19788 (N_19788,N_19556,N_19465);
xor U19789 (N_19789,N_19430,N_19544);
nand U19790 (N_19790,N_19434,N_19549);
nor U19791 (N_19791,N_19549,N_19553);
xnor U19792 (N_19792,N_19471,N_19478);
and U19793 (N_19793,N_19437,N_19519);
nor U19794 (N_19794,N_19505,N_19422);
xnor U19795 (N_19795,N_19442,N_19549);
and U19796 (N_19796,N_19506,N_19420);
nor U19797 (N_19797,N_19435,N_19411);
xor U19798 (N_19798,N_19517,N_19470);
nand U19799 (N_19799,N_19481,N_19588);
nor U19800 (N_19800,N_19693,N_19651);
nand U19801 (N_19801,N_19610,N_19712);
nor U19802 (N_19802,N_19751,N_19696);
nand U19803 (N_19803,N_19617,N_19749);
nand U19804 (N_19804,N_19704,N_19645);
nand U19805 (N_19805,N_19762,N_19646);
and U19806 (N_19806,N_19765,N_19622);
or U19807 (N_19807,N_19654,N_19690);
nand U19808 (N_19808,N_19675,N_19672);
xnor U19809 (N_19809,N_19640,N_19699);
or U19810 (N_19810,N_19630,N_19609);
xnor U19811 (N_19811,N_19717,N_19670);
nand U19812 (N_19812,N_19782,N_19629);
nor U19813 (N_19813,N_19603,N_19626);
nor U19814 (N_19814,N_19758,N_19618);
xnor U19815 (N_19815,N_19601,N_19748);
and U19816 (N_19816,N_19715,N_19708);
or U19817 (N_19817,N_19647,N_19679);
nor U19818 (N_19818,N_19607,N_19616);
or U19819 (N_19819,N_19697,N_19657);
nor U19820 (N_19820,N_19705,N_19784);
xor U19821 (N_19821,N_19727,N_19783);
or U19822 (N_19822,N_19786,N_19694);
nor U19823 (N_19823,N_19759,N_19706);
or U19824 (N_19824,N_19606,N_19678);
or U19825 (N_19825,N_19722,N_19775);
nand U19826 (N_19826,N_19650,N_19625);
xor U19827 (N_19827,N_19633,N_19767);
xor U19828 (N_19828,N_19683,N_19684);
nand U19829 (N_19829,N_19702,N_19663);
xor U19830 (N_19830,N_19720,N_19602);
nand U19831 (N_19831,N_19638,N_19725);
or U19832 (N_19832,N_19795,N_19777);
and U19833 (N_19833,N_19723,N_19792);
xor U19834 (N_19834,N_19692,N_19770);
xor U19835 (N_19835,N_19756,N_19773);
nor U19836 (N_19836,N_19644,N_19781);
nand U19837 (N_19837,N_19667,N_19774);
nand U19838 (N_19838,N_19769,N_19652);
xnor U19839 (N_19839,N_19760,N_19750);
nand U19840 (N_19840,N_19798,N_19674);
or U19841 (N_19841,N_19730,N_19639);
and U19842 (N_19842,N_19619,N_19662);
nor U19843 (N_19843,N_19738,N_19707);
and U19844 (N_19844,N_19643,N_19732);
nor U19845 (N_19845,N_19728,N_19649);
nor U19846 (N_19846,N_19666,N_19735);
xor U19847 (N_19847,N_19778,N_19772);
or U19848 (N_19848,N_19685,N_19604);
nand U19849 (N_19849,N_19658,N_19632);
nor U19850 (N_19850,N_19620,N_19641);
nor U19851 (N_19851,N_19761,N_19731);
nand U19852 (N_19852,N_19655,N_19710);
nand U19853 (N_19853,N_19743,N_19613);
and U19854 (N_19854,N_19789,N_19754);
xnor U19855 (N_19855,N_19611,N_19796);
and U19856 (N_19856,N_19739,N_19600);
and U19857 (N_19857,N_19745,N_19714);
and U19858 (N_19858,N_19788,N_19648);
and U19859 (N_19859,N_19768,N_19660);
nor U19860 (N_19860,N_19793,N_19744);
nor U19861 (N_19861,N_19713,N_19682);
and U19862 (N_19862,N_19680,N_19612);
or U19863 (N_19863,N_19665,N_19605);
xnor U19864 (N_19864,N_19716,N_19724);
and U19865 (N_19865,N_19791,N_19636);
nand U19866 (N_19866,N_19709,N_19623);
nor U19867 (N_19867,N_19780,N_19790);
and U19868 (N_19868,N_19741,N_19721);
nor U19869 (N_19869,N_19642,N_19676);
nand U19870 (N_19870,N_19747,N_19753);
and U19871 (N_19871,N_19763,N_19635);
xnor U19872 (N_19872,N_19797,N_19664);
and U19873 (N_19873,N_19737,N_19615);
nand U19874 (N_19874,N_19673,N_19746);
nor U19875 (N_19875,N_19757,N_19637);
xnor U19876 (N_19876,N_19718,N_19701);
or U19877 (N_19877,N_19733,N_19627);
nand U19878 (N_19878,N_19653,N_19688);
nor U19879 (N_19879,N_19711,N_19698);
and U19880 (N_19880,N_19669,N_19785);
nand U19881 (N_19881,N_19719,N_19787);
and U19882 (N_19882,N_19755,N_19668);
and U19883 (N_19883,N_19779,N_19621);
and U19884 (N_19884,N_19729,N_19736);
and U19885 (N_19885,N_19700,N_19799);
nor U19886 (N_19886,N_19687,N_19776);
or U19887 (N_19887,N_19764,N_19771);
nand U19888 (N_19888,N_19624,N_19628);
and U19889 (N_19889,N_19631,N_19691);
nand U19890 (N_19890,N_19656,N_19740);
or U19891 (N_19891,N_19742,N_19661);
and U19892 (N_19892,N_19681,N_19634);
xor U19893 (N_19893,N_19766,N_19671);
nand U19894 (N_19894,N_19686,N_19659);
and U19895 (N_19895,N_19608,N_19752);
or U19896 (N_19896,N_19726,N_19614);
and U19897 (N_19897,N_19703,N_19734);
and U19898 (N_19898,N_19677,N_19695);
xor U19899 (N_19899,N_19689,N_19794);
nand U19900 (N_19900,N_19648,N_19678);
nand U19901 (N_19901,N_19786,N_19759);
and U19902 (N_19902,N_19792,N_19662);
or U19903 (N_19903,N_19629,N_19640);
or U19904 (N_19904,N_19790,N_19665);
nand U19905 (N_19905,N_19696,N_19690);
xnor U19906 (N_19906,N_19670,N_19657);
and U19907 (N_19907,N_19787,N_19795);
nor U19908 (N_19908,N_19746,N_19611);
nand U19909 (N_19909,N_19769,N_19773);
or U19910 (N_19910,N_19640,N_19794);
and U19911 (N_19911,N_19704,N_19635);
xor U19912 (N_19912,N_19763,N_19765);
or U19913 (N_19913,N_19783,N_19611);
nand U19914 (N_19914,N_19656,N_19679);
or U19915 (N_19915,N_19684,N_19622);
nand U19916 (N_19916,N_19697,N_19797);
xnor U19917 (N_19917,N_19630,N_19602);
xnor U19918 (N_19918,N_19632,N_19787);
nand U19919 (N_19919,N_19696,N_19709);
nor U19920 (N_19920,N_19708,N_19636);
and U19921 (N_19921,N_19705,N_19727);
or U19922 (N_19922,N_19643,N_19702);
nand U19923 (N_19923,N_19749,N_19758);
and U19924 (N_19924,N_19705,N_19708);
and U19925 (N_19925,N_19733,N_19632);
nand U19926 (N_19926,N_19702,N_19721);
or U19927 (N_19927,N_19788,N_19631);
and U19928 (N_19928,N_19706,N_19739);
and U19929 (N_19929,N_19641,N_19792);
nor U19930 (N_19930,N_19742,N_19744);
xor U19931 (N_19931,N_19697,N_19631);
nor U19932 (N_19932,N_19691,N_19600);
nor U19933 (N_19933,N_19746,N_19608);
and U19934 (N_19934,N_19730,N_19668);
xnor U19935 (N_19935,N_19737,N_19664);
and U19936 (N_19936,N_19693,N_19714);
and U19937 (N_19937,N_19634,N_19784);
or U19938 (N_19938,N_19745,N_19775);
or U19939 (N_19939,N_19721,N_19684);
and U19940 (N_19940,N_19763,N_19764);
xor U19941 (N_19941,N_19799,N_19729);
nor U19942 (N_19942,N_19708,N_19724);
or U19943 (N_19943,N_19704,N_19772);
and U19944 (N_19944,N_19785,N_19703);
nand U19945 (N_19945,N_19650,N_19796);
or U19946 (N_19946,N_19791,N_19658);
nand U19947 (N_19947,N_19777,N_19670);
nor U19948 (N_19948,N_19786,N_19776);
and U19949 (N_19949,N_19792,N_19612);
and U19950 (N_19950,N_19739,N_19733);
nor U19951 (N_19951,N_19664,N_19769);
or U19952 (N_19952,N_19614,N_19646);
xnor U19953 (N_19953,N_19663,N_19784);
nand U19954 (N_19954,N_19769,N_19616);
xor U19955 (N_19955,N_19681,N_19622);
nor U19956 (N_19956,N_19706,N_19763);
nor U19957 (N_19957,N_19668,N_19742);
nand U19958 (N_19958,N_19713,N_19654);
nand U19959 (N_19959,N_19615,N_19783);
or U19960 (N_19960,N_19764,N_19663);
xnor U19961 (N_19961,N_19744,N_19708);
and U19962 (N_19962,N_19607,N_19601);
and U19963 (N_19963,N_19676,N_19769);
nor U19964 (N_19964,N_19761,N_19621);
and U19965 (N_19965,N_19671,N_19664);
or U19966 (N_19966,N_19714,N_19634);
xor U19967 (N_19967,N_19619,N_19718);
nor U19968 (N_19968,N_19643,N_19644);
xor U19969 (N_19969,N_19614,N_19766);
or U19970 (N_19970,N_19722,N_19679);
or U19971 (N_19971,N_19697,N_19620);
nor U19972 (N_19972,N_19645,N_19686);
and U19973 (N_19973,N_19635,N_19752);
nand U19974 (N_19974,N_19756,N_19795);
nand U19975 (N_19975,N_19618,N_19769);
nand U19976 (N_19976,N_19646,N_19603);
and U19977 (N_19977,N_19756,N_19648);
nand U19978 (N_19978,N_19671,N_19726);
nand U19979 (N_19979,N_19771,N_19607);
xor U19980 (N_19980,N_19615,N_19678);
or U19981 (N_19981,N_19734,N_19783);
nand U19982 (N_19982,N_19754,N_19693);
or U19983 (N_19983,N_19634,N_19617);
or U19984 (N_19984,N_19687,N_19734);
nor U19985 (N_19985,N_19651,N_19781);
xnor U19986 (N_19986,N_19700,N_19779);
or U19987 (N_19987,N_19659,N_19718);
nor U19988 (N_19988,N_19630,N_19792);
and U19989 (N_19989,N_19608,N_19734);
nand U19990 (N_19990,N_19641,N_19726);
or U19991 (N_19991,N_19756,N_19746);
or U19992 (N_19992,N_19774,N_19739);
and U19993 (N_19993,N_19793,N_19692);
or U19994 (N_19994,N_19791,N_19762);
nor U19995 (N_19995,N_19619,N_19601);
xnor U19996 (N_19996,N_19727,N_19623);
nor U19997 (N_19997,N_19695,N_19720);
and U19998 (N_19998,N_19655,N_19675);
or U19999 (N_19999,N_19706,N_19687);
or U20000 (N_20000,N_19867,N_19909);
and U20001 (N_20001,N_19969,N_19900);
nand U20002 (N_20002,N_19981,N_19899);
nor U20003 (N_20003,N_19870,N_19855);
and U20004 (N_20004,N_19943,N_19812);
xnor U20005 (N_20005,N_19828,N_19887);
nor U20006 (N_20006,N_19932,N_19888);
or U20007 (N_20007,N_19841,N_19930);
or U20008 (N_20008,N_19862,N_19941);
nand U20009 (N_20009,N_19956,N_19801);
and U20010 (N_20010,N_19991,N_19914);
nand U20011 (N_20011,N_19908,N_19924);
nand U20012 (N_20012,N_19989,N_19863);
nor U20013 (N_20013,N_19827,N_19800);
nor U20014 (N_20014,N_19815,N_19919);
nor U20015 (N_20015,N_19945,N_19940);
xnor U20016 (N_20016,N_19881,N_19944);
and U20017 (N_20017,N_19894,N_19869);
nand U20018 (N_20018,N_19835,N_19833);
or U20019 (N_20019,N_19830,N_19846);
and U20020 (N_20020,N_19880,N_19964);
nand U20021 (N_20021,N_19821,N_19977);
or U20022 (N_20022,N_19994,N_19813);
nor U20023 (N_20023,N_19839,N_19819);
or U20024 (N_20024,N_19885,N_19921);
and U20025 (N_20025,N_19875,N_19837);
and U20026 (N_20026,N_19906,N_19963);
or U20027 (N_20027,N_19953,N_19980);
xor U20028 (N_20028,N_19884,N_19952);
nand U20029 (N_20029,N_19999,N_19820);
or U20030 (N_20030,N_19893,N_19842);
nand U20031 (N_20031,N_19926,N_19849);
nor U20032 (N_20032,N_19942,N_19829);
nor U20033 (N_20033,N_19988,N_19861);
nor U20034 (N_20034,N_19911,N_19871);
or U20035 (N_20035,N_19928,N_19851);
nand U20036 (N_20036,N_19965,N_19915);
nor U20037 (N_20037,N_19973,N_19818);
xor U20038 (N_20038,N_19970,N_19986);
xnor U20039 (N_20039,N_19987,N_19810);
nor U20040 (N_20040,N_19975,N_19918);
nand U20041 (N_20041,N_19954,N_19803);
nor U20042 (N_20042,N_19805,N_19857);
or U20043 (N_20043,N_19934,N_19868);
or U20044 (N_20044,N_19901,N_19874);
nor U20045 (N_20045,N_19938,N_19967);
or U20046 (N_20046,N_19806,N_19825);
nand U20047 (N_20047,N_19990,N_19858);
and U20048 (N_20048,N_19895,N_19852);
or U20049 (N_20049,N_19834,N_19910);
and U20050 (N_20050,N_19878,N_19838);
xor U20051 (N_20051,N_19877,N_19896);
nand U20052 (N_20052,N_19984,N_19972);
or U20053 (N_20053,N_19971,N_19933);
nand U20054 (N_20054,N_19913,N_19974);
nor U20055 (N_20055,N_19843,N_19949);
xnor U20056 (N_20056,N_19985,N_19883);
or U20057 (N_20057,N_19951,N_19802);
or U20058 (N_20058,N_19922,N_19872);
nor U20059 (N_20059,N_19848,N_19866);
and U20060 (N_20060,N_19948,N_19923);
nand U20061 (N_20061,N_19936,N_19879);
xnor U20062 (N_20062,N_19889,N_19968);
and U20063 (N_20063,N_19959,N_19962);
nand U20064 (N_20064,N_19859,N_19860);
or U20065 (N_20065,N_19939,N_19840);
and U20066 (N_20066,N_19836,N_19876);
or U20067 (N_20067,N_19907,N_19935);
or U20068 (N_20068,N_19997,N_19904);
xor U20069 (N_20069,N_19998,N_19804);
or U20070 (N_20070,N_19957,N_19832);
xnor U20071 (N_20071,N_19854,N_19809);
nand U20072 (N_20072,N_19916,N_19864);
xnor U20073 (N_20073,N_19890,N_19978);
or U20074 (N_20074,N_19912,N_19950);
nor U20075 (N_20075,N_19897,N_19947);
and U20076 (N_20076,N_19822,N_19847);
nand U20077 (N_20077,N_19814,N_19873);
nor U20078 (N_20078,N_19845,N_19886);
nor U20079 (N_20079,N_19816,N_19853);
xor U20080 (N_20080,N_19931,N_19898);
and U20081 (N_20081,N_19937,N_19865);
and U20082 (N_20082,N_19917,N_19979);
nand U20083 (N_20083,N_19946,N_19927);
nor U20084 (N_20084,N_19955,N_19826);
or U20085 (N_20085,N_19856,N_19903);
nand U20086 (N_20086,N_19850,N_19831);
or U20087 (N_20087,N_19976,N_19996);
nand U20088 (N_20088,N_19811,N_19992);
and U20089 (N_20089,N_19824,N_19882);
and U20090 (N_20090,N_19995,N_19929);
and U20091 (N_20091,N_19817,N_19960);
nand U20092 (N_20092,N_19902,N_19958);
and U20093 (N_20093,N_19982,N_19823);
nand U20094 (N_20094,N_19993,N_19983);
or U20095 (N_20095,N_19966,N_19808);
xnor U20096 (N_20096,N_19905,N_19891);
nand U20097 (N_20097,N_19961,N_19920);
and U20098 (N_20098,N_19807,N_19892);
nor U20099 (N_20099,N_19925,N_19844);
and U20100 (N_20100,N_19951,N_19971);
nor U20101 (N_20101,N_19963,N_19929);
and U20102 (N_20102,N_19936,N_19846);
xnor U20103 (N_20103,N_19800,N_19998);
or U20104 (N_20104,N_19844,N_19815);
or U20105 (N_20105,N_19831,N_19893);
xor U20106 (N_20106,N_19962,N_19841);
or U20107 (N_20107,N_19918,N_19897);
nand U20108 (N_20108,N_19810,N_19867);
nor U20109 (N_20109,N_19806,N_19901);
and U20110 (N_20110,N_19940,N_19906);
nand U20111 (N_20111,N_19879,N_19871);
and U20112 (N_20112,N_19896,N_19848);
and U20113 (N_20113,N_19971,N_19804);
nor U20114 (N_20114,N_19994,N_19841);
nand U20115 (N_20115,N_19901,N_19974);
or U20116 (N_20116,N_19946,N_19891);
xor U20117 (N_20117,N_19873,N_19824);
or U20118 (N_20118,N_19860,N_19865);
xnor U20119 (N_20119,N_19855,N_19837);
or U20120 (N_20120,N_19881,N_19955);
nor U20121 (N_20121,N_19951,N_19960);
xnor U20122 (N_20122,N_19800,N_19826);
xnor U20123 (N_20123,N_19900,N_19958);
nand U20124 (N_20124,N_19807,N_19971);
nand U20125 (N_20125,N_19805,N_19839);
nand U20126 (N_20126,N_19858,N_19870);
and U20127 (N_20127,N_19862,N_19942);
or U20128 (N_20128,N_19822,N_19820);
and U20129 (N_20129,N_19835,N_19944);
and U20130 (N_20130,N_19850,N_19839);
nor U20131 (N_20131,N_19993,N_19818);
xnor U20132 (N_20132,N_19939,N_19946);
nor U20133 (N_20133,N_19896,N_19984);
nand U20134 (N_20134,N_19862,N_19964);
nand U20135 (N_20135,N_19856,N_19839);
or U20136 (N_20136,N_19919,N_19958);
or U20137 (N_20137,N_19885,N_19846);
xor U20138 (N_20138,N_19934,N_19904);
nand U20139 (N_20139,N_19861,N_19987);
nand U20140 (N_20140,N_19914,N_19997);
xnor U20141 (N_20141,N_19855,N_19809);
and U20142 (N_20142,N_19868,N_19905);
and U20143 (N_20143,N_19927,N_19925);
nand U20144 (N_20144,N_19838,N_19995);
or U20145 (N_20145,N_19876,N_19869);
or U20146 (N_20146,N_19976,N_19870);
xnor U20147 (N_20147,N_19972,N_19927);
nand U20148 (N_20148,N_19837,N_19808);
nor U20149 (N_20149,N_19805,N_19988);
and U20150 (N_20150,N_19978,N_19990);
xnor U20151 (N_20151,N_19951,N_19994);
nand U20152 (N_20152,N_19996,N_19948);
or U20153 (N_20153,N_19811,N_19983);
nor U20154 (N_20154,N_19979,N_19954);
xnor U20155 (N_20155,N_19919,N_19952);
and U20156 (N_20156,N_19831,N_19962);
nand U20157 (N_20157,N_19809,N_19813);
and U20158 (N_20158,N_19824,N_19914);
or U20159 (N_20159,N_19862,N_19917);
nand U20160 (N_20160,N_19995,N_19879);
nand U20161 (N_20161,N_19812,N_19926);
nor U20162 (N_20162,N_19956,N_19882);
nor U20163 (N_20163,N_19855,N_19930);
nor U20164 (N_20164,N_19960,N_19990);
xnor U20165 (N_20165,N_19868,N_19887);
nor U20166 (N_20166,N_19993,N_19821);
and U20167 (N_20167,N_19979,N_19902);
or U20168 (N_20168,N_19950,N_19988);
or U20169 (N_20169,N_19953,N_19818);
and U20170 (N_20170,N_19895,N_19812);
and U20171 (N_20171,N_19986,N_19923);
nand U20172 (N_20172,N_19834,N_19950);
xnor U20173 (N_20173,N_19810,N_19897);
nand U20174 (N_20174,N_19843,N_19959);
nor U20175 (N_20175,N_19962,N_19948);
xnor U20176 (N_20176,N_19906,N_19802);
xor U20177 (N_20177,N_19940,N_19806);
xnor U20178 (N_20178,N_19947,N_19969);
and U20179 (N_20179,N_19887,N_19911);
or U20180 (N_20180,N_19840,N_19960);
or U20181 (N_20181,N_19828,N_19821);
and U20182 (N_20182,N_19974,N_19803);
nand U20183 (N_20183,N_19986,N_19934);
xor U20184 (N_20184,N_19952,N_19851);
nand U20185 (N_20185,N_19906,N_19929);
or U20186 (N_20186,N_19879,N_19934);
or U20187 (N_20187,N_19867,N_19926);
or U20188 (N_20188,N_19913,N_19834);
nor U20189 (N_20189,N_19864,N_19820);
or U20190 (N_20190,N_19884,N_19885);
nor U20191 (N_20191,N_19865,N_19995);
and U20192 (N_20192,N_19854,N_19993);
xnor U20193 (N_20193,N_19921,N_19961);
and U20194 (N_20194,N_19823,N_19846);
xor U20195 (N_20195,N_19887,N_19912);
nor U20196 (N_20196,N_19958,N_19915);
nand U20197 (N_20197,N_19884,N_19899);
nor U20198 (N_20198,N_19881,N_19829);
or U20199 (N_20199,N_19980,N_19860);
xor U20200 (N_20200,N_20118,N_20001);
xor U20201 (N_20201,N_20096,N_20023);
nor U20202 (N_20202,N_20111,N_20193);
and U20203 (N_20203,N_20174,N_20100);
and U20204 (N_20204,N_20066,N_20139);
nor U20205 (N_20205,N_20172,N_20069);
and U20206 (N_20206,N_20058,N_20137);
nand U20207 (N_20207,N_20022,N_20005);
xor U20208 (N_20208,N_20013,N_20123);
nor U20209 (N_20209,N_20190,N_20038);
or U20210 (N_20210,N_20028,N_20093);
nand U20211 (N_20211,N_20018,N_20060);
or U20212 (N_20212,N_20188,N_20003);
and U20213 (N_20213,N_20162,N_20025);
and U20214 (N_20214,N_20113,N_20103);
and U20215 (N_20215,N_20009,N_20051);
xnor U20216 (N_20216,N_20032,N_20088);
nor U20217 (N_20217,N_20158,N_20065);
nand U20218 (N_20218,N_20068,N_20166);
nand U20219 (N_20219,N_20015,N_20160);
nand U20220 (N_20220,N_20143,N_20008);
xor U20221 (N_20221,N_20067,N_20136);
nand U20222 (N_20222,N_20191,N_20132);
or U20223 (N_20223,N_20052,N_20019);
or U20224 (N_20224,N_20178,N_20095);
xnor U20225 (N_20225,N_20129,N_20029);
nor U20226 (N_20226,N_20089,N_20194);
nand U20227 (N_20227,N_20034,N_20109);
and U20228 (N_20228,N_20037,N_20175);
xnor U20229 (N_20229,N_20061,N_20110);
nand U20230 (N_20230,N_20105,N_20185);
and U20231 (N_20231,N_20189,N_20036);
and U20232 (N_20232,N_20085,N_20176);
and U20233 (N_20233,N_20108,N_20041);
and U20234 (N_20234,N_20165,N_20184);
nor U20235 (N_20235,N_20048,N_20072);
nor U20236 (N_20236,N_20135,N_20117);
or U20237 (N_20237,N_20044,N_20039);
xor U20238 (N_20238,N_20074,N_20046);
xor U20239 (N_20239,N_20045,N_20027);
xnor U20240 (N_20240,N_20062,N_20186);
xor U20241 (N_20241,N_20002,N_20043);
xor U20242 (N_20242,N_20187,N_20170);
or U20243 (N_20243,N_20097,N_20076);
nor U20244 (N_20244,N_20196,N_20182);
and U20245 (N_20245,N_20083,N_20000);
nor U20246 (N_20246,N_20115,N_20177);
xor U20247 (N_20247,N_20198,N_20081);
nand U20248 (N_20248,N_20035,N_20133);
nor U20249 (N_20249,N_20112,N_20075);
xnor U20250 (N_20250,N_20114,N_20151);
and U20251 (N_20251,N_20050,N_20164);
and U20252 (N_20252,N_20126,N_20012);
xor U20253 (N_20253,N_20120,N_20159);
or U20254 (N_20254,N_20073,N_20121);
nand U20255 (N_20255,N_20130,N_20053);
or U20256 (N_20256,N_20004,N_20064);
or U20257 (N_20257,N_20195,N_20090);
nand U20258 (N_20258,N_20104,N_20150);
and U20259 (N_20259,N_20163,N_20007);
or U20260 (N_20260,N_20171,N_20059);
or U20261 (N_20261,N_20134,N_20128);
or U20262 (N_20262,N_20087,N_20055);
nor U20263 (N_20263,N_20071,N_20010);
and U20264 (N_20264,N_20124,N_20006);
and U20265 (N_20265,N_20183,N_20020);
and U20266 (N_20266,N_20017,N_20049);
xor U20267 (N_20267,N_20101,N_20122);
xnor U20268 (N_20268,N_20091,N_20127);
xnor U20269 (N_20269,N_20192,N_20156);
xor U20270 (N_20270,N_20078,N_20031);
nor U20271 (N_20271,N_20154,N_20197);
nor U20272 (N_20272,N_20116,N_20146);
xor U20273 (N_20273,N_20063,N_20054);
nor U20274 (N_20274,N_20016,N_20179);
xnor U20275 (N_20275,N_20107,N_20057);
nand U20276 (N_20276,N_20077,N_20153);
nand U20277 (N_20277,N_20094,N_20145);
and U20278 (N_20278,N_20033,N_20157);
and U20279 (N_20279,N_20161,N_20152);
nand U20280 (N_20280,N_20173,N_20099);
xor U20281 (N_20281,N_20011,N_20169);
xnor U20282 (N_20282,N_20080,N_20056);
and U20283 (N_20283,N_20168,N_20092);
or U20284 (N_20284,N_20047,N_20125);
xnor U20285 (N_20285,N_20106,N_20026);
nand U20286 (N_20286,N_20042,N_20030);
nor U20287 (N_20287,N_20014,N_20147);
xnor U20288 (N_20288,N_20119,N_20140);
xor U20289 (N_20289,N_20138,N_20141);
and U20290 (N_20290,N_20131,N_20142);
or U20291 (N_20291,N_20084,N_20102);
xor U20292 (N_20292,N_20024,N_20070);
and U20293 (N_20293,N_20180,N_20144);
nand U20294 (N_20294,N_20082,N_20086);
and U20295 (N_20295,N_20149,N_20181);
nand U20296 (N_20296,N_20098,N_20021);
xor U20297 (N_20297,N_20167,N_20148);
or U20298 (N_20298,N_20040,N_20199);
xor U20299 (N_20299,N_20155,N_20079);
xor U20300 (N_20300,N_20069,N_20081);
or U20301 (N_20301,N_20079,N_20000);
nand U20302 (N_20302,N_20013,N_20132);
xor U20303 (N_20303,N_20180,N_20168);
and U20304 (N_20304,N_20051,N_20046);
nor U20305 (N_20305,N_20084,N_20153);
xnor U20306 (N_20306,N_20098,N_20041);
nor U20307 (N_20307,N_20194,N_20185);
or U20308 (N_20308,N_20105,N_20035);
and U20309 (N_20309,N_20061,N_20106);
nand U20310 (N_20310,N_20141,N_20161);
xnor U20311 (N_20311,N_20172,N_20152);
or U20312 (N_20312,N_20029,N_20044);
or U20313 (N_20313,N_20022,N_20028);
nor U20314 (N_20314,N_20145,N_20185);
or U20315 (N_20315,N_20105,N_20126);
or U20316 (N_20316,N_20016,N_20152);
nor U20317 (N_20317,N_20016,N_20157);
and U20318 (N_20318,N_20119,N_20173);
or U20319 (N_20319,N_20134,N_20183);
nor U20320 (N_20320,N_20011,N_20076);
nor U20321 (N_20321,N_20166,N_20107);
xor U20322 (N_20322,N_20176,N_20105);
nand U20323 (N_20323,N_20198,N_20044);
or U20324 (N_20324,N_20132,N_20109);
and U20325 (N_20325,N_20156,N_20041);
or U20326 (N_20326,N_20008,N_20144);
or U20327 (N_20327,N_20023,N_20089);
and U20328 (N_20328,N_20072,N_20030);
nor U20329 (N_20329,N_20030,N_20049);
nor U20330 (N_20330,N_20029,N_20037);
nand U20331 (N_20331,N_20047,N_20122);
or U20332 (N_20332,N_20149,N_20055);
and U20333 (N_20333,N_20104,N_20048);
nand U20334 (N_20334,N_20096,N_20087);
xor U20335 (N_20335,N_20036,N_20197);
and U20336 (N_20336,N_20006,N_20090);
nor U20337 (N_20337,N_20107,N_20053);
or U20338 (N_20338,N_20071,N_20013);
xnor U20339 (N_20339,N_20190,N_20069);
nor U20340 (N_20340,N_20012,N_20166);
xor U20341 (N_20341,N_20089,N_20091);
nor U20342 (N_20342,N_20100,N_20007);
nand U20343 (N_20343,N_20115,N_20070);
nor U20344 (N_20344,N_20079,N_20125);
and U20345 (N_20345,N_20148,N_20073);
xor U20346 (N_20346,N_20139,N_20114);
xor U20347 (N_20347,N_20000,N_20137);
and U20348 (N_20348,N_20090,N_20169);
and U20349 (N_20349,N_20025,N_20029);
nand U20350 (N_20350,N_20138,N_20004);
nand U20351 (N_20351,N_20179,N_20071);
and U20352 (N_20352,N_20148,N_20003);
and U20353 (N_20353,N_20080,N_20162);
nand U20354 (N_20354,N_20008,N_20147);
nor U20355 (N_20355,N_20109,N_20103);
nor U20356 (N_20356,N_20195,N_20082);
xor U20357 (N_20357,N_20035,N_20020);
or U20358 (N_20358,N_20117,N_20177);
or U20359 (N_20359,N_20175,N_20084);
and U20360 (N_20360,N_20070,N_20179);
and U20361 (N_20361,N_20029,N_20193);
nand U20362 (N_20362,N_20018,N_20128);
nor U20363 (N_20363,N_20098,N_20026);
nand U20364 (N_20364,N_20098,N_20103);
nor U20365 (N_20365,N_20147,N_20005);
nor U20366 (N_20366,N_20079,N_20035);
or U20367 (N_20367,N_20166,N_20035);
and U20368 (N_20368,N_20122,N_20154);
nor U20369 (N_20369,N_20075,N_20093);
xor U20370 (N_20370,N_20005,N_20059);
or U20371 (N_20371,N_20181,N_20113);
xnor U20372 (N_20372,N_20191,N_20082);
nand U20373 (N_20373,N_20013,N_20130);
nor U20374 (N_20374,N_20080,N_20134);
or U20375 (N_20375,N_20076,N_20049);
and U20376 (N_20376,N_20054,N_20141);
and U20377 (N_20377,N_20062,N_20106);
or U20378 (N_20378,N_20105,N_20141);
or U20379 (N_20379,N_20153,N_20090);
nor U20380 (N_20380,N_20012,N_20146);
and U20381 (N_20381,N_20171,N_20144);
nor U20382 (N_20382,N_20114,N_20169);
xor U20383 (N_20383,N_20049,N_20047);
or U20384 (N_20384,N_20059,N_20118);
xnor U20385 (N_20385,N_20081,N_20151);
nor U20386 (N_20386,N_20098,N_20106);
and U20387 (N_20387,N_20127,N_20006);
xnor U20388 (N_20388,N_20098,N_20198);
xor U20389 (N_20389,N_20168,N_20108);
xor U20390 (N_20390,N_20140,N_20189);
nand U20391 (N_20391,N_20135,N_20177);
xor U20392 (N_20392,N_20044,N_20109);
nor U20393 (N_20393,N_20080,N_20159);
nor U20394 (N_20394,N_20176,N_20151);
xnor U20395 (N_20395,N_20133,N_20025);
and U20396 (N_20396,N_20136,N_20127);
or U20397 (N_20397,N_20189,N_20193);
nor U20398 (N_20398,N_20028,N_20197);
nor U20399 (N_20399,N_20020,N_20190);
nor U20400 (N_20400,N_20209,N_20336);
nand U20401 (N_20401,N_20384,N_20286);
xor U20402 (N_20402,N_20291,N_20344);
xnor U20403 (N_20403,N_20246,N_20276);
nor U20404 (N_20404,N_20362,N_20222);
xor U20405 (N_20405,N_20272,N_20357);
or U20406 (N_20406,N_20229,N_20201);
or U20407 (N_20407,N_20316,N_20275);
nand U20408 (N_20408,N_20278,N_20391);
nand U20409 (N_20409,N_20342,N_20393);
and U20410 (N_20410,N_20320,N_20345);
and U20411 (N_20411,N_20317,N_20343);
or U20412 (N_20412,N_20300,N_20376);
xor U20413 (N_20413,N_20254,N_20213);
nor U20414 (N_20414,N_20386,N_20240);
or U20415 (N_20415,N_20215,N_20328);
xnor U20416 (N_20416,N_20378,N_20238);
xnor U20417 (N_20417,N_20323,N_20263);
xnor U20418 (N_20418,N_20228,N_20292);
or U20419 (N_20419,N_20385,N_20324);
xnor U20420 (N_20420,N_20266,N_20383);
nor U20421 (N_20421,N_20258,N_20329);
nor U20422 (N_20422,N_20270,N_20368);
nand U20423 (N_20423,N_20299,N_20306);
and U20424 (N_20424,N_20371,N_20282);
xor U20425 (N_20425,N_20212,N_20369);
nor U20426 (N_20426,N_20231,N_20359);
xnor U20427 (N_20427,N_20287,N_20373);
and U20428 (N_20428,N_20330,N_20237);
or U20429 (N_20429,N_20250,N_20349);
nand U20430 (N_20430,N_20319,N_20236);
or U20431 (N_20431,N_20372,N_20308);
nand U20432 (N_20432,N_20200,N_20374);
or U20433 (N_20433,N_20239,N_20235);
nor U20434 (N_20434,N_20399,N_20252);
or U20435 (N_20435,N_20394,N_20234);
nor U20436 (N_20436,N_20367,N_20358);
and U20437 (N_20437,N_20283,N_20313);
and U20438 (N_20438,N_20261,N_20298);
nand U20439 (N_20439,N_20337,N_20353);
xnor U20440 (N_20440,N_20301,N_20225);
and U20441 (N_20441,N_20256,N_20363);
nand U20442 (N_20442,N_20351,N_20227);
nand U20443 (N_20443,N_20289,N_20294);
or U20444 (N_20444,N_20352,N_20346);
nor U20445 (N_20445,N_20271,N_20232);
nor U20446 (N_20446,N_20322,N_20377);
and U20447 (N_20447,N_20341,N_20249);
or U20448 (N_20448,N_20333,N_20284);
xnor U20449 (N_20449,N_20242,N_20302);
nor U20450 (N_20450,N_20366,N_20309);
xnor U20451 (N_20451,N_20260,N_20347);
and U20452 (N_20452,N_20327,N_20221);
xnor U20453 (N_20453,N_20395,N_20398);
or U20454 (N_20454,N_20279,N_20381);
nand U20455 (N_20455,N_20241,N_20390);
xnor U20456 (N_20456,N_20248,N_20223);
xor U20457 (N_20457,N_20233,N_20382);
xor U20458 (N_20458,N_20365,N_20207);
and U20459 (N_20459,N_20204,N_20206);
nor U20460 (N_20460,N_20257,N_20318);
or U20461 (N_20461,N_20334,N_20311);
nand U20462 (N_20462,N_20335,N_20296);
and U20463 (N_20463,N_20214,N_20304);
nor U20464 (N_20464,N_20332,N_20379);
or U20465 (N_20465,N_20217,N_20205);
and U20466 (N_20466,N_20265,N_20361);
and U20467 (N_20467,N_20211,N_20370);
or U20468 (N_20468,N_20244,N_20219);
and U20469 (N_20469,N_20354,N_20326);
xor U20470 (N_20470,N_20218,N_20312);
nor U20471 (N_20471,N_20277,N_20210);
and U20472 (N_20472,N_20307,N_20230);
nand U20473 (N_20473,N_20355,N_20387);
and U20474 (N_20474,N_20339,N_20295);
or U20475 (N_20475,N_20305,N_20290);
and U20476 (N_20476,N_20375,N_20356);
and U20477 (N_20477,N_20251,N_20338);
xnor U20478 (N_20478,N_20297,N_20285);
and U20479 (N_20479,N_20220,N_20288);
and U20480 (N_20480,N_20310,N_20267);
nand U20481 (N_20481,N_20247,N_20259);
xnor U20482 (N_20482,N_20303,N_20274);
or U20483 (N_20483,N_20331,N_20388);
nand U20484 (N_20484,N_20226,N_20280);
nor U20485 (N_20485,N_20380,N_20243);
and U20486 (N_20486,N_20321,N_20396);
nand U20487 (N_20487,N_20281,N_20245);
or U20488 (N_20488,N_20264,N_20253);
and U20489 (N_20489,N_20262,N_20350);
and U20490 (N_20490,N_20224,N_20315);
or U20491 (N_20491,N_20325,N_20392);
xnor U20492 (N_20492,N_20268,N_20360);
nand U20493 (N_20493,N_20314,N_20293);
xnor U20494 (N_20494,N_20389,N_20202);
and U20495 (N_20495,N_20340,N_20208);
or U20496 (N_20496,N_20397,N_20216);
or U20497 (N_20497,N_20348,N_20364);
nand U20498 (N_20498,N_20203,N_20273);
nor U20499 (N_20499,N_20269,N_20255);
xor U20500 (N_20500,N_20201,N_20254);
nand U20501 (N_20501,N_20325,N_20361);
and U20502 (N_20502,N_20264,N_20299);
and U20503 (N_20503,N_20374,N_20302);
nand U20504 (N_20504,N_20312,N_20234);
and U20505 (N_20505,N_20266,N_20321);
nand U20506 (N_20506,N_20246,N_20295);
or U20507 (N_20507,N_20267,N_20299);
or U20508 (N_20508,N_20354,N_20384);
nand U20509 (N_20509,N_20329,N_20293);
or U20510 (N_20510,N_20365,N_20348);
xnor U20511 (N_20511,N_20252,N_20354);
or U20512 (N_20512,N_20313,N_20334);
and U20513 (N_20513,N_20368,N_20306);
or U20514 (N_20514,N_20239,N_20321);
nand U20515 (N_20515,N_20299,N_20335);
nand U20516 (N_20516,N_20215,N_20204);
nand U20517 (N_20517,N_20378,N_20395);
or U20518 (N_20518,N_20209,N_20325);
nor U20519 (N_20519,N_20205,N_20248);
xor U20520 (N_20520,N_20275,N_20229);
xor U20521 (N_20521,N_20362,N_20313);
nand U20522 (N_20522,N_20246,N_20315);
and U20523 (N_20523,N_20225,N_20274);
nand U20524 (N_20524,N_20387,N_20395);
xnor U20525 (N_20525,N_20352,N_20215);
or U20526 (N_20526,N_20276,N_20273);
nand U20527 (N_20527,N_20366,N_20376);
nor U20528 (N_20528,N_20264,N_20222);
and U20529 (N_20529,N_20278,N_20395);
nand U20530 (N_20530,N_20331,N_20227);
nand U20531 (N_20531,N_20350,N_20357);
xor U20532 (N_20532,N_20278,N_20362);
nand U20533 (N_20533,N_20303,N_20392);
nand U20534 (N_20534,N_20297,N_20344);
and U20535 (N_20535,N_20220,N_20247);
and U20536 (N_20536,N_20316,N_20205);
or U20537 (N_20537,N_20305,N_20367);
and U20538 (N_20538,N_20311,N_20263);
nor U20539 (N_20539,N_20331,N_20399);
nor U20540 (N_20540,N_20326,N_20282);
or U20541 (N_20541,N_20221,N_20351);
xor U20542 (N_20542,N_20220,N_20230);
nor U20543 (N_20543,N_20293,N_20242);
and U20544 (N_20544,N_20224,N_20384);
and U20545 (N_20545,N_20322,N_20328);
nor U20546 (N_20546,N_20385,N_20335);
nand U20547 (N_20547,N_20200,N_20328);
nand U20548 (N_20548,N_20320,N_20247);
xnor U20549 (N_20549,N_20384,N_20232);
nor U20550 (N_20550,N_20310,N_20209);
or U20551 (N_20551,N_20312,N_20226);
nand U20552 (N_20552,N_20281,N_20377);
nor U20553 (N_20553,N_20386,N_20253);
nor U20554 (N_20554,N_20303,N_20351);
and U20555 (N_20555,N_20225,N_20263);
xnor U20556 (N_20556,N_20390,N_20353);
nand U20557 (N_20557,N_20251,N_20229);
and U20558 (N_20558,N_20231,N_20393);
or U20559 (N_20559,N_20289,N_20346);
xnor U20560 (N_20560,N_20238,N_20399);
xor U20561 (N_20561,N_20361,N_20305);
nor U20562 (N_20562,N_20327,N_20388);
and U20563 (N_20563,N_20359,N_20274);
or U20564 (N_20564,N_20343,N_20271);
or U20565 (N_20565,N_20366,N_20385);
nand U20566 (N_20566,N_20384,N_20395);
and U20567 (N_20567,N_20217,N_20227);
or U20568 (N_20568,N_20358,N_20369);
nand U20569 (N_20569,N_20329,N_20266);
or U20570 (N_20570,N_20205,N_20381);
xor U20571 (N_20571,N_20200,N_20277);
xnor U20572 (N_20572,N_20271,N_20244);
or U20573 (N_20573,N_20221,N_20324);
nor U20574 (N_20574,N_20214,N_20320);
nand U20575 (N_20575,N_20249,N_20354);
nand U20576 (N_20576,N_20387,N_20311);
nand U20577 (N_20577,N_20239,N_20325);
nor U20578 (N_20578,N_20210,N_20374);
nand U20579 (N_20579,N_20357,N_20377);
or U20580 (N_20580,N_20270,N_20226);
xnor U20581 (N_20581,N_20335,N_20339);
nand U20582 (N_20582,N_20254,N_20238);
and U20583 (N_20583,N_20299,N_20212);
nor U20584 (N_20584,N_20231,N_20249);
nand U20585 (N_20585,N_20212,N_20232);
xor U20586 (N_20586,N_20235,N_20243);
or U20587 (N_20587,N_20271,N_20345);
nand U20588 (N_20588,N_20353,N_20380);
nand U20589 (N_20589,N_20227,N_20393);
and U20590 (N_20590,N_20360,N_20381);
and U20591 (N_20591,N_20317,N_20371);
xnor U20592 (N_20592,N_20225,N_20332);
nor U20593 (N_20593,N_20208,N_20204);
or U20594 (N_20594,N_20371,N_20292);
nand U20595 (N_20595,N_20258,N_20365);
and U20596 (N_20596,N_20307,N_20210);
and U20597 (N_20597,N_20290,N_20257);
nand U20598 (N_20598,N_20248,N_20292);
xnor U20599 (N_20599,N_20303,N_20299);
xor U20600 (N_20600,N_20514,N_20579);
nor U20601 (N_20601,N_20558,N_20464);
nand U20602 (N_20602,N_20400,N_20582);
and U20603 (N_20603,N_20539,N_20478);
nor U20604 (N_20604,N_20541,N_20510);
or U20605 (N_20605,N_20475,N_20512);
nand U20606 (N_20606,N_20452,N_20440);
nor U20607 (N_20607,N_20405,N_20580);
xor U20608 (N_20608,N_20546,N_20474);
nor U20609 (N_20609,N_20410,N_20428);
or U20610 (N_20610,N_20492,N_20557);
xnor U20611 (N_20611,N_20457,N_20496);
nor U20612 (N_20612,N_20480,N_20447);
and U20613 (N_20613,N_20483,N_20519);
xnor U20614 (N_20614,N_20479,N_20565);
or U20615 (N_20615,N_20535,N_20592);
nand U20616 (N_20616,N_20571,N_20403);
nor U20617 (N_20617,N_20449,N_20598);
xor U20618 (N_20618,N_20431,N_20583);
nor U20619 (N_20619,N_20561,N_20578);
or U20620 (N_20620,N_20593,N_20529);
xor U20621 (N_20621,N_20499,N_20559);
xor U20622 (N_20622,N_20573,N_20581);
or U20623 (N_20623,N_20481,N_20502);
nor U20624 (N_20624,N_20443,N_20595);
and U20625 (N_20625,N_20442,N_20594);
or U20626 (N_20626,N_20459,N_20435);
or U20627 (N_20627,N_20513,N_20591);
or U20628 (N_20628,N_20586,N_20543);
nand U20629 (N_20629,N_20518,N_20425);
or U20630 (N_20630,N_20516,N_20532);
nand U20631 (N_20631,N_20528,N_20441);
and U20632 (N_20632,N_20491,N_20429);
xnor U20633 (N_20633,N_20527,N_20537);
and U20634 (N_20634,N_20501,N_20424);
nor U20635 (N_20635,N_20585,N_20488);
or U20636 (N_20636,N_20503,N_20420);
nor U20637 (N_20637,N_20453,N_20438);
nand U20638 (N_20638,N_20470,N_20576);
nor U20639 (N_20639,N_20515,N_20521);
nand U20640 (N_20640,N_20577,N_20551);
and U20641 (N_20641,N_20477,N_20404);
and U20642 (N_20642,N_20422,N_20590);
nand U20643 (N_20643,N_20427,N_20430);
and U20644 (N_20644,N_20506,N_20472);
xnor U20645 (N_20645,N_20432,N_20536);
nor U20646 (N_20646,N_20402,N_20460);
nand U20647 (N_20647,N_20486,N_20524);
and U20648 (N_20648,N_20493,N_20406);
nor U20649 (N_20649,N_20504,N_20560);
nand U20650 (N_20650,N_20531,N_20467);
nor U20651 (N_20651,N_20463,N_20553);
and U20652 (N_20652,N_20407,N_20497);
nand U20653 (N_20653,N_20434,N_20412);
or U20654 (N_20654,N_20451,N_20556);
or U20655 (N_20655,N_20542,N_20423);
or U20656 (N_20656,N_20584,N_20448);
xor U20657 (N_20657,N_20545,N_20525);
or U20658 (N_20658,N_20574,N_20476);
xnor U20659 (N_20659,N_20468,N_20462);
xor U20660 (N_20660,N_20439,N_20485);
nand U20661 (N_20661,N_20587,N_20526);
xor U20662 (N_20662,N_20437,N_20421);
or U20663 (N_20663,N_20550,N_20500);
nand U20664 (N_20664,N_20523,N_20401);
and U20665 (N_20665,N_20548,N_20409);
and U20666 (N_20666,N_20522,N_20456);
nor U20667 (N_20667,N_20552,N_20507);
nor U20668 (N_20668,N_20505,N_20446);
nor U20669 (N_20669,N_20597,N_20487);
nor U20670 (N_20670,N_20589,N_20569);
nor U20671 (N_20671,N_20540,N_20415);
xor U20672 (N_20672,N_20444,N_20414);
nor U20673 (N_20673,N_20436,N_20562);
or U20674 (N_20674,N_20461,N_20564);
xnor U20675 (N_20675,N_20419,N_20411);
or U20676 (N_20676,N_20567,N_20454);
nor U20677 (N_20677,N_20484,N_20555);
xnor U20678 (N_20678,N_20530,N_20575);
or U20679 (N_20679,N_20417,N_20413);
and U20680 (N_20680,N_20511,N_20520);
and U20681 (N_20681,N_20534,N_20418);
xnor U20682 (N_20682,N_20572,N_20509);
xnor U20683 (N_20683,N_20508,N_20469);
nand U20684 (N_20684,N_20588,N_20570);
and U20685 (N_20685,N_20466,N_20538);
and U20686 (N_20686,N_20426,N_20566);
or U20687 (N_20687,N_20489,N_20533);
and U20688 (N_20688,N_20596,N_20563);
nand U20689 (N_20689,N_20517,N_20458);
and U20690 (N_20690,N_20455,N_20473);
nor U20691 (N_20691,N_20568,N_20416);
nand U20692 (N_20692,N_20547,N_20554);
nor U20693 (N_20693,N_20494,N_20495);
nor U20694 (N_20694,N_20490,N_20433);
xor U20695 (N_20695,N_20549,N_20599);
or U20696 (N_20696,N_20498,N_20544);
nor U20697 (N_20697,N_20482,N_20450);
nor U20698 (N_20698,N_20445,N_20465);
xor U20699 (N_20699,N_20408,N_20471);
nand U20700 (N_20700,N_20596,N_20509);
nor U20701 (N_20701,N_20440,N_20589);
nor U20702 (N_20702,N_20539,N_20536);
nand U20703 (N_20703,N_20597,N_20516);
and U20704 (N_20704,N_20552,N_20426);
and U20705 (N_20705,N_20411,N_20541);
nand U20706 (N_20706,N_20427,N_20400);
and U20707 (N_20707,N_20512,N_20457);
and U20708 (N_20708,N_20570,N_20471);
or U20709 (N_20709,N_20561,N_20498);
and U20710 (N_20710,N_20498,N_20514);
nand U20711 (N_20711,N_20464,N_20478);
and U20712 (N_20712,N_20539,N_20449);
nand U20713 (N_20713,N_20475,N_20527);
nor U20714 (N_20714,N_20466,N_20543);
nor U20715 (N_20715,N_20436,N_20409);
and U20716 (N_20716,N_20575,N_20574);
and U20717 (N_20717,N_20486,N_20500);
xor U20718 (N_20718,N_20528,N_20402);
nor U20719 (N_20719,N_20515,N_20500);
or U20720 (N_20720,N_20578,N_20509);
nor U20721 (N_20721,N_20418,N_20480);
nor U20722 (N_20722,N_20569,N_20585);
xor U20723 (N_20723,N_20490,N_20562);
nand U20724 (N_20724,N_20549,N_20449);
or U20725 (N_20725,N_20549,N_20520);
and U20726 (N_20726,N_20542,N_20588);
nand U20727 (N_20727,N_20551,N_20428);
or U20728 (N_20728,N_20486,N_20588);
and U20729 (N_20729,N_20550,N_20429);
xnor U20730 (N_20730,N_20561,N_20433);
and U20731 (N_20731,N_20543,N_20528);
xnor U20732 (N_20732,N_20583,N_20465);
and U20733 (N_20733,N_20551,N_20430);
xnor U20734 (N_20734,N_20535,N_20568);
xor U20735 (N_20735,N_20579,N_20424);
or U20736 (N_20736,N_20595,N_20558);
nor U20737 (N_20737,N_20540,N_20560);
or U20738 (N_20738,N_20422,N_20461);
nand U20739 (N_20739,N_20554,N_20411);
or U20740 (N_20740,N_20556,N_20532);
and U20741 (N_20741,N_20431,N_20465);
nand U20742 (N_20742,N_20425,N_20439);
nor U20743 (N_20743,N_20563,N_20517);
xor U20744 (N_20744,N_20417,N_20568);
or U20745 (N_20745,N_20490,N_20542);
nor U20746 (N_20746,N_20544,N_20539);
nor U20747 (N_20747,N_20535,N_20482);
nand U20748 (N_20748,N_20563,N_20531);
nor U20749 (N_20749,N_20515,N_20470);
xnor U20750 (N_20750,N_20431,N_20459);
xor U20751 (N_20751,N_20551,N_20452);
nand U20752 (N_20752,N_20507,N_20467);
nor U20753 (N_20753,N_20598,N_20523);
xor U20754 (N_20754,N_20537,N_20425);
nor U20755 (N_20755,N_20596,N_20510);
xor U20756 (N_20756,N_20591,N_20550);
or U20757 (N_20757,N_20545,N_20508);
nor U20758 (N_20758,N_20508,N_20538);
xor U20759 (N_20759,N_20507,N_20483);
or U20760 (N_20760,N_20409,N_20527);
and U20761 (N_20761,N_20452,N_20572);
xnor U20762 (N_20762,N_20477,N_20501);
nand U20763 (N_20763,N_20418,N_20439);
nand U20764 (N_20764,N_20509,N_20543);
nor U20765 (N_20765,N_20534,N_20545);
or U20766 (N_20766,N_20469,N_20417);
xnor U20767 (N_20767,N_20474,N_20404);
nor U20768 (N_20768,N_20510,N_20528);
nand U20769 (N_20769,N_20440,N_20432);
xnor U20770 (N_20770,N_20467,N_20423);
nand U20771 (N_20771,N_20509,N_20409);
nor U20772 (N_20772,N_20434,N_20582);
xor U20773 (N_20773,N_20423,N_20538);
nand U20774 (N_20774,N_20425,N_20584);
nor U20775 (N_20775,N_20501,N_20572);
and U20776 (N_20776,N_20497,N_20511);
xor U20777 (N_20777,N_20464,N_20470);
or U20778 (N_20778,N_20479,N_20540);
or U20779 (N_20779,N_20449,N_20596);
xnor U20780 (N_20780,N_20436,N_20456);
or U20781 (N_20781,N_20441,N_20468);
xnor U20782 (N_20782,N_20505,N_20436);
and U20783 (N_20783,N_20587,N_20579);
or U20784 (N_20784,N_20460,N_20443);
or U20785 (N_20785,N_20491,N_20453);
xnor U20786 (N_20786,N_20573,N_20569);
and U20787 (N_20787,N_20426,N_20554);
nand U20788 (N_20788,N_20502,N_20524);
nor U20789 (N_20789,N_20462,N_20580);
or U20790 (N_20790,N_20432,N_20442);
nand U20791 (N_20791,N_20400,N_20460);
nand U20792 (N_20792,N_20547,N_20491);
or U20793 (N_20793,N_20540,N_20499);
or U20794 (N_20794,N_20455,N_20423);
or U20795 (N_20795,N_20531,N_20551);
or U20796 (N_20796,N_20470,N_20508);
and U20797 (N_20797,N_20425,N_20561);
nor U20798 (N_20798,N_20572,N_20536);
nor U20799 (N_20799,N_20450,N_20445);
nor U20800 (N_20800,N_20784,N_20686);
nor U20801 (N_20801,N_20648,N_20763);
or U20802 (N_20802,N_20681,N_20690);
nand U20803 (N_20803,N_20651,N_20682);
xnor U20804 (N_20804,N_20691,N_20720);
nor U20805 (N_20805,N_20748,N_20647);
or U20806 (N_20806,N_20676,N_20755);
nand U20807 (N_20807,N_20621,N_20660);
nor U20808 (N_20808,N_20782,N_20793);
xor U20809 (N_20809,N_20738,N_20638);
and U20810 (N_20810,N_20749,N_20732);
nand U20811 (N_20811,N_20769,N_20722);
and U20812 (N_20812,N_20635,N_20649);
nand U20813 (N_20813,N_20679,N_20778);
xnor U20814 (N_20814,N_20699,N_20600);
xnor U20815 (N_20815,N_20764,N_20637);
nand U20816 (N_20816,N_20689,N_20770);
xor U20817 (N_20817,N_20767,N_20771);
or U20818 (N_20818,N_20614,N_20716);
xnor U20819 (N_20819,N_20605,N_20612);
nand U20820 (N_20820,N_20628,N_20677);
or U20821 (N_20821,N_20733,N_20757);
and U20822 (N_20822,N_20643,N_20777);
xnor U20823 (N_20823,N_20646,N_20606);
xor U20824 (N_20824,N_20729,N_20795);
nand U20825 (N_20825,N_20725,N_20665);
or U20826 (N_20826,N_20797,N_20630);
or U20827 (N_20827,N_20659,N_20666);
nand U20828 (N_20828,N_20655,N_20693);
and U20829 (N_20829,N_20708,N_20611);
and U20830 (N_20830,N_20624,N_20712);
and U20831 (N_20831,N_20607,N_20785);
nor U20832 (N_20832,N_20616,N_20726);
nor U20833 (N_20833,N_20730,N_20696);
and U20834 (N_20834,N_20751,N_20758);
nor U20835 (N_20835,N_20762,N_20634);
and U20836 (N_20836,N_20645,N_20623);
or U20837 (N_20837,N_20791,N_20672);
or U20838 (N_20838,N_20740,N_20724);
nand U20839 (N_20839,N_20663,N_20629);
nand U20840 (N_20840,N_20713,N_20653);
or U20841 (N_20841,N_20664,N_20773);
nor U20842 (N_20842,N_20711,N_20687);
nand U20843 (N_20843,N_20756,N_20737);
nand U20844 (N_20844,N_20741,N_20669);
nor U20845 (N_20845,N_20619,N_20610);
and U20846 (N_20846,N_20717,N_20787);
and U20847 (N_20847,N_20746,N_20658);
or U20848 (N_20848,N_20745,N_20703);
nand U20849 (N_20849,N_20674,N_20657);
xnor U20850 (N_20850,N_20639,N_20794);
nand U20851 (N_20851,N_20707,N_20644);
xnor U20852 (N_20852,N_20620,N_20625);
and U20853 (N_20853,N_20661,N_20723);
or U20854 (N_20854,N_20705,N_20709);
nor U20855 (N_20855,N_20772,N_20673);
nor U20856 (N_20856,N_20678,N_20714);
xnor U20857 (N_20857,N_20759,N_20692);
or U20858 (N_20858,N_20671,N_20721);
xnor U20859 (N_20859,N_20750,N_20798);
xnor U20860 (N_20860,N_20731,N_20704);
or U20861 (N_20861,N_20615,N_20783);
xor U20862 (N_20862,N_20727,N_20761);
and U20863 (N_20863,N_20631,N_20608);
nor U20864 (N_20864,N_20662,N_20667);
nand U20865 (N_20865,N_20670,N_20719);
and U20866 (N_20866,N_20779,N_20701);
nor U20867 (N_20867,N_20744,N_20752);
and U20868 (N_20868,N_20753,N_20685);
xnor U20869 (N_20869,N_20640,N_20695);
xor U20870 (N_20870,N_20618,N_20710);
nand U20871 (N_20871,N_20796,N_20680);
nand U20872 (N_20872,N_20684,N_20668);
nor U20873 (N_20873,N_20775,N_20765);
nand U20874 (N_20874,N_20697,N_20736);
or U20875 (N_20875,N_20754,N_20786);
nand U20876 (N_20876,N_20715,N_20700);
xor U20877 (N_20877,N_20768,N_20742);
nand U20878 (N_20878,N_20788,N_20641);
nor U20879 (N_20879,N_20780,N_20718);
nand U20880 (N_20880,N_20632,N_20766);
nand U20881 (N_20881,N_20734,N_20603);
nand U20882 (N_20882,N_20602,N_20683);
nor U20883 (N_20883,N_20636,N_20656);
nand U20884 (N_20884,N_20789,N_20654);
nand U20885 (N_20885,N_20617,N_20698);
or U20886 (N_20886,N_20781,N_20774);
or U20887 (N_20887,N_20743,N_20622);
nand U20888 (N_20888,N_20702,N_20604);
xor U20889 (N_20889,N_20652,N_20650);
or U20890 (N_20890,N_20747,N_20675);
nand U20891 (N_20891,N_20790,N_20626);
xnor U20892 (N_20892,N_20735,N_20694);
xnor U20893 (N_20893,N_20627,N_20642);
and U20894 (N_20894,N_20792,N_20613);
xnor U20895 (N_20895,N_20633,N_20776);
or U20896 (N_20896,N_20706,N_20609);
nand U20897 (N_20897,N_20688,N_20739);
nand U20898 (N_20898,N_20728,N_20760);
or U20899 (N_20899,N_20601,N_20799);
nor U20900 (N_20900,N_20613,N_20623);
xor U20901 (N_20901,N_20630,N_20747);
or U20902 (N_20902,N_20793,N_20736);
xnor U20903 (N_20903,N_20615,N_20601);
or U20904 (N_20904,N_20690,N_20746);
nor U20905 (N_20905,N_20746,N_20618);
nand U20906 (N_20906,N_20731,N_20763);
nor U20907 (N_20907,N_20742,N_20719);
nor U20908 (N_20908,N_20760,N_20638);
nand U20909 (N_20909,N_20616,N_20754);
and U20910 (N_20910,N_20749,N_20692);
or U20911 (N_20911,N_20644,N_20716);
and U20912 (N_20912,N_20622,N_20795);
nand U20913 (N_20913,N_20740,N_20779);
or U20914 (N_20914,N_20623,N_20678);
or U20915 (N_20915,N_20798,N_20747);
xor U20916 (N_20916,N_20648,N_20752);
or U20917 (N_20917,N_20701,N_20681);
xor U20918 (N_20918,N_20774,N_20730);
xor U20919 (N_20919,N_20655,N_20678);
nand U20920 (N_20920,N_20615,N_20610);
xor U20921 (N_20921,N_20663,N_20794);
and U20922 (N_20922,N_20676,N_20750);
xnor U20923 (N_20923,N_20703,N_20626);
or U20924 (N_20924,N_20604,N_20775);
nand U20925 (N_20925,N_20619,N_20627);
xnor U20926 (N_20926,N_20654,N_20665);
xnor U20927 (N_20927,N_20641,N_20763);
and U20928 (N_20928,N_20760,N_20778);
nor U20929 (N_20929,N_20722,N_20682);
and U20930 (N_20930,N_20732,N_20646);
nor U20931 (N_20931,N_20774,N_20625);
nor U20932 (N_20932,N_20650,N_20714);
xor U20933 (N_20933,N_20744,N_20720);
nand U20934 (N_20934,N_20753,N_20734);
and U20935 (N_20935,N_20735,N_20795);
xnor U20936 (N_20936,N_20741,N_20770);
nand U20937 (N_20937,N_20728,N_20631);
nand U20938 (N_20938,N_20705,N_20701);
and U20939 (N_20939,N_20676,N_20629);
nor U20940 (N_20940,N_20646,N_20608);
or U20941 (N_20941,N_20630,N_20690);
xnor U20942 (N_20942,N_20768,N_20799);
or U20943 (N_20943,N_20660,N_20711);
nor U20944 (N_20944,N_20643,N_20734);
xnor U20945 (N_20945,N_20644,N_20621);
xnor U20946 (N_20946,N_20742,N_20741);
nand U20947 (N_20947,N_20739,N_20693);
xor U20948 (N_20948,N_20691,N_20687);
nand U20949 (N_20949,N_20782,N_20787);
xor U20950 (N_20950,N_20636,N_20757);
or U20951 (N_20951,N_20645,N_20780);
nor U20952 (N_20952,N_20714,N_20637);
nor U20953 (N_20953,N_20738,N_20602);
nor U20954 (N_20954,N_20729,N_20794);
and U20955 (N_20955,N_20737,N_20663);
or U20956 (N_20956,N_20703,N_20772);
nand U20957 (N_20957,N_20703,N_20708);
nand U20958 (N_20958,N_20647,N_20672);
nor U20959 (N_20959,N_20783,N_20617);
or U20960 (N_20960,N_20770,N_20610);
or U20961 (N_20961,N_20604,N_20792);
and U20962 (N_20962,N_20647,N_20747);
nand U20963 (N_20963,N_20610,N_20734);
nor U20964 (N_20964,N_20605,N_20780);
or U20965 (N_20965,N_20620,N_20747);
nand U20966 (N_20966,N_20750,N_20636);
nand U20967 (N_20967,N_20640,N_20602);
and U20968 (N_20968,N_20628,N_20758);
nor U20969 (N_20969,N_20607,N_20698);
and U20970 (N_20970,N_20669,N_20719);
nand U20971 (N_20971,N_20724,N_20647);
nor U20972 (N_20972,N_20729,N_20733);
nor U20973 (N_20973,N_20650,N_20611);
nand U20974 (N_20974,N_20693,N_20607);
nand U20975 (N_20975,N_20752,N_20746);
nand U20976 (N_20976,N_20735,N_20789);
nor U20977 (N_20977,N_20602,N_20721);
and U20978 (N_20978,N_20710,N_20624);
xor U20979 (N_20979,N_20795,N_20684);
or U20980 (N_20980,N_20650,N_20614);
and U20981 (N_20981,N_20637,N_20691);
and U20982 (N_20982,N_20758,N_20650);
xnor U20983 (N_20983,N_20772,N_20677);
nand U20984 (N_20984,N_20719,N_20629);
xnor U20985 (N_20985,N_20702,N_20779);
nor U20986 (N_20986,N_20685,N_20773);
nor U20987 (N_20987,N_20669,N_20673);
nand U20988 (N_20988,N_20654,N_20750);
nand U20989 (N_20989,N_20620,N_20736);
nand U20990 (N_20990,N_20718,N_20623);
nor U20991 (N_20991,N_20684,N_20765);
nand U20992 (N_20992,N_20605,N_20729);
nor U20993 (N_20993,N_20709,N_20726);
or U20994 (N_20994,N_20605,N_20678);
nor U20995 (N_20995,N_20665,N_20617);
or U20996 (N_20996,N_20611,N_20655);
nand U20997 (N_20997,N_20660,N_20664);
xnor U20998 (N_20998,N_20646,N_20760);
nand U20999 (N_20999,N_20743,N_20612);
xor U21000 (N_21000,N_20952,N_20958);
nand U21001 (N_21001,N_20947,N_20920);
nand U21002 (N_21002,N_20909,N_20933);
nor U21003 (N_21003,N_20995,N_20986);
nand U21004 (N_21004,N_20969,N_20837);
nor U21005 (N_21005,N_20859,N_20804);
nand U21006 (N_21006,N_20916,N_20882);
or U21007 (N_21007,N_20857,N_20993);
or U21008 (N_21008,N_20898,N_20824);
nor U21009 (N_21009,N_20818,N_20917);
nand U21010 (N_21010,N_20809,N_20904);
xnor U21011 (N_21011,N_20800,N_20825);
and U21012 (N_21012,N_20919,N_20862);
or U21013 (N_21013,N_20983,N_20937);
nor U21014 (N_21014,N_20901,N_20820);
or U21015 (N_21015,N_20812,N_20990);
or U21016 (N_21016,N_20959,N_20900);
nand U21017 (N_21017,N_20912,N_20830);
nor U21018 (N_21018,N_20902,N_20839);
xor U21019 (N_21019,N_20838,N_20895);
nor U21020 (N_21020,N_20842,N_20805);
nand U21021 (N_21021,N_20999,N_20935);
nor U21022 (N_21022,N_20954,N_20930);
and U21023 (N_21023,N_20946,N_20929);
xor U21024 (N_21024,N_20996,N_20973);
nor U21025 (N_21025,N_20994,N_20861);
nor U21026 (N_21026,N_20884,N_20876);
nand U21027 (N_21027,N_20807,N_20829);
nand U21028 (N_21028,N_20871,N_20803);
or U21029 (N_21029,N_20906,N_20892);
nand U21030 (N_21030,N_20915,N_20890);
nand U21031 (N_21031,N_20877,N_20921);
and U21032 (N_21032,N_20970,N_20887);
nand U21033 (N_21033,N_20950,N_20982);
and U21034 (N_21034,N_20963,N_20940);
or U21035 (N_21035,N_20886,N_20865);
and U21036 (N_21036,N_20891,N_20849);
nor U21037 (N_21037,N_20957,N_20932);
and U21038 (N_21038,N_20908,N_20945);
and U21039 (N_21039,N_20980,N_20855);
nor U21040 (N_21040,N_20948,N_20944);
and U21041 (N_21041,N_20971,N_20831);
nor U21042 (N_21042,N_20860,N_20905);
nand U21043 (N_21043,N_20863,N_20897);
and U21044 (N_21044,N_20806,N_20864);
xnor U21045 (N_21045,N_20956,N_20853);
xor U21046 (N_21046,N_20894,N_20850);
xnor U21047 (N_21047,N_20974,N_20813);
nand U21048 (N_21048,N_20827,N_20907);
xnor U21049 (N_21049,N_20832,N_20989);
nand U21050 (N_21050,N_20841,N_20997);
and U21051 (N_21051,N_20939,N_20815);
xnor U21052 (N_21052,N_20913,N_20873);
nand U21053 (N_21053,N_20979,N_20975);
nor U21054 (N_21054,N_20802,N_20869);
or U21055 (N_21055,N_20918,N_20936);
or U21056 (N_21056,N_20914,N_20903);
or U21057 (N_21057,N_20962,N_20835);
nor U21058 (N_21058,N_20927,N_20978);
xnor U21059 (N_21059,N_20981,N_20953);
nand U21060 (N_21060,N_20867,N_20972);
nand U21061 (N_21061,N_20987,N_20836);
xor U21062 (N_21062,N_20833,N_20931);
nand U21063 (N_21063,N_20883,N_20868);
nand U21064 (N_21064,N_20922,N_20885);
and U21065 (N_21065,N_20819,N_20880);
nand U21066 (N_21066,N_20888,N_20845);
xnor U21067 (N_21067,N_20872,N_20874);
nand U21068 (N_21068,N_20977,N_20928);
and U21069 (N_21069,N_20817,N_20961);
nand U21070 (N_21070,N_20960,N_20801);
nand U21071 (N_21071,N_20889,N_20878);
or U21072 (N_21072,N_20816,N_20828);
and U21073 (N_21073,N_20843,N_20847);
xor U21074 (N_21074,N_20964,N_20976);
nand U21075 (N_21075,N_20854,N_20879);
or U21076 (N_21076,N_20967,N_20893);
xor U21077 (N_21077,N_20814,N_20943);
or U21078 (N_21078,N_20984,N_20851);
nand U21079 (N_21079,N_20949,N_20941);
nand U21080 (N_21080,N_20966,N_20934);
nor U21081 (N_21081,N_20911,N_20992);
nor U21082 (N_21082,N_20808,N_20810);
xnor U21083 (N_21083,N_20991,N_20881);
xnor U21084 (N_21084,N_20858,N_20968);
nand U21085 (N_21085,N_20985,N_20923);
nor U21086 (N_21086,N_20925,N_20910);
and U21087 (N_21087,N_20844,N_20965);
nor U21088 (N_21088,N_20846,N_20998);
nand U21089 (N_21089,N_20899,N_20826);
nor U21090 (N_21090,N_20870,N_20924);
nor U21091 (N_21091,N_20834,N_20822);
and U21092 (N_21092,N_20823,N_20848);
and U21093 (N_21093,N_20821,N_20875);
and U21094 (N_21094,N_20896,N_20852);
xor U21095 (N_21095,N_20866,N_20942);
nor U21096 (N_21096,N_20811,N_20988);
nand U21097 (N_21097,N_20955,N_20840);
xor U21098 (N_21098,N_20926,N_20938);
nand U21099 (N_21099,N_20951,N_20856);
or U21100 (N_21100,N_20817,N_20815);
or U21101 (N_21101,N_20842,N_20950);
xor U21102 (N_21102,N_20964,N_20870);
xor U21103 (N_21103,N_20973,N_20892);
nor U21104 (N_21104,N_20817,N_20931);
nand U21105 (N_21105,N_20986,N_20820);
or U21106 (N_21106,N_20883,N_20967);
and U21107 (N_21107,N_20938,N_20853);
xnor U21108 (N_21108,N_20825,N_20909);
nand U21109 (N_21109,N_20959,N_20955);
or U21110 (N_21110,N_20868,N_20973);
nand U21111 (N_21111,N_20800,N_20898);
or U21112 (N_21112,N_20980,N_20833);
xor U21113 (N_21113,N_20955,N_20805);
xnor U21114 (N_21114,N_20954,N_20806);
and U21115 (N_21115,N_20822,N_20827);
nand U21116 (N_21116,N_20985,N_20894);
and U21117 (N_21117,N_20962,N_20846);
nor U21118 (N_21118,N_20920,N_20953);
xnor U21119 (N_21119,N_20923,N_20959);
and U21120 (N_21120,N_20930,N_20880);
and U21121 (N_21121,N_20858,N_20888);
and U21122 (N_21122,N_20902,N_20802);
xnor U21123 (N_21123,N_20976,N_20897);
and U21124 (N_21124,N_20904,N_20858);
xnor U21125 (N_21125,N_20881,N_20873);
xor U21126 (N_21126,N_20970,N_20938);
nor U21127 (N_21127,N_20820,N_20987);
nand U21128 (N_21128,N_20949,N_20807);
and U21129 (N_21129,N_20845,N_20963);
nor U21130 (N_21130,N_20922,N_20933);
or U21131 (N_21131,N_20812,N_20952);
or U21132 (N_21132,N_20950,N_20953);
nor U21133 (N_21133,N_20965,N_20843);
xor U21134 (N_21134,N_20830,N_20974);
and U21135 (N_21135,N_20921,N_20930);
nor U21136 (N_21136,N_20808,N_20984);
and U21137 (N_21137,N_20861,N_20801);
nand U21138 (N_21138,N_20973,N_20818);
nand U21139 (N_21139,N_20989,N_20877);
or U21140 (N_21140,N_20801,N_20885);
xnor U21141 (N_21141,N_20823,N_20871);
and U21142 (N_21142,N_20904,N_20981);
or U21143 (N_21143,N_20972,N_20891);
or U21144 (N_21144,N_20962,N_20967);
and U21145 (N_21145,N_20838,N_20816);
and U21146 (N_21146,N_20845,N_20890);
or U21147 (N_21147,N_20989,N_20998);
nor U21148 (N_21148,N_20847,N_20946);
xnor U21149 (N_21149,N_20960,N_20869);
and U21150 (N_21150,N_20851,N_20990);
xnor U21151 (N_21151,N_20892,N_20853);
nor U21152 (N_21152,N_20823,N_20997);
or U21153 (N_21153,N_20931,N_20946);
nand U21154 (N_21154,N_20875,N_20934);
nor U21155 (N_21155,N_20939,N_20919);
xor U21156 (N_21156,N_20842,N_20814);
xor U21157 (N_21157,N_20809,N_20836);
or U21158 (N_21158,N_20832,N_20967);
or U21159 (N_21159,N_20818,N_20924);
xnor U21160 (N_21160,N_20935,N_20915);
nor U21161 (N_21161,N_20923,N_20841);
nor U21162 (N_21162,N_20975,N_20856);
and U21163 (N_21163,N_20822,N_20813);
nor U21164 (N_21164,N_20976,N_20995);
and U21165 (N_21165,N_20936,N_20835);
xor U21166 (N_21166,N_20957,N_20905);
nor U21167 (N_21167,N_20854,N_20907);
and U21168 (N_21168,N_20888,N_20952);
and U21169 (N_21169,N_20809,N_20942);
or U21170 (N_21170,N_20926,N_20883);
xnor U21171 (N_21171,N_20955,N_20988);
nor U21172 (N_21172,N_20921,N_20910);
nor U21173 (N_21173,N_20825,N_20948);
or U21174 (N_21174,N_20915,N_20846);
nand U21175 (N_21175,N_20910,N_20820);
nand U21176 (N_21176,N_20957,N_20935);
or U21177 (N_21177,N_20892,N_20850);
nor U21178 (N_21178,N_20889,N_20974);
or U21179 (N_21179,N_20812,N_20865);
nor U21180 (N_21180,N_20911,N_20871);
xnor U21181 (N_21181,N_20998,N_20991);
or U21182 (N_21182,N_20913,N_20902);
or U21183 (N_21183,N_20954,N_20840);
or U21184 (N_21184,N_20845,N_20856);
or U21185 (N_21185,N_20839,N_20979);
xnor U21186 (N_21186,N_20990,N_20861);
or U21187 (N_21187,N_20876,N_20883);
nand U21188 (N_21188,N_20937,N_20884);
or U21189 (N_21189,N_20983,N_20813);
and U21190 (N_21190,N_20907,N_20848);
nor U21191 (N_21191,N_20951,N_20849);
xnor U21192 (N_21192,N_20928,N_20937);
xor U21193 (N_21193,N_20857,N_20879);
nor U21194 (N_21194,N_20922,N_20899);
or U21195 (N_21195,N_20924,N_20928);
nor U21196 (N_21196,N_20875,N_20939);
or U21197 (N_21197,N_20828,N_20973);
nor U21198 (N_21198,N_20975,N_20826);
and U21199 (N_21199,N_20919,N_20977);
nor U21200 (N_21200,N_21136,N_21053);
and U21201 (N_21201,N_21039,N_21092);
nand U21202 (N_21202,N_21001,N_21095);
and U21203 (N_21203,N_21189,N_21024);
nor U21204 (N_21204,N_21131,N_21052);
nand U21205 (N_21205,N_21132,N_21101);
or U21206 (N_21206,N_21094,N_21013);
nand U21207 (N_21207,N_21062,N_21076);
nor U21208 (N_21208,N_21198,N_21012);
nor U21209 (N_21209,N_21167,N_21086);
xor U21210 (N_21210,N_21152,N_21009);
xor U21211 (N_21211,N_21185,N_21058);
nor U21212 (N_21212,N_21111,N_21083);
nor U21213 (N_21213,N_21125,N_21133);
nor U21214 (N_21214,N_21134,N_21066);
xor U21215 (N_21215,N_21154,N_21044);
xnor U21216 (N_21216,N_21129,N_21141);
and U21217 (N_21217,N_21188,N_21192);
nor U21218 (N_21218,N_21117,N_21000);
and U21219 (N_21219,N_21183,N_21078);
xor U21220 (N_21220,N_21072,N_21156);
nor U21221 (N_21221,N_21075,N_21006);
or U21222 (N_21222,N_21182,N_21116);
or U21223 (N_21223,N_21140,N_21104);
and U21224 (N_21224,N_21080,N_21153);
xnor U21225 (N_21225,N_21191,N_21089);
nand U21226 (N_21226,N_21187,N_21130);
or U21227 (N_21227,N_21181,N_21081);
nand U21228 (N_21228,N_21020,N_21109);
or U21229 (N_21229,N_21060,N_21149);
nor U21230 (N_21230,N_21096,N_21110);
nor U21231 (N_21231,N_21157,N_21138);
nor U21232 (N_21232,N_21145,N_21139);
nor U21233 (N_21233,N_21033,N_21025);
or U21234 (N_21234,N_21023,N_21056);
or U21235 (N_21235,N_21151,N_21107);
nand U21236 (N_21236,N_21175,N_21073);
xnor U21237 (N_21237,N_21010,N_21160);
or U21238 (N_21238,N_21091,N_21158);
nand U21239 (N_21239,N_21035,N_21079);
xnor U21240 (N_21240,N_21098,N_21017);
nand U21241 (N_21241,N_21174,N_21124);
nand U21242 (N_21242,N_21047,N_21100);
xnor U21243 (N_21243,N_21041,N_21074);
nand U21244 (N_21244,N_21197,N_21128);
or U21245 (N_21245,N_21067,N_21176);
and U21246 (N_21246,N_21172,N_21122);
nand U21247 (N_21247,N_21199,N_21045);
xnor U21248 (N_21248,N_21150,N_21050);
xor U21249 (N_21249,N_21036,N_21088);
nand U21250 (N_21250,N_21071,N_21037);
or U21251 (N_21251,N_21031,N_21030);
nor U21252 (N_21252,N_21142,N_21126);
and U21253 (N_21253,N_21070,N_21105);
and U21254 (N_21254,N_21026,N_21097);
and U21255 (N_21255,N_21170,N_21195);
nor U21256 (N_21256,N_21169,N_21121);
or U21257 (N_21257,N_21190,N_21103);
or U21258 (N_21258,N_21148,N_21051);
nor U21259 (N_21259,N_21173,N_21042);
or U21260 (N_21260,N_21146,N_21108);
xnor U21261 (N_21261,N_21008,N_21038);
or U21262 (N_21262,N_21043,N_21165);
and U21263 (N_21263,N_21135,N_21163);
or U21264 (N_21264,N_21171,N_21159);
and U21265 (N_21265,N_21114,N_21179);
nor U21266 (N_21266,N_21049,N_21194);
xor U21267 (N_21267,N_21063,N_21028);
xnor U21268 (N_21268,N_21137,N_21143);
or U21269 (N_21269,N_21064,N_21155);
or U21270 (N_21270,N_21016,N_21102);
nand U21271 (N_21271,N_21048,N_21123);
or U21272 (N_21272,N_21082,N_21164);
and U21273 (N_21273,N_21004,N_21077);
nand U21274 (N_21274,N_21144,N_21115);
nand U21275 (N_21275,N_21018,N_21034);
xnor U21276 (N_21276,N_21120,N_21005);
and U21277 (N_21277,N_21068,N_21022);
or U21278 (N_21278,N_21055,N_21127);
nor U21279 (N_21279,N_21106,N_21166);
and U21280 (N_21280,N_21113,N_21011);
nor U21281 (N_21281,N_21040,N_21002);
or U21282 (N_21282,N_21046,N_21087);
xnor U21283 (N_21283,N_21093,N_21065);
or U21284 (N_21284,N_21090,N_21186);
and U21285 (N_21285,N_21014,N_21003);
nand U21286 (N_21286,N_21119,N_21084);
nor U21287 (N_21287,N_21054,N_21168);
xor U21288 (N_21288,N_21193,N_21029);
or U21289 (N_21289,N_21059,N_21032);
nor U21290 (N_21290,N_21015,N_21027);
nand U21291 (N_21291,N_21021,N_21099);
or U21292 (N_21292,N_21112,N_21184);
and U21293 (N_21293,N_21069,N_21180);
nand U21294 (N_21294,N_21007,N_21161);
xnor U21295 (N_21295,N_21118,N_21147);
nor U21296 (N_21296,N_21162,N_21019);
xnor U21297 (N_21297,N_21177,N_21057);
nor U21298 (N_21298,N_21178,N_21085);
nor U21299 (N_21299,N_21196,N_21061);
or U21300 (N_21300,N_21187,N_21175);
and U21301 (N_21301,N_21161,N_21058);
and U21302 (N_21302,N_21027,N_21142);
nand U21303 (N_21303,N_21116,N_21065);
or U21304 (N_21304,N_21134,N_21140);
or U21305 (N_21305,N_21065,N_21080);
nor U21306 (N_21306,N_21143,N_21020);
nor U21307 (N_21307,N_21030,N_21018);
xnor U21308 (N_21308,N_21038,N_21124);
and U21309 (N_21309,N_21191,N_21021);
nand U21310 (N_21310,N_21131,N_21066);
nor U21311 (N_21311,N_21156,N_21111);
and U21312 (N_21312,N_21180,N_21125);
nor U21313 (N_21313,N_21048,N_21178);
nor U21314 (N_21314,N_21005,N_21052);
nor U21315 (N_21315,N_21021,N_21039);
and U21316 (N_21316,N_21051,N_21034);
or U21317 (N_21317,N_21090,N_21028);
nand U21318 (N_21318,N_21020,N_21189);
nand U21319 (N_21319,N_21069,N_21083);
and U21320 (N_21320,N_21129,N_21084);
and U21321 (N_21321,N_21107,N_21116);
nor U21322 (N_21322,N_21027,N_21055);
nor U21323 (N_21323,N_21081,N_21133);
or U21324 (N_21324,N_21034,N_21123);
or U21325 (N_21325,N_21187,N_21106);
and U21326 (N_21326,N_21053,N_21161);
or U21327 (N_21327,N_21003,N_21053);
xnor U21328 (N_21328,N_21166,N_21128);
xnor U21329 (N_21329,N_21020,N_21065);
nor U21330 (N_21330,N_21170,N_21021);
and U21331 (N_21331,N_21134,N_21151);
xnor U21332 (N_21332,N_21125,N_21001);
xor U21333 (N_21333,N_21098,N_21143);
and U21334 (N_21334,N_21186,N_21058);
nor U21335 (N_21335,N_21129,N_21013);
and U21336 (N_21336,N_21134,N_21075);
nand U21337 (N_21337,N_21005,N_21114);
nand U21338 (N_21338,N_21093,N_21013);
or U21339 (N_21339,N_21049,N_21004);
nand U21340 (N_21340,N_21078,N_21021);
nand U21341 (N_21341,N_21100,N_21072);
nand U21342 (N_21342,N_21135,N_21104);
or U21343 (N_21343,N_21063,N_21020);
nor U21344 (N_21344,N_21186,N_21012);
nand U21345 (N_21345,N_21102,N_21046);
xnor U21346 (N_21346,N_21121,N_21120);
nand U21347 (N_21347,N_21184,N_21165);
nand U21348 (N_21348,N_21040,N_21105);
and U21349 (N_21349,N_21122,N_21033);
xnor U21350 (N_21350,N_21129,N_21115);
xnor U21351 (N_21351,N_21031,N_21119);
nand U21352 (N_21352,N_21008,N_21022);
or U21353 (N_21353,N_21016,N_21005);
or U21354 (N_21354,N_21183,N_21138);
or U21355 (N_21355,N_21037,N_21112);
xor U21356 (N_21356,N_21076,N_21067);
and U21357 (N_21357,N_21055,N_21138);
and U21358 (N_21358,N_21025,N_21140);
nand U21359 (N_21359,N_21037,N_21097);
nand U21360 (N_21360,N_21023,N_21130);
xor U21361 (N_21361,N_21057,N_21125);
nand U21362 (N_21362,N_21034,N_21033);
nor U21363 (N_21363,N_21134,N_21181);
xor U21364 (N_21364,N_21141,N_21162);
nand U21365 (N_21365,N_21090,N_21187);
nor U21366 (N_21366,N_21159,N_21031);
nor U21367 (N_21367,N_21039,N_21006);
and U21368 (N_21368,N_21075,N_21147);
and U21369 (N_21369,N_21026,N_21104);
nand U21370 (N_21370,N_21116,N_21129);
nor U21371 (N_21371,N_21116,N_21190);
nand U21372 (N_21372,N_21048,N_21031);
and U21373 (N_21373,N_21072,N_21163);
or U21374 (N_21374,N_21169,N_21082);
nor U21375 (N_21375,N_21068,N_21186);
nand U21376 (N_21376,N_21102,N_21170);
nor U21377 (N_21377,N_21014,N_21119);
nor U21378 (N_21378,N_21095,N_21036);
nor U21379 (N_21379,N_21068,N_21076);
nor U21380 (N_21380,N_21069,N_21138);
nand U21381 (N_21381,N_21031,N_21060);
xor U21382 (N_21382,N_21006,N_21167);
nand U21383 (N_21383,N_21161,N_21039);
xnor U21384 (N_21384,N_21044,N_21022);
xor U21385 (N_21385,N_21155,N_21195);
nand U21386 (N_21386,N_21053,N_21182);
nor U21387 (N_21387,N_21004,N_21057);
or U21388 (N_21388,N_21108,N_21041);
nor U21389 (N_21389,N_21113,N_21047);
nand U21390 (N_21390,N_21159,N_21041);
nor U21391 (N_21391,N_21011,N_21102);
or U21392 (N_21392,N_21087,N_21135);
xnor U21393 (N_21393,N_21099,N_21122);
xnor U21394 (N_21394,N_21134,N_21061);
and U21395 (N_21395,N_21188,N_21116);
or U21396 (N_21396,N_21080,N_21061);
xor U21397 (N_21397,N_21084,N_21016);
or U21398 (N_21398,N_21144,N_21036);
and U21399 (N_21399,N_21163,N_21006);
xnor U21400 (N_21400,N_21252,N_21239);
xnor U21401 (N_21401,N_21386,N_21201);
and U21402 (N_21402,N_21246,N_21249);
nor U21403 (N_21403,N_21248,N_21225);
nand U21404 (N_21404,N_21357,N_21266);
and U21405 (N_21405,N_21318,N_21341);
and U21406 (N_21406,N_21399,N_21378);
or U21407 (N_21407,N_21298,N_21307);
nor U21408 (N_21408,N_21329,N_21236);
nor U21409 (N_21409,N_21268,N_21370);
nor U21410 (N_21410,N_21313,N_21308);
or U21411 (N_21411,N_21243,N_21288);
and U21412 (N_21412,N_21227,N_21258);
xnor U21413 (N_21413,N_21398,N_21212);
nor U21414 (N_21414,N_21352,N_21218);
nand U21415 (N_21415,N_21397,N_21211);
nand U21416 (N_21416,N_21270,N_21247);
nor U21417 (N_21417,N_21337,N_21371);
nand U21418 (N_21418,N_21338,N_21328);
nor U21419 (N_21419,N_21215,N_21257);
nand U21420 (N_21420,N_21217,N_21299);
and U21421 (N_21421,N_21250,N_21204);
nor U21422 (N_21422,N_21346,N_21336);
or U21423 (N_21423,N_21222,N_21232);
and U21424 (N_21424,N_21332,N_21344);
nand U21425 (N_21425,N_21335,N_21278);
or U21426 (N_21426,N_21315,N_21210);
nor U21427 (N_21427,N_21368,N_21384);
and U21428 (N_21428,N_21383,N_21343);
and U21429 (N_21429,N_21291,N_21230);
nand U21430 (N_21430,N_21297,N_21234);
nor U21431 (N_21431,N_21260,N_21381);
xor U21432 (N_21432,N_21359,N_21231);
and U21433 (N_21433,N_21203,N_21327);
nor U21434 (N_21434,N_21382,N_21209);
and U21435 (N_21435,N_21285,N_21206);
xnor U21436 (N_21436,N_21290,N_21316);
nand U21437 (N_21437,N_21235,N_21224);
xnor U21438 (N_21438,N_21309,N_21342);
or U21439 (N_21439,N_21385,N_21275);
or U21440 (N_21440,N_21301,N_21241);
and U21441 (N_21441,N_21255,N_21366);
and U21442 (N_21442,N_21395,N_21334);
nor U21443 (N_21443,N_21281,N_21394);
or U21444 (N_21444,N_21393,N_21286);
or U21445 (N_21445,N_21311,N_21330);
nand U21446 (N_21446,N_21363,N_21277);
or U21447 (N_21447,N_21253,N_21279);
nand U21448 (N_21448,N_21282,N_21237);
nor U21449 (N_21449,N_21272,N_21353);
nor U21450 (N_21450,N_21347,N_21320);
xnor U21451 (N_21451,N_21223,N_21396);
xor U21452 (N_21452,N_21294,N_21333);
or U21453 (N_21453,N_21388,N_21207);
nor U21454 (N_21454,N_21391,N_21304);
xor U21455 (N_21455,N_21245,N_21273);
and U21456 (N_21456,N_21379,N_21295);
and U21457 (N_21457,N_21263,N_21375);
nand U21458 (N_21458,N_21303,N_21349);
nor U21459 (N_21459,N_21360,N_21305);
or U21460 (N_21460,N_21372,N_21262);
nor U21461 (N_21461,N_21221,N_21358);
and U21462 (N_21462,N_21254,N_21271);
nand U21463 (N_21463,N_21226,N_21233);
nor U21464 (N_21464,N_21373,N_21369);
or U21465 (N_21465,N_21259,N_21265);
xor U21466 (N_21466,N_21293,N_21300);
or U21467 (N_21467,N_21362,N_21280);
nand U21468 (N_21468,N_21242,N_21322);
nand U21469 (N_21469,N_21340,N_21216);
or U21470 (N_21470,N_21261,N_21377);
and U21471 (N_21471,N_21351,N_21365);
and U21472 (N_21472,N_21228,N_21376);
nor U21473 (N_21473,N_21380,N_21350);
nand U21474 (N_21474,N_21339,N_21264);
or U21475 (N_21475,N_21219,N_21345);
or U21476 (N_21476,N_21387,N_21367);
or U21477 (N_21477,N_21205,N_21356);
nand U21478 (N_21478,N_21251,N_21244);
xnor U21479 (N_21479,N_21287,N_21321);
or U21480 (N_21480,N_21326,N_21317);
and U21481 (N_21481,N_21213,N_21389);
nor U21482 (N_21482,N_21289,N_21283);
or U21483 (N_21483,N_21331,N_21240);
nand U21484 (N_21484,N_21323,N_21276);
nor U21485 (N_21485,N_21229,N_21296);
and U21486 (N_21486,N_21390,N_21312);
nand U21487 (N_21487,N_21200,N_21361);
xnor U21488 (N_21488,N_21214,N_21319);
and U21489 (N_21489,N_21364,N_21269);
or U21490 (N_21490,N_21355,N_21374);
or U21491 (N_21491,N_21392,N_21310);
xnor U21492 (N_21492,N_21220,N_21274);
xor U21493 (N_21493,N_21208,N_21238);
nor U21494 (N_21494,N_21325,N_21348);
nor U21495 (N_21495,N_21292,N_21306);
xor U21496 (N_21496,N_21256,N_21302);
or U21497 (N_21497,N_21284,N_21267);
or U21498 (N_21498,N_21324,N_21202);
and U21499 (N_21499,N_21314,N_21354);
or U21500 (N_21500,N_21219,N_21260);
and U21501 (N_21501,N_21365,N_21221);
nand U21502 (N_21502,N_21352,N_21324);
nor U21503 (N_21503,N_21354,N_21397);
xor U21504 (N_21504,N_21370,N_21305);
and U21505 (N_21505,N_21281,N_21354);
nand U21506 (N_21506,N_21296,N_21207);
or U21507 (N_21507,N_21323,N_21322);
nand U21508 (N_21508,N_21342,N_21369);
nand U21509 (N_21509,N_21211,N_21354);
xnor U21510 (N_21510,N_21227,N_21318);
nand U21511 (N_21511,N_21276,N_21266);
and U21512 (N_21512,N_21262,N_21395);
nor U21513 (N_21513,N_21220,N_21308);
and U21514 (N_21514,N_21280,N_21372);
and U21515 (N_21515,N_21283,N_21244);
or U21516 (N_21516,N_21214,N_21387);
nand U21517 (N_21517,N_21241,N_21262);
xor U21518 (N_21518,N_21294,N_21368);
nor U21519 (N_21519,N_21226,N_21333);
or U21520 (N_21520,N_21333,N_21220);
nand U21521 (N_21521,N_21326,N_21390);
nor U21522 (N_21522,N_21345,N_21321);
nor U21523 (N_21523,N_21234,N_21254);
nor U21524 (N_21524,N_21324,N_21380);
or U21525 (N_21525,N_21289,N_21204);
xor U21526 (N_21526,N_21318,N_21320);
nand U21527 (N_21527,N_21302,N_21365);
and U21528 (N_21528,N_21351,N_21336);
nor U21529 (N_21529,N_21300,N_21284);
nor U21530 (N_21530,N_21350,N_21353);
nand U21531 (N_21531,N_21204,N_21371);
nor U21532 (N_21532,N_21317,N_21267);
nand U21533 (N_21533,N_21295,N_21331);
and U21534 (N_21534,N_21270,N_21311);
and U21535 (N_21535,N_21356,N_21343);
or U21536 (N_21536,N_21209,N_21345);
xor U21537 (N_21537,N_21296,N_21365);
and U21538 (N_21538,N_21230,N_21268);
nand U21539 (N_21539,N_21349,N_21234);
and U21540 (N_21540,N_21386,N_21374);
or U21541 (N_21541,N_21351,N_21379);
or U21542 (N_21542,N_21323,N_21321);
nand U21543 (N_21543,N_21303,N_21390);
xnor U21544 (N_21544,N_21241,N_21268);
and U21545 (N_21545,N_21234,N_21278);
and U21546 (N_21546,N_21335,N_21398);
or U21547 (N_21547,N_21253,N_21312);
and U21548 (N_21548,N_21244,N_21385);
xor U21549 (N_21549,N_21259,N_21285);
nand U21550 (N_21550,N_21395,N_21372);
and U21551 (N_21551,N_21268,N_21310);
nand U21552 (N_21552,N_21219,N_21333);
nor U21553 (N_21553,N_21274,N_21308);
nor U21554 (N_21554,N_21248,N_21373);
xnor U21555 (N_21555,N_21289,N_21372);
or U21556 (N_21556,N_21387,N_21222);
nand U21557 (N_21557,N_21377,N_21225);
nor U21558 (N_21558,N_21232,N_21231);
xnor U21559 (N_21559,N_21339,N_21222);
nor U21560 (N_21560,N_21380,N_21236);
nand U21561 (N_21561,N_21339,N_21207);
or U21562 (N_21562,N_21254,N_21286);
nor U21563 (N_21563,N_21226,N_21394);
or U21564 (N_21564,N_21319,N_21249);
and U21565 (N_21565,N_21291,N_21377);
xnor U21566 (N_21566,N_21300,N_21389);
and U21567 (N_21567,N_21374,N_21340);
nand U21568 (N_21568,N_21361,N_21267);
nor U21569 (N_21569,N_21397,N_21361);
nor U21570 (N_21570,N_21315,N_21385);
xor U21571 (N_21571,N_21203,N_21336);
xor U21572 (N_21572,N_21388,N_21249);
nor U21573 (N_21573,N_21385,N_21316);
or U21574 (N_21574,N_21304,N_21363);
nand U21575 (N_21575,N_21224,N_21267);
nor U21576 (N_21576,N_21327,N_21319);
nor U21577 (N_21577,N_21283,N_21298);
nand U21578 (N_21578,N_21226,N_21288);
and U21579 (N_21579,N_21335,N_21342);
or U21580 (N_21580,N_21374,N_21296);
nand U21581 (N_21581,N_21237,N_21225);
or U21582 (N_21582,N_21260,N_21258);
or U21583 (N_21583,N_21212,N_21213);
nor U21584 (N_21584,N_21319,N_21331);
xnor U21585 (N_21585,N_21266,N_21234);
nand U21586 (N_21586,N_21320,N_21305);
nor U21587 (N_21587,N_21245,N_21364);
nor U21588 (N_21588,N_21322,N_21219);
nand U21589 (N_21589,N_21286,N_21296);
nor U21590 (N_21590,N_21251,N_21273);
or U21591 (N_21591,N_21281,N_21335);
nand U21592 (N_21592,N_21346,N_21242);
xor U21593 (N_21593,N_21342,N_21380);
and U21594 (N_21594,N_21373,N_21292);
nand U21595 (N_21595,N_21329,N_21321);
nor U21596 (N_21596,N_21343,N_21262);
nand U21597 (N_21597,N_21335,N_21294);
or U21598 (N_21598,N_21368,N_21207);
nor U21599 (N_21599,N_21398,N_21220);
nor U21600 (N_21600,N_21583,N_21523);
and U21601 (N_21601,N_21411,N_21501);
nor U21602 (N_21602,N_21592,N_21581);
or U21603 (N_21603,N_21496,N_21585);
and U21604 (N_21604,N_21446,N_21573);
xor U21605 (N_21605,N_21564,N_21415);
and U21606 (N_21606,N_21517,N_21545);
or U21607 (N_21607,N_21525,N_21463);
nor U21608 (N_21608,N_21559,N_21509);
and U21609 (N_21609,N_21563,N_21542);
xor U21610 (N_21610,N_21577,N_21457);
xor U21611 (N_21611,N_21543,N_21521);
nand U21612 (N_21612,N_21473,N_21534);
nor U21613 (N_21613,N_21492,N_21428);
and U21614 (N_21614,N_21491,N_21561);
and U21615 (N_21615,N_21567,N_21413);
nand U21616 (N_21616,N_21424,N_21423);
nand U21617 (N_21617,N_21589,N_21470);
nand U21618 (N_21618,N_21571,N_21579);
or U21619 (N_21619,N_21440,N_21429);
and U21620 (N_21620,N_21539,N_21497);
and U21621 (N_21621,N_21593,N_21481);
nor U21622 (N_21622,N_21519,N_21512);
xnor U21623 (N_21623,N_21547,N_21518);
nor U21624 (N_21624,N_21554,N_21529);
nor U21625 (N_21625,N_21430,N_21570);
xor U21626 (N_21626,N_21464,N_21505);
or U21627 (N_21627,N_21416,N_21449);
xor U21628 (N_21628,N_21439,N_21537);
xnor U21629 (N_21629,N_21520,N_21450);
or U21630 (N_21630,N_21405,N_21471);
nor U21631 (N_21631,N_21508,N_21466);
or U21632 (N_21632,N_21432,N_21469);
and U21633 (N_21633,N_21409,N_21498);
xnor U21634 (N_21634,N_21587,N_21533);
nor U21635 (N_21635,N_21414,N_21565);
nand U21636 (N_21636,N_21444,N_21455);
nor U21637 (N_21637,N_21524,N_21552);
or U21638 (N_21638,N_21553,N_21569);
and U21639 (N_21639,N_21532,N_21426);
nand U21640 (N_21640,N_21582,N_21419);
or U21641 (N_21641,N_21538,N_21541);
nand U21642 (N_21642,N_21502,N_21557);
xnor U21643 (N_21643,N_21477,N_21575);
and U21644 (N_21644,N_21462,N_21562);
or U21645 (N_21645,N_21596,N_21427);
or U21646 (N_21646,N_21443,N_21478);
nand U21647 (N_21647,N_21422,N_21506);
xnor U21648 (N_21648,N_21458,N_21550);
nor U21649 (N_21649,N_21510,N_21456);
or U21650 (N_21650,N_21504,N_21551);
or U21651 (N_21651,N_21438,N_21452);
or U21652 (N_21652,N_21467,N_21522);
and U21653 (N_21653,N_21485,N_21465);
nand U21654 (N_21654,N_21425,N_21560);
xnor U21655 (N_21655,N_21490,N_21487);
and U21656 (N_21656,N_21566,N_21459);
or U21657 (N_21657,N_21558,N_21453);
xor U21658 (N_21658,N_21420,N_21486);
nor U21659 (N_21659,N_21513,N_21507);
nor U21660 (N_21660,N_21590,N_21503);
nand U21661 (N_21661,N_21475,N_21500);
and U21662 (N_21662,N_21474,N_21499);
or U21663 (N_21663,N_21578,N_21454);
and U21664 (N_21664,N_21417,N_21514);
and U21665 (N_21665,N_21442,N_21536);
nor U21666 (N_21666,N_21403,N_21516);
xor U21667 (N_21667,N_21433,N_21540);
and U21668 (N_21668,N_21418,N_21594);
and U21669 (N_21669,N_21484,N_21435);
and U21670 (N_21670,N_21436,N_21407);
nand U21671 (N_21671,N_21580,N_21404);
and U21672 (N_21672,N_21568,N_21461);
nand U21673 (N_21673,N_21400,N_21599);
xnor U21674 (N_21674,N_21460,N_21493);
xor U21675 (N_21675,N_21526,N_21476);
nand U21676 (N_21676,N_21555,N_21406);
nor U21677 (N_21677,N_21494,N_21548);
nand U21678 (N_21678,N_21515,N_21483);
or U21679 (N_21679,N_21595,N_21488);
and U21680 (N_21680,N_21412,N_21401);
xnor U21681 (N_21681,N_21584,N_21597);
nand U21682 (N_21682,N_21586,N_21535);
xnor U21683 (N_21683,N_21511,N_21468);
nor U21684 (N_21684,N_21527,N_21588);
and U21685 (N_21685,N_21479,N_21556);
xnor U21686 (N_21686,N_21445,N_21528);
nor U21687 (N_21687,N_21408,N_21482);
and U21688 (N_21688,N_21437,N_21574);
nand U21689 (N_21689,N_21546,N_21431);
nor U21690 (N_21690,N_21576,N_21591);
nand U21691 (N_21691,N_21531,N_21448);
and U21692 (N_21692,N_21489,N_21549);
and U21693 (N_21693,N_21447,N_21451);
nand U21694 (N_21694,N_21421,N_21495);
or U21695 (N_21695,N_21480,N_21402);
and U21696 (N_21696,N_21434,N_21572);
or U21697 (N_21697,N_21472,N_21544);
xor U21698 (N_21698,N_21530,N_21441);
xor U21699 (N_21699,N_21598,N_21410);
nand U21700 (N_21700,N_21526,N_21458);
and U21701 (N_21701,N_21487,N_21515);
xor U21702 (N_21702,N_21407,N_21435);
or U21703 (N_21703,N_21442,N_21524);
or U21704 (N_21704,N_21584,N_21471);
xor U21705 (N_21705,N_21418,N_21593);
nand U21706 (N_21706,N_21581,N_21432);
xor U21707 (N_21707,N_21442,N_21552);
and U21708 (N_21708,N_21509,N_21535);
and U21709 (N_21709,N_21460,N_21495);
nor U21710 (N_21710,N_21533,N_21556);
xnor U21711 (N_21711,N_21576,N_21488);
xor U21712 (N_21712,N_21516,N_21541);
or U21713 (N_21713,N_21548,N_21482);
nor U21714 (N_21714,N_21455,N_21475);
and U21715 (N_21715,N_21532,N_21569);
xor U21716 (N_21716,N_21565,N_21541);
and U21717 (N_21717,N_21415,N_21529);
or U21718 (N_21718,N_21431,N_21539);
and U21719 (N_21719,N_21440,N_21583);
and U21720 (N_21720,N_21530,N_21474);
nand U21721 (N_21721,N_21440,N_21417);
and U21722 (N_21722,N_21411,N_21467);
xnor U21723 (N_21723,N_21554,N_21454);
and U21724 (N_21724,N_21407,N_21538);
or U21725 (N_21725,N_21540,N_21451);
xor U21726 (N_21726,N_21422,N_21477);
or U21727 (N_21727,N_21506,N_21589);
or U21728 (N_21728,N_21476,N_21449);
xnor U21729 (N_21729,N_21447,N_21575);
xnor U21730 (N_21730,N_21421,N_21441);
or U21731 (N_21731,N_21497,N_21544);
and U21732 (N_21732,N_21461,N_21548);
xor U21733 (N_21733,N_21428,N_21502);
nor U21734 (N_21734,N_21426,N_21544);
nor U21735 (N_21735,N_21439,N_21431);
or U21736 (N_21736,N_21478,N_21441);
xnor U21737 (N_21737,N_21524,N_21532);
nor U21738 (N_21738,N_21496,N_21499);
or U21739 (N_21739,N_21585,N_21469);
nand U21740 (N_21740,N_21472,N_21486);
and U21741 (N_21741,N_21435,N_21571);
or U21742 (N_21742,N_21570,N_21509);
nand U21743 (N_21743,N_21524,N_21582);
nor U21744 (N_21744,N_21410,N_21525);
nor U21745 (N_21745,N_21599,N_21438);
nand U21746 (N_21746,N_21521,N_21420);
xnor U21747 (N_21747,N_21403,N_21553);
xnor U21748 (N_21748,N_21473,N_21545);
nand U21749 (N_21749,N_21516,N_21450);
and U21750 (N_21750,N_21475,N_21488);
or U21751 (N_21751,N_21515,N_21431);
nor U21752 (N_21752,N_21400,N_21496);
or U21753 (N_21753,N_21516,N_21436);
xnor U21754 (N_21754,N_21580,N_21503);
xor U21755 (N_21755,N_21593,N_21419);
or U21756 (N_21756,N_21434,N_21480);
and U21757 (N_21757,N_21486,N_21454);
nor U21758 (N_21758,N_21552,N_21400);
and U21759 (N_21759,N_21424,N_21454);
and U21760 (N_21760,N_21454,N_21546);
xor U21761 (N_21761,N_21481,N_21495);
or U21762 (N_21762,N_21537,N_21585);
and U21763 (N_21763,N_21595,N_21591);
nand U21764 (N_21764,N_21539,N_21519);
and U21765 (N_21765,N_21409,N_21573);
or U21766 (N_21766,N_21563,N_21494);
nor U21767 (N_21767,N_21489,N_21566);
and U21768 (N_21768,N_21462,N_21597);
and U21769 (N_21769,N_21552,N_21419);
and U21770 (N_21770,N_21409,N_21407);
and U21771 (N_21771,N_21446,N_21531);
xnor U21772 (N_21772,N_21510,N_21462);
nor U21773 (N_21773,N_21414,N_21478);
nor U21774 (N_21774,N_21442,N_21561);
and U21775 (N_21775,N_21597,N_21567);
xnor U21776 (N_21776,N_21466,N_21563);
or U21777 (N_21777,N_21521,N_21578);
nor U21778 (N_21778,N_21502,N_21449);
nor U21779 (N_21779,N_21561,N_21477);
and U21780 (N_21780,N_21534,N_21486);
nand U21781 (N_21781,N_21563,N_21462);
or U21782 (N_21782,N_21402,N_21557);
nor U21783 (N_21783,N_21417,N_21510);
or U21784 (N_21784,N_21408,N_21428);
and U21785 (N_21785,N_21441,N_21419);
nor U21786 (N_21786,N_21591,N_21597);
nand U21787 (N_21787,N_21501,N_21589);
and U21788 (N_21788,N_21500,N_21410);
or U21789 (N_21789,N_21482,N_21544);
nor U21790 (N_21790,N_21406,N_21435);
and U21791 (N_21791,N_21449,N_21570);
or U21792 (N_21792,N_21418,N_21513);
or U21793 (N_21793,N_21591,N_21422);
xnor U21794 (N_21794,N_21417,N_21475);
nand U21795 (N_21795,N_21566,N_21462);
nor U21796 (N_21796,N_21596,N_21465);
and U21797 (N_21797,N_21528,N_21596);
nor U21798 (N_21798,N_21524,N_21429);
nor U21799 (N_21799,N_21406,N_21546);
nor U21800 (N_21800,N_21740,N_21755);
nand U21801 (N_21801,N_21639,N_21715);
nor U21802 (N_21802,N_21615,N_21719);
and U21803 (N_21803,N_21668,N_21735);
xor U21804 (N_21804,N_21741,N_21727);
nor U21805 (N_21805,N_21701,N_21638);
or U21806 (N_21806,N_21629,N_21779);
nor U21807 (N_21807,N_21770,N_21612);
or U21808 (N_21808,N_21603,N_21788);
xor U21809 (N_21809,N_21601,N_21757);
and U21810 (N_21810,N_21607,N_21653);
or U21811 (N_21811,N_21789,N_21768);
or U21812 (N_21812,N_21765,N_21797);
xnor U21813 (N_21813,N_21633,N_21763);
or U21814 (N_21814,N_21610,N_21764);
xor U21815 (N_21815,N_21739,N_21749);
or U21816 (N_21816,N_21743,N_21748);
or U21817 (N_21817,N_21664,N_21625);
nor U21818 (N_21818,N_21604,N_21717);
or U21819 (N_21819,N_21784,N_21661);
nor U21820 (N_21820,N_21760,N_21662);
nand U21821 (N_21821,N_21628,N_21677);
xnor U21822 (N_21822,N_21766,N_21796);
nand U21823 (N_21823,N_21746,N_21622);
or U21824 (N_21824,N_21754,N_21724);
nand U21825 (N_21825,N_21663,N_21713);
or U21826 (N_21826,N_21644,N_21613);
xor U21827 (N_21827,N_21708,N_21747);
nand U21828 (N_21828,N_21787,N_21620);
or U21829 (N_21829,N_21689,N_21790);
nand U21830 (N_21830,N_21720,N_21647);
xor U21831 (N_21831,N_21619,N_21753);
xor U21832 (N_21832,N_21710,N_21792);
xnor U21833 (N_21833,N_21736,N_21752);
nor U21834 (N_21834,N_21674,N_21687);
xnor U21835 (N_21835,N_21649,N_21667);
and U21836 (N_21836,N_21632,N_21617);
nand U21837 (N_21837,N_21775,N_21718);
or U21838 (N_21838,N_21680,N_21772);
nor U21839 (N_21839,N_21721,N_21682);
nand U21840 (N_21840,N_21780,N_21697);
or U21841 (N_21841,N_21616,N_21611);
and U21842 (N_21842,N_21636,N_21606);
and U21843 (N_21843,N_21703,N_21706);
or U21844 (N_21844,N_21675,N_21652);
nor U21845 (N_21845,N_21605,N_21669);
and U21846 (N_21846,N_21624,N_21737);
or U21847 (N_21847,N_21712,N_21695);
xor U21848 (N_21848,N_21691,N_21671);
or U21849 (N_21849,N_21781,N_21704);
xnor U21850 (N_21850,N_21783,N_21722);
xnor U21851 (N_21851,N_21778,N_21774);
and U21852 (N_21852,N_21609,N_21759);
or U21853 (N_21853,N_21693,N_21683);
and U21854 (N_21854,N_21696,N_21731);
or U21855 (N_21855,N_21690,N_21725);
and U21856 (N_21856,N_21685,N_21795);
or U21857 (N_21857,N_21621,N_21637);
and U21858 (N_21858,N_21631,N_21626);
nor U21859 (N_21859,N_21794,N_21635);
and U21860 (N_21860,N_21627,N_21751);
xor U21861 (N_21861,N_21769,N_21659);
nor U21862 (N_21862,N_21771,N_21634);
xor U21863 (N_21863,N_21732,N_21681);
nand U21864 (N_21864,N_21679,N_21726);
nand U21865 (N_21865,N_21694,N_21700);
xor U21866 (N_21866,N_21658,N_21729);
nor U21867 (N_21867,N_21767,N_21686);
nor U21868 (N_21868,N_21614,N_21643);
nor U21869 (N_21869,N_21738,N_21678);
nand U21870 (N_21870,N_21608,N_21782);
nand U21871 (N_21871,N_21761,N_21630);
nor U21872 (N_21872,N_21688,N_21707);
nor U21873 (N_21873,N_21657,N_21651);
or U21874 (N_21874,N_21734,N_21745);
nand U21875 (N_21875,N_21618,N_21776);
nor U21876 (N_21876,N_21750,N_21723);
or U21877 (N_21877,N_21709,N_21698);
and U21878 (N_21878,N_21762,N_21702);
xnor U21879 (N_21879,N_21623,N_21756);
xnor U21880 (N_21880,N_21600,N_21786);
and U21881 (N_21881,N_21670,N_21646);
or U21882 (N_21882,N_21730,N_21660);
or U21883 (N_21883,N_21673,N_21676);
or U21884 (N_21884,N_21602,N_21711);
nor U21885 (N_21885,N_21714,N_21650);
nand U21886 (N_21886,N_21793,N_21654);
xnor U21887 (N_21887,N_21641,N_21648);
and U21888 (N_21888,N_21655,N_21785);
and U21889 (N_21889,N_21798,N_21699);
nand U21890 (N_21890,N_21692,N_21656);
nor U21891 (N_21891,N_21716,N_21705);
xor U21892 (N_21892,N_21742,N_21645);
nand U21893 (N_21893,N_21666,N_21642);
and U21894 (N_21894,N_21777,N_21640);
xnor U21895 (N_21895,N_21791,N_21758);
nor U21896 (N_21896,N_21672,N_21684);
xor U21897 (N_21897,N_21773,N_21728);
and U21898 (N_21898,N_21744,N_21799);
nor U21899 (N_21899,N_21665,N_21733);
and U21900 (N_21900,N_21752,N_21627);
and U21901 (N_21901,N_21641,N_21681);
nand U21902 (N_21902,N_21763,N_21774);
and U21903 (N_21903,N_21654,N_21614);
or U21904 (N_21904,N_21727,N_21747);
and U21905 (N_21905,N_21604,N_21602);
and U21906 (N_21906,N_21756,N_21639);
nand U21907 (N_21907,N_21795,N_21600);
or U21908 (N_21908,N_21798,N_21759);
and U21909 (N_21909,N_21753,N_21670);
nand U21910 (N_21910,N_21611,N_21703);
or U21911 (N_21911,N_21771,N_21747);
nor U21912 (N_21912,N_21717,N_21749);
xor U21913 (N_21913,N_21694,N_21683);
or U21914 (N_21914,N_21745,N_21775);
or U21915 (N_21915,N_21761,N_21644);
xnor U21916 (N_21916,N_21639,N_21762);
nor U21917 (N_21917,N_21677,N_21648);
nor U21918 (N_21918,N_21629,N_21624);
and U21919 (N_21919,N_21615,N_21722);
and U21920 (N_21920,N_21632,N_21750);
nor U21921 (N_21921,N_21604,N_21780);
nor U21922 (N_21922,N_21602,N_21652);
xnor U21923 (N_21923,N_21683,N_21771);
and U21924 (N_21924,N_21771,N_21666);
nor U21925 (N_21925,N_21671,N_21641);
nor U21926 (N_21926,N_21612,N_21638);
and U21927 (N_21927,N_21643,N_21679);
nor U21928 (N_21928,N_21621,N_21702);
and U21929 (N_21929,N_21601,N_21772);
and U21930 (N_21930,N_21753,N_21761);
and U21931 (N_21931,N_21620,N_21606);
or U21932 (N_21932,N_21646,N_21716);
and U21933 (N_21933,N_21780,N_21644);
nand U21934 (N_21934,N_21612,N_21623);
nor U21935 (N_21935,N_21667,N_21797);
xor U21936 (N_21936,N_21755,N_21769);
and U21937 (N_21937,N_21740,N_21635);
nand U21938 (N_21938,N_21687,N_21701);
nor U21939 (N_21939,N_21706,N_21664);
xnor U21940 (N_21940,N_21784,N_21633);
nor U21941 (N_21941,N_21623,N_21795);
or U21942 (N_21942,N_21708,N_21777);
xor U21943 (N_21943,N_21715,N_21701);
xor U21944 (N_21944,N_21686,N_21637);
nor U21945 (N_21945,N_21646,N_21656);
and U21946 (N_21946,N_21715,N_21768);
nand U21947 (N_21947,N_21603,N_21664);
nand U21948 (N_21948,N_21763,N_21631);
nand U21949 (N_21949,N_21666,N_21784);
nand U21950 (N_21950,N_21722,N_21632);
or U21951 (N_21951,N_21772,N_21746);
xnor U21952 (N_21952,N_21686,N_21606);
or U21953 (N_21953,N_21676,N_21768);
nand U21954 (N_21954,N_21724,N_21675);
xor U21955 (N_21955,N_21637,N_21778);
xnor U21956 (N_21956,N_21653,N_21781);
or U21957 (N_21957,N_21758,N_21721);
or U21958 (N_21958,N_21769,N_21772);
nand U21959 (N_21959,N_21774,N_21730);
and U21960 (N_21960,N_21762,N_21697);
and U21961 (N_21961,N_21652,N_21727);
nand U21962 (N_21962,N_21608,N_21612);
and U21963 (N_21963,N_21724,N_21752);
nor U21964 (N_21964,N_21681,N_21728);
and U21965 (N_21965,N_21694,N_21715);
nand U21966 (N_21966,N_21697,N_21774);
nand U21967 (N_21967,N_21670,N_21767);
nand U21968 (N_21968,N_21782,N_21759);
or U21969 (N_21969,N_21694,N_21642);
xor U21970 (N_21970,N_21613,N_21719);
nor U21971 (N_21971,N_21701,N_21714);
and U21972 (N_21972,N_21728,N_21679);
or U21973 (N_21973,N_21734,N_21717);
nor U21974 (N_21974,N_21766,N_21680);
or U21975 (N_21975,N_21605,N_21698);
nand U21976 (N_21976,N_21765,N_21603);
xnor U21977 (N_21977,N_21684,N_21771);
or U21978 (N_21978,N_21630,N_21772);
or U21979 (N_21979,N_21761,N_21726);
xnor U21980 (N_21980,N_21684,N_21722);
or U21981 (N_21981,N_21632,N_21691);
xor U21982 (N_21982,N_21615,N_21752);
nor U21983 (N_21983,N_21627,N_21602);
or U21984 (N_21984,N_21705,N_21635);
nor U21985 (N_21985,N_21696,N_21776);
or U21986 (N_21986,N_21722,N_21777);
nand U21987 (N_21987,N_21753,N_21678);
and U21988 (N_21988,N_21780,N_21601);
and U21989 (N_21989,N_21619,N_21768);
or U21990 (N_21990,N_21696,N_21735);
nor U21991 (N_21991,N_21703,N_21601);
or U21992 (N_21992,N_21672,N_21630);
and U21993 (N_21993,N_21651,N_21640);
nand U21994 (N_21994,N_21714,N_21671);
or U21995 (N_21995,N_21789,N_21644);
or U21996 (N_21996,N_21784,N_21684);
xnor U21997 (N_21997,N_21613,N_21634);
nand U21998 (N_21998,N_21743,N_21655);
and U21999 (N_21999,N_21674,N_21769);
xor U22000 (N_22000,N_21878,N_21891);
or U22001 (N_22001,N_21928,N_21807);
and U22002 (N_22002,N_21905,N_21853);
xor U22003 (N_22003,N_21961,N_21808);
xor U22004 (N_22004,N_21993,N_21898);
and U22005 (N_22005,N_21942,N_21848);
or U22006 (N_22006,N_21900,N_21831);
xor U22007 (N_22007,N_21849,N_21906);
or U22008 (N_22008,N_21820,N_21802);
nor U22009 (N_22009,N_21913,N_21922);
and U22010 (N_22010,N_21924,N_21969);
xnor U22011 (N_22011,N_21865,N_21943);
nand U22012 (N_22012,N_21827,N_21862);
xor U22013 (N_22013,N_21896,N_21945);
xnor U22014 (N_22014,N_21954,N_21893);
nand U22015 (N_22015,N_21823,N_21971);
or U22016 (N_22016,N_21915,N_21956);
xnor U22017 (N_22017,N_21921,N_21814);
xnor U22018 (N_22018,N_21883,N_21816);
and U22019 (N_22019,N_21884,N_21938);
and U22020 (N_22020,N_21836,N_21851);
nand U22021 (N_22021,N_21977,N_21854);
nand U22022 (N_22022,N_21850,N_21813);
xnor U22023 (N_22023,N_21959,N_21970);
or U22024 (N_22024,N_21975,N_21890);
and U22025 (N_22025,N_21935,N_21840);
nor U22026 (N_22026,N_21958,N_21923);
nor U22027 (N_22027,N_21882,N_21837);
or U22028 (N_22028,N_21829,N_21978);
nor U22029 (N_22029,N_21887,N_21815);
and U22030 (N_22030,N_21952,N_21870);
nand U22031 (N_22031,N_21822,N_21819);
or U22032 (N_22032,N_21955,N_21858);
nand U22033 (N_22033,N_21903,N_21818);
nor U22034 (N_22034,N_21995,N_21902);
or U22035 (N_22035,N_21886,N_21981);
or U22036 (N_22036,N_21927,N_21801);
or U22037 (N_22037,N_21817,N_21987);
and U22038 (N_22038,N_21855,N_21907);
nand U22039 (N_22039,N_21830,N_21811);
xnor U22040 (N_22040,N_21868,N_21910);
nand U22041 (N_22041,N_21917,N_21992);
or U22042 (N_22042,N_21986,N_21843);
and U22043 (N_22043,N_21879,N_21991);
nand U22044 (N_22044,N_21967,N_21914);
nor U22045 (N_22045,N_21812,N_21965);
xor U22046 (N_22046,N_21957,N_21863);
and U22047 (N_22047,N_21940,N_21926);
and U22048 (N_22048,N_21835,N_21974);
nand U22049 (N_22049,N_21804,N_21916);
xnor U22050 (N_22050,N_21839,N_21859);
nor U22051 (N_22051,N_21976,N_21806);
nand U22052 (N_22052,N_21998,N_21983);
nand U22053 (N_22053,N_21885,N_21833);
nand U22054 (N_22054,N_21980,N_21908);
nand U22055 (N_22055,N_21845,N_21936);
nand U22056 (N_22056,N_21876,N_21857);
nor U22057 (N_22057,N_21824,N_21877);
and U22058 (N_22058,N_21918,N_21941);
nand U22059 (N_22059,N_21932,N_21925);
or U22060 (N_22060,N_21920,N_21989);
and U22061 (N_22061,N_21864,N_21964);
nor U22062 (N_22062,N_21994,N_21968);
nand U22063 (N_22063,N_21937,N_21825);
or U22064 (N_22064,N_21846,N_21985);
xnor U22065 (N_22065,N_21939,N_21996);
nand U22066 (N_22066,N_21904,N_21946);
xnor U22067 (N_22067,N_21805,N_21899);
and U22068 (N_22068,N_21966,N_21867);
or U22069 (N_22069,N_21872,N_21934);
nor U22070 (N_22070,N_21901,N_21875);
or U22071 (N_22071,N_21828,N_21892);
and U22072 (N_22072,N_21911,N_21947);
nor U22073 (N_22073,N_21832,N_21929);
and U22074 (N_22074,N_21953,N_21881);
nor U22075 (N_22075,N_21889,N_21931);
nand U22076 (N_22076,N_21861,N_21990);
nor U22077 (N_22077,N_21866,N_21897);
nand U22078 (N_22078,N_21856,N_21895);
xor U22079 (N_22079,N_21810,N_21852);
nor U22080 (N_22080,N_21860,N_21803);
xor U22081 (N_22081,N_21800,N_21841);
nor U22082 (N_22082,N_21909,N_21949);
or U22083 (N_22083,N_21979,N_21951);
or U22084 (N_22084,N_21888,N_21962);
nand U22085 (N_22085,N_21948,N_21944);
or U22086 (N_22086,N_21972,N_21873);
or U22087 (N_22087,N_21997,N_21930);
nand U22088 (N_22088,N_21821,N_21847);
or U22089 (N_22089,N_21988,N_21826);
and U22090 (N_22090,N_21933,N_21960);
nand U22091 (N_22091,N_21809,N_21982);
nand U22092 (N_22092,N_21874,N_21963);
or U22093 (N_22093,N_21894,N_21871);
nor U22094 (N_22094,N_21919,N_21912);
nor U22095 (N_22095,N_21984,N_21950);
nand U22096 (N_22096,N_21844,N_21869);
and U22097 (N_22097,N_21880,N_21838);
or U22098 (N_22098,N_21999,N_21834);
nand U22099 (N_22099,N_21973,N_21842);
and U22100 (N_22100,N_21886,N_21960);
nor U22101 (N_22101,N_21940,N_21977);
or U22102 (N_22102,N_21849,N_21870);
or U22103 (N_22103,N_21855,N_21974);
or U22104 (N_22104,N_21952,N_21815);
or U22105 (N_22105,N_21921,N_21948);
xnor U22106 (N_22106,N_21939,N_21956);
nand U22107 (N_22107,N_21850,N_21958);
or U22108 (N_22108,N_21911,N_21983);
nor U22109 (N_22109,N_21900,N_21905);
and U22110 (N_22110,N_21823,N_21861);
nor U22111 (N_22111,N_21933,N_21802);
or U22112 (N_22112,N_21808,N_21838);
nand U22113 (N_22113,N_21872,N_21958);
and U22114 (N_22114,N_21840,N_21868);
or U22115 (N_22115,N_21985,N_21834);
xor U22116 (N_22116,N_21867,N_21828);
nor U22117 (N_22117,N_21983,N_21846);
nand U22118 (N_22118,N_21924,N_21808);
xor U22119 (N_22119,N_21820,N_21859);
nor U22120 (N_22120,N_21844,N_21880);
nor U22121 (N_22121,N_21869,N_21905);
nand U22122 (N_22122,N_21919,N_21836);
or U22123 (N_22123,N_21987,N_21918);
nor U22124 (N_22124,N_21875,N_21816);
nor U22125 (N_22125,N_21932,N_21834);
and U22126 (N_22126,N_21807,N_21840);
nor U22127 (N_22127,N_21912,N_21967);
and U22128 (N_22128,N_21929,N_21802);
and U22129 (N_22129,N_21955,N_21802);
nand U22130 (N_22130,N_21829,N_21939);
nor U22131 (N_22131,N_21835,N_21814);
and U22132 (N_22132,N_21828,N_21804);
nand U22133 (N_22133,N_21974,N_21933);
or U22134 (N_22134,N_21992,N_21986);
nor U22135 (N_22135,N_21888,N_21926);
or U22136 (N_22136,N_21961,N_21921);
xnor U22137 (N_22137,N_21931,N_21907);
or U22138 (N_22138,N_21968,N_21854);
xor U22139 (N_22139,N_21972,N_21860);
xnor U22140 (N_22140,N_21830,N_21806);
nor U22141 (N_22141,N_21935,N_21835);
nor U22142 (N_22142,N_21831,N_21975);
nor U22143 (N_22143,N_21845,N_21956);
nand U22144 (N_22144,N_21848,N_21886);
nor U22145 (N_22145,N_21934,N_21865);
xor U22146 (N_22146,N_21896,N_21961);
nor U22147 (N_22147,N_21893,N_21957);
xor U22148 (N_22148,N_21896,N_21957);
nand U22149 (N_22149,N_21889,N_21853);
nor U22150 (N_22150,N_21862,N_21801);
or U22151 (N_22151,N_21902,N_21895);
or U22152 (N_22152,N_21850,N_21871);
and U22153 (N_22153,N_21978,N_21917);
xnor U22154 (N_22154,N_21802,N_21851);
and U22155 (N_22155,N_21872,N_21820);
nand U22156 (N_22156,N_21855,N_21808);
nand U22157 (N_22157,N_21942,N_21946);
nor U22158 (N_22158,N_21864,N_21841);
nand U22159 (N_22159,N_21988,N_21974);
nand U22160 (N_22160,N_21802,N_21937);
nor U22161 (N_22161,N_21923,N_21992);
or U22162 (N_22162,N_21805,N_21927);
or U22163 (N_22163,N_21841,N_21885);
nand U22164 (N_22164,N_21891,N_21966);
nor U22165 (N_22165,N_21871,N_21951);
or U22166 (N_22166,N_21980,N_21979);
nand U22167 (N_22167,N_21824,N_21999);
nor U22168 (N_22168,N_21982,N_21864);
nor U22169 (N_22169,N_21813,N_21964);
nor U22170 (N_22170,N_21900,N_21922);
nor U22171 (N_22171,N_21969,N_21908);
xnor U22172 (N_22172,N_21973,N_21832);
and U22173 (N_22173,N_21994,N_21846);
nand U22174 (N_22174,N_21960,N_21974);
xor U22175 (N_22175,N_21907,N_21820);
nand U22176 (N_22176,N_21817,N_21971);
and U22177 (N_22177,N_21827,N_21956);
and U22178 (N_22178,N_21886,N_21945);
or U22179 (N_22179,N_21807,N_21915);
and U22180 (N_22180,N_21914,N_21895);
and U22181 (N_22181,N_21903,N_21947);
or U22182 (N_22182,N_21994,N_21837);
or U22183 (N_22183,N_21904,N_21839);
or U22184 (N_22184,N_21963,N_21812);
or U22185 (N_22185,N_21907,N_21909);
and U22186 (N_22186,N_21848,N_21921);
xor U22187 (N_22187,N_21850,N_21866);
nor U22188 (N_22188,N_21951,N_21930);
nand U22189 (N_22189,N_21836,N_21806);
and U22190 (N_22190,N_21878,N_21873);
nand U22191 (N_22191,N_21825,N_21939);
or U22192 (N_22192,N_21948,N_21906);
nor U22193 (N_22193,N_21884,N_21882);
nand U22194 (N_22194,N_21826,N_21995);
and U22195 (N_22195,N_21897,N_21886);
and U22196 (N_22196,N_21821,N_21878);
nand U22197 (N_22197,N_21955,N_21974);
nand U22198 (N_22198,N_21924,N_21970);
xnor U22199 (N_22199,N_21854,N_21881);
nor U22200 (N_22200,N_22084,N_22152);
nor U22201 (N_22201,N_22009,N_22011);
and U22202 (N_22202,N_22001,N_22082);
nor U22203 (N_22203,N_22028,N_22147);
xor U22204 (N_22204,N_22135,N_22124);
nand U22205 (N_22205,N_22081,N_22062);
nor U22206 (N_22206,N_22179,N_22054);
nor U22207 (N_22207,N_22025,N_22101);
nor U22208 (N_22208,N_22137,N_22143);
nor U22209 (N_22209,N_22175,N_22131);
nand U22210 (N_22210,N_22037,N_22183);
nor U22211 (N_22211,N_22016,N_22058);
or U22212 (N_22212,N_22108,N_22076);
nor U22213 (N_22213,N_22048,N_22088);
and U22214 (N_22214,N_22004,N_22194);
nor U22215 (N_22215,N_22000,N_22046);
nand U22216 (N_22216,N_22130,N_22056);
xnor U22217 (N_22217,N_22049,N_22068);
nand U22218 (N_22218,N_22007,N_22167);
nor U22219 (N_22219,N_22010,N_22132);
nand U22220 (N_22220,N_22180,N_22107);
nand U22221 (N_22221,N_22191,N_22075);
nor U22222 (N_22222,N_22040,N_22050);
and U22223 (N_22223,N_22165,N_22109);
and U22224 (N_22224,N_22057,N_22142);
and U22225 (N_22225,N_22115,N_22185);
nor U22226 (N_22226,N_22012,N_22030);
and U22227 (N_22227,N_22117,N_22042);
xor U22228 (N_22228,N_22116,N_22177);
xor U22229 (N_22229,N_22083,N_22095);
xor U22230 (N_22230,N_22052,N_22174);
nor U22231 (N_22231,N_22077,N_22169);
nand U22232 (N_22232,N_22150,N_22158);
and U22233 (N_22233,N_22039,N_22035);
or U22234 (N_22234,N_22154,N_22188);
or U22235 (N_22235,N_22029,N_22125);
or U22236 (N_22236,N_22014,N_22178);
and U22237 (N_22237,N_22129,N_22079);
xnor U22238 (N_22238,N_22162,N_22120);
or U22239 (N_22239,N_22171,N_22078);
nand U22240 (N_22240,N_22148,N_22080);
xnor U22241 (N_22241,N_22060,N_22008);
nand U22242 (N_22242,N_22067,N_22114);
nand U22243 (N_22243,N_22098,N_22128);
or U22244 (N_22244,N_22156,N_22002);
nor U22245 (N_22245,N_22181,N_22161);
nor U22246 (N_22246,N_22089,N_22053);
nor U22247 (N_22247,N_22086,N_22036);
nand U22248 (N_22248,N_22100,N_22055);
or U22249 (N_22249,N_22112,N_22103);
nor U22250 (N_22250,N_22066,N_22034);
and U22251 (N_22251,N_22102,N_22106);
xor U22252 (N_22252,N_22122,N_22182);
nand U22253 (N_22253,N_22043,N_22155);
xor U22254 (N_22254,N_22099,N_22110);
xor U22255 (N_22255,N_22093,N_22087);
and U22256 (N_22256,N_22031,N_22196);
and U22257 (N_22257,N_22160,N_22006);
xnor U22258 (N_22258,N_22044,N_22134);
or U22259 (N_22259,N_22193,N_22097);
nor U22260 (N_22260,N_22070,N_22064);
nand U22261 (N_22261,N_22184,N_22092);
or U22262 (N_22262,N_22126,N_22198);
and U22263 (N_22263,N_22113,N_22013);
and U22264 (N_22264,N_22063,N_22111);
or U22265 (N_22265,N_22199,N_22020);
xor U22266 (N_22266,N_22003,N_22023);
nor U22267 (N_22267,N_22166,N_22173);
nor U22268 (N_22268,N_22026,N_22138);
xnor U22269 (N_22269,N_22176,N_22047);
nand U22270 (N_22270,N_22139,N_22061);
nor U22271 (N_22271,N_22159,N_22195);
and U22272 (N_22272,N_22065,N_22170);
nand U22273 (N_22273,N_22127,N_22038);
xnor U22274 (N_22274,N_22186,N_22071);
nor U22275 (N_22275,N_22051,N_22140);
nand U22276 (N_22276,N_22133,N_22073);
nand U22277 (N_22277,N_22172,N_22157);
or U22278 (N_22278,N_22024,N_22192);
nand U22279 (N_22279,N_22123,N_22119);
or U22280 (N_22280,N_22021,N_22027);
xnor U22281 (N_22281,N_22149,N_22197);
xnor U22282 (N_22282,N_22005,N_22164);
xor U22283 (N_22283,N_22104,N_22090);
and U22284 (N_22284,N_22105,N_22094);
or U22285 (N_22285,N_22187,N_22085);
nand U22286 (N_22286,N_22059,N_22033);
xnor U22287 (N_22287,N_22189,N_22069);
or U22288 (N_22288,N_22074,N_22144);
or U22289 (N_22289,N_22190,N_22136);
xnor U22290 (N_22290,N_22146,N_22091);
nand U22291 (N_22291,N_22141,N_22019);
nor U22292 (N_22292,N_22151,N_22072);
and U22293 (N_22293,N_22045,N_22153);
nand U22294 (N_22294,N_22015,N_22145);
xnor U22295 (N_22295,N_22041,N_22121);
xnor U22296 (N_22296,N_22017,N_22022);
nand U22297 (N_22297,N_22118,N_22096);
or U22298 (N_22298,N_22163,N_22018);
xor U22299 (N_22299,N_22032,N_22168);
and U22300 (N_22300,N_22108,N_22155);
or U22301 (N_22301,N_22169,N_22069);
nor U22302 (N_22302,N_22117,N_22035);
and U22303 (N_22303,N_22039,N_22196);
xnor U22304 (N_22304,N_22015,N_22068);
or U22305 (N_22305,N_22161,N_22124);
or U22306 (N_22306,N_22125,N_22016);
or U22307 (N_22307,N_22160,N_22090);
or U22308 (N_22308,N_22163,N_22130);
nor U22309 (N_22309,N_22064,N_22104);
xnor U22310 (N_22310,N_22047,N_22074);
nand U22311 (N_22311,N_22041,N_22003);
xor U22312 (N_22312,N_22079,N_22013);
or U22313 (N_22313,N_22194,N_22188);
and U22314 (N_22314,N_22148,N_22073);
xor U22315 (N_22315,N_22147,N_22086);
nand U22316 (N_22316,N_22045,N_22174);
or U22317 (N_22317,N_22069,N_22166);
nor U22318 (N_22318,N_22094,N_22146);
xor U22319 (N_22319,N_22037,N_22156);
nor U22320 (N_22320,N_22158,N_22106);
and U22321 (N_22321,N_22031,N_22074);
xor U22322 (N_22322,N_22195,N_22053);
nand U22323 (N_22323,N_22160,N_22159);
or U22324 (N_22324,N_22050,N_22014);
xnor U22325 (N_22325,N_22103,N_22101);
or U22326 (N_22326,N_22041,N_22036);
and U22327 (N_22327,N_22139,N_22088);
nor U22328 (N_22328,N_22017,N_22023);
and U22329 (N_22329,N_22082,N_22038);
and U22330 (N_22330,N_22183,N_22159);
xnor U22331 (N_22331,N_22029,N_22092);
xor U22332 (N_22332,N_22105,N_22108);
xnor U22333 (N_22333,N_22068,N_22121);
nand U22334 (N_22334,N_22154,N_22022);
xnor U22335 (N_22335,N_22138,N_22047);
or U22336 (N_22336,N_22029,N_22084);
or U22337 (N_22337,N_22031,N_22150);
and U22338 (N_22338,N_22035,N_22106);
and U22339 (N_22339,N_22186,N_22121);
and U22340 (N_22340,N_22056,N_22119);
and U22341 (N_22341,N_22087,N_22098);
nor U22342 (N_22342,N_22052,N_22046);
nor U22343 (N_22343,N_22020,N_22175);
and U22344 (N_22344,N_22105,N_22028);
nand U22345 (N_22345,N_22018,N_22070);
nor U22346 (N_22346,N_22021,N_22052);
xnor U22347 (N_22347,N_22191,N_22087);
or U22348 (N_22348,N_22056,N_22133);
xnor U22349 (N_22349,N_22166,N_22176);
xnor U22350 (N_22350,N_22129,N_22003);
and U22351 (N_22351,N_22058,N_22172);
nor U22352 (N_22352,N_22058,N_22009);
xnor U22353 (N_22353,N_22064,N_22198);
xor U22354 (N_22354,N_22135,N_22137);
nand U22355 (N_22355,N_22148,N_22030);
or U22356 (N_22356,N_22050,N_22098);
and U22357 (N_22357,N_22192,N_22018);
nand U22358 (N_22358,N_22000,N_22074);
and U22359 (N_22359,N_22129,N_22159);
xnor U22360 (N_22360,N_22109,N_22046);
xnor U22361 (N_22361,N_22173,N_22110);
nand U22362 (N_22362,N_22119,N_22138);
nand U22363 (N_22363,N_22076,N_22032);
xnor U22364 (N_22364,N_22147,N_22187);
nor U22365 (N_22365,N_22118,N_22084);
xnor U22366 (N_22366,N_22149,N_22126);
and U22367 (N_22367,N_22100,N_22173);
xor U22368 (N_22368,N_22101,N_22107);
xor U22369 (N_22369,N_22121,N_22008);
or U22370 (N_22370,N_22180,N_22018);
or U22371 (N_22371,N_22095,N_22059);
xnor U22372 (N_22372,N_22077,N_22134);
or U22373 (N_22373,N_22093,N_22003);
xnor U22374 (N_22374,N_22020,N_22030);
and U22375 (N_22375,N_22173,N_22122);
nand U22376 (N_22376,N_22081,N_22142);
nand U22377 (N_22377,N_22136,N_22059);
nand U22378 (N_22378,N_22197,N_22096);
nand U22379 (N_22379,N_22114,N_22123);
and U22380 (N_22380,N_22147,N_22082);
xor U22381 (N_22381,N_22097,N_22102);
or U22382 (N_22382,N_22098,N_22004);
and U22383 (N_22383,N_22005,N_22036);
nand U22384 (N_22384,N_22126,N_22182);
nor U22385 (N_22385,N_22049,N_22053);
nand U22386 (N_22386,N_22024,N_22185);
and U22387 (N_22387,N_22091,N_22193);
or U22388 (N_22388,N_22038,N_22087);
xnor U22389 (N_22389,N_22139,N_22104);
or U22390 (N_22390,N_22106,N_22164);
and U22391 (N_22391,N_22072,N_22021);
and U22392 (N_22392,N_22023,N_22020);
xor U22393 (N_22393,N_22006,N_22056);
nor U22394 (N_22394,N_22076,N_22118);
xor U22395 (N_22395,N_22085,N_22024);
xor U22396 (N_22396,N_22030,N_22061);
and U22397 (N_22397,N_22035,N_22122);
nand U22398 (N_22398,N_22168,N_22014);
nor U22399 (N_22399,N_22129,N_22157);
or U22400 (N_22400,N_22213,N_22363);
nor U22401 (N_22401,N_22340,N_22297);
or U22402 (N_22402,N_22316,N_22333);
and U22403 (N_22403,N_22269,N_22372);
and U22404 (N_22404,N_22380,N_22231);
xnor U22405 (N_22405,N_22391,N_22229);
xnor U22406 (N_22406,N_22225,N_22344);
nor U22407 (N_22407,N_22280,N_22302);
xnor U22408 (N_22408,N_22322,N_22392);
or U22409 (N_22409,N_22334,N_22375);
or U22410 (N_22410,N_22346,N_22202);
and U22411 (N_22411,N_22318,N_22367);
and U22412 (N_22412,N_22287,N_22365);
or U22413 (N_22413,N_22312,N_22289);
or U22414 (N_22414,N_22324,N_22376);
xor U22415 (N_22415,N_22219,N_22249);
nand U22416 (N_22416,N_22321,N_22248);
xnor U22417 (N_22417,N_22212,N_22320);
and U22418 (N_22418,N_22329,N_22224);
nand U22419 (N_22419,N_22327,N_22371);
nor U22420 (N_22420,N_22236,N_22209);
nand U22421 (N_22421,N_22382,N_22298);
or U22422 (N_22422,N_22360,N_22331);
xor U22423 (N_22423,N_22345,N_22221);
nor U22424 (N_22424,N_22305,N_22241);
xnor U22425 (N_22425,N_22238,N_22352);
xor U22426 (N_22426,N_22342,N_22338);
nand U22427 (N_22427,N_22273,N_22210);
or U22428 (N_22428,N_22390,N_22336);
nor U22429 (N_22429,N_22330,N_22315);
and U22430 (N_22430,N_22310,N_22240);
nor U22431 (N_22431,N_22239,N_22245);
nor U22432 (N_22432,N_22286,N_22265);
xnor U22433 (N_22433,N_22208,N_22351);
or U22434 (N_22434,N_22203,N_22296);
nand U22435 (N_22435,N_22207,N_22230);
nand U22436 (N_22436,N_22319,N_22260);
and U22437 (N_22437,N_22341,N_22254);
nor U22438 (N_22438,N_22317,N_22226);
nor U22439 (N_22439,N_22200,N_22282);
xnor U22440 (N_22440,N_22301,N_22303);
xnor U22441 (N_22441,N_22311,N_22350);
xnor U22442 (N_22442,N_22362,N_22252);
xnor U22443 (N_22443,N_22393,N_22357);
and U22444 (N_22444,N_22270,N_22272);
or U22445 (N_22445,N_22274,N_22227);
xor U22446 (N_22446,N_22250,N_22204);
nand U22447 (N_22447,N_22355,N_22228);
nand U22448 (N_22448,N_22397,N_22294);
or U22449 (N_22449,N_22271,N_22242);
nand U22450 (N_22450,N_22379,N_22394);
nor U22451 (N_22451,N_22278,N_22347);
nand U22452 (N_22452,N_22262,N_22358);
and U22453 (N_22453,N_22205,N_22284);
or U22454 (N_22454,N_22281,N_22247);
and U22455 (N_22455,N_22220,N_22313);
and U22456 (N_22456,N_22368,N_22256);
nand U22457 (N_22457,N_22218,N_22261);
nor U22458 (N_22458,N_22323,N_22361);
or U22459 (N_22459,N_22325,N_22383);
nand U22460 (N_22460,N_22388,N_22237);
nand U22461 (N_22461,N_22257,N_22216);
and U22462 (N_22462,N_22214,N_22335);
xor U22463 (N_22463,N_22263,N_22279);
or U22464 (N_22464,N_22277,N_22292);
nor U22465 (N_22465,N_22255,N_22217);
or U22466 (N_22466,N_22285,N_22246);
and U22467 (N_22467,N_22337,N_22253);
nor U22468 (N_22468,N_22307,N_22243);
and U22469 (N_22469,N_22399,N_22251);
nand U22470 (N_22470,N_22332,N_22314);
or U22471 (N_22471,N_22374,N_22306);
xor U22472 (N_22472,N_22309,N_22385);
or U22473 (N_22473,N_22267,N_22395);
xnor U22474 (N_22474,N_22258,N_22364);
and U22475 (N_22475,N_22398,N_22396);
xnor U22476 (N_22476,N_22222,N_22201);
nand U22477 (N_22477,N_22378,N_22328);
or U22478 (N_22478,N_22386,N_22343);
or U22479 (N_22479,N_22232,N_22300);
nor U22480 (N_22480,N_22373,N_22264);
nand U22481 (N_22481,N_22291,N_22366);
nand U22482 (N_22482,N_22370,N_22359);
or U22483 (N_22483,N_22215,N_22211);
nor U22484 (N_22484,N_22295,N_22381);
nor U22485 (N_22485,N_22235,N_22259);
nand U22486 (N_22486,N_22293,N_22244);
and U22487 (N_22487,N_22384,N_22353);
xor U22488 (N_22488,N_22348,N_22304);
nand U22489 (N_22489,N_22288,N_22369);
and U22490 (N_22490,N_22266,N_22349);
or U22491 (N_22491,N_22233,N_22299);
xnor U22492 (N_22492,N_22339,N_22354);
or U22493 (N_22493,N_22223,N_22377);
nand U22494 (N_22494,N_22234,N_22275);
nor U22495 (N_22495,N_22389,N_22268);
xor U22496 (N_22496,N_22276,N_22283);
xor U22497 (N_22497,N_22206,N_22308);
xor U22498 (N_22498,N_22290,N_22326);
and U22499 (N_22499,N_22356,N_22387);
or U22500 (N_22500,N_22205,N_22219);
nand U22501 (N_22501,N_22293,N_22332);
and U22502 (N_22502,N_22351,N_22389);
xor U22503 (N_22503,N_22242,N_22308);
and U22504 (N_22504,N_22228,N_22314);
xnor U22505 (N_22505,N_22314,N_22355);
or U22506 (N_22506,N_22362,N_22275);
nand U22507 (N_22507,N_22247,N_22250);
nor U22508 (N_22508,N_22203,N_22378);
nand U22509 (N_22509,N_22256,N_22278);
nand U22510 (N_22510,N_22222,N_22252);
nor U22511 (N_22511,N_22269,N_22209);
and U22512 (N_22512,N_22278,N_22355);
xor U22513 (N_22513,N_22221,N_22397);
or U22514 (N_22514,N_22215,N_22370);
nor U22515 (N_22515,N_22249,N_22381);
nand U22516 (N_22516,N_22224,N_22332);
nor U22517 (N_22517,N_22393,N_22228);
nor U22518 (N_22518,N_22250,N_22220);
nor U22519 (N_22519,N_22226,N_22243);
nand U22520 (N_22520,N_22391,N_22201);
nor U22521 (N_22521,N_22360,N_22264);
nand U22522 (N_22522,N_22220,N_22273);
or U22523 (N_22523,N_22348,N_22275);
or U22524 (N_22524,N_22212,N_22374);
xor U22525 (N_22525,N_22368,N_22318);
and U22526 (N_22526,N_22241,N_22355);
nand U22527 (N_22527,N_22311,N_22298);
nand U22528 (N_22528,N_22303,N_22270);
xnor U22529 (N_22529,N_22242,N_22309);
nand U22530 (N_22530,N_22206,N_22332);
nand U22531 (N_22531,N_22392,N_22389);
nor U22532 (N_22532,N_22305,N_22281);
nand U22533 (N_22533,N_22263,N_22388);
nand U22534 (N_22534,N_22379,N_22282);
or U22535 (N_22535,N_22386,N_22247);
nor U22536 (N_22536,N_22281,N_22230);
nand U22537 (N_22537,N_22345,N_22249);
or U22538 (N_22538,N_22233,N_22395);
xor U22539 (N_22539,N_22255,N_22207);
nor U22540 (N_22540,N_22363,N_22392);
nand U22541 (N_22541,N_22263,N_22291);
nor U22542 (N_22542,N_22280,N_22206);
and U22543 (N_22543,N_22354,N_22206);
nand U22544 (N_22544,N_22315,N_22284);
or U22545 (N_22545,N_22383,N_22269);
nand U22546 (N_22546,N_22273,N_22256);
xor U22547 (N_22547,N_22347,N_22365);
nand U22548 (N_22548,N_22283,N_22316);
nand U22549 (N_22549,N_22319,N_22399);
or U22550 (N_22550,N_22285,N_22343);
or U22551 (N_22551,N_22218,N_22250);
and U22552 (N_22552,N_22316,N_22263);
nor U22553 (N_22553,N_22382,N_22297);
or U22554 (N_22554,N_22364,N_22319);
and U22555 (N_22555,N_22281,N_22246);
and U22556 (N_22556,N_22241,N_22201);
nand U22557 (N_22557,N_22364,N_22327);
nand U22558 (N_22558,N_22204,N_22303);
and U22559 (N_22559,N_22385,N_22355);
nand U22560 (N_22560,N_22203,N_22316);
nand U22561 (N_22561,N_22347,N_22264);
and U22562 (N_22562,N_22215,N_22295);
and U22563 (N_22563,N_22347,N_22265);
and U22564 (N_22564,N_22342,N_22276);
or U22565 (N_22565,N_22331,N_22329);
xnor U22566 (N_22566,N_22358,N_22384);
xor U22567 (N_22567,N_22223,N_22396);
or U22568 (N_22568,N_22236,N_22344);
nor U22569 (N_22569,N_22392,N_22398);
nor U22570 (N_22570,N_22338,N_22216);
xor U22571 (N_22571,N_22208,N_22337);
xnor U22572 (N_22572,N_22345,N_22394);
or U22573 (N_22573,N_22302,N_22225);
nor U22574 (N_22574,N_22233,N_22223);
nand U22575 (N_22575,N_22245,N_22225);
nand U22576 (N_22576,N_22372,N_22397);
xor U22577 (N_22577,N_22216,N_22387);
nand U22578 (N_22578,N_22328,N_22219);
nor U22579 (N_22579,N_22369,N_22282);
nor U22580 (N_22580,N_22224,N_22278);
nand U22581 (N_22581,N_22376,N_22301);
nor U22582 (N_22582,N_22287,N_22350);
nor U22583 (N_22583,N_22241,N_22393);
nand U22584 (N_22584,N_22333,N_22268);
nand U22585 (N_22585,N_22307,N_22205);
nor U22586 (N_22586,N_22299,N_22262);
or U22587 (N_22587,N_22298,N_22295);
nor U22588 (N_22588,N_22290,N_22330);
and U22589 (N_22589,N_22341,N_22359);
nand U22590 (N_22590,N_22276,N_22310);
xor U22591 (N_22591,N_22226,N_22398);
or U22592 (N_22592,N_22268,N_22213);
nand U22593 (N_22593,N_22359,N_22354);
nand U22594 (N_22594,N_22384,N_22348);
or U22595 (N_22595,N_22323,N_22397);
or U22596 (N_22596,N_22371,N_22339);
nor U22597 (N_22597,N_22393,N_22284);
nor U22598 (N_22598,N_22230,N_22321);
and U22599 (N_22599,N_22354,N_22255);
or U22600 (N_22600,N_22478,N_22403);
nand U22601 (N_22601,N_22518,N_22490);
and U22602 (N_22602,N_22412,N_22417);
nor U22603 (N_22603,N_22553,N_22545);
or U22604 (N_22604,N_22581,N_22585);
nand U22605 (N_22605,N_22400,N_22498);
nor U22606 (N_22606,N_22512,N_22415);
xor U22607 (N_22607,N_22431,N_22413);
nand U22608 (N_22608,N_22586,N_22452);
nand U22609 (N_22609,N_22589,N_22508);
nor U22610 (N_22610,N_22582,N_22594);
nand U22611 (N_22611,N_22410,N_22556);
and U22612 (N_22612,N_22476,N_22570);
and U22613 (N_22613,N_22475,N_22566);
xnor U22614 (N_22614,N_22466,N_22447);
xor U22615 (N_22615,N_22569,N_22554);
nand U22616 (N_22616,N_22536,N_22481);
xor U22617 (N_22617,N_22456,N_22494);
or U22618 (N_22618,N_22437,N_22474);
or U22619 (N_22619,N_22416,N_22561);
nor U22620 (N_22620,N_22493,N_22500);
and U22621 (N_22621,N_22441,N_22537);
nor U22622 (N_22622,N_22522,N_22596);
xnor U22623 (N_22623,N_22408,N_22461);
nand U22624 (N_22624,N_22547,N_22515);
or U22625 (N_22625,N_22434,N_22588);
or U22626 (N_22626,N_22517,N_22409);
nor U22627 (N_22627,N_22531,N_22445);
nand U22628 (N_22628,N_22563,N_22442);
and U22629 (N_22629,N_22446,N_22577);
nand U22630 (N_22630,N_22425,N_22485);
nand U22631 (N_22631,N_22533,N_22489);
xor U22632 (N_22632,N_22497,N_22454);
and U22633 (N_22633,N_22443,N_22573);
nor U22634 (N_22634,N_22579,N_22543);
or U22635 (N_22635,N_22571,N_22469);
or U22636 (N_22636,N_22495,N_22590);
and U22637 (N_22637,N_22513,N_22457);
nand U22638 (N_22638,N_22502,N_22482);
nor U22639 (N_22639,N_22555,N_22486);
xnor U22640 (N_22640,N_22432,N_22421);
xor U22641 (N_22641,N_22453,N_22424);
nand U22642 (N_22642,N_22503,N_22578);
or U22643 (N_22643,N_22575,N_22455);
nor U22644 (N_22644,N_22529,N_22551);
or U22645 (N_22645,N_22567,N_22507);
and U22646 (N_22646,N_22464,N_22414);
xor U22647 (N_22647,N_22562,N_22524);
xnor U22648 (N_22648,N_22587,N_22418);
and U22649 (N_22649,N_22574,N_22560);
nor U22650 (N_22650,N_22439,N_22584);
or U22651 (N_22651,N_22467,N_22460);
nor U22652 (N_22652,N_22451,N_22528);
and U22653 (N_22653,N_22406,N_22458);
or U22654 (N_22654,N_22568,N_22423);
nand U22655 (N_22655,N_22595,N_22462);
xnor U22656 (N_22656,N_22420,N_22565);
and U22657 (N_22657,N_22510,N_22572);
and U22658 (N_22658,N_22550,N_22549);
nand U22659 (N_22659,N_22411,N_22558);
nand U22660 (N_22660,N_22520,N_22534);
nor U22661 (N_22661,N_22435,N_22598);
and U22662 (N_22662,N_22592,N_22473);
or U22663 (N_22663,N_22516,N_22433);
nand U22664 (N_22664,N_22430,N_22527);
and U22665 (N_22665,N_22404,N_22505);
nor U22666 (N_22666,N_22491,N_22405);
xor U22667 (N_22667,N_22407,N_22487);
nor U22668 (N_22668,N_22580,N_22402);
xor U22669 (N_22669,N_22422,N_22479);
xnor U22670 (N_22670,N_22465,N_22484);
xor U22671 (N_22671,N_22544,N_22535);
nand U22672 (N_22672,N_22429,N_22576);
nand U22673 (N_22673,N_22428,N_22591);
xor U22674 (N_22674,N_22444,N_22564);
or U22675 (N_22675,N_22538,N_22559);
nor U22676 (N_22676,N_22448,N_22427);
nand U22677 (N_22677,N_22480,N_22532);
nor U22678 (N_22678,N_22540,N_22548);
nor U22679 (N_22679,N_22468,N_22521);
nor U22680 (N_22680,N_22470,N_22599);
nor U22681 (N_22681,N_22511,N_22463);
or U22682 (N_22682,N_22552,N_22436);
xnor U22683 (N_22683,N_22501,N_22526);
xor U22684 (N_22684,N_22514,N_22471);
or U22685 (N_22685,N_22546,N_22504);
nand U22686 (N_22686,N_22438,N_22597);
and U22687 (N_22687,N_22499,N_22492);
nand U22688 (N_22688,N_22530,N_22519);
or U22689 (N_22689,N_22426,N_22472);
or U22690 (N_22690,N_22583,N_22593);
nand U22691 (N_22691,N_22496,N_22506);
nand U22692 (N_22692,N_22539,N_22401);
xor U22693 (N_22693,N_22450,N_22488);
and U22694 (N_22694,N_22483,N_22440);
nor U22695 (N_22695,N_22419,N_22459);
and U22696 (N_22696,N_22509,N_22523);
and U22697 (N_22697,N_22542,N_22525);
nand U22698 (N_22698,N_22449,N_22541);
xnor U22699 (N_22699,N_22477,N_22557);
nand U22700 (N_22700,N_22497,N_22514);
nor U22701 (N_22701,N_22574,N_22479);
or U22702 (N_22702,N_22572,N_22597);
or U22703 (N_22703,N_22508,N_22501);
nand U22704 (N_22704,N_22571,N_22412);
nand U22705 (N_22705,N_22560,N_22415);
xnor U22706 (N_22706,N_22484,N_22570);
and U22707 (N_22707,N_22436,N_22476);
and U22708 (N_22708,N_22591,N_22498);
nor U22709 (N_22709,N_22479,N_22487);
or U22710 (N_22710,N_22486,N_22540);
and U22711 (N_22711,N_22580,N_22413);
and U22712 (N_22712,N_22402,N_22520);
nand U22713 (N_22713,N_22556,N_22545);
xnor U22714 (N_22714,N_22510,N_22438);
or U22715 (N_22715,N_22579,N_22444);
and U22716 (N_22716,N_22502,N_22520);
nor U22717 (N_22717,N_22408,N_22594);
and U22718 (N_22718,N_22559,N_22452);
xnor U22719 (N_22719,N_22579,N_22408);
and U22720 (N_22720,N_22479,N_22409);
nor U22721 (N_22721,N_22446,N_22561);
or U22722 (N_22722,N_22507,N_22524);
nand U22723 (N_22723,N_22462,N_22493);
xnor U22724 (N_22724,N_22519,N_22501);
nand U22725 (N_22725,N_22593,N_22433);
or U22726 (N_22726,N_22586,N_22406);
or U22727 (N_22727,N_22420,N_22558);
xnor U22728 (N_22728,N_22520,N_22595);
or U22729 (N_22729,N_22491,N_22587);
and U22730 (N_22730,N_22488,N_22533);
and U22731 (N_22731,N_22430,N_22585);
nand U22732 (N_22732,N_22512,N_22573);
or U22733 (N_22733,N_22446,N_22481);
nor U22734 (N_22734,N_22528,N_22490);
nand U22735 (N_22735,N_22483,N_22461);
and U22736 (N_22736,N_22579,N_22566);
xnor U22737 (N_22737,N_22427,N_22482);
nor U22738 (N_22738,N_22460,N_22557);
and U22739 (N_22739,N_22483,N_22587);
or U22740 (N_22740,N_22501,N_22515);
or U22741 (N_22741,N_22534,N_22591);
nor U22742 (N_22742,N_22550,N_22552);
nand U22743 (N_22743,N_22400,N_22521);
and U22744 (N_22744,N_22499,N_22509);
nor U22745 (N_22745,N_22546,N_22563);
xor U22746 (N_22746,N_22422,N_22526);
xor U22747 (N_22747,N_22482,N_22589);
and U22748 (N_22748,N_22448,N_22458);
xor U22749 (N_22749,N_22511,N_22538);
or U22750 (N_22750,N_22571,N_22425);
xor U22751 (N_22751,N_22533,N_22540);
nand U22752 (N_22752,N_22410,N_22588);
and U22753 (N_22753,N_22473,N_22542);
nor U22754 (N_22754,N_22497,N_22484);
and U22755 (N_22755,N_22589,N_22580);
and U22756 (N_22756,N_22447,N_22476);
nand U22757 (N_22757,N_22475,N_22599);
and U22758 (N_22758,N_22453,N_22543);
xor U22759 (N_22759,N_22525,N_22509);
xnor U22760 (N_22760,N_22526,N_22481);
nor U22761 (N_22761,N_22498,N_22444);
xor U22762 (N_22762,N_22400,N_22476);
nor U22763 (N_22763,N_22436,N_22491);
and U22764 (N_22764,N_22472,N_22571);
and U22765 (N_22765,N_22414,N_22405);
nor U22766 (N_22766,N_22429,N_22552);
or U22767 (N_22767,N_22454,N_22513);
xor U22768 (N_22768,N_22434,N_22554);
nor U22769 (N_22769,N_22585,N_22495);
or U22770 (N_22770,N_22574,N_22449);
or U22771 (N_22771,N_22559,N_22403);
nand U22772 (N_22772,N_22546,N_22594);
nor U22773 (N_22773,N_22495,N_22542);
and U22774 (N_22774,N_22518,N_22405);
nand U22775 (N_22775,N_22458,N_22461);
nor U22776 (N_22776,N_22413,N_22485);
nor U22777 (N_22777,N_22531,N_22529);
nor U22778 (N_22778,N_22469,N_22589);
and U22779 (N_22779,N_22425,N_22508);
nor U22780 (N_22780,N_22466,N_22426);
nor U22781 (N_22781,N_22520,N_22596);
or U22782 (N_22782,N_22548,N_22416);
nor U22783 (N_22783,N_22589,N_22517);
xor U22784 (N_22784,N_22453,N_22503);
xnor U22785 (N_22785,N_22482,N_22440);
or U22786 (N_22786,N_22506,N_22509);
or U22787 (N_22787,N_22535,N_22566);
and U22788 (N_22788,N_22431,N_22488);
nor U22789 (N_22789,N_22424,N_22558);
or U22790 (N_22790,N_22457,N_22576);
xor U22791 (N_22791,N_22518,N_22548);
and U22792 (N_22792,N_22457,N_22540);
nand U22793 (N_22793,N_22412,N_22544);
nor U22794 (N_22794,N_22525,N_22408);
and U22795 (N_22795,N_22534,N_22564);
and U22796 (N_22796,N_22495,N_22559);
and U22797 (N_22797,N_22598,N_22404);
nor U22798 (N_22798,N_22578,N_22488);
nor U22799 (N_22799,N_22420,N_22568);
xor U22800 (N_22800,N_22616,N_22752);
nor U22801 (N_22801,N_22617,N_22639);
xor U22802 (N_22802,N_22736,N_22675);
or U22803 (N_22803,N_22691,N_22648);
and U22804 (N_22804,N_22710,N_22660);
nand U22805 (N_22805,N_22677,N_22731);
and U22806 (N_22806,N_22608,N_22738);
or U22807 (N_22807,N_22681,N_22605);
xor U22808 (N_22808,N_22651,N_22729);
nand U22809 (N_22809,N_22601,N_22786);
xnor U22810 (N_22810,N_22743,N_22694);
or U22811 (N_22811,N_22705,N_22603);
nor U22812 (N_22812,N_22636,N_22781);
xnor U22813 (N_22813,N_22655,N_22707);
and U22814 (N_22814,N_22645,N_22600);
nor U22815 (N_22815,N_22700,N_22610);
and U22816 (N_22816,N_22785,N_22627);
nor U22817 (N_22817,N_22638,N_22757);
and U22818 (N_22818,N_22673,N_22719);
or U22819 (N_22819,N_22614,N_22797);
or U22820 (N_22820,N_22630,N_22782);
nor U22821 (N_22821,N_22754,N_22606);
nor U22822 (N_22822,N_22733,N_22658);
or U22823 (N_22823,N_22696,N_22748);
and U22824 (N_22824,N_22634,N_22721);
nand U22825 (N_22825,N_22724,N_22667);
and U22826 (N_22826,N_22794,N_22779);
nand U22827 (N_22827,N_22650,N_22625);
nor U22828 (N_22828,N_22713,N_22626);
or U22829 (N_22829,N_22697,N_22756);
nor U22830 (N_22830,N_22602,N_22720);
nor U22831 (N_22831,N_22665,N_22780);
nor U22832 (N_22832,N_22722,N_22760);
nor U22833 (N_22833,N_22633,N_22726);
xnor U22834 (N_22834,N_22747,N_22799);
or U22835 (N_22835,N_22755,N_22668);
xor U22836 (N_22836,N_22611,N_22764);
xor U22837 (N_22837,N_22787,N_22690);
or U22838 (N_22838,N_22661,N_22604);
xor U22839 (N_22839,N_22740,N_22678);
or U22840 (N_22840,N_22663,N_22659);
nand U22841 (N_22841,N_22615,N_22620);
xor U22842 (N_22842,N_22766,N_22687);
nand U22843 (N_22843,N_22749,N_22623);
nor U22844 (N_22844,N_22784,N_22763);
and U22845 (N_22845,N_22772,N_22709);
and U22846 (N_22846,N_22684,N_22708);
and U22847 (N_22847,N_22621,N_22717);
nand U22848 (N_22848,N_22613,N_22783);
and U22849 (N_22849,N_22618,N_22657);
nor U22850 (N_22850,N_22656,N_22649);
and U22851 (N_22851,N_22742,N_22622);
or U22852 (N_22852,N_22686,N_22664);
and U22853 (N_22853,N_22695,N_22685);
or U22854 (N_22854,N_22632,N_22641);
xor U22855 (N_22855,N_22716,N_22728);
or U22856 (N_22856,N_22727,N_22771);
and U22857 (N_22857,N_22778,N_22777);
nand U22858 (N_22858,N_22741,N_22790);
and U22859 (N_22859,N_22635,N_22746);
nand U22860 (N_22860,N_22624,N_22789);
and U22861 (N_22861,N_22793,N_22737);
xnor U22862 (N_22862,N_22699,N_22672);
xnor U22863 (N_22863,N_22765,N_22642);
nor U22864 (N_22864,N_22739,N_22674);
and U22865 (N_22865,N_22683,N_22770);
or U22866 (N_22866,N_22671,N_22706);
nor U22867 (N_22867,N_22703,N_22725);
or U22868 (N_22868,N_22776,N_22669);
and U22869 (N_22869,N_22612,N_22732);
or U22870 (N_22870,N_22775,N_22734);
or U22871 (N_22871,N_22792,N_22682);
or U22872 (N_22872,N_22744,N_22640);
or U22873 (N_22873,N_22718,N_22712);
nor U22874 (N_22874,N_22619,N_22735);
and U22875 (N_22875,N_22628,N_22670);
and U22876 (N_22876,N_22761,N_22796);
and U22877 (N_22877,N_22769,N_22704);
nand U22878 (N_22878,N_22689,N_22688);
xnor U22879 (N_22879,N_22750,N_22654);
or U22880 (N_22880,N_22759,N_22774);
nand U22881 (N_22881,N_22767,N_22676);
or U22882 (N_22882,N_22631,N_22788);
and U22883 (N_22883,N_22773,N_22652);
or U22884 (N_22884,N_22791,N_22653);
xnor U22885 (N_22885,N_22753,N_22730);
and U22886 (N_22886,N_22607,N_22711);
or U22887 (N_22887,N_22702,N_22680);
and U22888 (N_22888,N_22679,N_22723);
nor U22889 (N_22889,N_22758,N_22662);
xnor U22890 (N_22890,N_22701,N_22698);
xnor U22891 (N_22891,N_22629,N_22692);
nor U22892 (N_22892,N_22609,N_22647);
and U22893 (N_22893,N_22643,N_22768);
or U22894 (N_22894,N_22714,N_22646);
xor U22895 (N_22895,N_22715,N_22798);
nand U22896 (N_22896,N_22745,N_22762);
nand U22897 (N_22897,N_22751,N_22795);
nand U22898 (N_22898,N_22637,N_22644);
or U22899 (N_22899,N_22693,N_22666);
nand U22900 (N_22900,N_22737,N_22603);
or U22901 (N_22901,N_22774,N_22766);
and U22902 (N_22902,N_22706,N_22767);
and U22903 (N_22903,N_22706,N_22781);
or U22904 (N_22904,N_22794,N_22699);
and U22905 (N_22905,N_22795,N_22614);
nor U22906 (N_22906,N_22621,N_22716);
nand U22907 (N_22907,N_22663,N_22796);
or U22908 (N_22908,N_22792,N_22629);
or U22909 (N_22909,N_22769,N_22674);
nand U22910 (N_22910,N_22797,N_22675);
nor U22911 (N_22911,N_22725,N_22609);
and U22912 (N_22912,N_22798,N_22683);
or U22913 (N_22913,N_22617,N_22683);
and U22914 (N_22914,N_22733,N_22742);
nor U22915 (N_22915,N_22617,N_22714);
nand U22916 (N_22916,N_22767,N_22722);
or U22917 (N_22917,N_22658,N_22695);
and U22918 (N_22918,N_22671,N_22684);
xnor U22919 (N_22919,N_22741,N_22630);
and U22920 (N_22920,N_22607,N_22633);
nor U22921 (N_22921,N_22635,N_22655);
and U22922 (N_22922,N_22605,N_22644);
xor U22923 (N_22923,N_22678,N_22674);
nor U22924 (N_22924,N_22673,N_22641);
or U22925 (N_22925,N_22725,N_22702);
and U22926 (N_22926,N_22694,N_22614);
and U22927 (N_22927,N_22702,N_22733);
or U22928 (N_22928,N_22644,N_22755);
nor U22929 (N_22929,N_22615,N_22675);
or U22930 (N_22930,N_22768,N_22645);
nor U22931 (N_22931,N_22607,N_22618);
and U22932 (N_22932,N_22620,N_22699);
and U22933 (N_22933,N_22614,N_22793);
nand U22934 (N_22934,N_22688,N_22637);
and U22935 (N_22935,N_22610,N_22640);
xnor U22936 (N_22936,N_22741,N_22693);
nand U22937 (N_22937,N_22751,N_22623);
or U22938 (N_22938,N_22680,N_22705);
and U22939 (N_22939,N_22613,N_22781);
nor U22940 (N_22940,N_22754,N_22621);
nor U22941 (N_22941,N_22761,N_22654);
or U22942 (N_22942,N_22626,N_22706);
nor U22943 (N_22943,N_22783,N_22667);
nor U22944 (N_22944,N_22685,N_22652);
nand U22945 (N_22945,N_22765,N_22762);
nor U22946 (N_22946,N_22769,N_22696);
xor U22947 (N_22947,N_22695,N_22764);
or U22948 (N_22948,N_22642,N_22780);
xor U22949 (N_22949,N_22769,N_22709);
nand U22950 (N_22950,N_22635,N_22607);
or U22951 (N_22951,N_22665,N_22649);
or U22952 (N_22952,N_22792,N_22785);
nand U22953 (N_22953,N_22727,N_22656);
and U22954 (N_22954,N_22684,N_22702);
or U22955 (N_22955,N_22644,N_22688);
nand U22956 (N_22956,N_22683,N_22727);
nand U22957 (N_22957,N_22615,N_22608);
xor U22958 (N_22958,N_22788,N_22778);
nand U22959 (N_22959,N_22656,N_22762);
nand U22960 (N_22960,N_22734,N_22646);
xnor U22961 (N_22961,N_22791,N_22689);
and U22962 (N_22962,N_22664,N_22633);
xnor U22963 (N_22963,N_22635,N_22761);
nor U22964 (N_22964,N_22614,N_22732);
or U22965 (N_22965,N_22604,N_22653);
nand U22966 (N_22966,N_22689,N_22771);
nand U22967 (N_22967,N_22726,N_22634);
nor U22968 (N_22968,N_22682,N_22645);
or U22969 (N_22969,N_22652,N_22742);
xnor U22970 (N_22970,N_22725,N_22745);
xnor U22971 (N_22971,N_22756,N_22719);
nor U22972 (N_22972,N_22680,N_22772);
xnor U22973 (N_22973,N_22649,N_22788);
or U22974 (N_22974,N_22670,N_22650);
xnor U22975 (N_22975,N_22638,N_22700);
xnor U22976 (N_22976,N_22745,N_22651);
xor U22977 (N_22977,N_22707,N_22731);
nand U22978 (N_22978,N_22736,N_22731);
nand U22979 (N_22979,N_22783,N_22693);
nor U22980 (N_22980,N_22631,N_22746);
xnor U22981 (N_22981,N_22724,N_22741);
xor U22982 (N_22982,N_22713,N_22753);
or U22983 (N_22983,N_22754,N_22604);
and U22984 (N_22984,N_22673,N_22707);
and U22985 (N_22985,N_22754,N_22655);
xor U22986 (N_22986,N_22725,N_22784);
nand U22987 (N_22987,N_22665,N_22640);
or U22988 (N_22988,N_22664,N_22698);
nand U22989 (N_22989,N_22699,N_22718);
nand U22990 (N_22990,N_22651,N_22734);
xnor U22991 (N_22991,N_22777,N_22640);
or U22992 (N_22992,N_22642,N_22758);
and U22993 (N_22993,N_22719,N_22675);
xnor U22994 (N_22994,N_22794,N_22791);
xor U22995 (N_22995,N_22741,N_22667);
nor U22996 (N_22996,N_22755,N_22761);
nor U22997 (N_22997,N_22729,N_22614);
nor U22998 (N_22998,N_22768,N_22672);
xnor U22999 (N_22999,N_22671,N_22679);
nor U23000 (N_23000,N_22865,N_22819);
xnor U23001 (N_23001,N_22999,N_22876);
xor U23002 (N_23002,N_22996,N_22880);
or U23003 (N_23003,N_22981,N_22831);
nand U23004 (N_23004,N_22830,N_22821);
nor U23005 (N_23005,N_22995,N_22861);
nor U23006 (N_23006,N_22839,N_22976);
or U23007 (N_23007,N_22935,N_22939);
or U23008 (N_23008,N_22825,N_22900);
xnor U23009 (N_23009,N_22911,N_22932);
nor U23010 (N_23010,N_22841,N_22930);
nor U23011 (N_23011,N_22970,N_22853);
xnor U23012 (N_23012,N_22804,N_22964);
nor U23013 (N_23013,N_22848,N_22815);
xnor U23014 (N_23014,N_22800,N_22901);
nor U23015 (N_23015,N_22884,N_22818);
and U23016 (N_23016,N_22951,N_22855);
or U23017 (N_23017,N_22802,N_22857);
or U23018 (N_23018,N_22994,N_22931);
or U23019 (N_23019,N_22806,N_22927);
xor U23020 (N_23020,N_22950,N_22858);
and U23021 (N_23021,N_22974,N_22875);
nor U23022 (N_23022,N_22835,N_22902);
or U23023 (N_23023,N_22938,N_22953);
nand U23024 (N_23024,N_22898,N_22895);
xnor U23025 (N_23025,N_22940,N_22822);
and U23026 (N_23026,N_22920,N_22984);
and U23027 (N_23027,N_22879,N_22922);
and U23028 (N_23028,N_22980,N_22917);
nand U23029 (N_23029,N_22811,N_22833);
and U23030 (N_23030,N_22892,N_22993);
nor U23031 (N_23031,N_22870,N_22842);
xnor U23032 (N_23032,N_22838,N_22967);
or U23033 (N_23033,N_22828,N_22867);
nand U23034 (N_23034,N_22992,N_22918);
xnor U23035 (N_23035,N_22899,N_22873);
and U23036 (N_23036,N_22845,N_22891);
or U23037 (N_23037,N_22947,N_22864);
xnor U23038 (N_23038,N_22926,N_22913);
and U23039 (N_23039,N_22943,N_22933);
nor U23040 (N_23040,N_22937,N_22854);
nor U23041 (N_23041,N_22890,N_22960);
or U23042 (N_23042,N_22908,N_22972);
xor U23043 (N_23043,N_22924,N_22897);
nor U23044 (N_23044,N_22881,N_22948);
xor U23045 (N_23045,N_22871,N_22836);
and U23046 (N_23046,N_22820,N_22945);
nand U23047 (N_23047,N_22962,N_22889);
and U23048 (N_23048,N_22847,N_22949);
and U23049 (N_23049,N_22987,N_22921);
nor U23050 (N_23050,N_22968,N_22837);
nand U23051 (N_23051,N_22843,N_22934);
xor U23052 (N_23052,N_22966,N_22941);
or U23053 (N_23053,N_22963,N_22827);
nand U23054 (N_23054,N_22975,N_22810);
nand U23055 (N_23055,N_22872,N_22869);
xor U23056 (N_23056,N_22813,N_22958);
and U23057 (N_23057,N_22936,N_22840);
xnor U23058 (N_23058,N_22803,N_22971);
and U23059 (N_23059,N_22979,N_22894);
and U23060 (N_23060,N_22834,N_22801);
nor U23061 (N_23061,N_22978,N_22832);
xor U23062 (N_23062,N_22903,N_22849);
nand U23063 (N_23063,N_22859,N_22956);
and U23064 (N_23064,N_22977,N_22883);
nor U23065 (N_23065,N_22905,N_22896);
nand U23066 (N_23066,N_22997,N_22805);
nor U23067 (N_23067,N_22816,N_22959);
and U23068 (N_23068,N_22906,N_22928);
xor U23069 (N_23069,N_22916,N_22874);
or U23070 (N_23070,N_22965,N_22985);
or U23071 (N_23071,N_22946,N_22860);
and U23072 (N_23072,N_22808,N_22929);
and U23073 (N_23073,N_22912,N_22893);
and U23074 (N_23074,N_22983,N_22907);
nor U23075 (N_23075,N_22851,N_22923);
and U23076 (N_23076,N_22925,N_22807);
nand U23077 (N_23077,N_22868,N_22882);
nand U23078 (N_23078,N_22988,N_22910);
and U23079 (N_23079,N_22990,N_22852);
and U23080 (N_23080,N_22904,N_22850);
and U23081 (N_23081,N_22824,N_22846);
and U23082 (N_23082,N_22955,N_22919);
nand U23083 (N_23083,N_22812,N_22844);
nor U23084 (N_23084,N_22989,N_22973);
and U23085 (N_23085,N_22914,N_22969);
xnor U23086 (N_23086,N_22952,N_22866);
nor U23087 (N_23087,N_22885,N_22877);
or U23088 (N_23088,N_22942,N_22863);
nand U23089 (N_23089,N_22915,N_22878);
nand U23090 (N_23090,N_22909,N_22856);
and U23091 (N_23091,N_22823,N_22957);
and U23092 (N_23092,N_22888,N_22991);
nor U23093 (N_23093,N_22944,N_22829);
nor U23094 (N_23094,N_22998,N_22817);
nor U23095 (N_23095,N_22982,N_22826);
xor U23096 (N_23096,N_22886,N_22809);
nand U23097 (N_23097,N_22954,N_22814);
xnor U23098 (N_23098,N_22961,N_22986);
nand U23099 (N_23099,N_22862,N_22887);
and U23100 (N_23100,N_22920,N_22898);
nor U23101 (N_23101,N_22804,N_22874);
xnor U23102 (N_23102,N_22981,N_22838);
and U23103 (N_23103,N_22891,N_22812);
nand U23104 (N_23104,N_22942,N_22864);
nor U23105 (N_23105,N_22974,N_22991);
and U23106 (N_23106,N_22913,N_22932);
or U23107 (N_23107,N_22911,N_22816);
or U23108 (N_23108,N_22861,N_22940);
and U23109 (N_23109,N_22800,N_22893);
and U23110 (N_23110,N_22897,N_22902);
and U23111 (N_23111,N_22926,N_22994);
or U23112 (N_23112,N_22922,N_22917);
nor U23113 (N_23113,N_22988,N_22920);
nor U23114 (N_23114,N_22879,N_22971);
nor U23115 (N_23115,N_22830,N_22876);
and U23116 (N_23116,N_22875,N_22890);
or U23117 (N_23117,N_22857,N_22826);
and U23118 (N_23118,N_22986,N_22890);
nor U23119 (N_23119,N_22818,N_22861);
nor U23120 (N_23120,N_22817,N_22852);
or U23121 (N_23121,N_22968,N_22910);
nand U23122 (N_23122,N_22947,N_22830);
nor U23123 (N_23123,N_22829,N_22999);
nand U23124 (N_23124,N_22807,N_22954);
xnor U23125 (N_23125,N_22862,N_22924);
nor U23126 (N_23126,N_22848,N_22875);
and U23127 (N_23127,N_22854,N_22892);
and U23128 (N_23128,N_22886,N_22844);
and U23129 (N_23129,N_22951,N_22961);
xor U23130 (N_23130,N_22839,N_22916);
xor U23131 (N_23131,N_22905,N_22926);
xnor U23132 (N_23132,N_22873,N_22931);
nand U23133 (N_23133,N_22991,N_22816);
or U23134 (N_23134,N_22803,N_22930);
nand U23135 (N_23135,N_22866,N_22937);
and U23136 (N_23136,N_22841,N_22806);
nor U23137 (N_23137,N_22819,N_22848);
and U23138 (N_23138,N_22893,N_22824);
xor U23139 (N_23139,N_22870,N_22864);
nor U23140 (N_23140,N_22907,N_22853);
and U23141 (N_23141,N_22941,N_22994);
and U23142 (N_23142,N_22878,N_22929);
nand U23143 (N_23143,N_22963,N_22923);
or U23144 (N_23144,N_22905,N_22954);
nand U23145 (N_23145,N_22997,N_22905);
nand U23146 (N_23146,N_22920,N_22936);
xnor U23147 (N_23147,N_22892,N_22804);
xnor U23148 (N_23148,N_22981,N_22918);
xor U23149 (N_23149,N_22980,N_22896);
nor U23150 (N_23150,N_22947,N_22802);
xor U23151 (N_23151,N_22810,N_22988);
xnor U23152 (N_23152,N_22805,N_22942);
or U23153 (N_23153,N_22999,N_22996);
nor U23154 (N_23154,N_22929,N_22902);
and U23155 (N_23155,N_22931,N_22937);
or U23156 (N_23156,N_22833,N_22956);
or U23157 (N_23157,N_22991,N_22936);
and U23158 (N_23158,N_22984,N_22818);
xnor U23159 (N_23159,N_22811,N_22858);
or U23160 (N_23160,N_22938,N_22921);
xnor U23161 (N_23161,N_22812,N_22926);
xor U23162 (N_23162,N_22959,N_22935);
xnor U23163 (N_23163,N_22947,N_22921);
nor U23164 (N_23164,N_22892,N_22991);
and U23165 (N_23165,N_22909,N_22945);
and U23166 (N_23166,N_22960,N_22905);
nand U23167 (N_23167,N_22876,N_22814);
nor U23168 (N_23168,N_22951,N_22904);
and U23169 (N_23169,N_22899,N_22963);
and U23170 (N_23170,N_22914,N_22963);
or U23171 (N_23171,N_22831,N_22979);
nand U23172 (N_23172,N_22847,N_22939);
and U23173 (N_23173,N_22854,N_22996);
nand U23174 (N_23174,N_22936,N_22919);
xor U23175 (N_23175,N_22807,N_22936);
nor U23176 (N_23176,N_22852,N_22811);
or U23177 (N_23177,N_22818,N_22837);
and U23178 (N_23178,N_22958,N_22881);
or U23179 (N_23179,N_22800,N_22962);
or U23180 (N_23180,N_22816,N_22831);
nand U23181 (N_23181,N_22881,N_22957);
xor U23182 (N_23182,N_22866,N_22998);
and U23183 (N_23183,N_22838,N_22800);
or U23184 (N_23184,N_22878,N_22938);
xor U23185 (N_23185,N_22859,N_22909);
or U23186 (N_23186,N_22860,N_22925);
xnor U23187 (N_23187,N_22963,N_22897);
xor U23188 (N_23188,N_22933,N_22905);
or U23189 (N_23189,N_22952,N_22902);
or U23190 (N_23190,N_22902,N_22963);
xor U23191 (N_23191,N_22937,N_22842);
nor U23192 (N_23192,N_22812,N_22927);
or U23193 (N_23193,N_22812,N_22958);
xor U23194 (N_23194,N_22906,N_22808);
or U23195 (N_23195,N_22846,N_22919);
nand U23196 (N_23196,N_22837,N_22819);
xor U23197 (N_23197,N_22864,N_22805);
nor U23198 (N_23198,N_22839,N_22902);
or U23199 (N_23199,N_22821,N_22838);
xnor U23200 (N_23200,N_23148,N_23080);
nand U23201 (N_23201,N_23081,N_23175);
or U23202 (N_23202,N_23180,N_23100);
nand U23203 (N_23203,N_23197,N_23031);
or U23204 (N_23204,N_23196,N_23154);
nor U23205 (N_23205,N_23063,N_23064);
or U23206 (N_23206,N_23158,N_23141);
xor U23207 (N_23207,N_23007,N_23094);
xnor U23208 (N_23208,N_23005,N_23170);
nor U23209 (N_23209,N_23190,N_23042);
nor U23210 (N_23210,N_23013,N_23161);
and U23211 (N_23211,N_23126,N_23073);
or U23212 (N_23212,N_23066,N_23095);
and U23213 (N_23213,N_23118,N_23183);
nand U23214 (N_23214,N_23068,N_23167);
or U23215 (N_23215,N_23146,N_23039);
nor U23216 (N_23216,N_23150,N_23016);
or U23217 (N_23217,N_23067,N_23113);
and U23218 (N_23218,N_23033,N_23134);
nand U23219 (N_23219,N_23105,N_23090);
nand U23220 (N_23220,N_23050,N_23179);
nand U23221 (N_23221,N_23143,N_23117);
nor U23222 (N_23222,N_23120,N_23099);
xor U23223 (N_23223,N_23124,N_23145);
nand U23224 (N_23224,N_23054,N_23109);
or U23225 (N_23225,N_23058,N_23025);
or U23226 (N_23226,N_23135,N_23041);
xnor U23227 (N_23227,N_23168,N_23122);
xnor U23228 (N_23228,N_23087,N_23053);
nor U23229 (N_23229,N_23102,N_23116);
nand U23230 (N_23230,N_23075,N_23159);
xnor U23231 (N_23231,N_23079,N_23106);
xnor U23232 (N_23232,N_23115,N_23009);
nand U23233 (N_23233,N_23026,N_23084);
or U23234 (N_23234,N_23028,N_23037);
and U23235 (N_23235,N_23089,N_23119);
nand U23236 (N_23236,N_23078,N_23070);
or U23237 (N_23237,N_23011,N_23131);
or U23238 (N_23238,N_23128,N_23055);
nand U23239 (N_23239,N_23085,N_23108);
and U23240 (N_23240,N_23022,N_23166);
or U23241 (N_23241,N_23060,N_23072);
and U23242 (N_23242,N_23097,N_23133);
nand U23243 (N_23243,N_23047,N_23049);
or U23244 (N_23244,N_23151,N_23184);
nand U23245 (N_23245,N_23069,N_23176);
nand U23246 (N_23246,N_23110,N_23012);
and U23247 (N_23247,N_23173,N_23125);
nor U23248 (N_23248,N_23149,N_23027);
and U23249 (N_23249,N_23059,N_23144);
and U23250 (N_23250,N_23169,N_23040);
xnor U23251 (N_23251,N_23136,N_23017);
nand U23252 (N_23252,N_23130,N_23043);
nand U23253 (N_23253,N_23199,N_23062);
nand U23254 (N_23254,N_23061,N_23123);
nand U23255 (N_23255,N_23103,N_23098);
nand U23256 (N_23256,N_23091,N_23004);
and U23257 (N_23257,N_23019,N_23164);
nand U23258 (N_23258,N_23153,N_23138);
nor U23259 (N_23259,N_23194,N_23142);
and U23260 (N_23260,N_23077,N_23181);
nor U23261 (N_23261,N_23003,N_23147);
xnor U23262 (N_23262,N_23177,N_23046);
nor U23263 (N_23263,N_23178,N_23185);
xor U23264 (N_23264,N_23023,N_23000);
nand U23265 (N_23265,N_23056,N_23076);
or U23266 (N_23266,N_23140,N_23018);
nor U23267 (N_23267,N_23074,N_23065);
and U23268 (N_23268,N_23052,N_23034);
or U23269 (N_23269,N_23030,N_23157);
xor U23270 (N_23270,N_23189,N_23048);
and U23271 (N_23271,N_23127,N_23051);
or U23272 (N_23272,N_23156,N_23163);
or U23273 (N_23273,N_23015,N_23137);
nor U23274 (N_23274,N_23086,N_23191);
nor U23275 (N_23275,N_23032,N_23107);
xor U23276 (N_23276,N_23193,N_23024);
or U23277 (N_23277,N_23171,N_23008);
nand U23278 (N_23278,N_23198,N_23083);
and U23279 (N_23279,N_23014,N_23021);
or U23280 (N_23280,N_23038,N_23035);
or U23281 (N_23281,N_23001,N_23088);
or U23282 (N_23282,N_23162,N_23045);
nor U23283 (N_23283,N_23186,N_23036);
nand U23284 (N_23284,N_23111,N_23188);
or U23285 (N_23285,N_23101,N_23029);
and U23286 (N_23286,N_23182,N_23192);
or U23287 (N_23287,N_23071,N_23132);
nor U23288 (N_23288,N_23152,N_23093);
and U23289 (N_23289,N_23121,N_23044);
nand U23290 (N_23290,N_23187,N_23010);
nor U23291 (N_23291,N_23195,N_23139);
nand U23292 (N_23292,N_23155,N_23112);
nor U23293 (N_23293,N_23082,N_23057);
nand U23294 (N_23294,N_23114,N_23020);
nand U23295 (N_23295,N_23174,N_23172);
or U23296 (N_23296,N_23092,N_23006);
nand U23297 (N_23297,N_23002,N_23160);
or U23298 (N_23298,N_23104,N_23165);
and U23299 (N_23299,N_23096,N_23129);
and U23300 (N_23300,N_23141,N_23154);
or U23301 (N_23301,N_23055,N_23000);
and U23302 (N_23302,N_23140,N_23001);
nand U23303 (N_23303,N_23038,N_23157);
and U23304 (N_23304,N_23076,N_23080);
or U23305 (N_23305,N_23042,N_23067);
nor U23306 (N_23306,N_23016,N_23042);
or U23307 (N_23307,N_23148,N_23097);
or U23308 (N_23308,N_23059,N_23150);
nand U23309 (N_23309,N_23157,N_23004);
or U23310 (N_23310,N_23108,N_23121);
nand U23311 (N_23311,N_23046,N_23118);
nand U23312 (N_23312,N_23101,N_23043);
xor U23313 (N_23313,N_23158,N_23166);
nor U23314 (N_23314,N_23188,N_23103);
or U23315 (N_23315,N_23032,N_23137);
nand U23316 (N_23316,N_23054,N_23175);
nand U23317 (N_23317,N_23074,N_23053);
and U23318 (N_23318,N_23170,N_23136);
and U23319 (N_23319,N_23014,N_23166);
nor U23320 (N_23320,N_23148,N_23049);
nand U23321 (N_23321,N_23199,N_23118);
or U23322 (N_23322,N_23067,N_23184);
xnor U23323 (N_23323,N_23109,N_23173);
and U23324 (N_23324,N_23130,N_23127);
nand U23325 (N_23325,N_23007,N_23153);
nand U23326 (N_23326,N_23078,N_23083);
and U23327 (N_23327,N_23036,N_23127);
nand U23328 (N_23328,N_23123,N_23137);
or U23329 (N_23329,N_23150,N_23006);
xor U23330 (N_23330,N_23156,N_23161);
xnor U23331 (N_23331,N_23015,N_23063);
or U23332 (N_23332,N_23128,N_23157);
or U23333 (N_23333,N_23184,N_23061);
xnor U23334 (N_23334,N_23063,N_23005);
nand U23335 (N_23335,N_23141,N_23145);
and U23336 (N_23336,N_23180,N_23012);
nor U23337 (N_23337,N_23079,N_23063);
nand U23338 (N_23338,N_23116,N_23170);
or U23339 (N_23339,N_23074,N_23154);
nand U23340 (N_23340,N_23114,N_23123);
or U23341 (N_23341,N_23155,N_23140);
nand U23342 (N_23342,N_23074,N_23187);
nor U23343 (N_23343,N_23120,N_23105);
nand U23344 (N_23344,N_23129,N_23156);
and U23345 (N_23345,N_23118,N_23069);
nand U23346 (N_23346,N_23044,N_23168);
or U23347 (N_23347,N_23188,N_23115);
xnor U23348 (N_23348,N_23048,N_23129);
nand U23349 (N_23349,N_23003,N_23192);
nand U23350 (N_23350,N_23134,N_23074);
or U23351 (N_23351,N_23031,N_23010);
nand U23352 (N_23352,N_23102,N_23065);
nand U23353 (N_23353,N_23057,N_23075);
and U23354 (N_23354,N_23055,N_23065);
xor U23355 (N_23355,N_23125,N_23113);
and U23356 (N_23356,N_23151,N_23074);
xor U23357 (N_23357,N_23093,N_23192);
or U23358 (N_23358,N_23132,N_23064);
xnor U23359 (N_23359,N_23177,N_23023);
nand U23360 (N_23360,N_23080,N_23190);
xnor U23361 (N_23361,N_23090,N_23053);
nor U23362 (N_23362,N_23007,N_23171);
nor U23363 (N_23363,N_23128,N_23161);
or U23364 (N_23364,N_23117,N_23099);
and U23365 (N_23365,N_23000,N_23085);
and U23366 (N_23366,N_23103,N_23191);
nor U23367 (N_23367,N_23128,N_23126);
or U23368 (N_23368,N_23147,N_23177);
and U23369 (N_23369,N_23064,N_23116);
xor U23370 (N_23370,N_23023,N_23086);
nand U23371 (N_23371,N_23093,N_23080);
and U23372 (N_23372,N_23001,N_23097);
nor U23373 (N_23373,N_23066,N_23051);
xnor U23374 (N_23374,N_23148,N_23016);
xor U23375 (N_23375,N_23100,N_23151);
or U23376 (N_23376,N_23013,N_23182);
nor U23377 (N_23377,N_23117,N_23024);
xor U23378 (N_23378,N_23199,N_23009);
or U23379 (N_23379,N_23164,N_23047);
nor U23380 (N_23380,N_23144,N_23156);
and U23381 (N_23381,N_23062,N_23169);
and U23382 (N_23382,N_23049,N_23106);
or U23383 (N_23383,N_23199,N_23100);
and U23384 (N_23384,N_23033,N_23008);
xnor U23385 (N_23385,N_23104,N_23019);
nor U23386 (N_23386,N_23134,N_23191);
nand U23387 (N_23387,N_23146,N_23199);
xor U23388 (N_23388,N_23111,N_23110);
and U23389 (N_23389,N_23079,N_23199);
or U23390 (N_23390,N_23146,N_23111);
or U23391 (N_23391,N_23082,N_23019);
nand U23392 (N_23392,N_23110,N_23142);
or U23393 (N_23393,N_23013,N_23191);
nor U23394 (N_23394,N_23164,N_23012);
nor U23395 (N_23395,N_23134,N_23071);
xor U23396 (N_23396,N_23198,N_23095);
nor U23397 (N_23397,N_23185,N_23018);
nand U23398 (N_23398,N_23140,N_23077);
xnor U23399 (N_23399,N_23107,N_23010);
nor U23400 (N_23400,N_23359,N_23242);
and U23401 (N_23401,N_23391,N_23286);
nand U23402 (N_23402,N_23282,N_23250);
nor U23403 (N_23403,N_23275,N_23293);
and U23404 (N_23404,N_23396,N_23279);
or U23405 (N_23405,N_23301,N_23256);
and U23406 (N_23406,N_23292,N_23270);
and U23407 (N_23407,N_23268,N_23325);
or U23408 (N_23408,N_23376,N_23343);
xnor U23409 (N_23409,N_23361,N_23351);
and U23410 (N_23410,N_23373,N_23360);
and U23411 (N_23411,N_23375,N_23260);
or U23412 (N_23412,N_23399,N_23271);
nor U23413 (N_23413,N_23228,N_23245);
nor U23414 (N_23414,N_23384,N_23357);
xnor U23415 (N_23415,N_23202,N_23305);
or U23416 (N_23416,N_23322,N_23394);
and U23417 (N_23417,N_23297,N_23265);
xnor U23418 (N_23418,N_23267,N_23206);
and U23419 (N_23419,N_23365,N_23362);
nor U23420 (N_23420,N_23230,N_23253);
nor U23421 (N_23421,N_23304,N_23319);
or U23422 (N_23422,N_23390,N_23214);
and U23423 (N_23423,N_23278,N_23353);
nor U23424 (N_23424,N_23312,N_23371);
nor U23425 (N_23425,N_23204,N_23283);
xor U23426 (N_23426,N_23231,N_23246);
nor U23427 (N_23427,N_23328,N_23382);
nand U23428 (N_23428,N_23272,N_23316);
or U23429 (N_23429,N_23273,N_23342);
or U23430 (N_23430,N_23281,N_23317);
and U23431 (N_23431,N_23233,N_23350);
or U23432 (N_23432,N_23257,N_23363);
xor U23433 (N_23433,N_23315,N_23240);
nor U23434 (N_23434,N_23220,N_23326);
or U23435 (N_23435,N_23381,N_23300);
and U23436 (N_23436,N_23338,N_23303);
xor U23437 (N_23437,N_23336,N_23333);
nor U23438 (N_23438,N_23366,N_23380);
nor U23439 (N_23439,N_23308,N_23311);
and U23440 (N_23440,N_23244,N_23236);
or U23441 (N_23441,N_23263,N_23234);
nand U23442 (N_23442,N_23252,N_23295);
nor U23443 (N_23443,N_23280,N_23367);
xnor U23444 (N_23444,N_23335,N_23290);
and U23445 (N_23445,N_23393,N_23229);
xor U23446 (N_23446,N_23217,N_23392);
nor U23447 (N_23447,N_23370,N_23212);
xor U23448 (N_23448,N_23216,N_23299);
nor U23449 (N_23449,N_23337,N_23309);
xor U23450 (N_23450,N_23235,N_23302);
nand U23451 (N_23451,N_23369,N_23332);
and U23452 (N_23452,N_23398,N_23219);
or U23453 (N_23453,N_23383,N_23203);
and U23454 (N_23454,N_23347,N_23288);
and U23455 (N_23455,N_23354,N_23324);
and U23456 (N_23456,N_23227,N_23205);
and U23457 (N_23457,N_23243,N_23339);
nand U23458 (N_23458,N_23291,N_23298);
xnor U23459 (N_23459,N_23372,N_23387);
and U23460 (N_23460,N_23284,N_23241);
nand U23461 (N_23461,N_23379,N_23331);
and U23462 (N_23462,N_23251,N_23277);
nand U23463 (N_23463,N_23222,N_23248);
nor U23464 (N_23464,N_23237,N_23346);
or U23465 (N_23465,N_23294,N_23218);
or U23466 (N_23466,N_23340,N_23395);
nand U23467 (N_23467,N_23254,N_23258);
and U23468 (N_23468,N_23223,N_23388);
nand U23469 (N_23469,N_23289,N_23262);
or U23470 (N_23470,N_23374,N_23314);
or U23471 (N_23471,N_23352,N_23356);
nand U23472 (N_23472,N_23385,N_23378);
nor U23473 (N_23473,N_23221,N_23323);
or U23474 (N_23474,N_23261,N_23349);
nand U23475 (N_23475,N_23239,N_23226);
and U23476 (N_23476,N_23318,N_23276);
xor U23477 (N_23477,N_23274,N_23264);
xor U23478 (N_23478,N_23341,N_23306);
and U23479 (N_23479,N_23210,N_23334);
nor U23480 (N_23480,N_23255,N_23329);
nand U23481 (N_23481,N_23201,N_23330);
nor U23482 (N_23482,N_23377,N_23327);
nand U23483 (N_23483,N_23320,N_23213);
and U23484 (N_23484,N_23287,N_23296);
nand U23485 (N_23485,N_23208,N_23238);
nor U23486 (N_23486,N_23200,N_23364);
nand U23487 (N_23487,N_23249,N_23345);
and U23488 (N_23488,N_23259,N_23348);
or U23489 (N_23489,N_23247,N_23344);
nor U23490 (N_23490,N_23269,N_23389);
nor U23491 (N_23491,N_23368,N_23207);
xnor U23492 (N_23492,N_23225,N_23355);
nand U23493 (N_23493,N_23358,N_23397);
xor U23494 (N_23494,N_23224,N_23285);
xnor U23495 (N_23495,N_23266,N_23215);
and U23496 (N_23496,N_23307,N_23232);
nand U23497 (N_23497,N_23211,N_23386);
nor U23498 (N_23498,N_23209,N_23313);
xor U23499 (N_23499,N_23321,N_23310);
nor U23500 (N_23500,N_23275,N_23338);
xnor U23501 (N_23501,N_23369,N_23208);
or U23502 (N_23502,N_23245,N_23279);
nand U23503 (N_23503,N_23396,N_23262);
and U23504 (N_23504,N_23211,N_23259);
nand U23505 (N_23505,N_23230,N_23305);
or U23506 (N_23506,N_23217,N_23260);
or U23507 (N_23507,N_23393,N_23345);
or U23508 (N_23508,N_23295,N_23259);
nor U23509 (N_23509,N_23353,N_23316);
nor U23510 (N_23510,N_23250,N_23286);
and U23511 (N_23511,N_23358,N_23324);
xnor U23512 (N_23512,N_23272,N_23366);
nor U23513 (N_23513,N_23216,N_23233);
nor U23514 (N_23514,N_23322,N_23269);
nand U23515 (N_23515,N_23312,N_23215);
xor U23516 (N_23516,N_23300,N_23327);
nand U23517 (N_23517,N_23298,N_23386);
xor U23518 (N_23518,N_23252,N_23348);
nand U23519 (N_23519,N_23393,N_23293);
nor U23520 (N_23520,N_23383,N_23298);
or U23521 (N_23521,N_23263,N_23303);
xnor U23522 (N_23522,N_23275,N_23369);
or U23523 (N_23523,N_23234,N_23232);
nor U23524 (N_23524,N_23242,N_23262);
and U23525 (N_23525,N_23327,N_23347);
nand U23526 (N_23526,N_23389,N_23347);
nor U23527 (N_23527,N_23342,N_23365);
or U23528 (N_23528,N_23358,N_23310);
nand U23529 (N_23529,N_23222,N_23365);
or U23530 (N_23530,N_23392,N_23283);
xor U23531 (N_23531,N_23234,N_23337);
nand U23532 (N_23532,N_23253,N_23211);
or U23533 (N_23533,N_23346,N_23399);
nand U23534 (N_23534,N_23374,N_23321);
xnor U23535 (N_23535,N_23202,N_23330);
xor U23536 (N_23536,N_23309,N_23212);
nand U23537 (N_23537,N_23347,N_23383);
and U23538 (N_23538,N_23391,N_23377);
nor U23539 (N_23539,N_23327,N_23255);
nor U23540 (N_23540,N_23313,N_23224);
and U23541 (N_23541,N_23375,N_23372);
xnor U23542 (N_23542,N_23288,N_23256);
nor U23543 (N_23543,N_23220,N_23245);
nand U23544 (N_23544,N_23275,N_23289);
nand U23545 (N_23545,N_23385,N_23379);
and U23546 (N_23546,N_23201,N_23229);
and U23547 (N_23547,N_23239,N_23222);
and U23548 (N_23548,N_23348,N_23339);
and U23549 (N_23549,N_23241,N_23291);
or U23550 (N_23550,N_23227,N_23233);
and U23551 (N_23551,N_23250,N_23245);
nor U23552 (N_23552,N_23260,N_23280);
xor U23553 (N_23553,N_23209,N_23391);
and U23554 (N_23554,N_23319,N_23345);
nor U23555 (N_23555,N_23216,N_23267);
xnor U23556 (N_23556,N_23287,N_23304);
nand U23557 (N_23557,N_23345,N_23328);
nor U23558 (N_23558,N_23338,N_23382);
or U23559 (N_23559,N_23273,N_23275);
or U23560 (N_23560,N_23345,N_23333);
xor U23561 (N_23561,N_23341,N_23217);
nor U23562 (N_23562,N_23200,N_23306);
and U23563 (N_23563,N_23308,N_23227);
xnor U23564 (N_23564,N_23318,N_23339);
nand U23565 (N_23565,N_23319,N_23305);
nand U23566 (N_23566,N_23218,N_23247);
or U23567 (N_23567,N_23340,N_23234);
or U23568 (N_23568,N_23211,N_23329);
and U23569 (N_23569,N_23249,N_23383);
nor U23570 (N_23570,N_23213,N_23201);
or U23571 (N_23571,N_23314,N_23343);
or U23572 (N_23572,N_23349,N_23365);
or U23573 (N_23573,N_23253,N_23296);
nor U23574 (N_23574,N_23348,N_23263);
xnor U23575 (N_23575,N_23312,N_23350);
nor U23576 (N_23576,N_23258,N_23263);
or U23577 (N_23577,N_23277,N_23267);
xnor U23578 (N_23578,N_23371,N_23360);
and U23579 (N_23579,N_23252,N_23372);
nand U23580 (N_23580,N_23353,N_23212);
and U23581 (N_23581,N_23294,N_23238);
or U23582 (N_23582,N_23335,N_23209);
nand U23583 (N_23583,N_23379,N_23212);
nor U23584 (N_23584,N_23234,N_23328);
and U23585 (N_23585,N_23397,N_23264);
or U23586 (N_23586,N_23217,N_23331);
and U23587 (N_23587,N_23329,N_23339);
nand U23588 (N_23588,N_23298,N_23232);
xor U23589 (N_23589,N_23322,N_23278);
nand U23590 (N_23590,N_23293,N_23239);
xnor U23591 (N_23591,N_23356,N_23376);
xor U23592 (N_23592,N_23396,N_23294);
nand U23593 (N_23593,N_23258,N_23300);
xnor U23594 (N_23594,N_23302,N_23257);
and U23595 (N_23595,N_23345,N_23254);
and U23596 (N_23596,N_23224,N_23216);
nand U23597 (N_23597,N_23379,N_23252);
and U23598 (N_23598,N_23245,N_23314);
nand U23599 (N_23599,N_23216,N_23381);
xor U23600 (N_23600,N_23466,N_23559);
xor U23601 (N_23601,N_23522,N_23549);
or U23602 (N_23602,N_23592,N_23573);
xor U23603 (N_23603,N_23595,N_23515);
or U23604 (N_23604,N_23531,N_23408);
and U23605 (N_23605,N_23550,N_23547);
or U23606 (N_23606,N_23441,N_23470);
and U23607 (N_23607,N_23539,N_23589);
and U23608 (N_23608,N_23434,N_23501);
or U23609 (N_23609,N_23579,N_23502);
and U23610 (N_23610,N_23425,N_23472);
nand U23611 (N_23611,N_23513,N_23505);
nor U23612 (N_23612,N_23536,N_23553);
nand U23613 (N_23613,N_23458,N_23524);
and U23614 (N_23614,N_23542,N_23416);
and U23615 (N_23615,N_23431,N_23599);
or U23616 (N_23616,N_23422,N_23528);
xnor U23617 (N_23617,N_23444,N_23473);
xor U23618 (N_23618,N_23421,N_23529);
xor U23619 (N_23619,N_23429,N_23534);
or U23620 (N_23620,N_23450,N_23488);
xor U23621 (N_23621,N_23455,N_23483);
xor U23622 (N_23622,N_23413,N_23499);
nor U23623 (N_23623,N_23479,N_23403);
and U23624 (N_23624,N_23525,N_23457);
xor U23625 (N_23625,N_23497,N_23538);
nor U23626 (N_23626,N_23535,N_23411);
nor U23627 (N_23627,N_23548,N_23576);
nand U23628 (N_23628,N_23404,N_23566);
nand U23629 (N_23629,N_23495,N_23467);
nor U23630 (N_23630,N_23494,N_23582);
nand U23631 (N_23631,N_23406,N_23509);
nor U23632 (N_23632,N_23516,N_23555);
xnor U23633 (N_23633,N_23591,N_23463);
xnor U23634 (N_23634,N_23527,N_23593);
nor U23635 (N_23635,N_23504,N_23514);
nand U23636 (N_23636,N_23506,N_23445);
or U23637 (N_23637,N_23478,N_23546);
or U23638 (N_23638,N_23480,N_23462);
xor U23639 (N_23639,N_23405,N_23432);
nor U23640 (N_23640,N_23552,N_23428);
and U23641 (N_23641,N_23482,N_23437);
nor U23642 (N_23642,N_23453,N_23436);
and U23643 (N_23643,N_23551,N_23448);
or U23644 (N_23644,N_23414,N_23451);
xnor U23645 (N_23645,N_23517,N_23430);
nor U23646 (N_23646,N_23400,N_23597);
nand U23647 (N_23647,N_23409,N_23433);
nand U23648 (N_23648,N_23561,N_23490);
nand U23649 (N_23649,N_23401,N_23540);
or U23650 (N_23650,N_23440,N_23521);
xnor U23651 (N_23651,N_23484,N_23447);
nand U23652 (N_23652,N_23465,N_23565);
nand U23653 (N_23653,N_23586,N_23438);
and U23654 (N_23654,N_23557,N_23503);
xor U23655 (N_23655,N_23496,N_23512);
xnor U23656 (N_23656,N_23412,N_23491);
or U23657 (N_23657,N_23489,N_23474);
or U23658 (N_23658,N_23485,N_23454);
xor U23659 (N_23659,N_23571,N_23584);
nand U23660 (N_23660,N_23459,N_23475);
nand U23661 (N_23661,N_23456,N_23569);
nor U23662 (N_23662,N_23520,N_23507);
nand U23663 (N_23663,N_23424,N_23594);
or U23664 (N_23664,N_23543,N_23446);
xor U23665 (N_23665,N_23581,N_23427);
xnor U23666 (N_23666,N_23533,N_23588);
xnor U23667 (N_23667,N_23574,N_23460);
xor U23668 (N_23668,N_23598,N_23452);
or U23669 (N_23669,N_23410,N_23402);
or U23670 (N_23670,N_23498,N_23461);
nor U23671 (N_23671,N_23541,N_23449);
and U23672 (N_23672,N_23580,N_23519);
nand U23673 (N_23673,N_23419,N_23596);
nor U23674 (N_23674,N_23492,N_23423);
and U23675 (N_23675,N_23439,N_23426);
nand U23676 (N_23676,N_23523,N_23563);
nor U23677 (N_23677,N_23558,N_23567);
and U23678 (N_23678,N_23477,N_23511);
or U23679 (N_23679,N_23476,N_23518);
nor U23680 (N_23680,N_23545,N_23487);
nor U23681 (N_23681,N_23443,N_23417);
and U23682 (N_23682,N_23570,N_23510);
nor U23683 (N_23683,N_23481,N_23407);
and U23684 (N_23684,N_23554,N_23585);
xnor U23685 (N_23685,N_23500,N_23572);
or U23686 (N_23686,N_23578,N_23556);
and U23687 (N_23687,N_23486,N_23508);
and U23688 (N_23688,N_23587,N_23526);
xor U23689 (N_23689,N_23420,N_23575);
or U23690 (N_23690,N_23415,N_23493);
nand U23691 (N_23691,N_23442,N_23532);
or U23692 (N_23692,N_23418,N_23471);
and U23693 (N_23693,N_23537,N_23468);
and U23694 (N_23694,N_23562,N_23469);
xor U23695 (N_23695,N_23583,N_23564);
or U23696 (N_23696,N_23464,N_23544);
and U23697 (N_23697,N_23577,N_23590);
nor U23698 (N_23698,N_23560,N_23435);
and U23699 (N_23699,N_23568,N_23530);
and U23700 (N_23700,N_23585,N_23545);
nor U23701 (N_23701,N_23550,N_23421);
xor U23702 (N_23702,N_23468,N_23551);
xnor U23703 (N_23703,N_23523,N_23570);
or U23704 (N_23704,N_23569,N_23447);
or U23705 (N_23705,N_23412,N_23502);
xor U23706 (N_23706,N_23555,N_23467);
or U23707 (N_23707,N_23503,N_23407);
nand U23708 (N_23708,N_23407,N_23530);
or U23709 (N_23709,N_23564,N_23518);
or U23710 (N_23710,N_23573,N_23439);
and U23711 (N_23711,N_23570,N_23509);
nor U23712 (N_23712,N_23541,N_23484);
xnor U23713 (N_23713,N_23453,N_23416);
nand U23714 (N_23714,N_23475,N_23572);
nand U23715 (N_23715,N_23579,N_23592);
and U23716 (N_23716,N_23531,N_23456);
xor U23717 (N_23717,N_23505,N_23536);
and U23718 (N_23718,N_23493,N_23514);
nand U23719 (N_23719,N_23468,N_23439);
and U23720 (N_23720,N_23513,N_23481);
xnor U23721 (N_23721,N_23544,N_23401);
nand U23722 (N_23722,N_23410,N_23479);
nor U23723 (N_23723,N_23482,N_23549);
nand U23724 (N_23724,N_23570,N_23459);
nand U23725 (N_23725,N_23546,N_23453);
xnor U23726 (N_23726,N_23443,N_23403);
nand U23727 (N_23727,N_23489,N_23558);
or U23728 (N_23728,N_23449,N_23443);
or U23729 (N_23729,N_23404,N_23463);
nor U23730 (N_23730,N_23423,N_23558);
nor U23731 (N_23731,N_23579,N_23460);
nor U23732 (N_23732,N_23405,N_23583);
and U23733 (N_23733,N_23533,N_23552);
xor U23734 (N_23734,N_23531,N_23565);
or U23735 (N_23735,N_23409,N_23450);
and U23736 (N_23736,N_23486,N_23595);
and U23737 (N_23737,N_23431,N_23477);
xnor U23738 (N_23738,N_23511,N_23588);
nand U23739 (N_23739,N_23407,N_23540);
or U23740 (N_23740,N_23437,N_23487);
and U23741 (N_23741,N_23512,N_23582);
and U23742 (N_23742,N_23401,N_23472);
and U23743 (N_23743,N_23542,N_23507);
xnor U23744 (N_23744,N_23484,N_23477);
or U23745 (N_23745,N_23419,N_23464);
or U23746 (N_23746,N_23485,N_23523);
and U23747 (N_23747,N_23572,N_23496);
xnor U23748 (N_23748,N_23473,N_23443);
or U23749 (N_23749,N_23487,N_23567);
or U23750 (N_23750,N_23510,N_23488);
and U23751 (N_23751,N_23432,N_23437);
or U23752 (N_23752,N_23561,N_23452);
xnor U23753 (N_23753,N_23588,N_23516);
and U23754 (N_23754,N_23443,N_23421);
and U23755 (N_23755,N_23544,N_23490);
nand U23756 (N_23756,N_23447,N_23479);
or U23757 (N_23757,N_23409,N_23571);
or U23758 (N_23758,N_23469,N_23550);
or U23759 (N_23759,N_23415,N_23558);
nand U23760 (N_23760,N_23408,N_23560);
nand U23761 (N_23761,N_23568,N_23523);
or U23762 (N_23762,N_23430,N_23500);
xnor U23763 (N_23763,N_23508,N_23582);
nand U23764 (N_23764,N_23590,N_23422);
nor U23765 (N_23765,N_23440,N_23525);
xnor U23766 (N_23766,N_23404,N_23416);
nand U23767 (N_23767,N_23420,N_23597);
nor U23768 (N_23768,N_23406,N_23505);
or U23769 (N_23769,N_23436,N_23439);
or U23770 (N_23770,N_23575,N_23576);
nor U23771 (N_23771,N_23421,N_23479);
xor U23772 (N_23772,N_23534,N_23489);
nand U23773 (N_23773,N_23422,N_23575);
xor U23774 (N_23774,N_23554,N_23512);
nor U23775 (N_23775,N_23479,N_23476);
nand U23776 (N_23776,N_23534,N_23542);
xor U23777 (N_23777,N_23501,N_23431);
or U23778 (N_23778,N_23580,N_23400);
or U23779 (N_23779,N_23475,N_23430);
or U23780 (N_23780,N_23438,N_23454);
and U23781 (N_23781,N_23432,N_23542);
or U23782 (N_23782,N_23566,N_23462);
nor U23783 (N_23783,N_23453,N_23427);
xnor U23784 (N_23784,N_23416,N_23418);
and U23785 (N_23785,N_23534,N_23516);
nand U23786 (N_23786,N_23502,N_23407);
xor U23787 (N_23787,N_23506,N_23534);
or U23788 (N_23788,N_23410,N_23565);
nor U23789 (N_23789,N_23485,N_23555);
and U23790 (N_23790,N_23511,N_23487);
nor U23791 (N_23791,N_23403,N_23496);
xor U23792 (N_23792,N_23562,N_23491);
or U23793 (N_23793,N_23423,N_23509);
nand U23794 (N_23794,N_23494,N_23414);
nand U23795 (N_23795,N_23585,N_23537);
and U23796 (N_23796,N_23527,N_23443);
xor U23797 (N_23797,N_23463,N_23503);
nor U23798 (N_23798,N_23566,N_23430);
nor U23799 (N_23799,N_23576,N_23413);
xnor U23800 (N_23800,N_23724,N_23758);
and U23801 (N_23801,N_23773,N_23701);
and U23802 (N_23802,N_23763,N_23780);
nor U23803 (N_23803,N_23761,N_23746);
xor U23804 (N_23804,N_23656,N_23669);
xor U23805 (N_23805,N_23700,N_23796);
or U23806 (N_23806,N_23781,N_23732);
and U23807 (N_23807,N_23650,N_23689);
nor U23808 (N_23808,N_23606,N_23742);
and U23809 (N_23809,N_23767,N_23659);
or U23810 (N_23810,N_23671,N_23768);
nand U23811 (N_23811,N_23697,N_23641);
or U23812 (N_23812,N_23640,N_23653);
xor U23813 (N_23813,N_23764,N_23645);
or U23814 (N_23814,N_23605,N_23691);
and U23815 (N_23815,N_23617,N_23782);
and U23816 (N_23816,N_23699,N_23642);
nand U23817 (N_23817,N_23733,N_23721);
or U23818 (N_23818,N_23667,N_23756);
nor U23819 (N_23819,N_23647,N_23709);
and U23820 (N_23820,N_23658,N_23603);
nand U23821 (N_23821,N_23692,N_23620);
and U23822 (N_23822,N_23661,N_23744);
and U23823 (N_23823,N_23706,N_23655);
nor U23824 (N_23824,N_23696,N_23779);
xnor U23825 (N_23825,N_23720,N_23619);
or U23826 (N_23826,N_23678,N_23601);
nor U23827 (N_23827,N_23795,N_23688);
or U23828 (N_23828,N_23797,N_23725);
nor U23829 (N_23829,N_23679,N_23654);
nand U23830 (N_23830,N_23784,N_23638);
nand U23831 (N_23831,N_23712,N_23684);
or U23832 (N_23832,N_23713,N_23668);
nor U23833 (N_23833,N_23672,N_23718);
or U23834 (N_23834,N_23786,N_23651);
or U23835 (N_23835,N_23778,N_23687);
nor U23836 (N_23836,N_23757,N_23792);
xor U23837 (N_23837,N_23707,N_23785);
nand U23838 (N_23838,N_23600,N_23755);
nand U23839 (N_23839,N_23680,N_23693);
or U23840 (N_23840,N_23739,N_23788);
xor U23841 (N_23841,N_23636,N_23698);
nand U23842 (N_23842,N_23793,N_23783);
nand U23843 (N_23843,N_23631,N_23618);
and U23844 (N_23844,N_23694,N_23625);
xnor U23845 (N_23845,N_23607,N_23611);
or U23846 (N_23846,N_23633,N_23787);
xor U23847 (N_23847,N_23754,N_23677);
and U23848 (N_23848,N_23676,N_23657);
and U23849 (N_23849,N_23740,N_23634);
nor U23850 (N_23850,N_23751,N_23644);
nor U23851 (N_23851,N_23705,N_23753);
nand U23852 (N_23852,N_23708,N_23730);
nand U23853 (N_23853,N_23735,N_23776);
nor U23854 (N_23854,N_23772,N_23704);
nand U23855 (N_23855,N_23789,N_23799);
or U23856 (N_23856,N_23609,N_23649);
xor U23857 (N_23857,N_23723,N_23662);
and U23858 (N_23858,N_23711,N_23775);
or U23859 (N_23859,N_23760,N_23612);
and U23860 (N_23860,N_23726,N_23748);
nor U23861 (N_23861,N_23635,N_23727);
nor U23862 (N_23862,N_23627,N_23621);
and U23863 (N_23863,N_23769,N_23614);
and U23864 (N_23864,N_23664,N_23695);
and U23865 (N_23865,N_23719,N_23683);
nor U23866 (N_23866,N_23728,N_23717);
xnor U23867 (N_23867,N_23613,N_23710);
xor U23868 (N_23868,N_23674,N_23798);
and U23869 (N_23869,N_23629,N_23745);
nand U23870 (N_23870,N_23630,N_23731);
or U23871 (N_23871,N_23670,N_23703);
xnor U23872 (N_23872,N_23643,N_23616);
nand U23873 (N_23873,N_23759,N_23652);
nand U23874 (N_23874,N_23646,N_23666);
nand U23875 (N_23875,N_23622,N_23663);
xor U23876 (N_23876,N_23660,N_23615);
nand U23877 (N_23877,N_23682,N_23604);
or U23878 (N_23878,N_23637,N_23624);
or U23879 (N_23879,N_23743,N_23602);
nand U23880 (N_23880,N_23749,N_23648);
xnor U23881 (N_23881,N_23716,N_23722);
or U23882 (N_23882,N_23752,N_23771);
xnor U23883 (N_23883,N_23690,N_23777);
xor U23884 (N_23884,N_23794,N_23736);
and U23885 (N_23885,N_23610,N_23608);
xnor U23886 (N_23886,N_23762,N_23702);
nand U23887 (N_23887,N_23626,N_23774);
nand U23888 (N_23888,N_23734,N_23685);
nor U23889 (N_23889,N_23665,N_23686);
xnor U23890 (N_23890,N_23623,N_23715);
xnor U23891 (N_23891,N_23738,N_23765);
or U23892 (N_23892,N_23628,N_23729);
nor U23893 (N_23893,N_23632,N_23747);
nor U23894 (N_23894,N_23791,N_23639);
and U23895 (N_23895,N_23675,N_23681);
nand U23896 (N_23896,N_23766,N_23770);
nor U23897 (N_23897,N_23714,N_23673);
xnor U23898 (N_23898,N_23750,N_23790);
nor U23899 (N_23899,N_23737,N_23741);
nor U23900 (N_23900,N_23645,N_23696);
and U23901 (N_23901,N_23796,N_23638);
nor U23902 (N_23902,N_23650,N_23663);
and U23903 (N_23903,N_23723,N_23632);
nand U23904 (N_23904,N_23752,N_23782);
or U23905 (N_23905,N_23616,N_23654);
nor U23906 (N_23906,N_23609,N_23630);
and U23907 (N_23907,N_23797,N_23784);
and U23908 (N_23908,N_23735,N_23662);
nor U23909 (N_23909,N_23786,N_23635);
xor U23910 (N_23910,N_23716,N_23611);
or U23911 (N_23911,N_23645,N_23745);
or U23912 (N_23912,N_23780,N_23791);
nor U23913 (N_23913,N_23731,N_23658);
xnor U23914 (N_23914,N_23693,N_23786);
nor U23915 (N_23915,N_23666,N_23644);
and U23916 (N_23916,N_23702,N_23740);
nand U23917 (N_23917,N_23678,N_23711);
and U23918 (N_23918,N_23607,N_23723);
nand U23919 (N_23919,N_23737,N_23727);
or U23920 (N_23920,N_23657,N_23778);
and U23921 (N_23921,N_23681,N_23621);
nor U23922 (N_23922,N_23699,N_23698);
and U23923 (N_23923,N_23670,N_23702);
xnor U23924 (N_23924,N_23601,N_23648);
or U23925 (N_23925,N_23704,N_23612);
nor U23926 (N_23926,N_23796,N_23791);
nand U23927 (N_23927,N_23665,N_23729);
xor U23928 (N_23928,N_23689,N_23684);
and U23929 (N_23929,N_23767,N_23657);
or U23930 (N_23930,N_23695,N_23625);
or U23931 (N_23931,N_23601,N_23609);
xnor U23932 (N_23932,N_23685,N_23699);
nand U23933 (N_23933,N_23750,N_23625);
nand U23934 (N_23934,N_23794,N_23615);
and U23935 (N_23935,N_23722,N_23682);
or U23936 (N_23936,N_23640,N_23654);
and U23937 (N_23937,N_23687,N_23641);
or U23938 (N_23938,N_23733,N_23620);
nor U23939 (N_23939,N_23766,N_23650);
xnor U23940 (N_23940,N_23760,N_23775);
xnor U23941 (N_23941,N_23622,N_23686);
nor U23942 (N_23942,N_23763,N_23648);
or U23943 (N_23943,N_23622,N_23643);
nand U23944 (N_23944,N_23720,N_23763);
and U23945 (N_23945,N_23726,N_23781);
or U23946 (N_23946,N_23799,N_23723);
nor U23947 (N_23947,N_23786,N_23722);
xor U23948 (N_23948,N_23647,N_23737);
or U23949 (N_23949,N_23610,N_23647);
and U23950 (N_23950,N_23688,N_23755);
and U23951 (N_23951,N_23793,N_23673);
nor U23952 (N_23952,N_23759,N_23795);
nor U23953 (N_23953,N_23663,N_23641);
and U23954 (N_23954,N_23669,N_23602);
nand U23955 (N_23955,N_23638,N_23762);
nand U23956 (N_23956,N_23699,N_23682);
or U23957 (N_23957,N_23650,N_23658);
xnor U23958 (N_23958,N_23783,N_23753);
nor U23959 (N_23959,N_23784,N_23717);
or U23960 (N_23960,N_23750,N_23609);
nor U23961 (N_23961,N_23656,N_23759);
nand U23962 (N_23962,N_23761,N_23783);
nor U23963 (N_23963,N_23782,N_23625);
and U23964 (N_23964,N_23652,N_23657);
nand U23965 (N_23965,N_23724,N_23765);
xor U23966 (N_23966,N_23638,N_23785);
or U23967 (N_23967,N_23611,N_23712);
or U23968 (N_23968,N_23689,N_23696);
xnor U23969 (N_23969,N_23648,N_23709);
nand U23970 (N_23970,N_23631,N_23606);
nand U23971 (N_23971,N_23648,N_23652);
or U23972 (N_23972,N_23768,N_23616);
nor U23973 (N_23973,N_23632,N_23709);
xnor U23974 (N_23974,N_23647,N_23700);
xor U23975 (N_23975,N_23722,N_23638);
nor U23976 (N_23976,N_23633,N_23655);
nand U23977 (N_23977,N_23724,N_23757);
nor U23978 (N_23978,N_23605,N_23643);
nor U23979 (N_23979,N_23630,N_23685);
nor U23980 (N_23980,N_23793,N_23688);
or U23981 (N_23981,N_23785,N_23773);
and U23982 (N_23982,N_23627,N_23648);
xnor U23983 (N_23983,N_23703,N_23626);
nand U23984 (N_23984,N_23646,N_23699);
xor U23985 (N_23985,N_23657,N_23600);
and U23986 (N_23986,N_23668,N_23707);
nor U23987 (N_23987,N_23736,N_23610);
and U23988 (N_23988,N_23732,N_23762);
or U23989 (N_23989,N_23630,N_23755);
xor U23990 (N_23990,N_23760,N_23742);
and U23991 (N_23991,N_23618,N_23626);
and U23992 (N_23992,N_23603,N_23613);
nand U23993 (N_23993,N_23789,N_23656);
nor U23994 (N_23994,N_23745,N_23703);
xor U23995 (N_23995,N_23604,N_23624);
or U23996 (N_23996,N_23740,N_23707);
xor U23997 (N_23997,N_23757,N_23745);
and U23998 (N_23998,N_23637,N_23744);
and U23999 (N_23999,N_23799,N_23660);
xor U24000 (N_24000,N_23941,N_23993);
nor U24001 (N_24001,N_23892,N_23837);
xor U24002 (N_24002,N_23970,N_23909);
nand U24003 (N_24003,N_23836,N_23829);
or U24004 (N_24004,N_23895,N_23844);
nor U24005 (N_24005,N_23897,N_23808);
xnor U24006 (N_24006,N_23992,N_23854);
nor U24007 (N_24007,N_23918,N_23804);
and U24008 (N_24008,N_23974,N_23818);
or U24009 (N_24009,N_23870,N_23891);
nand U24010 (N_24010,N_23972,N_23811);
or U24011 (N_24011,N_23874,N_23817);
nand U24012 (N_24012,N_23981,N_23957);
or U24013 (N_24013,N_23894,N_23979);
nor U24014 (N_24014,N_23871,N_23821);
or U24015 (N_24015,N_23819,N_23907);
xnor U24016 (N_24016,N_23991,N_23872);
and U24017 (N_24017,N_23868,N_23947);
nor U24018 (N_24018,N_23880,N_23826);
and U24019 (N_24019,N_23916,N_23859);
or U24020 (N_24020,N_23848,N_23980);
nand U24021 (N_24021,N_23852,N_23824);
nand U24022 (N_24022,N_23961,N_23948);
nor U24023 (N_24023,N_23904,N_23830);
and U24024 (N_24024,N_23926,N_23955);
or U24025 (N_24025,N_23885,N_23806);
and U24026 (N_24026,N_23813,N_23967);
nand U24027 (N_24027,N_23828,N_23949);
xor U24028 (N_24028,N_23915,N_23919);
and U24029 (N_24029,N_23896,N_23944);
nor U24030 (N_24030,N_23985,N_23914);
nand U24031 (N_24031,N_23984,N_23803);
or U24032 (N_24032,N_23936,N_23827);
nand U24033 (N_24033,N_23958,N_23878);
nor U24034 (N_24034,N_23853,N_23900);
nor U24035 (N_24035,N_23997,N_23903);
or U24036 (N_24036,N_23969,N_23884);
nand U24037 (N_24037,N_23950,N_23986);
xnor U24038 (N_24038,N_23939,N_23906);
and U24039 (N_24039,N_23883,N_23932);
or U24040 (N_24040,N_23959,N_23876);
xnor U24041 (N_24041,N_23809,N_23893);
or U24042 (N_24042,N_23954,N_23801);
and U24043 (N_24043,N_23987,N_23898);
nor U24044 (N_24044,N_23822,N_23882);
or U24045 (N_24045,N_23945,N_23825);
or U24046 (N_24046,N_23942,N_23847);
nor U24047 (N_24047,N_23940,N_23911);
or U24048 (N_24048,N_23865,N_23839);
nor U24049 (N_24049,N_23965,N_23927);
xnor U24050 (N_24050,N_23857,N_23976);
or U24051 (N_24051,N_23973,N_23858);
nor U24052 (N_24052,N_23856,N_23938);
nand U24053 (N_24053,N_23962,N_23937);
xor U24054 (N_24054,N_23953,N_23866);
and U24055 (N_24055,N_23995,N_23802);
or U24056 (N_24056,N_23823,N_23929);
nand U24057 (N_24057,N_23816,N_23846);
nor U24058 (N_24058,N_23861,N_23901);
or U24059 (N_24059,N_23989,N_23815);
xnor U24060 (N_24060,N_23849,N_23908);
xor U24061 (N_24061,N_23998,N_23964);
nor U24062 (N_24062,N_23943,N_23913);
and U24063 (N_24063,N_23843,N_23982);
and U24064 (N_24064,N_23842,N_23931);
nand U24065 (N_24065,N_23851,N_23833);
and U24066 (N_24066,N_23838,N_23978);
and U24067 (N_24067,N_23820,N_23888);
nand U24068 (N_24068,N_23923,N_23924);
nand U24069 (N_24069,N_23890,N_23887);
nor U24070 (N_24070,N_23905,N_23863);
nand U24071 (N_24071,N_23867,N_23886);
nand U24072 (N_24072,N_23850,N_23988);
nand U24073 (N_24073,N_23934,N_23832);
and U24074 (N_24074,N_23855,N_23935);
or U24075 (N_24075,N_23917,N_23831);
or U24076 (N_24076,N_23860,N_23800);
nand U24077 (N_24077,N_23971,N_23946);
xnor U24078 (N_24078,N_23902,N_23994);
nand U24079 (N_24079,N_23841,N_23960);
xor U24080 (N_24080,N_23810,N_23862);
nor U24081 (N_24081,N_23968,N_23990);
nor U24082 (N_24082,N_23952,N_23996);
nand U24083 (N_24083,N_23899,N_23873);
xor U24084 (N_24084,N_23966,N_23933);
nand U24085 (N_24085,N_23812,N_23875);
xor U24086 (N_24086,N_23889,N_23928);
or U24087 (N_24087,N_23845,N_23956);
and U24088 (N_24088,N_23910,N_23951);
or U24089 (N_24089,N_23877,N_23881);
or U24090 (N_24090,N_23834,N_23805);
xor U24091 (N_24091,N_23835,N_23977);
nor U24092 (N_24092,N_23879,N_23930);
nand U24093 (N_24093,N_23864,N_23807);
and U24094 (N_24094,N_23814,N_23912);
and U24095 (N_24095,N_23975,N_23963);
or U24096 (N_24096,N_23921,N_23925);
xor U24097 (N_24097,N_23920,N_23983);
xnor U24098 (N_24098,N_23922,N_23999);
nand U24099 (N_24099,N_23840,N_23869);
xor U24100 (N_24100,N_23809,N_23917);
xnor U24101 (N_24101,N_23849,N_23942);
and U24102 (N_24102,N_23867,N_23940);
nor U24103 (N_24103,N_23890,N_23929);
xor U24104 (N_24104,N_23862,N_23819);
xnor U24105 (N_24105,N_23861,N_23909);
nand U24106 (N_24106,N_23948,N_23890);
nor U24107 (N_24107,N_23862,N_23976);
xnor U24108 (N_24108,N_23915,N_23861);
and U24109 (N_24109,N_23825,N_23858);
nor U24110 (N_24110,N_23826,N_23901);
nor U24111 (N_24111,N_23985,N_23956);
or U24112 (N_24112,N_23811,N_23913);
xnor U24113 (N_24113,N_23930,N_23946);
nor U24114 (N_24114,N_23916,N_23918);
nor U24115 (N_24115,N_23892,N_23895);
or U24116 (N_24116,N_23882,N_23814);
or U24117 (N_24117,N_23990,N_23849);
nand U24118 (N_24118,N_23829,N_23996);
nand U24119 (N_24119,N_23973,N_23869);
xnor U24120 (N_24120,N_23839,N_23996);
or U24121 (N_24121,N_23965,N_23883);
nor U24122 (N_24122,N_23942,N_23854);
and U24123 (N_24123,N_23831,N_23863);
or U24124 (N_24124,N_23829,N_23854);
or U24125 (N_24125,N_23883,N_23917);
xnor U24126 (N_24126,N_23857,N_23822);
xnor U24127 (N_24127,N_23833,N_23814);
xnor U24128 (N_24128,N_23808,N_23902);
or U24129 (N_24129,N_23933,N_23863);
nor U24130 (N_24130,N_23874,N_23809);
nor U24131 (N_24131,N_23965,N_23945);
nand U24132 (N_24132,N_23808,N_23909);
xor U24133 (N_24133,N_23969,N_23881);
or U24134 (N_24134,N_23811,N_23870);
and U24135 (N_24135,N_23933,N_23819);
and U24136 (N_24136,N_23952,N_23880);
or U24137 (N_24137,N_23883,N_23890);
nor U24138 (N_24138,N_23908,N_23906);
or U24139 (N_24139,N_23813,N_23831);
xor U24140 (N_24140,N_23810,N_23832);
and U24141 (N_24141,N_23815,N_23833);
nor U24142 (N_24142,N_23969,N_23883);
and U24143 (N_24143,N_23925,N_23918);
nand U24144 (N_24144,N_23966,N_23821);
and U24145 (N_24145,N_23994,N_23855);
nand U24146 (N_24146,N_23807,N_23939);
nand U24147 (N_24147,N_23923,N_23959);
xnor U24148 (N_24148,N_23801,N_23979);
xor U24149 (N_24149,N_23923,N_23870);
xor U24150 (N_24150,N_23810,N_23942);
or U24151 (N_24151,N_23934,N_23865);
nor U24152 (N_24152,N_23994,N_23896);
or U24153 (N_24153,N_23857,N_23845);
nand U24154 (N_24154,N_23815,N_23976);
or U24155 (N_24155,N_23991,N_23974);
nor U24156 (N_24156,N_23946,N_23947);
and U24157 (N_24157,N_23844,N_23827);
nor U24158 (N_24158,N_23969,N_23830);
xnor U24159 (N_24159,N_23886,N_23936);
xor U24160 (N_24160,N_23876,N_23996);
or U24161 (N_24161,N_23930,N_23884);
xor U24162 (N_24162,N_23963,N_23840);
xor U24163 (N_24163,N_23973,N_23890);
nor U24164 (N_24164,N_23963,N_23842);
or U24165 (N_24165,N_23896,N_23986);
nand U24166 (N_24166,N_23994,N_23845);
xnor U24167 (N_24167,N_23852,N_23814);
and U24168 (N_24168,N_23911,N_23839);
or U24169 (N_24169,N_23822,N_23993);
nor U24170 (N_24170,N_23885,N_23904);
or U24171 (N_24171,N_23928,N_23837);
nor U24172 (N_24172,N_23918,N_23885);
xor U24173 (N_24173,N_23837,N_23920);
nand U24174 (N_24174,N_23931,N_23999);
nor U24175 (N_24175,N_23906,N_23936);
nor U24176 (N_24176,N_23946,N_23852);
xor U24177 (N_24177,N_23868,N_23931);
xor U24178 (N_24178,N_23853,N_23877);
xor U24179 (N_24179,N_23808,N_23945);
or U24180 (N_24180,N_23946,N_23863);
xor U24181 (N_24181,N_23823,N_23992);
and U24182 (N_24182,N_23961,N_23859);
or U24183 (N_24183,N_23920,N_23958);
xnor U24184 (N_24184,N_23828,N_23929);
nand U24185 (N_24185,N_23858,N_23917);
xnor U24186 (N_24186,N_23853,N_23983);
nand U24187 (N_24187,N_23863,N_23917);
and U24188 (N_24188,N_23999,N_23840);
or U24189 (N_24189,N_23971,N_23855);
and U24190 (N_24190,N_23824,N_23925);
nand U24191 (N_24191,N_23901,N_23809);
and U24192 (N_24192,N_23991,N_23997);
xnor U24193 (N_24193,N_23916,N_23942);
or U24194 (N_24194,N_23847,N_23866);
and U24195 (N_24195,N_23951,N_23918);
nor U24196 (N_24196,N_23982,N_23986);
and U24197 (N_24197,N_23967,N_23832);
nand U24198 (N_24198,N_23908,N_23937);
or U24199 (N_24199,N_23979,N_23950);
xnor U24200 (N_24200,N_24084,N_24174);
xnor U24201 (N_24201,N_24081,N_24004);
and U24202 (N_24202,N_24070,N_24112);
nor U24203 (N_24203,N_24137,N_24005);
nor U24204 (N_24204,N_24063,N_24140);
xnor U24205 (N_24205,N_24092,N_24051);
nand U24206 (N_24206,N_24022,N_24017);
and U24207 (N_24207,N_24189,N_24043);
xnor U24208 (N_24208,N_24050,N_24044);
nor U24209 (N_24209,N_24149,N_24127);
xor U24210 (N_24210,N_24024,N_24011);
nor U24211 (N_24211,N_24030,N_24179);
or U24212 (N_24212,N_24150,N_24012);
nor U24213 (N_24213,N_24072,N_24001);
nor U24214 (N_24214,N_24083,N_24034);
xnor U24215 (N_24215,N_24154,N_24058);
or U24216 (N_24216,N_24136,N_24059);
and U24217 (N_24217,N_24052,N_24124);
and U24218 (N_24218,N_24060,N_24000);
or U24219 (N_24219,N_24135,N_24057);
nor U24220 (N_24220,N_24039,N_24199);
nor U24221 (N_24221,N_24141,N_24076);
nor U24222 (N_24222,N_24156,N_24187);
nor U24223 (N_24223,N_24089,N_24148);
nor U24224 (N_24224,N_24131,N_24080);
nor U24225 (N_24225,N_24153,N_24097);
or U24226 (N_24226,N_24191,N_24013);
and U24227 (N_24227,N_24099,N_24133);
xnor U24228 (N_24228,N_24096,N_24082);
xor U24229 (N_24229,N_24014,N_24079);
xnor U24230 (N_24230,N_24125,N_24122);
nand U24231 (N_24231,N_24177,N_24031);
and U24232 (N_24232,N_24173,N_24067);
xor U24233 (N_24233,N_24075,N_24061);
xor U24234 (N_24234,N_24164,N_24002);
xnor U24235 (N_24235,N_24123,N_24049);
nor U24236 (N_24236,N_24016,N_24100);
and U24237 (N_24237,N_24032,N_24129);
nor U24238 (N_24238,N_24180,N_24026);
nand U24239 (N_24239,N_24066,N_24168);
and U24240 (N_24240,N_24071,N_24006);
xor U24241 (N_24241,N_24197,N_24144);
xor U24242 (N_24242,N_24166,N_24165);
nor U24243 (N_24243,N_24036,N_24118);
nand U24244 (N_24244,N_24183,N_24160);
nand U24245 (N_24245,N_24078,N_24065);
and U24246 (N_24246,N_24119,N_24158);
nor U24247 (N_24247,N_24198,N_24151);
xor U24248 (N_24248,N_24105,N_24155);
nand U24249 (N_24249,N_24116,N_24181);
xor U24250 (N_24250,N_24117,N_24064);
and U24251 (N_24251,N_24020,N_24093);
xor U24252 (N_24252,N_24161,N_24028);
xor U24253 (N_24253,N_24040,N_24037);
nor U24254 (N_24254,N_24101,N_24106);
and U24255 (N_24255,N_24132,N_24015);
nor U24256 (N_24256,N_24169,N_24053);
nor U24257 (N_24257,N_24029,N_24171);
nor U24258 (N_24258,N_24062,N_24188);
xnor U24259 (N_24259,N_24054,N_24033);
nand U24260 (N_24260,N_24073,N_24107);
nand U24261 (N_24261,N_24069,N_24134);
xnor U24262 (N_24262,N_24115,N_24055);
or U24263 (N_24263,N_24120,N_24194);
or U24264 (N_24264,N_24159,N_24121);
nor U24265 (N_24265,N_24139,N_24027);
nand U24266 (N_24266,N_24138,N_24186);
nand U24267 (N_24267,N_24196,N_24172);
xnor U24268 (N_24268,N_24085,N_24023);
nor U24269 (N_24269,N_24042,N_24007);
xor U24270 (N_24270,N_24077,N_24088);
nand U24271 (N_24271,N_24047,N_24086);
nor U24272 (N_24272,N_24103,N_24095);
nor U24273 (N_24273,N_24091,N_24175);
and U24274 (N_24274,N_24048,N_24162);
or U24275 (N_24275,N_24157,N_24046);
nor U24276 (N_24276,N_24182,N_24094);
and U24277 (N_24277,N_24190,N_24192);
nand U24278 (N_24278,N_24074,N_24090);
nor U24279 (N_24279,N_24143,N_24111);
nor U24280 (N_24280,N_24145,N_24184);
nor U24281 (N_24281,N_24018,N_24068);
nor U24282 (N_24282,N_24009,N_24113);
or U24283 (N_24283,N_24041,N_24008);
and U24284 (N_24284,N_24170,N_24021);
and U24285 (N_24285,N_24146,N_24163);
nor U24286 (N_24286,N_24010,N_24176);
or U24287 (N_24287,N_24025,N_24108);
and U24288 (N_24288,N_24126,N_24114);
xor U24289 (N_24289,N_24130,N_24142);
and U24290 (N_24290,N_24110,N_24195);
or U24291 (N_24291,N_24019,N_24128);
nor U24292 (N_24292,N_24152,N_24167);
or U24293 (N_24293,N_24102,N_24147);
and U24294 (N_24294,N_24087,N_24193);
nor U24295 (N_24295,N_24098,N_24109);
and U24296 (N_24296,N_24056,N_24035);
or U24297 (N_24297,N_24178,N_24003);
or U24298 (N_24298,N_24185,N_24038);
xnor U24299 (N_24299,N_24104,N_24045);
nor U24300 (N_24300,N_24107,N_24097);
nand U24301 (N_24301,N_24111,N_24014);
nor U24302 (N_24302,N_24048,N_24190);
and U24303 (N_24303,N_24146,N_24119);
nand U24304 (N_24304,N_24062,N_24117);
and U24305 (N_24305,N_24110,N_24038);
xor U24306 (N_24306,N_24095,N_24074);
nand U24307 (N_24307,N_24107,N_24085);
xnor U24308 (N_24308,N_24099,N_24141);
nor U24309 (N_24309,N_24012,N_24044);
or U24310 (N_24310,N_24024,N_24081);
or U24311 (N_24311,N_24185,N_24094);
or U24312 (N_24312,N_24100,N_24138);
nor U24313 (N_24313,N_24163,N_24071);
xor U24314 (N_24314,N_24045,N_24037);
or U24315 (N_24315,N_24033,N_24031);
nor U24316 (N_24316,N_24128,N_24176);
nand U24317 (N_24317,N_24139,N_24029);
and U24318 (N_24318,N_24106,N_24116);
nor U24319 (N_24319,N_24019,N_24094);
nand U24320 (N_24320,N_24128,N_24056);
nand U24321 (N_24321,N_24089,N_24002);
nand U24322 (N_24322,N_24064,N_24078);
or U24323 (N_24323,N_24071,N_24090);
xor U24324 (N_24324,N_24019,N_24194);
and U24325 (N_24325,N_24071,N_24182);
nor U24326 (N_24326,N_24109,N_24186);
nor U24327 (N_24327,N_24128,N_24107);
nor U24328 (N_24328,N_24113,N_24144);
and U24329 (N_24329,N_24048,N_24050);
nor U24330 (N_24330,N_24058,N_24110);
or U24331 (N_24331,N_24145,N_24199);
nand U24332 (N_24332,N_24094,N_24159);
nand U24333 (N_24333,N_24068,N_24072);
xnor U24334 (N_24334,N_24198,N_24073);
nand U24335 (N_24335,N_24131,N_24123);
and U24336 (N_24336,N_24188,N_24190);
nor U24337 (N_24337,N_24027,N_24018);
xor U24338 (N_24338,N_24180,N_24194);
or U24339 (N_24339,N_24038,N_24190);
nand U24340 (N_24340,N_24021,N_24116);
and U24341 (N_24341,N_24108,N_24039);
nor U24342 (N_24342,N_24011,N_24173);
nand U24343 (N_24343,N_24145,N_24071);
and U24344 (N_24344,N_24035,N_24129);
nor U24345 (N_24345,N_24196,N_24128);
and U24346 (N_24346,N_24176,N_24184);
nor U24347 (N_24347,N_24168,N_24051);
xor U24348 (N_24348,N_24124,N_24158);
and U24349 (N_24349,N_24132,N_24089);
nor U24350 (N_24350,N_24006,N_24138);
and U24351 (N_24351,N_24070,N_24113);
nor U24352 (N_24352,N_24174,N_24167);
nand U24353 (N_24353,N_24072,N_24134);
and U24354 (N_24354,N_24098,N_24177);
nand U24355 (N_24355,N_24136,N_24033);
or U24356 (N_24356,N_24008,N_24104);
or U24357 (N_24357,N_24076,N_24179);
nor U24358 (N_24358,N_24172,N_24067);
nand U24359 (N_24359,N_24065,N_24175);
xor U24360 (N_24360,N_24156,N_24030);
nand U24361 (N_24361,N_24060,N_24007);
or U24362 (N_24362,N_24055,N_24011);
or U24363 (N_24363,N_24018,N_24011);
nand U24364 (N_24364,N_24192,N_24042);
or U24365 (N_24365,N_24111,N_24049);
and U24366 (N_24366,N_24186,N_24018);
nand U24367 (N_24367,N_24077,N_24185);
nand U24368 (N_24368,N_24136,N_24077);
nand U24369 (N_24369,N_24186,N_24058);
and U24370 (N_24370,N_24118,N_24196);
and U24371 (N_24371,N_24182,N_24118);
nor U24372 (N_24372,N_24147,N_24043);
and U24373 (N_24373,N_24005,N_24180);
and U24374 (N_24374,N_24066,N_24110);
and U24375 (N_24375,N_24019,N_24048);
or U24376 (N_24376,N_24140,N_24146);
or U24377 (N_24377,N_24199,N_24105);
nor U24378 (N_24378,N_24083,N_24194);
or U24379 (N_24379,N_24103,N_24099);
and U24380 (N_24380,N_24101,N_24186);
and U24381 (N_24381,N_24180,N_24000);
or U24382 (N_24382,N_24027,N_24056);
nand U24383 (N_24383,N_24014,N_24054);
nor U24384 (N_24384,N_24036,N_24046);
or U24385 (N_24385,N_24176,N_24145);
and U24386 (N_24386,N_24130,N_24065);
nor U24387 (N_24387,N_24041,N_24037);
or U24388 (N_24388,N_24176,N_24144);
or U24389 (N_24389,N_24126,N_24025);
xnor U24390 (N_24390,N_24001,N_24146);
or U24391 (N_24391,N_24023,N_24140);
nand U24392 (N_24392,N_24022,N_24106);
nand U24393 (N_24393,N_24194,N_24163);
or U24394 (N_24394,N_24004,N_24150);
nor U24395 (N_24395,N_24054,N_24083);
or U24396 (N_24396,N_24148,N_24080);
nand U24397 (N_24397,N_24110,N_24064);
nor U24398 (N_24398,N_24153,N_24016);
and U24399 (N_24399,N_24190,N_24005);
xnor U24400 (N_24400,N_24271,N_24351);
nor U24401 (N_24401,N_24326,N_24329);
xnor U24402 (N_24402,N_24284,N_24259);
or U24403 (N_24403,N_24219,N_24260);
nor U24404 (N_24404,N_24321,N_24339);
nor U24405 (N_24405,N_24308,N_24281);
and U24406 (N_24406,N_24222,N_24305);
or U24407 (N_24407,N_24244,N_24338);
nand U24408 (N_24408,N_24393,N_24320);
nor U24409 (N_24409,N_24379,N_24212);
xor U24410 (N_24410,N_24235,N_24388);
and U24411 (N_24411,N_24263,N_24210);
xor U24412 (N_24412,N_24395,N_24389);
nor U24413 (N_24413,N_24289,N_24291);
nor U24414 (N_24414,N_24360,N_24256);
nand U24415 (N_24415,N_24361,N_24334);
nand U24416 (N_24416,N_24253,N_24322);
nand U24417 (N_24417,N_24343,N_24348);
nor U24418 (N_24418,N_24382,N_24228);
nand U24419 (N_24419,N_24397,N_24297);
or U24420 (N_24420,N_24215,N_24302);
or U24421 (N_24421,N_24243,N_24312);
nand U24422 (N_24422,N_24333,N_24349);
nor U24423 (N_24423,N_24276,N_24331);
nor U24424 (N_24424,N_24304,N_24300);
nor U24425 (N_24425,N_24265,N_24267);
nand U24426 (N_24426,N_24399,N_24218);
and U24427 (N_24427,N_24209,N_24207);
and U24428 (N_24428,N_24232,N_24238);
nor U24429 (N_24429,N_24272,N_24341);
or U24430 (N_24430,N_24396,N_24342);
and U24431 (N_24431,N_24234,N_24377);
and U24432 (N_24432,N_24248,N_24231);
nor U24433 (N_24433,N_24319,N_24298);
and U24434 (N_24434,N_24293,N_24290);
nor U24435 (N_24435,N_24310,N_24373);
nor U24436 (N_24436,N_24328,N_24296);
xor U24437 (N_24437,N_24223,N_24340);
and U24438 (N_24438,N_24239,N_24372);
nor U24439 (N_24439,N_24346,N_24200);
or U24440 (N_24440,N_24229,N_24285);
nor U24441 (N_24441,N_24268,N_24345);
nor U24442 (N_24442,N_24287,N_24230);
nand U24443 (N_24443,N_24286,N_24390);
and U24444 (N_24444,N_24315,N_24227);
nand U24445 (N_24445,N_24236,N_24357);
nand U24446 (N_24446,N_24262,N_24362);
nand U24447 (N_24447,N_24208,N_24366);
nor U24448 (N_24448,N_24278,N_24233);
xnor U24449 (N_24449,N_24280,N_24358);
nor U24450 (N_24450,N_24213,N_24269);
and U24451 (N_24451,N_24385,N_24214);
and U24452 (N_24452,N_24299,N_24306);
and U24453 (N_24453,N_24275,N_24337);
nand U24454 (N_24454,N_24283,N_24344);
and U24455 (N_24455,N_24317,N_24225);
or U24456 (N_24456,N_24277,N_24381);
and U24457 (N_24457,N_24250,N_24355);
nor U24458 (N_24458,N_24318,N_24398);
nor U24459 (N_24459,N_24336,N_24217);
nand U24460 (N_24460,N_24350,N_24258);
xnor U24461 (N_24461,N_24363,N_24384);
nand U24462 (N_24462,N_24356,N_24303);
nand U24463 (N_24463,N_24245,N_24392);
and U24464 (N_24464,N_24380,N_24279);
nor U24465 (N_24465,N_24220,N_24216);
and U24466 (N_24466,N_24224,N_24365);
and U24467 (N_24467,N_24391,N_24257);
nor U24468 (N_24468,N_24364,N_24307);
and U24469 (N_24469,N_24252,N_24387);
or U24470 (N_24470,N_24367,N_24242);
nor U24471 (N_24471,N_24274,N_24335);
nor U24472 (N_24472,N_24203,N_24394);
nand U24473 (N_24473,N_24347,N_24266);
nand U24474 (N_24474,N_24288,N_24264);
nand U24475 (N_24475,N_24255,N_24202);
nand U24476 (N_24476,N_24226,N_24301);
xnor U24477 (N_24477,N_24327,N_24251);
or U24478 (N_24478,N_24352,N_24374);
nor U24479 (N_24479,N_24370,N_24292);
or U24480 (N_24480,N_24237,N_24311);
nand U24481 (N_24481,N_24254,N_24383);
nor U24482 (N_24482,N_24201,N_24294);
or U24483 (N_24483,N_24309,N_24324);
nor U24484 (N_24484,N_24204,N_24295);
nand U24485 (N_24485,N_24247,N_24221);
or U24486 (N_24486,N_24206,N_24325);
nor U24487 (N_24487,N_24316,N_24282);
or U24488 (N_24488,N_24241,N_24270);
and U24489 (N_24489,N_24368,N_24246);
and U24490 (N_24490,N_24261,N_24205);
or U24491 (N_24491,N_24376,N_24240);
and U24492 (N_24492,N_24371,N_24359);
or U24493 (N_24493,N_24353,N_24314);
nand U24494 (N_24494,N_24332,N_24211);
or U24495 (N_24495,N_24273,N_24386);
nor U24496 (N_24496,N_24330,N_24378);
or U24497 (N_24497,N_24375,N_24369);
nand U24498 (N_24498,N_24354,N_24313);
and U24499 (N_24499,N_24249,N_24323);
nor U24500 (N_24500,N_24311,N_24280);
or U24501 (N_24501,N_24360,N_24205);
xnor U24502 (N_24502,N_24265,N_24347);
or U24503 (N_24503,N_24356,N_24241);
and U24504 (N_24504,N_24364,N_24313);
xor U24505 (N_24505,N_24302,N_24256);
or U24506 (N_24506,N_24293,N_24204);
and U24507 (N_24507,N_24235,N_24383);
or U24508 (N_24508,N_24238,N_24369);
and U24509 (N_24509,N_24359,N_24252);
nand U24510 (N_24510,N_24297,N_24351);
and U24511 (N_24511,N_24240,N_24293);
xor U24512 (N_24512,N_24319,N_24326);
xnor U24513 (N_24513,N_24327,N_24208);
nor U24514 (N_24514,N_24225,N_24324);
or U24515 (N_24515,N_24368,N_24317);
nor U24516 (N_24516,N_24347,N_24390);
or U24517 (N_24517,N_24309,N_24320);
nand U24518 (N_24518,N_24216,N_24343);
and U24519 (N_24519,N_24237,N_24203);
nand U24520 (N_24520,N_24364,N_24219);
and U24521 (N_24521,N_24227,N_24265);
nand U24522 (N_24522,N_24349,N_24371);
nor U24523 (N_24523,N_24381,N_24292);
nor U24524 (N_24524,N_24339,N_24324);
or U24525 (N_24525,N_24289,N_24299);
and U24526 (N_24526,N_24343,N_24388);
xor U24527 (N_24527,N_24255,N_24317);
and U24528 (N_24528,N_24333,N_24245);
xnor U24529 (N_24529,N_24368,N_24301);
or U24530 (N_24530,N_24315,N_24346);
and U24531 (N_24531,N_24380,N_24271);
nand U24532 (N_24532,N_24321,N_24311);
and U24533 (N_24533,N_24238,N_24353);
and U24534 (N_24534,N_24275,N_24386);
and U24535 (N_24535,N_24302,N_24232);
nor U24536 (N_24536,N_24226,N_24349);
and U24537 (N_24537,N_24353,N_24351);
or U24538 (N_24538,N_24371,N_24221);
nand U24539 (N_24539,N_24344,N_24398);
and U24540 (N_24540,N_24342,N_24267);
or U24541 (N_24541,N_24208,N_24234);
nor U24542 (N_24542,N_24316,N_24230);
or U24543 (N_24543,N_24239,N_24280);
xnor U24544 (N_24544,N_24270,N_24227);
and U24545 (N_24545,N_24238,N_24224);
xor U24546 (N_24546,N_24226,N_24286);
or U24547 (N_24547,N_24261,N_24393);
and U24548 (N_24548,N_24260,N_24233);
nand U24549 (N_24549,N_24348,N_24304);
xnor U24550 (N_24550,N_24341,N_24298);
xor U24551 (N_24551,N_24329,N_24389);
or U24552 (N_24552,N_24358,N_24337);
nor U24553 (N_24553,N_24270,N_24399);
and U24554 (N_24554,N_24292,N_24344);
xnor U24555 (N_24555,N_24281,N_24212);
and U24556 (N_24556,N_24316,N_24235);
xor U24557 (N_24557,N_24383,N_24262);
nor U24558 (N_24558,N_24228,N_24270);
nand U24559 (N_24559,N_24311,N_24248);
xor U24560 (N_24560,N_24259,N_24223);
and U24561 (N_24561,N_24350,N_24363);
nor U24562 (N_24562,N_24247,N_24369);
and U24563 (N_24563,N_24353,N_24372);
nand U24564 (N_24564,N_24333,N_24283);
xnor U24565 (N_24565,N_24244,N_24380);
or U24566 (N_24566,N_24386,N_24242);
nand U24567 (N_24567,N_24234,N_24274);
and U24568 (N_24568,N_24365,N_24350);
nand U24569 (N_24569,N_24353,N_24398);
or U24570 (N_24570,N_24386,N_24317);
xnor U24571 (N_24571,N_24256,N_24260);
nor U24572 (N_24572,N_24291,N_24378);
nor U24573 (N_24573,N_24271,N_24241);
nor U24574 (N_24574,N_24353,N_24315);
xor U24575 (N_24575,N_24373,N_24319);
nor U24576 (N_24576,N_24389,N_24375);
or U24577 (N_24577,N_24226,N_24309);
and U24578 (N_24578,N_24289,N_24257);
nand U24579 (N_24579,N_24314,N_24348);
or U24580 (N_24580,N_24210,N_24339);
or U24581 (N_24581,N_24304,N_24206);
or U24582 (N_24582,N_24268,N_24260);
or U24583 (N_24583,N_24265,N_24208);
nor U24584 (N_24584,N_24206,N_24342);
or U24585 (N_24585,N_24388,N_24330);
nand U24586 (N_24586,N_24342,N_24258);
and U24587 (N_24587,N_24296,N_24342);
or U24588 (N_24588,N_24379,N_24248);
or U24589 (N_24589,N_24336,N_24388);
nor U24590 (N_24590,N_24305,N_24396);
nand U24591 (N_24591,N_24357,N_24361);
or U24592 (N_24592,N_24381,N_24328);
nand U24593 (N_24593,N_24216,N_24212);
and U24594 (N_24594,N_24211,N_24216);
nand U24595 (N_24595,N_24311,N_24345);
xor U24596 (N_24596,N_24252,N_24315);
and U24597 (N_24597,N_24395,N_24328);
nor U24598 (N_24598,N_24360,N_24237);
or U24599 (N_24599,N_24374,N_24285);
and U24600 (N_24600,N_24439,N_24504);
or U24601 (N_24601,N_24453,N_24524);
nor U24602 (N_24602,N_24516,N_24596);
nand U24603 (N_24603,N_24530,N_24514);
and U24604 (N_24604,N_24484,N_24488);
and U24605 (N_24605,N_24507,N_24492);
xor U24606 (N_24606,N_24464,N_24442);
and U24607 (N_24607,N_24526,N_24546);
xnor U24608 (N_24608,N_24558,N_24440);
xnor U24609 (N_24609,N_24433,N_24496);
xor U24610 (N_24610,N_24432,N_24460);
nor U24611 (N_24611,N_24584,N_24500);
or U24612 (N_24612,N_24580,N_24571);
and U24613 (N_24613,N_24474,N_24578);
and U24614 (N_24614,N_24407,N_24446);
or U24615 (N_24615,N_24489,N_24557);
nor U24616 (N_24616,N_24417,N_24473);
xor U24617 (N_24617,N_24490,N_24475);
or U24618 (N_24618,N_24517,N_24503);
or U24619 (N_24619,N_24538,N_24477);
or U24620 (N_24620,N_24468,N_24494);
or U24621 (N_24621,N_24561,N_24569);
xnor U24622 (N_24622,N_24497,N_24411);
nand U24623 (N_24623,N_24427,N_24556);
or U24624 (N_24624,N_24586,N_24532);
nor U24625 (N_24625,N_24552,N_24574);
nand U24626 (N_24626,N_24450,N_24413);
nor U24627 (N_24627,N_24531,N_24520);
xor U24628 (N_24628,N_24593,N_24548);
and U24629 (N_24629,N_24588,N_24577);
nand U24630 (N_24630,N_24592,N_24563);
and U24631 (N_24631,N_24438,N_24521);
nand U24632 (N_24632,N_24452,N_24581);
nor U24633 (N_24633,N_24481,N_24567);
nand U24634 (N_24634,N_24410,N_24466);
xnor U24635 (N_24635,N_24583,N_24443);
xor U24636 (N_24636,N_24595,N_24591);
nand U24637 (N_24637,N_24576,N_24467);
nor U24638 (N_24638,N_24506,N_24406);
or U24639 (N_24639,N_24568,N_24445);
and U24640 (N_24640,N_24478,N_24560);
and U24641 (N_24641,N_24415,N_24599);
nor U24642 (N_24642,N_24405,N_24476);
nand U24643 (N_24643,N_24543,N_24470);
or U24644 (N_24644,N_24454,N_24551);
xor U24645 (N_24645,N_24545,N_24422);
and U24646 (N_24646,N_24431,N_24429);
nor U24647 (N_24647,N_24508,N_24434);
and U24648 (N_24648,N_24501,N_24585);
nor U24649 (N_24649,N_24455,N_24573);
xor U24650 (N_24650,N_24562,N_24502);
nor U24651 (N_24651,N_24553,N_24419);
xnor U24652 (N_24652,N_24550,N_24483);
nor U24653 (N_24653,N_24533,N_24401);
or U24654 (N_24654,N_24426,N_24491);
or U24655 (N_24655,N_24510,N_24527);
and U24656 (N_24656,N_24570,N_24424);
nand U24657 (N_24657,N_24547,N_24572);
xor U24658 (N_24658,N_24536,N_24498);
and U24659 (N_24659,N_24400,N_24589);
nand U24660 (N_24660,N_24493,N_24512);
nand U24661 (N_24661,N_24441,N_24487);
and U24662 (N_24662,N_24435,N_24482);
and U24663 (N_24663,N_24461,N_24403);
and U24664 (N_24664,N_24554,N_24540);
and U24665 (N_24665,N_24449,N_24518);
nor U24666 (N_24666,N_24402,N_24505);
xnor U24667 (N_24667,N_24539,N_24587);
or U24668 (N_24668,N_24541,N_24418);
nor U24669 (N_24669,N_24404,N_24421);
or U24670 (N_24670,N_24519,N_24447);
or U24671 (N_24671,N_24409,N_24448);
and U24672 (N_24672,N_24451,N_24416);
nor U24673 (N_24673,N_24597,N_24480);
and U24674 (N_24674,N_24499,N_24479);
nor U24675 (N_24675,N_24575,N_24457);
nor U24676 (N_24676,N_24428,N_24456);
or U24677 (N_24677,N_24528,N_24436);
nand U24678 (N_24678,N_24486,N_24515);
and U24679 (N_24679,N_24559,N_24529);
and U24680 (N_24680,N_24472,N_24523);
or U24681 (N_24681,N_24590,N_24469);
or U24682 (N_24682,N_24579,N_24471);
and U24683 (N_24683,N_24511,N_24495);
nor U24684 (N_24684,N_24444,N_24463);
nor U24685 (N_24685,N_24408,N_24423);
nand U24686 (N_24686,N_24458,N_24535);
nand U24687 (N_24687,N_24549,N_24594);
and U24688 (N_24688,N_24420,N_24465);
nor U24689 (N_24689,N_24509,N_24425);
xor U24690 (N_24690,N_24412,N_24414);
nor U24691 (N_24691,N_24566,N_24555);
or U24692 (N_24692,N_24525,N_24544);
nor U24693 (N_24693,N_24542,N_24462);
xnor U24694 (N_24694,N_24513,N_24437);
nor U24695 (N_24695,N_24565,N_24485);
and U24696 (N_24696,N_24537,N_24522);
nor U24697 (N_24697,N_24564,N_24459);
nand U24698 (N_24698,N_24598,N_24582);
xor U24699 (N_24699,N_24534,N_24430);
and U24700 (N_24700,N_24503,N_24413);
and U24701 (N_24701,N_24576,N_24406);
nand U24702 (N_24702,N_24472,N_24475);
or U24703 (N_24703,N_24437,N_24462);
nor U24704 (N_24704,N_24407,N_24588);
nand U24705 (N_24705,N_24500,N_24589);
nand U24706 (N_24706,N_24540,N_24491);
or U24707 (N_24707,N_24527,N_24490);
nand U24708 (N_24708,N_24434,N_24563);
nand U24709 (N_24709,N_24442,N_24449);
or U24710 (N_24710,N_24541,N_24548);
or U24711 (N_24711,N_24498,N_24538);
nand U24712 (N_24712,N_24541,N_24495);
nand U24713 (N_24713,N_24556,N_24482);
or U24714 (N_24714,N_24538,N_24438);
nand U24715 (N_24715,N_24556,N_24432);
nor U24716 (N_24716,N_24564,N_24478);
xor U24717 (N_24717,N_24529,N_24480);
xnor U24718 (N_24718,N_24565,N_24589);
nand U24719 (N_24719,N_24586,N_24418);
xnor U24720 (N_24720,N_24400,N_24427);
and U24721 (N_24721,N_24513,N_24546);
nor U24722 (N_24722,N_24527,N_24597);
and U24723 (N_24723,N_24568,N_24479);
and U24724 (N_24724,N_24548,N_24536);
nor U24725 (N_24725,N_24483,N_24538);
and U24726 (N_24726,N_24490,N_24552);
nor U24727 (N_24727,N_24471,N_24442);
or U24728 (N_24728,N_24468,N_24514);
or U24729 (N_24729,N_24486,N_24491);
or U24730 (N_24730,N_24541,N_24470);
nor U24731 (N_24731,N_24402,N_24498);
xnor U24732 (N_24732,N_24485,N_24493);
or U24733 (N_24733,N_24442,N_24437);
nor U24734 (N_24734,N_24561,N_24498);
or U24735 (N_24735,N_24507,N_24545);
nor U24736 (N_24736,N_24480,N_24586);
and U24737 (N_24737,N_24533,N_24442);
nor U24738 (N_24738,N_24463,N_24421);
nand U24739 (N_24739,N_24476,N_24450);
nor U24740 (N_24740,N_24574,N_24429);
nand U24741 (N_24741,N_24479,N_24590);
xnor U24742 (N_24742,N_24569,N_24586);
nand U24743 (N_24743,N_24445,N_24475);
nor U24744 (N_24744,N_24463,N_24476);
or U24745 (N_24745,N_24429,N_24427);
or U24746 (N_24746,N_24467,N_24508);
nand U24747 (N_24747,N_24483,N_24506);
nor U24748 (N_24748,N_24535,N_24524);
nand U24749 (N_24749,N_24413,N_24553);
nor U24750 (N_24750,N_24578,N_24526);
or U24751 (N_24751,N_24471,N_24480);
and U24752 (N_24752,N_24461,N_24491);
nor U24753 (N_24753,N_24570,N_24477);
nand U24754 (N_24754,N_24470,N_24526);
and U24755 (N_24755,N_24559,N_24482);
and U24756 (N_24756,N_24538,N_24514);
xnor U24757 (N_24757,N_24426,N_24536);
nor U24758 (N_24758,N_24534,N_24575);
or U24759 (N_24759,N_24422,N_24521);
nand U24760 (N_24760,N_24588,N_24464);
nand U24761 (N_24761,N_24586,N_24578);
or U24762 (N_24762,N_24480,N_24590);
xnor U24763 (N_24763,N_24472,N_24562);
nand U24764 (N_24764,N_24464,N_24519);
nand U24765 (N_24765,N_24567,N_24427);
and U24766 (N_24766,N_24558,N_24485);
nand U24767 (N_24767,N_24556,N_24542);
or U24768 (N_24768,N_24557,N_24536);
or U24769 (N_24769,N_24550,N_24491);
xnor U24770 (N_24770,N_24525,N_24553);
or U24771 (N_24771,N_24544,N_24542);
or U24772 (N_24772,N_24482,N_24587);
nand U24773 (N_24773,N_24509,N_24560);
nand U24774 (N_24774,N_24493,N_24435);
xor U24775 (N_24775,N_24464,N_24433);
and U24776 (N_24776,N_24433,N_24446);
nand U24777 (N_24777,N_24572,N_24554);
and U24778 (N_24778,N_24588,N_24423);
and U24779 (N_24779,N_24524,N_24435);
nor U24780 (N_24780,N_24549,N_24582);
and U24781 (N_24781,N_24460,N_24475);
nor U24782 (N_24782,N_24431,N_24436);
nand U24783 (N_24783,N_24473,N_24561);
nor U24784 (N_24784,N_24449,N_24560);
nor U24785 (N_24785,N_24536,N_24528);
nor U24786 (N_24786,N_24563,N_24523);
nand U24787 (N_24787,N_24594,N_24479);
nand U24788 (N_24788,N_24407,N_24526);
nand U24789 (N_24789,N_24564,N_24476);
xor U24790 (N_24790,N_24556,N_24562);
nor U24791 (N_24791,N_24448,N_24491);
xnor U24792 (N_24792,N_24526,N_24549);
xor U24793 (N_24793,N_24565,N_24425);
xor U24794 (N_24794,N_24582,N_24517);
xnor U24795 (N_24795,N_24408,N_24518);
nor U24796 (N_24796,N_24572,N_24510);
xnor U24797 (N_24797,N_24491,N_24505);
or U24798 (N_24798,N_24451,N_24591);
nor U24799 (N_24799,N_24521,N_24558);
nor U24800 (N_24800,N_24670,N_24682);
xor U24801 (N_24801,N_24667,N_24724);
nand U24802 (N_24802,N_24617,N_24662);
and U24803 (N_24803,N_24638,N_24679);
nor U24804 (N_24804,N_24629,N_24661);
or U24805 (N_24805,N_24614,N_24630);
xor U24806 (N_24806,N_24770,N_24793);
xor U24807 (N_24807,N_24720,N_24694);
or U24808 (N_24808,N_24717,N_24751);
xnor U24809 (N_24809,N_24719,N_24772);
or U24810 (N_24810,N_24708,N_24603);
and U24811 (N_24811,N_24792,N_24650);
and U24812 (N_24812,N_24785,N_24652);
nand U24813 (N_24813,N_24733,N_24780);
nand U24814 (N_24814,N_24731,N_24659);
nand U24815 (N_24815,N_24636,N_24711);
nand U24816 (N_24816,N_24695,N_24728);
nor U24817 (N_24817,N_24737,N_24705);
or U24818 (N_24818,N_24746,N_24699);
nand U24819 (N_24819,N_24658,N_24759);
nor U24820 (N_24820,N_24620,N_24796);
xor U24821 (N_24821,N_24660,N_24762);
xnor U24822 (N_24822,N_24697,N_24788);
and U24823 (N_24823,N_24797,N_24721);
nor U24824 (N_24824,N_24714,N_24752);
nor U24825 (N_24825,N_24778,N_24726);
nand U24826 (N_24826,N_24691,N_24609);
xor U24827 (N_24827,N_24791,N_24651);
nand U24828 (N_24828,N_24698,N_24753);
or U24829 (N_24829,N_24602,N_24637);
and U24830 (N_24830,N_24730,N_24775);
or U24831 (N_24831,N_24795,N_24649);
nor U24832 (N_24832,N_24779,N_24668);
or U24833 (N_24833,N_24718,N_24703);
nor U24834 (N_24834,N_24712,N_24756);
nand U24835 (N_24835,N_24757,N_24601);
and U24836 (N_24836,N_24615,N_24610);
xor U24837 (N_24837,N_24623,N_24642);
nand U24838 (N_24838,N_24787,N_24639);
nand U24839 (N_24839,N_24624,N_24777);
and U24840 (N_24840,N_24789,N_24631);
nand U24841 (N_24841,N_24635,N_24776);
nand U24842 (N_24842,N_24687,N_24755);
nand U24843 (N_24843,N_24600,N_24771);
and U24844 (N_24844,N_24673,N_24713);
or U24845 (N_24845,N_24680,N_24655);
and U24846 (N_24846,N_24736,N_24641);
and U24847 (N_24847,N_24765,N_24754);
or U24848 (N_24848,N_24743,N_24773);
nand U24849 (N_24849,N_24625,N_24611);
nand U24850 (N_24850,N_24786,N_24716);
nor U24851 (N_24851,N_24616,N_24783);
and U24852 (N_24852,N_24738,N_24799);
nand U24853 (N_24853,N_24729,N_24790);
nor U24854 (N_24854,N_24696,N_24760);
and U24855 (N_24855,N_24798,N_24607);
and U24856 (N_24856,N_24690,N_24782);
and U24857 (N_24857,N_24741,N_24683);
nor U24858 (N_24858,N_24722,N_24707);
or U24859 (N_24859,N_24669,N_24622);
nand U24860 (N_24860,N_24763,N_24676);
xnor U24861 (N_24861,N_24732,N_24628);
and U24862 (N_24862,N_24640,N_24633);
or U24863 (N_24863,N_24723,N_24604);
or U24864 (N_24864,N_24747,N_24685);
nor U24865 (N_24865,N_24727,N_24768);
and U24866 (N_24866,N_24774,N_24619);
xor U24867 (N_24867,N_24794,N_24688);
nand U24868 (N_24868,N_24704,N_24643);
nor U24869 (N_24869,N_24613,N_24644);
nor U24870 (N_24870,N_24608,N_24648);
or U24871 (N_24871,N_24761,N_24671);
nor U24872 (N_24872,N_24663,N_24645);
or U24873 (N_24873,N_24769,N_24664);
and U24874 (N_24874,N_24689,N_24748);
xnor U24875 (N_24875,N_24646,N_24742);
xor U24876 (N_24876,N_24626,N_24740);
nand U24877 (N_24877,N_24710,N_24709);
and U24878 (N_24878,N_24605,N_24693);
or U24879 (N_24879,N_24654,N_24735);
nand U24880 (N_24880,N_24715,N_24672);
or U24881 (N_24881,N_24749,N_24634);
nand U24882 (N_24882,N_24781,N_24657);
and U24883 (N_24883,N_24686,N_24675);
and U24884 (N_24884,N_24678,N_24665);
nand U24885 (N_24885,N_24758,N_24684);
nor U24886 (N_24886,N_24692,N_24744);
nor U24887 (N_24887,N_24647,N_24700);
or U24888 (N_24888,N_24612,N_24745);
nand U24889 (N_24889,N_24666,N_24674);
nand U24890 (N_24890,N_24702,N_24677);
nand U24891 (N_24891,N_24766,N_24725);
and U24892 (N_24892,N_24618,N_24627);
nand U24893 (N_24893,N_24621,N_24701);
and U24894 (N_24894,N_24767,N_24739);
and U24895 (N_24895,N_24706,N_24656);
nand U24896 (N_24896,N_24681,N_24632);
xnor U24897 (N_24897,N_24606,N_24734);
or U24898 (N_24898,N_24653,N_24750);
and U24899 (N_24899,N_24764,N_24784);
and U24900 (N_24900,N_24781,N_24765);
or U24901 (N_24901,N_24795,N_24757);
nand U24902 (N_24902,N_24661,N_24682);
nand U24903 (N_24903,N_24679,N_24774);
xor U24904 (N_24904,N_24762,N_24671);
xor U24905 (N_24905,N_24762,N_24782);
and U24906 (N_24906,N_24651,N_24711);
nor U24907 (N_24907,N_24653,N_24711);
nor U24908 (N_24908,N_24712,N_24623);
nor U24909 (N_24909,N_24777,N_24760);
xor U24910 (N_24910,N_24699,N_24638);
and U24911 (N_24911,N_24747,N_24612);
and U24912 (N_24912,N_24649,N_24683);
nand U24913 (N_24913,N_24622,N_24785);
nand U24914 (N_24914,N_24611,N_24698);
nor U24915 (N_24915,N_24640,N_24791);
nand U24916 (N_24916,N_24667,N_24790);
or U24917 (N_24917,N_24767,N_24664);
nor U24918 (N_24918,N_24784,N_24718);
and U24919 (N_24919,N_24608,N_24602);
xor U24920 (N_24920,N_24762,N_24798);
xor U24921 (N_24921,N_24628,N_24756);
and U24922 (N_24922,N_24787,N_24743);
xor U24923 (N_24923,N_24660,N_24716);
nor U24924 (N_24924,N_24686,N_24775);
xor U24925 (N_24925,N_24703,N_24773);
xor U24926 (N_24926,N_24688,N_24695);
or U24927 (N_24927,N_24696,N_24668);
and U24928 (N_24928,N_24763,N_24783);
nand U24929 (N_24929,N_24628,N_24778);
nand U24930 (N_24930,N_24671,N_24736);
xor U24931 (N_24931,N_24719,N_24779);
or U24932 (N_24932,N_24608,N_24691);
nor U24933 (N_24933,N_24724,N_24737);
or U24934 (N_24934,N_24649,N_24741);
and U24935 (N_24935,N_24671,N_24793);
xnor U24936 (N_24936,N_24664,N_24631);
nand U24937 (N_24937,N_24608,N_24745);
nand U24938 (N_24938,N_24633,N_24705);
nor U24939 (N_24939,N_24653,N_24605);
xnor U24940 (N_24940,N_24694,N_24644);
or U24941 (N_24941,N_24603,N_24760);
nand U24942 (N_24942,N_24621,N_24742);
nand U24943 (N_24943,N_24730,N_24627);
nor U24944 (N_24944,N_24625,N_24646);
nor U24945 (N_24945,N_24699,N_24663);
nor U24946 (N_24946,N_24710,N_24673);
nand U24947 (N_24947,N_24781,N_24628);
xnor U24948 (N_24948,N_24705,N_24776);
and U24949 (N_24949,N_24610,N_24674);
nor U24950 (N_24950,N_24664,N_24630);
nor U24951 (N_24951,N_24717,N_24731);
and U24952 (N_24952,N_24662,N_24770);
xor U24953 (N_24953,N_24696,N_24697);
xor U24954 (N_24954,N_24723,N_24771);
or U24955 (N_24955,N_24697,N_24707);
or U24956 (N_24956,N_24772,N_24796);
and U24957 (N_24957,N_24714,N_24742);
and U24958 (N_24958,N_24618,N_24686);
and U24959 (N_24959,N_24651,N_24670);
xnor U24960 (N_24960,N_24763,N_24718);
nor U24961 (N_24961,N_24750,N_24784);
xnor U24962 (N_24962,N_24784,N_24786);
or U24963 (N_24963,N_24688,N_24716);
nor U24964 (N_24964,N_24731,N_24782);
xor U24965 (N_24965,N_24652,N_24677);
or U24966 (N_24966,N_24642,N_24707);
and U24967 (N_24967,N_24743,N_24789);
xnor U24968 (N_24968,N_24751,N_24709);
and U24969 (N_24969,N_24777,N_24629);
nand U24970 (N_24970,N_24616,N_24623);
or U24971 (N_24971,N_24677,N_24602);
or U24972 (N_24972,N_24659,N_24761);
or U24973 (N_24973,N_24797,N_24781);
nor U24974 (N_24974,N_24762,N_24709);
and U24975 (N_24975,N_24762,N_24659);
nand U24976 (N_24976,N_24621,N_24640);
nor U24977 (N_24977,N_24793,N_24718);
xor U24978 (N_24978,N_24672,N_24666);
nand U24979 (N_24979,N_24720,N_24697);
or U24980 (N_24980,N_24797,N_24749);
and U24981 (N_24981,N_24765,N_24746);
and U24982 (N_24982,N_24755,N_24757);
or U24983 (N_24983,N_24633,N_24615);
xnor U24984 (N_24984,N_24722,N_24746);
xnor U24985 (N_24985,N_24672,N_24643);
or U24986 (N_24986,N_24652,N_24751);
nand U24987 (N_24987,N_24738,N_24773);
nor U24988 (N_24988,N_24680,N_24692);
xor U24989 (N_24989,N_24714,N_24648);
nand U24990 (N_24990,N_24721,N_24690);
nand U24991 (N_24991,N_24685,N_24774);
or U24992 (N_24992,N_24627,N_24672);
and U24993 (N_24993,N_24609,N_24653);
nand U24994 (N_24994,N_24657,N_24662);
or U24995 (N_24995,N_24697,N_24771);
or U24996 (N_24996,N_24630,N_24701);
and U24997 (N_24997,N_24621,N_24685);
and U24998 (N_24998,N_24785,N_24631);
nand U24999 (N_24999,N_24653,N_24634);
xor UO_0 (O_0,N_24877,N_24829);
nand UO_1 (O_1,N_24804,N_24890);
nor UO_2 (O_2,N_24876,N_24874);
nor UO_3 (O_3,N_24937,N_24850);
nor UO_4 (O_4,N_24925,N_24853);
xor UO_5 (O_5,N_24900,N_24983);
or UO_6 (O_6,N_24950,N_24940);
nand UO_7 (O_7,N_24898,N_24966);
or UO_8 (O_8,N_24843,N_24864);
xnor UO_9 (O_9,N_24916,N_24969);
xor UO_10 (O_10,N_24817,N_24986);
nor UO_11 (O_11,N_24857,N_24888);
xnor UO_12 (O_12,N_24845,N_24926);
or UO_13 (O_13,N_24944,N_24987);
nand UO_14 (O_14,N_24998,N_24825);
nand UO_15 (O_15,N_24931,N_24828);
xor UO_16 (O_16,N_24820,N_24912);
and UO_17 (O_17,N_24805,N_24847);
nand UO_18 (O_18,N_24884,N_24835);
xor UO_19 (O_19,N_24826,N_24899);
or UO_20 (O_20,N_24985,N_24870);
xnor UO_21 (O_21,N_24967,N_24852);
nor UO_22 (O_22,N_24975,N_24891);
and UO_23 (O_23,N_24801,N_24895);
or UO_24 (O_24,N_24956,N_24973);
or UO_25 (O_25,N_24911,N_24863);
and UO_26 (O_26,N_24968,N_24907);
and UO_27 (O_27,N_24980,N_24892);
xor UO_28 (O_28,N_24803,N_24909);
xnor UO_29 (O_29,N_24903,N_24812);
nor UO_30 (O_30,N_24851,N_24988);
and UO_31 (O_31,N_24800,N_24878);
and UO_32 (O_32,N_24977,N_24929);
nor UO_33 (O_33,N_24855,N_24994);
and UO_34 (O_34,N_24936,N_24894);
or UO_35 (O_35,N_24930,N_24955);
or UO_36 (O_36,N_24919,N_24871);
or UO_37 (O_37,N_24979,N_24808);
or UO_38 (O_38,N_24984,N_24814);
nand UO_39 (O_39,N_24844,N_24954);
and UO_40 (O_40,N_24952,N_24861);
and UO_41 (O_41,N_24971,N_24862);
nand UO_42 (O_42,N_24906,N_24881);
and UO_43 (O_43,N_24920,N_24962);
nand UO_44 (O_44,N_24993,N_24941);
xor UO_45 (O_45,N_24875,N_24872);
and UO_46 (O_46,N_24982,N_24886);
and UO_47 (O_47,N_24905,N_24992);
and UO_48 (O_48,N_24913,N_24841);
nor UO_49 (O_49,N_24928,N_24959);
and UO_50 (O_50,N_24945,N_24946);
or UO_51 (O_51,N_24932,N_24818);
xor UO_52 (O_52,N_24951,N_24823);
xor UO_53 (O_53,N_24961,N_24976);
and UO_54 (O_54,N_24918,N_24834);
and UO_55 (O_55,N_24939,N_24824);
xor UO_56 (O_56,N_24990,N_24873);
nor UO_57 (O_57,N_24908,N_24883);
xnor UO_58 (O_58,N_24849,N_24947);
xnor UO_59 (O_59,N_24810,N_24949);
and UO_60 (O_60,N_24815,N_24974);
or UO_61 (O_61,N_24963,N_24921);
nor UO_62 (O_62,N_24989,N_24830);
nand UO_63 (O_63,N_24901,N_24904);
and UO_64 (O_64,N_24867,N_24933);
xnor UO_65 (O_65,N_24816,N_24923);
and UO_66 (O_66,N_24811,N_24910);
and UO_67 (O_67,N_24965,N_24943);
or UO_68 (O_68,N_24914,N_24869);
xnor UO_69 (O_69,N_24935,N_24832);
xnor UO_70 (O_70,N_24836,N_24822);
and UO_71 (O_71,N_24934,N_24897);
xnor UO_72 (O_72,N_24999,N_24893);
xnor UO_73 (O_73,N_24831,N_24879);
and UO_74 (O_74,N_24865,N_24837);
nand UO_75 (O_75,N_24880,N_24866);
xor UO_76 (O_76,N_24848,N_24885);
nor UO_77 (O_77,N_24991,N_24809);
nor UO_78 (O_78,N_24927,N_24889);
nor UO_79 (O_79,N_24802,N_24819);
nand UO_80 (O_80,N_24938,N_24896);
or UO_81 (O_81,N_24806,N_24838);
nand UO_82 (O_82,N_24924,N_24922);
nor UO_83 (O_83,N_24960,N_24917);
nor UO_84 (O_84,N_24981,N_24840);
or UO_85 (O_85,N_24996,N_24978);
nand UO_86 (O_86,N_24972,N_24942);
nor UO_87 (O_87,N_24854,N_24807);
xnor UO_88 (O_88,N_24957,N_24915);
xnor UO_89 (O_89,N_24821,N_24948);
xnor UO_90 (O_90,N_24953,N_24887);
nand UO_91 (O_91,N_24856,N_24859);
and UO_92 (O_92,N_24958,N_24964);
xnor UO_93 (O_93,N_24860,N_24813);
and UO_94 (O_94,N_24827,N_24842);
nand UO_95 (O_95,N_24902,N_24882);
xor UO_96 (O_96,N_24997,N_24858);
or UO_97 (O_97,N_24839,N_24833);
and UO_98 (O_98,N_24868,N_24995);
xor UO_99 (O_99,N_24846,N_24970);
xnor UO_100 (O_100,N_24942,N_24977);
xor UO_101 (O_101,N_24867,N_24967);
nand UO_102 (O_102,N_24955,N_24839);
and UO_103 (O_103,N_24813,N_24873);
or UO_104 (O_104,N_24961,N_24828);
nor UO_105 (O_105,N_24854,N_24976);
nor UO_106 (O_106,N_24800,N_24847);
nand UO_107 (O_107,N_24954,N_24872);
nand UO_108 (O_108,N_24880,N_24833);
and UO_109 (O_109,N_24853,N_24830);
nor UO_110 (O_110,N_24942,N_24828);
nand UO_111 (O_111,N_24892,N_24853);
xnor UO_112 (O_112,N_24942,N_24805);
nand UO_113 (O_113,N_24814,N_24936);
and UO_114 (O_114,N_24873,N_24870);
xnor UO_115 (O_115,N_24993,N_24939);
xnor UO_116 (O_116,N_24901,N_24948);
xor UO_117 (O_117,N_24906,N_24997);
nand UO_118 (O_118,N_24915,N_24821);
nor UO_119 (O_119,N_24880,N_24825);
or UO_120 (O_120,N_24827,N_24922);
nand UO_121 (O_121,N_24825,N_24983);
and UO_122 (O_122,N_24919,N_24838);
or UO_123 (O_123,N_24839,N_24919);
nand UO_124 (O_124,N_24997,N_24970);
xnor UO_125 (O_125,N_24932,N_24979);
or UO_126 (O_126,N_24842,N_24961);
xor UO_127 (O_127,N_24818,N_24994);
nand UO_128 (O_128,N_24830,N_24931);
xnor UO_129 (O_129,N_24847,N_24872);
or UO_130 (O_130,N_24982,N_24932);
or UO_131 (O_131,N_24823,N_24895);
or UO_132 (O_132,N_24812,N_24910);
or UO_133 (O_133,N_24812,N_24832);
nor UO_134 (O_134,N_24891,N_24811);
nor UO_135 (O_135,N_24875,N_24811);
nand UO_136 (O_136,N_24887,N_24908);
and UO_137 (O_137,N_24951,N_24922);
nor UO_138 (O_138,N_24873,N_24842);
xor UO_139 (O_139,N_24966,N_24820);
xor UO_140 (O_140,N_24938,N_24829);
or UO_141 (O_141,N_24888,N_24818);
nor UO_142 (O_142,N_24984,N_24818);
nand UO_143 (O_143,N_24969,N_24802);
nand UO_144 (O_144,N_24814,N_24989);
nand UO_145 (O_145,N_24867,N_24957);
and UO_146 (O_146,N_24822,N_24919);
nand UO_147 (O_147,N_24873,N_24821);
and UO_148 (O_148,N_24995,N_24926);
xnor UO_149 (O_149,N_24847,N_24989);
and UO_150 (O_150,N_24856,N_24936);
nand UO_151 (O_151,N_24933,N_24847);
nor UO_152 (O_152,N_24836,N_24811);
xor UO_153 (O_153,N_24800,N_24825);
nand UO_154 (O_154,N_24894,N_24994);
xnor UO_155 (O_155,N_24844,N_24920);
or UO_156 (O_156,N_24825,N_24925);
and UO_157 (O_157,N_24926,N_24997);
nor UO_158 (O_158,N_24980,N_24974);
and UO_159 (O_159,N_24896,N_24873);
and UO_160 (O_160,N_24940,N_24907);
nand UO_161 (O_161,N_24891,N_24951);
xor UO_162 (O_162,N_24935,N_24986);
and UO_163 (O_163,N_24804,N_24841);
or UO_164 (O_164,N_24934,N_24826);
nor UO_165 (O_165,N_24932,N_24845);
nand UO_166 (O_166,N_24908,N_24854);
and UO_167 (O_167,N_24844,N_24955);
and UO_168 (O_168,N_24974,N_24826);
nor UO_169 (O_169,N_24885,N_24886);
and UO_170 (O_170,N_24846,N_24926);
and UO_171 (O_171,N_24807,N_24846);
or UO_172 (O_172,N_24912,N_24959);
xnor UO_173 (O_173,N_24870,N_24992);
and UO_174 (O_174,N_24895,N_24821);
nand UO_175 (O_175,N_24958,N_24903);
xor UO_176 (O_176,N_24992,N_24908);
nand UO_177 (O_177,N_24955,N_24854);
xor UO_178 (O_178,N_24863,N_24978);
nor UO_179 (O_179,N_24886,N_24828);
nand UO_180 (O_180,N_24974,N_24932);
nor UO_181 (O_181,N_24872,N_24857);
or UO_182 (O_182,N_24826,N_24952);
nor UO_183 (O_183,N_24879,N_24986);
or UO_184 (O_184,N_24953,N_24851);
nor UO_185 (O_185,N_24850,N_24897);
nand UO_186 (O_186,N_24929,N_24829);
and UO_187 (O_187,N_24940,N_24994);
and UO_188 (O_188,N_24843,N_24965);
xor UO_189 (O_189,N_24919,N_24896);
and UO_190 (O_190,N_24988,N_24916);
or UO_191 (O_191,N_24880,N_24828);
and UO_192 (O_192,N_24961,N_24964);
xnor UO_193 (O_193,N_24956,N_24938);
or UO_194 (O_194,N_24935,N_24833);
and UO_195 (O_195,N_24839,N_24869);
and UO_196 (O_196,N_24857,N_24922);
nor UO_197 (O_197,N_24846,N_24808);
or UO_198 (O_198,N_24850,N_24921);
xnor UO_199 (O_199,N_24864,N_24816);
or UO_200 (O_200,N_24819,N_24919);
or UO_201 (O_201,N_24866,N_24833);
nor UO_202 (O_202,N_24944,N_24964);
and UO_203 (O_203,N_24896,N_24887);
nand UO_204 (O_204,N_24866,N_24911);
xor UO_205 (O_205,N_24864,N_24819);
and UO_206 (O_206,N_24941,N_24807);
or UO_207 (O_207,N_24913,N_24957);
nand UO_208 (O_208,N_24820,N_24916);
and UO_209 (O_209,N_24899,N_24860);
nand UO_210 (O_210,N_24828,N_24837);
nand UO_211 (O_211,N_24818,N_24846);
nand UO_212 (O_212,N_24973,N_24941);
nand UO_213 (O_213,N_24850,N_24853);
or UO_214 (O_214,N_24958,N_24834);
or UO_215 (O_215,N_24854,N_24806);
and UO_216 (O_216,N_24836,N_24929);
and UO_217 (O_217,N_24815,N_24824);
or UO_218 (O_218,N_24984,N_24967);
and UO_219 (O_219,N_24804,N_24840);
xor UO_220 (O_220,N_24819,N_24983);
nand UO_221 (O_221,N_24978,N_24899);
and UO_222 (O_222,N_24991,N_24811);
and UO_223 (O_223,N_24800,N_24892);
nor UO_224 (O_224,N_24899,N_24999);
and UO_225 (O_225,N_24846,N_24874);
and UO_226 (O_226,N_24914,N_24905);
nor UO_227 (O_227,N_24807,N_24837);
xnor UO_228 (O_228,N_24926,N_24928);
nor UO_229 (O_229,N_24994,N_24975);
nand UO_230 (O_230,N_24861,N_24956);
nor UO_231 (O_231,N_24815,N_24867);
nor UO_232 (O_232,N_24821,N_24998);
nor UO_233 (O_233,N_24957,N_24829);
nand UO_234 (O_234,N_24866,N_24952);
xor UO_235 (O_235,N_24854,N_24929);
and UO_236 (O_236,N_24815,N_24950);
and UO_237 (O_237,N_24830,N_24835);
xnor UO_238 (O_238,N_24825,N_24979);
or UO_239 (O_239,N_24842,N_24839);
nor UO_240 (O_240,N_24874,N_24969);
and UO_241 (O_241,N_24990,N_24835);
and UO_242 (O_242,N_24852,N_24805);
and UO_243 (O_243,N_24966,N_24810);
nor UO_244 (O_244,N_24989,N_24984);
or UO_245 (O_245,N_24887,N_24806);
nand UO_246 (O_246,N_24938,N_24970);
nor UO_247 (O_247,N_24899,N_24904);
or UO_248 (O_248,N_24959,N_24984);
nand UO_249 (O_249,N_24852,N_24846);
and UO_250 (O_250,N_24921,N_24919);
or UO_251 (O_251,N_24920,N_24972);
nor UO_252 (O_252,N_24986,N_24996);
and UO_253 (O_253,N_24948,N_24977);
nor UO_254 (O_254,N_24902,N_24994);
and UO_255 (O_255,N_24978,N_24853);
nor UO_256 (O_256,N_24970,N_24829);
or UO_257 (O_257,N_24827,N_24884);
xor UO_258 (O_258,N_24912,N_24855);
and UO_259 (O_259,N_24933,N_24882);
and UO_260 (O_260,N_24870,N_24970);
nor UO_261 (O_261,N_24834,N_24971);
nand UO_262 (O_262,N_24976,N_24998);
nor UO_263 (O_263,N_24878,N_24828);
or UO_264 (O_264,N_24928,N_24937);
and UO_265 (O_265,N_24919,N_24836);
nand UO_266 (O_266,N_24892,N_24810);
nand UO_267 (O_267,N_24996,N_24851);
and UO_268 (O_268,N_24966,N_24983);
nand UO_269 (O_269,N_24946,N_24870);
nand UO_270 (O_270,N_24891,N_24884);
xor UO_271 (O_271,N_24934,N_24879);
or UO_272 (O_272,N_24810,N_24945);
or UO_273 (O_273,N_24881,N_24934);
nand UO_274 (O_274,N_24953,N_24916);
xnor UO_275 (O_275,N_24869,N_24857);
nor UO_276 (O_276,N_24863,N_24837);
nand UO_277 (O_277,N_24947,N_24943);
and UO_278 (O_278,N_24921,N_24923);
and UO_279 (O_279,N_24931,N_24891);
or UO_280 (O_280,N_24881,N_24945);
or UO_281 (O_281,N_24865,N_24993);
xnor UO_282 (O_282,N_24920,N_24816);
and UO_283 (O_283,N_24924,N_24842);
and UO_284 (O_284,N_24879,N_24808);
or UO_285 (O_285,N_24980,N_24967);
and UO_286 (O_286,N_24911,N_24842);
xnor UO_287 (O_287,N_24963,N_24945);
and UO_288 (O_288,N_24825,N_24999);
nand UO_289 (O_289,N_24944,N_24933);
nor UO_290 (O_290,N_24850,N_24839);
and UO_291 (O_291,N_24984,N_24864);
nor UO_292 (O_292,N_24856,N_24815);
or UO_293 (O_293,N_24837,N_24810);
nor UO_294 (O_294,N_24901,N_24955);
xnor UO_295 (O_295,N_24978,N_24802);
nand UO_296 (O_296,N_24928,N_24995);
and UO_297 (O_297,N_24944,N_24886);
xor UO_298 (O_298,N_24817,N_24922);
or UO_299 (O_299,N_24993,N_24948);
nor UO_300 (O_300,N_24918,N_24889);
nand UO_301 (O_301,N_24800,N_24924);
xnor UO_302 (O_302,N_24921,N_24827);
xor UO_303 (O_303,N_24835,N_24814);
nor UO_304 (O_304,N_24970,N_24975);
xor UO_305 (O_305,N_24851,N_24812);
xnor UO_306 (O_306,N_24845,N_24817);
nor UO_307 (O_307,N_24813,N_24915);
or UO_308 (O_308,N_24840,N_24913);
nor UO_309 (O_309,N_24872,N_24826);
or UO_310 (O_310,N_24884,N_24974);
nand UO_311 (O_311,N_24994,N_24830);
and UO_312 (O_312,N_24949,N_24804);
or UO_313 (O_313,N_24965,N_24881);
nand UO_314 (O_314,N_24884,N_24875);
and UO_315 (O_315,N_24843,N_24916);
nor UO_316 (O_316,N_24802,N_24891);
nor UO_317 (O_317,N_24997,N_24940);
nand UO_318 (O_318,N_24910,N_24997);
xnor UO_319 (O_319,N_24861,N_24968);
nor UO_320 (O_320,N_24827,N_24969);
and UO_321 (O_321,N_24989,N_24907);
nor UO_322 (O_322,N_24995,N_24977);
nand UO_323 (O_323,N_24843,N_24898);
and UO_324 (O_324,N_24946,N_24882);
or UO_325 (O_325,N_24925,N_24944);
and UO_326 (O_326,N_24965,N_24851);
xor UO_327 (O_327,N_24944,N_24939);
nor UO_328 (O_328,N_24938,N_24815);
or UO_329 (O_329,N_24990,N_24815);
nor UO_330 (O_330,N_24972,N_24957);
and UO_331 (O_331,N_24955,N_24888);
nand UO_332 (O_332,N_24990,N_24845);
and UO_333 (O_333,N_24911,N_24929);
nor UO_334 (O_334,N_24852,N_24832);
and UO_335 (O_335,N_24804,N_24964);
and UO_336 (O_336,N_24958,N_24844);
nand UO_337 (O_337,N_24883,N_24891);
nor UO_338 (O_338,N_24927,N_24862);
nor UO_339 (O_339,N_24900,N_24988);
nand UO_340 (O_340,N_24833,N_24908);
nand UO_341 (O_341,N_24800,N_24802);
nand UO_342 (O_342,N_24870,N_24988);
nand UO_343 (O_343,N_24925,N_24843);
nand UO_344 (O_344,N_24892,N_24829);
nor UO_345 (O_345,N_24917,N_24805);
and UO_346 (O_346,N_24927,N_24897);
or UO_347 (O_347,N_24881,N_24980);
xnor UO_348 (O_348,N_24965,N_24976);
nor UO_349 (O_349,N_24893,N_24835);
xnor UO_350 (O_350,N_24855,N_24862);
and UO_351 (O_351,N_24902,N_24935);
xnor UO_352 (O_352,N_24956,N_24933);
xor UO_353 (O_353,N_24935,N_24942);
nand UO_354 (O_354,N_24850,N_24962);
xor UO_355 (O_355,N_24920,N_24979);
nor UO_356 (O_356,N_24893,N_24952);
and UO_357 (O_357,N_24998,N_24868);
or UO_358 (O_358,N_24975,N_24972);
nor UO_359 (O_359,N_24959,N_24966);
or UO_360 (O_360,N_24810,N_24898);
nor UO_361 (O_361,N_24889,N_24871);
or UO_362 (O_362,N_24813,N_24830);
xor UO_363 (O_363,N_24915,N_24978);
nor UO_364 (O_364,N_24964,N_24858);
xnor UO_365 (O_365,N_24865,N_24876);
and UO_366 (O_366,N_24846,N_24975);
and UO_367 (O_367,N_24932,N_24994);
xnor UO_368 (O_368,N_24985,N_24993);
nand UO_369 (O_369,N_24923,N_24830);
nor UO_370 (O_370,N_24920,N_24945);
and UO_371 (O_371,N_24886,N_24865);
nand UO_372 (O_372,N_24846,N_24820);
nand UO_373 (O_373,N_24986,N_24972);
and UO_374 (O_374,N_24837,N_24919);
xor UO_375 (O_375,N_24914,N_24976);
nand UO_376 (O_376,N_24921,N_24967);
or UO_377 (O_377,N_24909,N_24949);
nand UO_378 (O_378,N_24839,N_24819);
and UO_379 (O_379,N_24894,N_24837);
xor UO_380 (O_380,N_24988,N_24847);
nor UO_381 (O_381,N_24834,N_24973);
xor UO_382 (O_382,N_24903,N_24996);
xnor UO_383 (O_383,N_24908,N_24851);
nand UO_384 (O_384,N_24878,N_24886);
and UO_385 (O_385,N_24857,N_24809);
nor UO_386 (O_386,N_24961,N_24956);
or UO_387 (O_387,N_24903,N_24945);
xnor UO_388 (O_388,N_24826,N_24896);
xnor UO_389 (O_389,N_24933,N_24968);
xor UO_390 (O_390,N_24879,N_24963);
nor UO_391 (O_391,N_24817,N_24934);
and UO_392 (O_392,N_24944,N_24897);
nand UO_393 (O_393,N_24889,N_24999);
nor UO_394 (O_394,N_24838,N_24844);
or UO_395 (O_395,N_24910,N_24891);
and UO_396 (O_396,N_24845,N_24922);
xor UO_397 (O_397,N_24957,N_24835);
nor UO_398 (O_398,N_24940,N_24931);
nor UO_399 (O_399,N_24884,N_24919);
nand UO_400 (O_400,N_24823,N_24820);
nand UO_401 (O_401,N_24800,N_24920);
nand UO_402 (O_402,N_24906,N_24823);
and UO_403 (O_403,N_24948,N_24932);
xor UO_404 (O_404,N_24964,N_24864);
and UO_405 (O_405,N_24810,N_24934);
or UO_406 (O_406,N_24855,N_24835);
nand UO_407 (O_407,N_24821,N_24986);
and UO_408 (O_408,N_24927,N_24893);
nor UO_409 (O_409,N_24841,N_24825);
nor UO_410 (O_410,N_24928,N_24903);
xor UO_411 (O_411,N_24995,N_24969);
xnor UO_412 (O_412,N_24921,N_24809);
nand UO_413 (O_413,N_24872,N_24858);
and UO_414 (O_414,N_24919,N_24918);
nor UO_415 (O_415,N_24836,N_24966);
nand UO_416 (O_416,N_24990,N_24961);
xor UO_417 (O_417,N_24871,N_24887);
and UO_418 (O_418,N_24930,N_24895);
nor UO_419 (O_419,N_24953,N_24920);
nand UO_420 (O_420,N_24942,N_24974);
nand UO_421 (O_421,N_24949,N_24863);
or UO_422 (O_422,N_24851,N_24991);
or UO_423 (O_423,N_24993,N_24802);
and UO_424 (O_424,N_24844,N_24965);
nor UO_425 (O_425,N_24954,N_24826);
and UO_426 (O_426,N_24879,N_24973);
xnor UO_427 (O_427,N_24805,N_24938);
nand UO_428 (O_428,N_24832,N_24918);
and UO_429 (O_429,N_24812,N_24999);
nor UO_430 (O_430,N_24965,N_24914);
and UO_431 (O_431,N_24997,N_24823);
and UO_432 (O_432,N_24960,N_24951);
and UO_433 (O_433,N_24824,N_24910);
xnor UO_434 (O_434,N_24932,N_24895);
nand UO_435 (O_435,N_24891,N_24835);
nand UO_436 (O_436,N_24913,N_24810);
or UO_437 (O_437,N_24853,N_24890);
nand UO_438 (O_438,N_24930,N_24972);
or UO_439 (O_439,N_24804,N_24905);
and UO_440 (O_440,N_24846,N_24877);
and UO_441 (O_441,N_24832,N_24848);
nor UO_442 (O_442,N_24943,N_24986);
or UO_443 (O_443,N_24838,N_24837);
xor UO_444 (O_444,N_24921,N_24801);
and UO_445 (O_445,N_24888,N_24902);
or UO_446 (O_446,N_24882,N_24871);
xor UO_447 (O_447,N_24821,N_24906);
nor UO_448 (O_448,N_24938,N_24806);
and UO_449 (O_449,N_24842,N_24875);
and UO_450 (O_450,N_24811,N_24935);
nand UO_451 (O_451,N_24828,N_24846);
nor UO_452 (O_452,N_24824,N_24919);
or UO_453 (O_453,N_24846,N_24974);
nand UO_454 (O_454,N_24832,N_24855);
xor UO_455 (O_455,N_24835,N_24874);
xnor UO_456 (O_456,N_24815,N_24988);
and UO_457 (O_457,N_24843,N_24871);
nand UO_458 (O_458,N_24803,N_24949);
nor UO_459 (O_459,N_24992,N_24875);
nor UO_460 (O_460,N_24816,N_24903);
nor UO_461 (O_461,N_24982,N_24945);
or UO_462 (O_462,N_24929,N_24865);
nand UO_463 (O_463,N_24923,N_24961);
xnor UO_464 (O_464,N_24924,N_24961);
nor UO_465 (O_465,N_24818,N_24831);
or UO_466 (O_466,N_24850,N_24847);
nand UO_467 (O_467,N_24942,N_24879);
nor UO_468 (O_468,N_24962,N_24890);
xnor UO_469 (O_469,N_24812,N_24898);
and UO_470 (O_470,N_24978,N_24864);
or UO_471 (O_471,N_24976,N_24881);
nand UO_472 (O_472,N_24911,N_24925);
nand UO_473 (O_473,N_24980,N_24800);
xor UO_474 (O_474,N_24906,N_24828);
and UO_475 (O_475,N_24886,N_24837);
nor UO_476 (O_476,N_24945,N_24965);
nand UO_477 (O_477,N_24805,N_24843);
xnor UO_478 (O_478,N_24858,N_24919);
xnor UO_479 (O_479,N_24805,N_24839);
or UO_480 (O_480,N_24873,N_24913);
xor UO_481 (O_481,N_24893,N_24972);
nor UO_482 (O_482,N_24831,N_24807);
nor UO_483 (O_483,N_24899,N_24956);
nor UO_484 (O_484,N_24937,N_24851);
xnor UO_485 (O_485,N_24976,N_24852);
nor UO_486 (O_486,N_24915,N_24853);
and UO_487 (O_487,N_24998,N_24990);
nor UO_488 (O_488,N_24931,N_24880);
or UO_489 (O_489,N_24931,N_24919);
and UO_490 (O_490,N_24811,N_24950);
or UO_491 (O_491,N_24926,N_24924);
or UO_492 (O_492,N_24823,N_24928);
nand UO_493 (O_493,N_24954,N_24912);
nand UO_494 (O_494,N_24873,N_24993);
or UO_495 (O_495,N_24914,N_24885);
nand UO_496 (O_496,N_24943,N_24910);
xor UO_497 (O_497,N_24919,N_24823);
nor UO_498 (O_498,N_24910,N_24848);
xor UO_499 (O_499,N_24948,N_24935);
nor UO_500 (O_500,N_24890,N_24845);
xnor UO_501 (O_501,N_24890,N_24819);
xor UO_502 (O_502,N_24864,N_24968);
nand UO_503 (O_503,N_24921,N_24840);
and UO_504 (O_504,N_24894,N_24931);
nor UO_505 (O_505,N_24959,N_24872);
nor UO_506 (O_506,N_24986,N_24874);
nand UO_507 (O_507,N_24997,N_24983);
nand UO_508 (O_508,N_24931,N_24930);
xor UO_509 (O_509,N_24881,N_24984);
nand UO_510 (O_510,N_24810,N_24863);
nand UO_511 (O_511,N_24926,N_24823);
or UO_512 (O_512,N_24893,N_24934);
or UO_513 (O_513,N_24891,N_24990);
and UO_514 (O_514,N_24839,N_24851);
and UO_515 (O_515,N_24854,N_24883);
and UO_516 (O_516,N_24899,N_24927);
xor UO_517 (O_517,N_24947,N_24855);
and UO_518 (O_518,N_24883,N_24920);
nor UO_519 (O_519,N_24856,N_24971);
nand UO_520 (O_520,N_24996,N_24871);
nor UO_521 (O_521,N_24921,N_24981);
or UO_522 (O_522,N_24988,N_24820);
xor UO_523 (O_523,N_24878,N_24817);
xor UO_524 (O_524,N_24926,N_24800);
or UO_525 (O_525,N_24961,N_24839);
nor UO_526 (O_526,N_24847,N_24934);
nand UO_527 (O_527,N_24884,N_24988);
and UO_528 (O_528,N_24934,N_24941);
nor UO_529 (O_529,N_24898,N_24900);
xnor UO_530 (O_530,N_24808,N_24943);
nand UO_531 (O_531,N_24939,N_24925);
or UO_532 (O_532,N_24881,N_24949);
or UO_533 (O_533,N_24834,N_24929);
nor UO_534 (O_534,N_24839,N_24809);
and UO_535 (O_535,N_24856,N_24946);
xor UO_536 (O_536,N_24854,N_24824);
xnor UO_537 (O_537,N_24934,N_24976);
nor UO_538 (O_538,N_24974,N_24921);
and UO_539 (O_539,N_24826,N_24972);
xnor UO_540 (O_540,N_24905,N_24909);
nand UO_541 (O_541,N_24971,N_24932);
and UO_542 (O_542,N_24856,N_24843);
nor UO_543 (O_543,N_24848,N_24986);
xor UO_544 (O_544,N_24828,N_24812);
nor UO_545 (O_545,N_24947,N_24925);
and UO_546 (O_546,N_24822,N_24906);
nor UO_547 (O_547,N_24859,N_24942);
nand UO_548 (O_548,N_24860,N_24846);
xor UO_549 (O_549,N_24820,N_24942);
nor UO_550 (O_550,N_24890,N_24987);
or UO_551 (O_551,N_24826,N_24864);
xor UO_552 (O_552,N_24860,N_24946);
nand UO_553 (O_553,N_24906,N_24907);
or UO_554 (O_554,N_24811,N_24815);
and UO_555 (O_555,N_24887,N_24951);
nand UO_556 (O_556,N_24933,N_24830);
nor UO_557 (O_557,N_24932,N_24950);
nand UO_558 (O_558,N_24957,N_24848);
or UO_559 (O_559,N_24877,N_24800);
or UO_560 (O_560,N_24902,N_24895);
and UO_561 (O_561,N_24811,N_24986);
or UO_562 (O_562,N_24941,N_24914);
nor UO_563 (O_563,N_24953,N_24882);
nand UO_564 (O_564,N_24809,N_24897);
nor UO_565 (O_565,N_24998,N_24920);
nor UO_566 (O_566,N_24943,N_24933);
xnor UO_567 (O_567,N_24973,N_24979);
or UO_568 (O_568,N_24918,N_24902);
and UO_569 (O_569,N_24884,N_24856);
nor UO_570 (O_570,N_24982,N_24854);
nor UO_571 (O_571,N_24835,N_24937);
xor UO_572 (O_572,N_24840,N_24898);
nand UO_573 (O_573,N_24860,N_24843);
nor UO_574 (O_574,N_24828,N_24945);
or UO_575 (O_575,N_24926,N_24831);
or UO_576 (O_576,N_24885,N_24994);
nor UO_577 (O_577,N_24923,N_24871);
nand UO_578 (O_578,N_24996,N_24864);
and UO_579 (O_579,N_24898,N_24825);
nor UO_580 (O_580,N_24917,N_24882);
nor UO_581 (O_581,N_24851,N_24825);
nand UO_582 (O_582,N_24835,N_24837);
nor UO_583 (O_583,N_24965,N_24941);
xor UO_584 (O_584,N_24992,N_24984);
xor UO_585 (O_585,N_24831,N_24984);
nor UO_586 (O_586,N_24883,N_24870);
nand UO_587 (O_587,N_24814,N_24815);
or UO_588 (O_588,N_24806,N_24918);
nor UO_589 (O_589,N_24813,N_24952);
nand UO_590 (O_590,N_24900,N_24920);
or UO_591 (O_591,N_24867,N_24851);
and UO_592 (O_592,N_24945,N_24952);
nor UO_593 (O_593,N_24826,N_24985);
nor UO_594 (O_594,N_24846,N_24956);
nor UO_595 (O_595,N_24838,N_24917);
and UO_596 (O_596,N_24831,N_24966);
and UO_597 (O_597,N_24934,N_24894);
xor UO_598 (O_598,N_24878,N_24852);
nand UO_599 (O_599,N_24801,N_24950);
xnor UO_600 (O_600,N_24844,N_24877);
nand UO_601 (O_601,N_24906,N_24864);
and UO_602 (O_602,N_24805,N_24950);
and UO_603 (O_603,N_24803,N_24850);
or UO_604 (O_604,N_24887,N_24936);
or UO_605 (O_605,N_24816,N_24971);
xor UO_606 (O_606,N_24949,N_24833);
or UO_607 (O_607,N_24945,N_24862);
or UO_608 (O_608,N_24804,N_24844);
or UO_609 (O_609,N_24956,N_24910);
nand UO_610 (O_610,N_24938,N_24823);
nand UO_611 (O_611,N_24827,N_24950);
nor UO_612 (O_612,N_24933,N_24883);
nand UO_613 (O_613,N_24865,N_24981);
or UO_614 (O_614,N_24842,N_24991);
and UO_615 (O_615,N_24913,N_24892);
or UO_616 (O_616,N_24977,N_24978);
or UO_617 (O_617,N_24801,N_24994);
xor UO_618 (O_618,N_24938,N_24964);
nand UO_619 (O_619,N_24889,N_24973);
and UO_620 (O_620,N_24911,N_24940);
or UO_621 (O_621,N_24947,N_24971);
or UO_622 (O_622,N_24905,N_24941);
xnor UO_623 (O_623,N_24826,N_24980);
nand UO_624 (O_624,N_24977,N_24987);
or UO_625 (O_625,N_24946,N_24938);
nand UO_626 (O_626,N_24869,N_24942);
or UO_627 (O_627,N_24875,N_24944);
xnor UO_628 (O_628,N_24912,N_24853);
xor UO_629 (O_629,N_24991,N_24983);
and UO_630 (O_630,N_24996,N_24832);
and UO_631 (O_631,N_24835,N_24817);
nand UO_632 (O_632,N_24923,N_24998);
or UO_633 (O_633,N_24833,N_24806);
nor UO_634 (O_634,N_24966,N_24953);
and UO_635 (O_635,N_24915,N_24958);
nor UO_636 (O_636,N_24952,N_24894);
nor UO_637 (O_637,N_24999,N_24926);
nand UO_638 (O_638,N_24924,N_24822);
nand UO_639 (O_639,N_24825,N_24927);
nand UO_640 (O_640,N_24973,N_24924);
or UO_641 (O_641,N_24879,N_24939);
nor UO_642 (O_642,N_24909,N_24872);
nand UO_643 (O_643,N_24981,N_24836);
nor UO_644 (O_644,N_24845,N_24900);
and UO_645 (O_645,N_24839,N_24830);
and UO_646 (O_646,N_24854,N_24811);
and UO_647 (O_647,N_24900,N_24903);
and UO_648 (O_648,N_24997,N_24957);
nand UO_649 (O_649,N_24840,N_24887);
and UO_650 (O_650,N_24929,N_24909);
nand UO_651 (O_651,N_24880,N_24976);
xnor UO_652 (O_652,N_24904,N_24873);
or UO_653 (O_653,N_24924,N_24943);
or UO_654 (O_654,N_24933,N_24914);
nor UO_655 (O_655,N_24886,N_24983);
or UO_656 (O_656,N_24879,N_24983);
nor UO_657 (O_657,N_24841,N_24960);
and UO_658 (O_658,N_24966,N_24825);
and UO_659 (O_659,N_24933,N_24906);
or UO_660 (O_660,N_24992,N_24961);
and UO_661 (O_661,N_24978,N_24872);
xor UO_662 (O_662,N_24888,N_24844);
nand UO_663 (O_663,N_24935,N_24937);
or UO_664 (O_664,N_24888,N_24945);
nand UO_665 (O_665,N_24878,N_24832);
xor UO_666 (O_666,N_24960,N_24893);
and UO_667 (O_667,N_24802,N_24873);
nand UO_668 (O_668,N_24863,N_24977);
xor UO_669 (O_669,N_24901,N_24890);
and UO_670 (O_670,N_24899,N_24892);
xnor UO_671 (O_671,N_24891,N_24925);
nand UO_672 (O_672,N_24934,N_24956);
xor UO_673 (O_673,N_24979,N_24996);
and UO_674 (O_674,N_24839,N_24938);
or UO_675 (O_675,N_24841,N_24930);
or UO_676 (O_676,N_24974,N_24938);
xor UO_677 (O_677,N_24935,N_24880);
or UO_678 (O_678,N_24891,N_24842);
and UO_679 (O_679,N_24948,N_24988);
nor UO_680 (O_680,N_24850,N_24819);
xor UO_681 (O_681,N_24832,N_24991);
nor UO_682 (O_682,N_24810,N_24816);
nand UO_683 (O_683,N_24986,N_24926);
nand UO_684 (O_684,N_24875,N_24928);
xnor UO_685 (O_685,N_24978,N_24873);
nand UO_686 (O_686,N_24815,N_24821);
xnor UO_687 (O_687,N_24866,N_24829);
xnor UO_688 (O_688,N_24871,N_24840);
or UO_689 (O_689,N_24936,N_24886);
nand UO_690 (O_690,N_24831,N_24917);
or UO_691 (O_691,N_24915,N_24859);
and UO_692 (O_692,N_24900,N_24818);
xnor UO_693 (O_693,N_24883,N_24939);
nor UO_694 (O_694,N_24909,N_24953);
xor UO_695 (O_695,N_24869,N_24825);
and UO_696 (O_696,N_24802,N_24880);
and UO_697 (O_697,N_24940,N_24981);
and UO_698 (O_698,N_24853,N_24887);
nor UO_699 (O_699,N_24977,N_24985);
and UO_700 (O_700,N_24910,N_24880);
nor UO_701 (O_701,N_24812,N_24876);
xor UO_702 (O_702,N_24882,N_24833);
nand UO_703 (O_703,N_24912,N_24916);
or UO_704 (O_704,N_24907,N_24891);
xnor UO_705 (O_705,N_24859,N_24801);
nor UO_706 (O_706,N_24979,N_24911);
and UO_707 (O_707,N_24811,N_24826);
or UO_708 (O_708,N_24973,N_24880);
nand UO_709 (O_709,N_24944,N_24982);
and UO_710 (O_710,N_24831,N_24902);
xor UO_711 (O_711,N_24887,N_24802);
or UO_712 (O_712,N_24997,N_24886);
and UO_713 (O_713,N_24855,N_24963);
or UO_714 (O_714,N_24807,N_24975);
or UO_715 (O_715,N_24806,N_24965);
nor UO_716 (O_716,N_24802,N_24870);
or UO_717 (O_717,N_24925,N_24873);
or UO_718 (O_718,N_24863,N_24927);
nand UO_719 (O_719,N_24880,N_24984);
nand UO_720 (O_720,N_24847,N_24927);
or UO_721 (O_721,N_24890,N_24850);
and UO_722 (O_722,N_24923,N_24847);
and UO_723 (O_723,N_24867,N_24910);
or UO_724 (O_724,N_24913,N_24900);
nor UO_725 (O_725,N_24979,N_24831);
nand UO_726 (O_726,N_24976,N_24943);
nor UO_727 (O_727,N_24909,N_24837);
nand UO_728 (O_728,N_24998,N_24978);
or UO_729 (O_729,N_24909,N_24908);
xor UO_730 (O_730,N_24850,N_24979);
or UO_731 (O_731,N_24898,N_24896);
and UO_732 (O_732,N_24909,N_24917);
nor UO_733 (O_733,N_24970,N_24991);
nor UO_734 (O_734,N_24949,N_24892);
or UO_735 (O_735,N_24871,N_24932);
xnor UO_736 (O_736,N_24874,N_24910);
xnor UO_737 (O_737,N_24812,N_24836);
xnor UO_738 (O_738,N_24820,N_24896);
nand UO_739 (O_739,N_24917,N_24839);
and UO_740 (O_740,N_24898,N_24905);
xor UO_741 (O_741,N_24860,N_24851);
xnor UO_742 (O_742,N_24900,N_24941);
or UO_743 (O_743,N_24845,N_24852);
and UO_744 (O_744,N_24835,N_24946);
and UO_745 (O_745,N_24875,N_24858);
or UO_746 (O_746,N_24955,N_24887);
and UO_747 (O_747,N_24848,N_24970);
nand UO_748 (O_748,N_24985,N_24875);
nor UO_749 (O_749,N_24841,N_24892);
or UO_750 (O_750,N_24851,N_24832);
nand UO_751 (O_751,N_24840,N_24962);
or UO_752 (O_752,N_24919,N_24848);
nor UO_753 (O_753,N_24823,N_24840);
and UO_754 (O_754,N_24897,N_24906);
xnor UO_755 (O_755,N_24854,N_24931);
nor UO_756 (O_756,N_24849,N_24822);
xnor UO_757 (O_757,N_24878,N_24816);
or UO_758 (O_758,N_24818,N_24920);
or UO_759 (O_759,N_24923,N_24972);
or UO_760 (O_760,N_24825,N_24937);
nand UO_761 (O_761,N_24917,N_24856);
or UO_762 (O_762,N_24824,N_24989);
and UO_763 (O_763,N_24984,N_24980);
nand UO_764 (O_764,N_24927,N_24905);
nor UO_765 (O_765,N_24876,N_24914);
nor UO_766 (O_766,N_24812,N_24859);
nor UO_767 (O_767,N_24844,N_24987);
nand UO_768 (O_768,N_24915,N_24960);
or UO_769 (O_769,N_24918,N_24881);
and UO_770 (O_770,N_24895,N_24815);
nand UO_771 (O_771,N_24927,N_24900);
and UO_772 (O_772,N_24887,N_24922);
or UO_773 (O_773,N_24800,N_24991);
nand UO_774 (O_774,N_24954,N_24949);
xnor UO_775 (O_775,N_24953,N_24945);
xor UO_776 (O_776,N_24892,N_24882);
and UO_777 (O_777,N_24995,N_24844);
nand UO_778 (O_778,N_24967,N_24898);
nor UO_779 (O_779,N_24808,N_24871);
xnor UO_780 (O_780,N_24925,N_24874);
and UO_781 (O_781,N_24831,N_24801);
xor UO_782 (O_782,N_24807,N_24942);
xor UO_783 (O_783,N_24855,N_24989);
nand UO_784 (O_784,N_24818,N_24860);
or UO_785 (O_785,N_24874,N_24871);
xnor UO_786 (O_786,N_24923,N_24813);
or UO_787 (O_787,N_24894,N_24811);
xor UO_788 (O_788,N_24992,N_24878);
xor UO_789 (O_789,N_24936,N_24921);
xor UO_790 (O_790,N_24818,N_24967);
and UO_791 (O_791,N_24981,N_24999);
nor UO_792 (O_792,N_24800,N_24928);
and UO_793 (O_793,N_24905,N_24966);
and UO_794 (O_794,N_24873,N_24936);
nand UO_795 (O_795,N_24818,N_24848);
or UO_796 (O_796,N_24901,N_24935);
xor UO_797 (O_797,N_24971,N_24861);
xnor UO_798 (O_798,N_24913,N_24925);
or UO_799 (O_799,N_24955,N_24847);
nand UO_800 (O_800,N_24927,N_24932);
or UO_801 (O_801,N_24887,N_24983);
and UO_802 (O_802,N_24928,N_24811);
nand UO_803 (O_803,N_24811,N_24904);
nor UO_804 (O_804,N_24967,N_24920);
and UO_805 (O_805,N_24804,N_24942);
and UO_806 (O_806,N_24831,N_24830);
nand UO_807 (O_807,N_24826,N_24923);
xnor UO_808 (O_808,N_24952,N_24833);
and UO_809 (O_809,N_24884,N_24834);
nor UO_810 (O_810,N_24861,N_24815);
xnor UO_811 (O_811,N_24982,N_24947);
nand UO_812 (O_812,N_24837,N_24890);
nand UO_813 (O_813,N_24861,N_24914);
nand UO_814 (O_814,N_24826,N_24994);
or UO_815 (O_815,N_24914,N_24917);
or UO_816 (O_816,N_24981,N_24953);
or UO_817 (O_817,N_24817,N_24833);
and UO_818 (O_818,N_24802,N_24811);
and UO_819 (O_819,N_24908,N_24947);
and UO_820 (O_820,N_24863,N_24806);
nor UO_821 (O_821,N_24852,N_24962);
and UO_822 (O_822,N_24840,N_24806);
xor UO_823 (O_823,N_24942,N_24991);
xnor UO_824 (O_824,N_24970,N_24961);
or UO_825 (O_825,N_24890,N_24802);
or UO_826 (O_826,N_24991,N_24893);
nor UO_827 (O_827,N_24904,N_24887);
or UO_828 (O_828,N_24834,N_24874);
nor UO_829 (O_829,N_24844,N_24993);
xor UO_830 (O_830,N_24843,N_24967);
xnor UO_831 (O_831,N_24852,N_24865);
nor UO_832 (O_832,N_24955,N_24867);
xor UO_833 (O_833,N_24898,N_24858);
and UO_834 (O_834,N_24907,N_24841);
xor UO_835 (O_835,N_24816,N_24818);
and UO_836 (O_836,N_24925,N_24970);
xor UO_837 (O_837,N_24805,N_24910);
xnor UO_838 (O_838,N_24928,N_24971);
and UO_839 (O_839,N_24823,N_24989);
xnor UO_840 (O_840,N_24875,N_24963);
xor UO_841 (O_841,N_24938,N_24942);
and UO_842 (O_842,N_24906,N_24954);
nand UO_843 (O_843,N_24905,N_24895);
or UO_844 (O_844,N_24965,N_24807);
nor UO_845 (O_845,N_24981,N_24980);
or UO_846 (O_846,N_24816,N_24917);
nor UO_847 (O_847,N_24991,N_24926);
or UO_848 (O_848,N_24945,N_24928);
or UO_849 (O_849,N_24930,N_24952);
or UO_850 (O_850,N_24918,N_24815);
nand UO_851 (O_851,N_24833,N_24931);
and UO_852 (O_852,N_24993,N_24935);
and UO_853 (O_853,N_24894,N_24928);
nor UO_854 (O_854,N_24850,N_24940);
xor UO_855 (O_855,N_24872,N_24967);
nor UO_856 (O_856,N_24924,N_24999);
xor UO_857 (O_857,N_24816,N_24866);
nand UO_858 (O_858,N_24846,N_24916);
nand UO_859 (O_859,N_24843,N_24928);
or UO_860 (O_860,N_24834,N_24858);
or UO_861 (O_861,N_24878,N_24928);
nor UO_862 (O_862,N_24817,N_24987);
xor UO_863 (O_863,N_24893,N_24993);
xnor UO_864 (O_864,N_24997,N_24981);
nor UO_865 (O_865,N_24906,N_24826);
nor UO_866 (O_866,N_24852,N_24949);
xor UO_867 (O_867,N_24998,N_24910);
or UO_868 (O_868,N_24870,N_24876);
and UO_869 (O_869,N_24920,N_24806);
nor UO_870 (O_870,N_24973,N_24895);
nand UO_871 (O_871,N_24842,N_24870);
and UO_872 (O_872,N_24952,N_24834);
xor UO_873 (O_873,N_24908,N_24826);
nor UO_874 (O_874,N_24850,N_24918);
or UO_875 (O_875,N_24953,N_24922);
nand UO_876 (O_876,N_24900,N_24999);
nand UO_877 (O_877,N_24978,N_24940);
nor UO_878 (O_878,N_24960,N_24838);
nand UO_879 (O_879,N_24961,N_24860);
xor UO_880 (O_880,N_24930,N_24855);
xnor UO_881 (O_881,N_24940,N_24815);
nand UO_882 (O_882,N_24974,N_24843);
nor UO_883 (O_883,N_24848,N_24974);
nor UO_884 (O_884,N_24866,N_24922);
or UO_885 (O_885,N_24971,N_24984);
nand UO_886 (O_886,N_24892,N_24957);
and UO_887 (O_887,N_24925,N_24858);
nand UO_888 (O_888,N_24949,N_24889);
nor UO_889 (O_889,N_24905,N_24946);
nor UO_890 (O_890,N_24800,N_24969);
nor UO_891 (O_891,N_24834,N_24953);
and UO_892 (O_892,N_24952,N_24814);
or UO_893 (O_893,N_24917,N_24886);
nor UO_894 (O_894,N_24912,N_24854);
nor UO_895 (O_895,N_24823,N_24937);
or UO_896 (O_896,N_24922,N_24909);
and UO_897 (O_897,N_24980,N_24880);
nand UO_898 (O_898,N_24853,N_24859);
or UO_899 (O_899,N_24818,N_24995);
or UO_900 (O_900,N_24994,N_24903);
and UO_901 (O_901,N_24867,N_24865);
or UO_902 (O_902,N_24887,N_24804);
nand UO_903 (O_903,N_24850,N_24965);
xnor UO_904 (O_904,N_24986,N_24870);
nand UO_905 (O_905,N_24833,N_24948);
and UO_906 (O_906,N_24805,N_24925);
nand UO_907 (O_907,N_24926,N_24966);
xnor UO_908 (O_908,N_24834,N_24949);
and UO_909 (O_909,N_24827,N_24826);
xnor UO_910 (O_910,N_24819,N_24964);
xnor UO_911 (O_911,N_24852,N_24816);
xor UO_912 (O_912,N_24841,N_24912);
xnor UO_913 (O_913,N_24827,N_24803);
or UO_914 (O_914,N_24839,N_24853);
or UO_915 (O_915,N_24922,N_24852);
and UO_916 (O_916,N_24904,N_24884);
xor UO_917 (O_917,N_24894,N_24814);
xor UO_918 (O_918,N_24881,N_24931);
xnor UO_919 (O_919,N_24963,N_24950);
nor UO_920 (O_920,N_24933,N_24952);
xnor UO_921 (O_921,N_24942,N_24851);
or UO_922 (O_922,N_24877,N_24810);
nand UO_923 (O_923,N_24879,N_24953);
nand UO_924 (O_924,N_24828,N_24856);
nand UO_925 (O_925,N_24824,N_24980);
or UO_926 (O_926,N_24858,N_24982);
or UO_927 (O_927,N_24921,N_24823);
and UO_928 (O_928,N_24965,N_24978);
xor UO_929 (O_929,N_24897,N_24992);
and UO_930 (O_930,N_24820,N_24986);
xnor UO_931 (O_931,N_24853,N_24814);
xor UO_932 (O_932,N_24854,N_24896);
nor UO_933 (O_933,N_24830,N_24804);
nand UO_934 (O_934,N_24895,N_24873);
nand UO_935 (O_935,N_24954,N_24997);
nor UO_936 (O_936,N_24883,N_24813);
and UO_937 (O_937,N_24844,N_24895);
nor UO_938 (O_938,N_24959,N_24851);
nand UO_939 (O_939,N_24956,N_24907);
nand UO_940 (O_940,N_24840,N_24919);
and UO_941 (O_941,N_24925,N_24926);
xnor UO_942 (O_942,N_24925,N_24897);
nor UO_943 (O_943,N_24900,N_24986);
and UO_944 (O_944,N_24868,N_24854);
xor UO_945 (O_945,N_24933,N_24911);
nor UO_946 (O_946,N_24809,N_24924);
and UO_947 (O_947,N_24829,N_24869);
nor UO_948 (O_948,N_24811,N_24865);
xnor UO_949 (O_949,N_24964,N_24811);
and UO_950 (O_950,N_24977,N_24859);
and UO_951 (O_951,N_24907,N_24843);
nand UO_952 (O_952,N_24830,N_24862);
nor UO_953 (O_953,N_24951,N_24913);
xor UO_954 (O_954,N_24824,N_24846);
and UO_955 (O_955,N_24817,N_24873);
xnor UO_956 (O_956,N_24852,N_24974);
or UO_957 (O_957,N_24930,N_24848);
or UO_958 (O_958,N_24823,N_24970);
and UO_959 (O_959,N_24988,N_24938);
nand UO_960 (O_960,N_24903,N_24978);
nor UO_961 (O_961,N_24879,N_24884);
xnor UO_962 (O_962,N_24936,N_24864);
or UO_963 (O_963,N_24865,N_24909);
xor UO_964 (O_964,N_24808,N_24901);
nor UO_965 (O_965,N_24830,N_24915);
nor UO_966 (O_966,N_24841,N_24844);
nor UO_967 (O_967,N_24936,N_24915);
xor UO_968 (O_968,N_24974,N_24809);
nand UO_969 (O_969,N_24990,N_24818);
or UO_970 (O_970,N_24800,N_24871);
xor UO_971 (O_971,N_24903,N_24986);
nand UO_972 (O_972,N_24879,N_24883);
or UO_973 (O_973,N_24960,N_24806);
nand UO_974 (O_974,N_24843,N_24906);
nand UO_975 (O_975,N_24886,N_24957);
xor UO_976 (O_976,N_24990,N_24900);
and UO_977 (O_977,N_24866,N_24839);
nor UO_978 (O_978,N_24808,N_24926);
and UO_979 (O_979,N_24889,N_24956);
nor UO_980 (O_980,N_24918,N_24811);
or UO_981 (O_981,N_24923,N_24986);
nand UO_982 (O_982,N_24884,N_24994);
nor UO_983 (O_983,N_24843,N_24886);
and UO_984 (O_984,N_24814,N_24930);
nand UO_985 (O_985,N_24885,N_24801);
and UO_986 (O_986,N_24997,N_24819);
xor UO_987 (O_987,N_24849,N_24882);
xnor UO_988 (O_988,N_24871,N_24878);
xnor UO_989 (O_989,N_24868,N_24876);
and UO_990 (O_990,N_24981,N_24824);
nor UO_991 (O_991,N_24937,N_24967);
or UO_992 (O_992,N_24916,N_24809);
or UO_993 (O_993,N_24901,N_24978);
and UO_994 (O_994,N_24846,N_24841);
nor UO_995 (O_995,N_24932,N_24812);
nand UO_996 (O_996,N_24876,N_24978);
or UO_997 (O_997,N_24991,N_24838);
or UO_998 (O_998,N_24971,N_24840);
nand UO_999 (O_999,N_24920,N_24866);
nor UO_1000 (O_1000,N_24918,N_24972);
and UO_1001 (O_1001,N_24821,N_24802);
and UO_1002 (O_1002,N_24965,N_24916);
and UO_1003 (O_1003,N_24951,N_24910);
xor UO_1004 (O_1004,N_24835,N_24892);
nand UO_1005 (O_1005,N_24999,N_24950);
or UO_1006 (O_1006,N_24920,N_24830);
nand UO_1007 (O_1007,N_24864,N_24835);
nand UO_1008 (O_1008,N_24861,N_24822);
xor UO_1009 (O_1009,N_24852,N_24835);
xnor UO_1010 (O_1010,N_24940,N_24830);
nand UO_1011 (O_1011,N_24905,N_24818);
xor UO_1012 (O_1012,N_24832,N_24951);
xnor UO_1013 (O_1013,N_24987,N_24813);
xnor UO_1014 (O_1014,N_24947,N_24865);
or UO_1015 (O_1015,N_24994,N_24971);
and UO_1016 (O_1016,N_24871,N_24895);
nor UO_1017 (O_1017,N_24886,N_24849);
and UO_1018 (O_1018,N_24850,N_24947);
nor UO_1019 (O_1019,N_24895,N_24961);
xnor UO_1020 (O_1020,N_24986,N_24818);
xnor UO_1021 (O_1021,N_24888,N_24904);
xnor UO_1022 (O_1022,N_24890,N_24904);
and UO_1023 (O_1023,N_24922,N_24802);
and UO_1024 (O_1024,N_24905,N_24987);
and UO_1025 (O_1025,N_24834,N_24864);
nand UO_1026 (O_1026,N_24993,N_24849);
nor UO_1027 (O_1027,N_24943,N_24903);
and UO_1028 (O_1028,N_24978,N_24890);
and UO_1029 (O_1029,N_24847,N_24991);
xor UO_1030 (O_1030,N_24815,N_24822);
nor UO_1031 (O_1031,N_24905,N_24867);
nand UO_1032 (O_1032,N_24987,N_24815);
nand UO_1033 (O_1033,N_24863,N_24931);
and UO_1034 (O_1034,N_24965,N_24954);
xor UO_1035 (O_1035,N_24981,N_24895);
nand UO_1036 (O_1036,N_24927,N_24936);
or UO_1037 (O_1037,N_24813,N_24985);
and UO_1038 (O_1038,N_24957,N_24971);
xor UO_1039 (O_1039,N_24842,N_24996);
or UO_1040 (O_1040,N_24880,N_24967);
and UO_1041 (O_1041,N_24838,N_24873);
nand UO_1042 (O_1042,N_24820,N_24968);
xnor UO_1043 (O_1043,N_24946,N_24816);
or UO_1044 (O_1044,N_24935,N_24820);
xor UO_1045 (O_1045,N_24885,N_24903);
and UO_1046 (O_1046,N_24944,N_24992);
and UO_1047 (O_1047,N_24850,N_24981);
or UO_1048 (O_1048,N_24839,N_24829);
or UO_1049 (O_1049,N_24823,N_24950);
xor UO_1050 (O_1050,N_24988,N_24907);
or UO_1051 (O_1051,N_24997,N_24900);
and UO_1052 (O_1052,N_24842,N_24942);
and UO_1053 (O_1053,N_24958,N_24860);
xor UO_1054 (O_1054,N_24851,N_24993);
xor UO_1055 (O_1055,N_24895,N_24899);
or UO_1056 (O_1056,N_24977,N_24941);
or UO_1057 (O_1057,N_24911,N_24881);
and UO_1058 (O_1058,N_24972,N_24883);
or UO_1059 (O_1059,N_24981,N_24843);
and UO_1060 (O_1060,N_24812,N_24850);
xor UO_1061 (O_1061,N_24837,N_24815);
nor UO_1062 (O_1062,N_24871,N_24804);
nand UO_1063 (O_1063,N_24942,N_24855);
nor UO_1064 (O_1064,N_24962,N_24961);
nand UO_1065 (O_1065,N_24867,N_24984);
and UO_1066 (O_1066,N_24992,N_24890);
and UO_1067 (O_1067,N_24868,N_24958);
nand UO_1068 (O_1068,N_24856,N_24912);
and UO_1069 (O_1069,N_24819,N_24897);
xnor UO_1070 (O_1070,N_24897,N_24998);
nor UO_1071 (O_1071,N_24917,N_24934);
nand UO_1072 (O_1072,N_24950,N_24922);
or UO_1073 (O_1073,N_24851,N_24980);
and UO_1074 (O_1074,N_24895,N_24993);
xnor UO_1075 (O_1075,N_24886,N_24972);
xnor UO_1076 (O_1076,N_24958,N_24938);
xor UO_1077 (O_1077,N_24961,N_24936);
xor UO_1078 (O_1078,N_24831,N_24919);
and UO_1079 (O_1079,N_24929,N_24978);
and UO_1080 (O_1080,N_24993,N_24807);
nor UO_1081 (O_1081,N_24956,N_24901);
xnor UO_1082 (O_1082,N_24897,N_24831);
nand UO_1083 (O_1083,N_24840,N_24878);
xor UO_1084 (O_1084,N_24853,N_24961);
nor UO_1085 (O_1085,N_24871,N_24841);
nand UO_1086 (O_1086,N_24953,N_24855);
and UO_1087 (O_1087,N_24839,N_24823);
or UO_1088 (O_1088,N_24862,N_24952);
nor UO_1089 (O_1089,N_24926,N_24844);
or UO_1090 (O_1090,N_24813,N_24887);
and UO_1091 (O_1091,N_24941,N_24819);
or UO_1092 (O_1092,N_24842,N_24896);
and UO_1093 (O_1093,N_24887,N_24926);
xor UO_1094 (O_1094,N_24887,N_24915);
or UO_1095 (O_1095,N_24884,N_24957);
or UO_1096 (O_1096,N_24820,N_24841);
xnor UO_1097 (O_1097,N_24892,N_24944);
and UO_1098 (O_1098,N_24975,N_24849);
nor UO_1099 (O_1099,N_24984,N_24918);
and UO_1100 (O_1100,N_24838,N_24867);
nand UO_1101 (O_1101,N_24837,N_24880);
nor UO_1102 (O_1102,N_24981,N_24916);
or UO_1103 (O_1103,N_24813,N_24978);
xnor UO_1104 (O_1104,N_24946,N_24943);
and UO_1105 (O_1105,N_24929,N_24845);
or UO_1106 (O_1106,N_24968,N_24970);
and UO_1107 (O_1107,N_24851,N_24915);
or UO_1108 (O_1108,N_24991,N_24997);
xnor UO_1109 (O_1109,N_24900,N_24812);
and UO_1110 (O_1110,N_24859,N_24928);
nand UO_1111 (O_1111,N_24845,N_24918);
xnor UO_1112 (O_1112,N_24834,N_24954);
and UO_1113 (O_1113,N_24878,N_24951);
nor UO_1114 (O_1114,N_24895,N_24965);
and UO_1115 (O_1115,N_24895,N_24928);
xor UO_1116 (O_1116,N_24911,N_24896);
nor UO_1117 (O_1117,N_24859,N_24959);
or UO_1118 (O_1118,N_24940,N_24917);
xnor UO_1119 (O_1119,N_24982,N_24920);
nor UO_1120 (O_1120,N_24807,N_24948);
xor UO_1121 (O_1121,N_24906,N_24938);
xor UO_1122 (O_1122,N_24850,N_24988);
nand UO_1123 (O_1123,N_24938,N_24887);
or UO_1124 (O_1124,N_24871,N_24823);
or UO_1125 (O_1125,N_24842,N_24841);
xor UO_1126 (O_1126,N_24825,N_24818);
xnor UO_1127 (O_1127,N_24892,N_24875);
and UO_1128 (O_1128,N_24976,N_24820);
nor UO_1129 (O_1129,N_24909,N_24840);
nor UO_1130 (O_1130,N_24862,N_24932);
nand UO_1131 (O_1131,N_24958,N_24939);
xnor UO_1132 (O_1132,N_24948,N_24816);
nor UO_1133 (O_1133,N_24868,N_24899);
nor UO_1134 (O_1134,N_24832,N_24807);
nand UO_1135 (O_1135,N_24856,N_24830);
and UO_1136 (O_1136,N_24826,N_24893);
nand UO_1137 (O_1137,N_24908,N_24846);
nor UO_1138 (O_1138,N_24920,N_24973);
nand UO_1139 (O_1139,N_24874,N_24920);
and UO_1140 (O_1140,N_24840,N_24819);
xor UO_1141 (O_1141,N_24832,N_24821);
nor UO_1142 (O_1142,N_24996,N_24867);
or UO_1143 (O_1143,N_24815,N_24849);
nor UO_1144 (O_1144,N_24905,N_24924);
xnor UO_1145 (O_1145,N_24810,N_24909);
nor UO_1146 (O_1146,N_24917,N_24875);
or UO_1147 (O_1147,N_24824,N_24804);
or UO_1148 (O_1148,N_24867,N_24962);
or UO_1149 (O_1149,N_24918,N_24801);
xor UO_1150 (O_1150,N_24825,N_24823);
or UO_1151 (O_1151,N_24996,N_24857);
nor UO_1152 (O_1152,N_24893,N_24856);
nand UO_1153 (O_1153,N_24898,N_24875);
or UO_1154 (O_1154,N_24879,N_24970);
xor UO_1155 (O_1155,N_24971,N_24833);
nand UO_1156 (O_1156,N_24846,N_24812);
nor UO_1157 (O_1157,N_24930,N_24933);
or UO_1158 (O_1158,N_24970,N_24902);
xnor UO_1159 (O_1159,N_24975,N_24973);
and UO_1160 (O_1160,N_24960,N_24955);
nor UO_1161 (O_1161,N_24954,N_24953);
or UO_1162 (O_1162,N_24875,N_24941);
and UO_1163 (O_1163,N_24995,N_24975);
nor UO_1164 (O_1164,N_24927,N_24964);
nor UO_1165 (O_1165,N_24856,N_24986);
and UO_1166 (O_1166,N_24833,N_24962);
and UO_1167 (O_1167,N_24850,N_24892);
xor UO_1168 (O_1168,N_24823,N_24822);
nand UO_1169 (O_1169,N_24839,N_24826);
xnor UO_1170 (O_1170,N_24994,N_24808);
nand UO_1171 (O_1171,N_24850,N_24809);
or UO_1172 (O_1172,N_24844,N_24974);
and UO_1173 (O_1173,N_24940,N_24958);
nand UO_1174 (O_1174,N_24818,N_24962);
nand UO_1175 (O_1175,N_24854,N_24964);
nand UO_1176 (O_1176,N_24854,N_24989);
nor UO_1177 (O_1177,N_24838,N_24819);
xor UO_1178 (O_1178,N_24943,N_24922);
xor UO_1179 (O_1179,N_24945,N_24910);
or UO_1180 (O_1180,N_24801,N_24872);
nand UO_1181 (O_1181,N_24931,N_24862);
nor UO_1182 (O_1182,N_24830,N_24849);
nor UO_1183 (O_1183,N_24910,N_24898);
or UO_1184 (O_1184,N_24935,N_24998);
and UO_1185 (O_1185,N_24863,N_24964);
nor UO_1186 (O_1186,N_24951,N_24930);
and UO_1187 (O_1187,N_24989,N_24813);
or UO_1188 (O_1188,N_24840,N_24892);
and UO_1189 (O_1189,N_24802,N_24923);
xor UO_1190 (O_1190,N_24977,N_24900);
nand UO_1191 (O_1191,N_24875,N_24986);
or UO_1192 (O_1192,N_24907,N_24858);
xor UO_1193 (O_1193,N_24865,N_24952);
and UO_1194 (O_1194,N_24955,N_24972);
xor UO_1195 (O_1195,N_24877,N_24926);
nor UO_1196 (O_1196,N_24939,N_24960);
nand UO_1197 (O_1197,N_24848,N_24935);
nor UO_1198 (O_1198,N_24849,N_24916);
nand UO_1199 (O_1199,N_24858,N_24915);
or UO_1200 (O_1200,N_24969,N_24925);
nand UO_1201 (O_1201,N_24859,N_24930);
and UO_1202 (O_1202,N_24987,N_24955);
nand UO_1203 (O_1203,N_24936,N_24960);
or UO_1204 (O_1204,N_24842,N_24815);
and UO_1205 (O_1205,N_24805,N_24802);
xnor UO_1206 (O_1206,N_24829,N_24945);
and UO_1207 (O_1207,N_24896,N_24876);
and UO_1208 (O_1208,N_24895,N_24988);
nand UO_1209 (O_1209,N_24859,N_24913);
nand UO_1210 (O_1210,N_24870,N_24931);
nor UO_1211 (O_1211,N_24815,N_24979);
nand UO_1212 (O_1212,N_24926,N_24836);
and UO_1213 (O_1213,N_24816,N_24831);
nand UO_1214 (O_1214,N_24983,N_24842);
or UO_1215 (O_1215,N_24991,N_24930);
nor UO_1216 (O_1216,N_24951,N_24926);
or UO_1217 (O_1217,N_24964,N_24835);
or UO_1218 (O_1218,N_24902,N_24965);
nor UO_1219 (O_1219,N_24989,N_24827);
xor UO_1220 (O_1220,N_24852,N_24822);
and UO_1221 (O_1221,N_24998,N_24885);
nand UO_1222 (O_1222,N_24802,N_24905);
or UO_1223 (O_1223,N_24827,N_24805);
nor UO_1224 (O_1224,N_24880,N_24856);
xnor UO_1225 (O_1225,N_24831,N_24804);
nand UO_1226 (O_1226,N_24943,N_24972);
nor UO_1227 (O_1227,N_24982,N_24809);
nand UO_1228 (O_1228,N_24804,N_24899);
nand UO_1229 (O_1229,N_24889,N_24863);
nor UO_1230 (O_1230,N_24826,N_24943);
nand UO_1231 (O_1231,N_24997,N_24874);
nor UO_1232 (O_1232,N_24877,N_24801);
and UO_1233 (O_1233,N_24958,N_24804);
and UO_1234 (O_1234,N_24997,N_24840);
or UO_1235 (O_1235,N_24815,N_24912);
or UO_1236 (O_1236,N_24981,N_24986);
nand UO_1237 (O_1237,N_24995,N_24880);
nor UO_1238 (O_1238,N_24978,N_24860);
and UO_1239 (O_1239,N_24895,N_24999);
and UO_1240 (O_1240,N_24817,N_24843);
nand UO_1241 (O_1241,N_24959,N_24828);
and UO_1242 (O_1242,N_24847,N_24911);
and UO_1243 (O_1243,N_24818,N_24941);
xnor UO_1244 (O_1244,N_24830,N_24909);
nor UO_1245 (O_1245,N_24958,N_24816);
nor UO_1246 (O_1246,N_24866,N_24962);
and UO_1247 (O_1247,N_24819,N_24873);
xor UO_1248 (O_1248,N_24925,N_24811);
nor UO_1249 (O_1249,N_24860,N_24927);
and UO_1250 (O_1250,N_24956,N_24818);
nor UO_1251 (O_1251,N_24879,N_24918);
and UO_1252 (O_1252,N_24968,N_24916);
nor UO_1253 (O_1253,N_24802,N_24828);
or UO_1254 (O_1254,N_24833,N_24887);
nand UO_1255 (O_1255,N_24855,N_24987);
xnor UO_1256 (O_1256,N_24863,N_24920);
nand UO_1257 (O_1257,N_24862,N_24852);
or UO_1258 (O_1258,N_24839,N_24834);
xnor UO_1259 (O_1259,N_24938,N_24801);
xor UO_1260 (O_1260,N_24855,N_24840);
xor UO_1261 (O_1261,N_24866,N_24855);
nand UO_1262 (O_1262,N_24850,N_24810);
xnor UO_1263 (O_1263,N_24878,N_24869);
or UO_1264 (O_1264,N_24876,N_24969);
nor UO_1265 (O_1265,N_24812,N_24942);
nand UO_1266 (O_1266,N_24830,N_24894);
and UO_1267 (O_1267,N_24984,N_24840);
or UO_1268 (O_1268,N_24899,N_24909);
nand UO_1269 (O_1269,N_24818,N_24899);
nand UO_1270 (O_1270,N_24830,N_24885);
and UO_1271 (O_1271,N_24869,N_24836);
nor UO_1272 (O_1272,N_24916,N_24997);
nand UO_1273 (O_1273,N_24873,N_24866);
xnor UO_1274 (O_1274,N_24979,N_24823);
xor UO_1275 (O_1275,N_24972,N_24953);
xnor UO_1276 (O_1276,N_24805,N_24858);
nor UO_1277 (O_1277,N_24802,N_24846);
nor UO_1278 (O_1278,N_24898,N_24941);
nor UO_1279 (O_1279,N_24812,N_24977);
or UO_1280 (O_1280,N_24914,N_24902);
or UO_1281 (O_1281,N_24951,N_24940);
nand UO_1282 (O_1282,N_24831,N_24808);
xnor UO_1283 (O_1283,N_24880,N_24846);
xor UO_1284 (O_1284,N_24997,N_24808);
and UO_1285 (O_1285,N_24947,N_24883);
or UO_1286 (O_1286,N_24996,N_24846);
or UO_1287 (O_1287,N_24871,N_24941);
nor UO_1288 (O_1288,N_24873,N_24989);
and UO_1289 (O_1289,N_24991,N_24820);
xnor UO_1290 (O_1290,N_24941,N_24858);
or UO_1291 (O_1291,N_24819,N_24938);
nor UO_1292 (O_1292,N_24813,N_24840);
nor UO_1293 (O_1293,N_24988,N_24848);
xnor UO_1294 (O_1294,N_24993,N_24826);
and UO_1295 (O_1295,N_24999,N_24978);
nor UO_1296 (O_1296,N_24805,N_24831);
and UO_1297 (O_1297,N_24934,N_24944);
nor UO_1298 (O_1298,N_24891,N_24813);
nor UO_1299 (O_1299,N_24834,N_24939);
or UO_1300 (O_1300,N_24842,N_24848);
or UO_1301 (O_1301,N_24809,N_24955);
or UO_1302 (O_1302,N_24973,N_24829);
nand UO_1303 (O_1303,N_24883,N_24867);
nor UO_1304 (O_1304,N_24973,N_24926);
xnor UO_1305 (O_1305,N_24844,N_24915);
xnor UO_1306 (O_1306,N_24912,N_24836);
xor UO_1307 (O_1307,N_24955,N_24820);
nand UO_1308 (O_1308,N_24925,N_24951);
xnor UO_1309 (O_1309,N_24979,N_24809);
nor UO_1310 (O_1310,N_24962,N_24941);
or UO_1311 (O_1311,N_24970,N_24867);
or UO_1312 (O_1312,N_24887,N_24959);
nand UO_1313 (O_1313,N_24908,N_24885);
or UO_1314 (O_1314,N_24997,N_24920);
or UO_1315 (O_1315,N_24970,N_24952);
or UO_1316 (O_1316,N_24961,N_24912);
nand UO_1317 (O_1317,N_24855,N_24937);
and UO_1318 (O_1318,N_24831,N_24997);
xor UO_1319 (O_1319,N_24966,N_24918);
or UO_1320 (O_1320,N_24907,N_24945);
and UO_1321 (O_1321,N_24981,N_24933);
xnor UO_1322 (O_1322,N_24976,N_24878);
xnor UO_1323 (O_1323,N_24933,N_24935);
nand UO_1324 (O_1324,N_24828,N_24891);
and UO_1325 (O_1325,N_24825,N_24848);
nand UO_1326 (O_1326,N_24816,N_24999);
nor UO_1327 (O_1327,N_24943,N_24897);
nor UO_1328 (O_1328,N_24824,N_24933);
xor UO_1329 (O_1329,N_24833,N_24901);
xor UO_1330 (O_1330,N_24883,N_24838);
and UO_1331 (O_1331,N_24844,N_24882);
and UO_1332 (O_1332,N_24975,N_24991);
nor UO_1333 (O_1333,N_24907,N_24993);
xor UO_1334 (O_1334,N_24885,N_24839);
and UO_1335 (O_1335,N_24872,N_24855);
nor UO_1336 (O_1336,N_24871,N_24931);
xor UO_1337 (O_1337,N_24863,N_24963);
and UO_1338 (O_1338,N_24885,N_24812);
nand UO_1339 (O_1339,N_24876,N_24861);
nand UO_1340 (O_1340,N_24841,N_24937);
xnor UO_1341 (O_1341,N_24928,N_24850);
xnor UO_1342 (O_1342,N_24993,N_24808);
xor UO_1343 (O_1343,N_24885,N_24968);
nor UO_1344 (O_1344,N_24954,N_24990);
xor UO_1345 (O_1345,N_24888,N_24833);
nand UO_1346 (O_1346,N_24875,N_24829);
nor UO_1347 (O_1347,N_24930,N_24965);
xnor UO_1348 (O_1348,N_24997,N_24973);
xor UO_1349 (O_1349,N_24800,N_24837);
nor UO_1350 (O_1350,N_24823,N_24940);
and UO_1351 (O_1351,N_24841,N_24829);
and UO_1352 (O_1352,N_24856,N_24962);
nor UO_1353 (O_1353,N_24945,N_24884);
xnor UO_1354 (O_1354,N_24964,N_24998);
and UO_1355 (O_1355,N_24946,N_24930);
nand UO_1356 (O_1356,N_24881,N_24919);
xor UO_1357 (O_1357,N_24803,N_24852);
and UO_1358 (O_1358,N_24976,N_24883);
and UO_1359 (O_1359,N_24913,N_24846);
nor UO_1360 (O_1360,N_24819,N_24910);
or UO_1361 (O_1361,N_24980,N_24901);
nor UO_1362 (O_1362,N_24873,N_24906);
and UO_1363 (O_1363,N_24898,N_24866);
or UO_1364 (O_1364,N_24857,N_24847);
or UO_1365 (O_1365,N_24883,N_24978);
and UO_1366 (O_1366,N_24861,N_24811);
nor UO_1367 (O_1367,N_24845,N_24848);
xnor UO_1368 (O_1368,N_24909,N_24805);
nor UO_1369 (O_1369,N_24917,N_24947);
nor UO_1370 (O_1370,N_24842,N_24853);
nor UO_1371 (O_1371,N_24901,N_24868);
nand UO_1372 (O_1372,N_24956,N_24952);
nor UO_1373 (O_1373,N_24992,N_24958);
nor UO_1374 (O_1374,N_24818,N_24927);
and UO_1375 (O_1375,N_24885,N_24869);
or UO_1376 (O_1376,N_24827,N_24811);
and UO_1377 (O_1377,N_24823,N_24925);
and UO_1378 (O_1378,N_24852,N_24964);
nor UO_1379 (O_1379,N_24879,N_24989);
or UO_1380 (O_1380,N_24984,N_24872);
nand UO_1381 (O_1381,N_24911,N_24935);
nor UO_1382 (O_1382,N_24800,N_24884);
or UO_1383 (O_1383,N_24911,N_24841);
and UO_1384 (O_1384,N_24845,N_24984);
xnor UO_1385 (O_1385,N_24804,N_24896);
nor UO_1386 (O_1386,N_24849,N_24874);
nor UO_1387 (O_1387,N_24842,N_24966);
xnor UO_1388 (O_1388,N_24880,N_24968);
or UO_1389 (O_1389,N_24927,N_24970);
and UO_1390 (O_1390,N_24968,N_24894);
and UO_1391 (O_1391,N_24834,N_24849);
nor UO_1392 (O_1392,N_24904,N_24801);
or UO_1393 (O_1393,N_24815,N_24903);
nand UO_1394 (O_1394,N_24842,N_24953);
nand UO_1395 (O_1395,N_24959,N_24868);
nor UO_1396 (O_1396,N_24818,N_24983);
nor UO_1397 (O_1397,N_24853,N_24863);
nand UO_1398 (O_1398,N_24828,N_24850);
nand UO_1399 (O_1399,N_24955,N_24877);
nor UO_1400 (O_1400,N_24955,N_24840);
or UO_1401 (O_1401,N_24911,N_24878);
or UO_1402 (O_1402,N_24882,N_24830);
or UO_1403 (O_1403,N_24912,N_24921);
nand UO_1404 (O_1404,N_24883,N_24912);
xor UO_1405 (O_1405,N_24918,N_24962);
or UO_1406 (O_1406,N_24963,N_24989);
nand UO_1407 (O_1407,N_24845,N_24850);
and UO_1408 (O_1408,N_24995,N_24816);
nor UO_1409 (O_1409,N_24996,N_24812);
nand UO_1410 (O_1410,N_24965,N_24836);
nor UO_1411 (O_1411,N_24984,N_24907);
nor UO_1412 (O_1412,N_24801,N_24900);
and UO_1413 (O_1413,N_24806,N_24878);
nor UO_1414 (O_1414,N_24996,N_24974);
and UO_1415 (O_1415,N_24871,N_24901);
nor UO_1416 (O_1416,N_24960,N_24959);
xor UO_1417 (O_1417,N_24882,N_24847);
and UO_1418 (O_1418,N_24908,N_24886);
nand UO_1419 (O_1419,N_24844,N_24910);
or UO_1420 (O_1420,N_24868,N_24955);
xor UO_1421 (O_1421,N_24911,N_24856);
and UO_1422 (O_1422,N_24877,N_24862);
nand UO_1423 (O_1423,N_24950,N_24951);
and UO_1424 (O_1424,N_24827,N_24857);
and UO_1425 (O_1425,N_24960,N_24935);
nor UO_1426 (O_1426,N_24805,N_24860);
or UO_1427 (O_1427,N_24962,N_24801);
nor UO_1428 (O_1428,N_24830,N_24960);
xor UO_1429 (O_1429,N_24982,N_24801);
and UO_1430 (O_1430,N_24939,N_24969);
xnor UO_1431 (O_1431,N_24923,N_24974);
and UO_1432 (O_1432,N_24918,N_24940);
nor UO_1433 (O_1433,N_24950,N_24871);
nor UO_1434 (O_1434,N_24818,N_24922);
or UO_1435 (O_1435,N_24912,N_24971);
nor UO_1436 (O_1436,N_24854,N_24867);
nand UO_1437 (O_1437,N_24977,N_24966);
nand UO_1438 (O_1438,N_24877,N_24966);
nor UO_1439 (O_1439,N_24943,N_24814);
and UO_1440 (O_1440,N_24849,N_24832);
and UO_1441 (O_1441,N_24817,N_24888);
nor UO_1442 (O_1442,N_24956,N_24991);
and UO_1443 (O_1443,N_24937,N_24933);
xnor UO_1444 (O_1444,N_24857,N_24873);
nand UO_1445 (O_1445,N_24884,N_24981);
nor UO_1446 (O_1446,N_24957,N_24812);
or UO_1447 (O_1447,N_24989,N_24844);
or UO_1448 (O_1448,N_24939,N_24835);
xnor UO_1449 (O_1449,N_24908,N_24878);
and UO_1450 (O_1450,N_24835,N_24940);
nor UO_1451 (O_1451,N_24950,N_24850);
nor UO_1452 (O_1452,N_24887,N_24832);
and UO_1453 (O_1453,N_24970,N_24939);
or UO_1454 (O_1454,N_24988,N_24866);
nor UO_1455 (O_1455,N_24984,N_24863);
or UO_1456 (O_1456,N_24959,N_24902);
nor UO_1457 (O_1457,N_24862,N_24900);
xnor UO_1458 (O_1458,N_24928,N_24952);
and UO_1459 (O_1459,N_24951,N_24886);
xor UO_1460 (O_1460,N_24816,N_24892);
nand UO_1461 (O_1461,N_24996,N_24823);
and UO_1462 (O_1462,N_24832,N_24963);
and UO_1463 (O_1463,N_24822,N_24831);
nor UO_1464 (O_1464,N_24991,N_24998);
or UO_1465 (O_1465,N_24950,N_24909);
and UO_1466 (O_1466,N_24953,N_24805);
nand UO_1467 (O_1467,N_24878,N_24838);
and UO_1468 (O_1468,N_24962,N_24986);
nor UO_1469 (O_1469,N_24876,N_24907);
or UO_1470 (O_1470,N_24813,N_24818);
nand UO_1471 (O_1471,N_24834,N_24823);
xor UO_1472 (O_1472,N_24871,N_24818);
and UO_1473 (O_1473,N_24861,N_24850);
or UO_1474 (O_1474,N_24815,N_24924);
or UO_1475 (O_1475,N_24829,N_24944);
and UO_1476 (O_1476,N_24924,N_24891);
or UO_1477 (O_1477,N_24971,N_24814);
and UO_1478 (O_1478,N_24812,N_24825);
xor UO_1479 (O_1479,N_24890,N_24897);
nor UO_1480 (O_1480,N_24883,N_24914);
xor UO_1481 (O_1481,N_24974,N_24860);
or UO_1482 (O_1482,N_24813,N_24974);
nand UO_1483 (O_1483,N_24897,N_24952);
nor UO_1484 (O_1484,N_24917,N_24936);
nor UO_1485 (O_1485,N_24814,N_24864);
or UO_1486 (O_1486,N_24851,N_24823);
or UO_1487 (O_1487,N_24917,N_24954);
and UO_1488 (O_1488,N_24817,N_24852);
and UO_1489 (O_1489,N_24999,N_24991);
nor UO_1490 (O_1490,N_24866,N_24814);
nor UO_1491 (O_1491,N_24994,N_24825);
and UO_1492 (O_1492,N_24991,N_24878);
and UO_1493 (O_1493,N_24950,N_24875);
nand UO_1494 (O_1494,N_24971,N_24895);
nor UO_1495 (O_1495,N_24879,N_24825);
and UO_1496 (O_1496,N_24861,N_24800);
xnor UO_1497 (O_1497,N_24972,N_24941);
and UO_1498 (O_1498,N_24964,N_24842);
nand UO_1499 (O_1499,N_24916,N_24935);
and UO_1500 (O_1500,N_24969,N_24814);
and UO_1501 (O_1501,N_24853,N_24861);
and UO_1502 (O_1502,N_24930,N_24823);
xor UO_1503 (O_1503,N_24899,N_24847);
nor UO_1504 (O_1504,N_24856,N_24889);
xnor UO_1505 (O_1505,N_24868,N_24931);
or UO_1506 (O_1506,N_24968,N_24892);
xnor UO_1507 (O_1507,N_24875,N_24859);
or UO_1508 (O_1508,N_24830,N_24911);
xnor UO_1509 (O_1509,N_24970,N_24909);
xor UO_1510 (O_1510,N_24919,N_24954);
nand UO_1511 (O_1511,N_24862,N_24985);
and UO_1512 (O_1512,N_24968,N_24852);
nor UO_1513 (O_1513,N_24872,N_24990);
xnor UO_1514 (O_1514,N_24928,N_24877);
nand UO_1515 (O_1515,N_24927,N_24954);
nand UO_1516 (O_1516,N_24913,N_24854);
xor UO_1517 (O_1517,N_24878,N_24895);
or UO_1518 (O_1518,N_24973,N_24821);
nand UO_1519 (O_1519,N_24911,N_24941);
xnor UO_1520 (O_1520,N_24801,N_24847);
xnor UO_1521 (O_1521,N_24996,N_24887);
nand UO_1522 (O_1522,N_24941,N_24882);
nor UO_1523 (O_1523,N_24801,N_24866);
or UO_1524 (O_1524,N_24877,N_24843);
nor UO_1525 (O_1525,N_24944,N_24927);
xor UO_1526 (O_1526,N_24821,N_24955);
xnor UO_1527 (O_1527,N_24894,N_24802);
or UO_1528 (O_1528,N_24865,N_24988);
nor UO_1529 (O_1529,N_24968,N_24840);
or UO_1530 (O_1530,N_24956,N_24954);
and UO_1531 (O_1531,N_24925,N_24937);
xnor UO_1532 (O_1532,N_24872,N_24815);
nor UO_1533 (O_1533,N_24838,N_24801);
and UO_1534 (O_1534,N_24898,N_24904);
or UO_1535 (O_1535,N_24966,N_24970);
and UO_1536 (O_1536,N_24914,N_24915);
and UO_1537 (O_1537,N_24957,N_24897);
or UO_1538 (O_1538,N_24888,N_24933);
nor UO_1539 (O_1539,N_24979,N_24828);
and UO_1540 (O_1540,N_24988,N_24940);
nor UO_1541 (O_1541,N_24890,N_24923);
nand UO_1542 (O_1542,N_24849,N_24918);
xnor UO_1543 (O_1543,N_24937,N_24997);
xnor UO_1544 (O_1544,N_24924,N_24871);
nor UO_1545 (O_1545,N_24907,N_24974);
or UO_1546 (O_1546,N_24906,N_24937);
xnor UO_1547 (O_1547,N_24825,N_24933);
and UO_1548 (O_1548,N_24971,N_24842);
nor UO_1549 (O_1549,N_24851,N_24971);
xor UO_1550 (O_1550,N_24868,N_24904);
xnor UO_1551 (O_1551,N_24898,N_24838);
or UO_1552 (O_1552,N_24933,N_24803);
or UO_1553 (O_1553,N_24883,N_24821);
nor UO_1554 (O_1554,N_24816,N_24930);
nand UO_1555 (O_1555,N_24811,N_24999);
nor UO_1556 (O_1556,N_24845,N_24954);
nand UO_1557 (O_1557,N_24824,N_24945);
nor UO_1558 (O_1558,N_24927,N_24826);
nor UO_1559 (O_1559,N_24820,N_24832);
xor UO_1560 (O_1560,N_24931,N_24895);
nor UO_1561 (O_1561,N_24982,N_24864);
nor UO_1562 (O_1562,N_24833,N_24912);
or UO_1563 (O_1563,N_24821,N_24851);
xnor UO_1564 (O_1564,N_24992,N_24997);
and UO_1565 (O_1565,N_24811,N_24824);
or UO_1566 (O_1566,N_24893,N_24917);
nor UO_1567 (O_1567,N_24998,N_24968);
or UO_1568 (O_1568,N_24910,N_24834);
xnor UO_1569 (O_1569,N_24971,N_24909);
xor UO_1570 (O_1570,N_24808,N_24959);
nand UO_1571 (O_1571,N_24912,N_24852);
nand UO_1572 (O_1572,N_24813,N_24833);
xnor UO_1573 (O_1573,N_24912,N_24943);
xnor UO_1574 (O_1574,N_24874,N_24836);
nand UO_1575 (O_1575,N_24815,N_24855);
xor UO_1576 (O_1576,N_24894,N_24912);
or UO_1577 (O_1577,N_24940,N_24883);
or UO_1578 (O_1578,N_24956,N_24816);
nor UO_1579 (O_1579,N_24869,N_24813);
or UO_1580 (O_1580,N_24874,N_24861);
or UO_1581 (O_1581,N_24904,N_24891);
nand UO_1582 (O_1582,N_24814,N_24977);
or UO_1583 (O_1583,N_24981,N_24957);
or UO_1584 (O_1584,N_24938,N_24991);
nor UO_1585 (O_1585,N_24993,N_24803);
and UO_1586 (O_1586,N_24944,N_24849);
nand UO_1587 (O_1587,N_24844,N_24944);
nand UO_1588 (O_1588,N_24867,N_24816);
nand UO_1589 (O_1589,N_24908,N_24920);
nand UO_1590 (O_1590,N_24850,N_24880);
nand UO_1591 (O_1591,N_24861,N_24814);
xnor UO_1592 (O_1592,N_24931,N_24887);
nor UO_1593 (O_1593,N_24846,N_24899);
nand UO_1594 (O_1594,N_24985,N_24916);
and UO_1595 (O_1595,N_24856,N_24901);
nor UO_1596 (O_1596,N_24835,N_24849);
xor UO_1597 (O_1597,N_24818,N_24838);
and UO_1598 (O_1598,N_24847,N_24996);
nand UO_1599 (O_1599,N_24888,N_24921);
xnor UO_1600 (O_1600,N_24935,N_24965);
and UO_1601 (O_1601,N_24971,N_24911);
xnor UO_1602 (O_1602,N_24868,N_24953);
and UO_1603 (O_1603,N_24867,N_24812);
or UO_1604 (O_1604,N_24806,N_24973);
nor UO_1605 (O_1605,N_24907,N_24865);
xor UO_1606 (O_1606,N_24834,N_24944);
or UO_1607 (O_1607,N_24946,N_24981);
and UO_1608 (O_1608,N_24804,N_24900);
nor UO_1609 (O_1609,N_24890,N_24941);
nand UO_1610 (O_1610,N_24809,N_24963);
and UO_1611 (O_1611,N_24988,N_24905);
xor UO_1612 (O_1612,N_24850,N_24837);
nor UO_1613 (O_1613,N_24925,N_24804);
nor UO_1614 (O_1614,N_24947,N_24817);
or UO_1615 (O_1615,N_24814,N_24932);
nor UO_1616 (O_1616,N_24867,N_24849);
or UO_1617 (O_1617,N_24890,N_24936);
and UO_1618 (O_1618,N_24959,N_24883);
or UO_1619 (O_1619,N_24931,N_24844);
nand UO_1620 (O_1620,N_24936,N_24877);
nand UO_1621 (O_1621,N_24911,N_24966);
or UO_1622 (O_1622,N_24824,N_24904);
nand UO_1623 (O_1623,N_24862,N_24917);
nand UO_1624 (O_1624,N_24889,N_24928);
or UO_1625 (O_1625,N_24889,N_24905);
nand UO_1626 (O_1626,N_24832,N_24947);
or UO_1627 (O_1627,N_24929,N_24870);
nand UO_1628 (O_1628,N_24972,N_24977);
and UO_1629 (O_1629,N_24930,N_24984);
nor UO_1630 (O_1630,N_24956,N_24815);
xnor UO_1631 (O_1631,N_24962,N_24969);
xnor UO_1632 (O_1632,N_24930,N_24809);
nor UO_1633 (O_1633,N_24811,N_24872);
nand UO_1634 (O_1634,N_24963,N_24906);
nand UO_1635 (O_1635,N_24874,N_24855);
nand UO_1636 (O_1636,N_24892,N_24836);
and UO_1637 (O_1637,N_24911,N_24922);
nor UO_1638 (O_1638,N_24916,N_24957);
xor UO_1639 (O_1639,N_24802,N_24906);
and UO_1640 (O_1640,N_24915,N_24954);
nor UO_1641 (O_1641,N_24940,N_24936);
xor UO_1642 (O_1642,N_24993,N_24910);
and UO_1643 (O_1643,N_24992,N_24947);
and UO_1644 (O_1644,N_24984,N_24922);
nor UO_1645 (O_1645,N_24946,N_24956);
nor UO_1646 (O_1646,N_24881,N_24956);
and UO_1647 (O_1647,N_24977,N_24971);
xor UO_1648 (O_1648,N_24872,N_24912);
nor UO_1649 (O_1649,N_24911,N_24920);
and UO_1650 (O_1650,N_24880,N_24920);
nand UO_1651 (O_1651,N_24861,N_24962);
nand UO_1652 (O_1652,N_24802,N_24983);
or UO_1653 (O_1653,N_24940,N_24908);
xnor UO_1654 (O_1654,N_24804,N_24952);
xor UO_1655 (O_1655,N_24936,N_24984);
xor UO_1656 (O_1656,N_24938,N_24881);
nor UO_1657 (O_1657,N_24930,N_24919);
xnor UO_1658 (O_1658,N_24882,N_24978);
xor UO_1659 (O_1659,N_24953,N_24931);
or UO_1660 (O_1660,N_24862,N_24874);
xnor UO_1661 (O_1661,N_24867,N_24969);
xnor UO_1662 (O_1662,N_24868,N_24972);
and UO_1663 (O_1663,N_24971,N_24876);
and UO_1664 (O_1664,N_24983,N_24800);
and UO_1665 (O_1665,N_24905,N_24810);
or UO_1666 (O_1666,N_24945,N_24866);
nor UO_1667 (O_1667,N_24951,N_24974);
xnor UO_1668 (O_1668,N_24816,N_24908);
or UO_1669 (O_1669,N_24913,N_24881);
nor UO_1670 (O_1670,N_24870,N_24964);
xnor UO_1671 (O_1671,N_24841,N_24914);
xnor UO_1672 (O_1672,N_24935,N_24976);
xor UO_1673 (O_1673,N_24971,N_24879);
and UO_1674 (O_1674,N_24845,N_24843);
and UO_1675 (O_1675,N_24925,N_24927);
xnor UO_1676 (O_1676,N_24851,N_24885);
nand UO_1677 (O_1677,N_24808,N_24965);
nor UO_1678 (O_1678,N_24907,N_24852);
xnor UO_1679 (O_1679,N_24949,N_24921);
nor UO_1680 (O_1680,N_24916,N_24818);
and UO_1681 (O_1681,N_24804,N_24878);
or UO_1682 (O_1682,N_24968,N_24973);
nor UO_1683 (O_1683,N_24932,N_24841);
nand UO_1684 (O_1684,N_24972,N_24956);
nor UO_1685 (O_1685,N_24841,N_24908);
nand UO_1686 (O_1686,N_24808,N_24866);
or UO_1687 (O_1687,N_24827,N_24978);
nor UO_1688 (O_1688,N_24974,N_24872);
and UO_1689 (O_1689,N_24879,N_24914);
or UO_1690 (O_1690,N_24807,N_24913);
xor UO_1691 (O_1691,N_24952,N_24929);
xor UO_1692 (O_1692,N_24844,N_24807);
nand UO_1693 (O_1693,N_24867,N_24992);
and UO_1694 (O_1694,N_24914,N_24863);
nand UO_1695 (O_1695,N_24841,N_24856);
or UO_1696 (O_1696,N_24872,N_24995);
and UO_1697 (O_1697,N_24881,N_24974);
xnor UO_1698 (O_1698,N_24839,N_24855);
nor UO_1699 (O_1699,N_24804,N_24943);
nor UO_1700 (O_1700,N_24966,N_24851);
or UO_1701 (O_1701,N_24920,N_24934);
and UO_1702 (O_1702,N_24940,N_24987);
nor UO_1703 (O_1703,N_24922,N_24853);
and UO_1704 (O_1704,N_24879,N_24935);
or UO_1705 (O_1705,N_24957,N_24950);
or UO_1706 (O_1706,N_24808,N_24857);
nand UO_1707 (O_1707,N_24981,N_24958);
xor UO_1708 (O_1708,N_24953,N_24921);
xor UO_1709 (O_1709,N_24942,N_24832);
nand UO_1710 (O_1710,N_24978,N_24968);
or UO_1711 (O_1711,N_24839,N_24951);
and UO_1712 (O_1712,N_24867,N_24926);
and UO_1713 (O_1713,N_24838,N_24852);
nand UO_1714 (O_1714,N_24881,N_24986);
xnor UO_1715 (O_1715,N_24842,N_24935);
nand UO_1716 (O_1716,N_24835,N_24982);
nor UO_1717 (O_1717,N_24993,N_24913);
nand UO_1718 (O_1718,N_24897,N_24995);
xor UO_1719 (O_1719,N_24910,N_24875);
nand UO_1720 (O_1720,N_24809,N_24989);
nor UO_1721 (O_1721,N_24992,N_24933);
and UO_1722 (O_1722,N_24945,N_24972);
xnor UO_1723 (O_1723,N_24998,N_24818);
or UO_1724 (O_1724,N_24846,N_24937);
nand UO_1725 (O_1725,N_24926,N_24884);
nand UO_1726 (O_1726,N_24938,N_24924);
or UO_1727 (O_1727,N_24853,N_24876);
and UO_1728 (O_1728,N_24880,N_24818);
and UO_1729 (O_1729,N_24821,N_24992);
nor UO_1730 (O_1730,N_24832,N_24983);
and UO_1731 (O_1731,N_24984,N_24817);
or UO_1732 (O_1732,N_24929,N_24901);
or UO_1733 (O_1733,N_24828,N_24996);
xor UO_1734 (O_1734,N_24931,N_24857);
nor UO_1735 (O_1735,N_24922,N_24968);
nor UO_1736 (O_1736,N_24947,N_24989);
xnor UO_1737 (O_1737,N_24916,N_24834);
nand UO_1738 (O_1738,N_24882,N_24843);
xor UO_1739 (O_1739,N_24881,N_24879);
nor UO_1740 (O_1740,N_24884,N_24901);
or UO_1741 (O_1741,N_24927,N_24824);
nor UO_1742 (O_1742,N_24902,N_24884);
xnor UO_1743 (O_1743,N_24827,N_24945);
or UO_1744 (O_1744,N_24861,N_24870);
nand UO_1745 (O_1745,N_24884,N_24927);
nand UO_1746 (O_1746,N_24873,N_24956);
or UO_1747 (O_1747,N_24823,N_24955);
and UO_1748 (O_1748,N_24818,N_24978);
and UO_1749 (O_1749,N_24824,N_24870);
nor UO_1750 (O_1750,N_24843,N_24952);
and UO_1751 (O_1751,N_24887,N_24933);
nor UO_1752 (O_1752,N_24832,N_24959);
nor UO_1753 (O_1753,N_24883,N_24946);
xnor UO_1754 (O_1754,N_24810,N_24800);
and UO_1755 (O_1755,N_24869,N_24956);
and UO_1756 (O_1756,N_24820,N_24842);
or UO_1757 (O_1757,N_24818,N_24849);
xor UO_1758 (O_1758,N_24888,N_24836);
xor UO_1759 (O_1759,N_24965,N_24959);
xnor UO_1760 (O_1760,N_24911,N_24943);
and UO_1761 (O_1761,N_24931,N_24910);
nand UO_1762 (O_1762,N_24871,N_24850);
nor UO_1763 (O_1763,N_24887,N_24889);
or UO_1764 (O_1764,N_24985,N_24814);
nor UO_1765 (O_1765,N_24919,N_24901);
or UO_1766 (O_1766,N_24830,N_24893);
xnor UO_1767 (O_1767,N_24898,N_24950);
nand UO_1768 (O_1768,N_24828,N_24969);
or UO_1769 (O_1769,N_24837,N_24862);
nor UO_1770 (O_1770,N_24984,N_24874);
nand UO_1771 (O_1771,N_24993,N_24861);
xor UO_1772 (O_1772,N_24937,N_24888);
nor UO_1773 (O_1773,N_24974,N_24917);
or UO_1774 (O_1774,N_24853,N_24844);
nor UO_1775 (O_1775,N_24997,N_24974);
or UO_1776 (O_1776,N_24900,N_24932);
and UO_1777 (O_1777,N_24966,N_24909);
and UO_1778 (O_1778,N_24899,N_24993);
nor UO_1779 (O_1779,N_24914,N_24954);
nor UO_1780 (O_1780,N_24831,N_24866);
xnor UO_1781 (O_1781,N_24940,N_24971);
or UO_1782 (O_1782,N_24824,N_24853);
nor UO_1783 (O_1783,N_24995,N_24829);
and UO_1784 (O_1784,N_24832,N_24927);
or UO_1785 (O_1785,N_24936,N_24840);
nor UO_1786 (O_1786,N_24828,N_24885);
or UO_1787 (O_1787,N_24888,N_24915);
and UO_1788 (O_1788,N_24843,N_24841);
or UO_1789 (O_1789,N_24894,N_24949);
xor UO_1790 (O_1790,N_24946,N_24895);
and UO_1791 (O_1791,N_24944,N_24970);
nand UO_1792 (O_1792,N_24932,N_24838);
and UO_1793 (O_1793,N_24914,N_24875);
and UO_1794 (O_1794,N_24931,N_24899);
nor UO_1795 (O_1795,N_24853,N_24878);
or UO_1796 (O_1796,N_24859,N_24837);
and UO_1797 (O_1797,N_24935,N_24802);
nor UO_1798 (O_1798,N_24851,N_24870);
or UO_1799 (O_1799,N_24889,N_24952);
nor UO_1800 (O_1800,N_24929,N_24826);
xnor UO_1801 (O_1801,N_24948,N_24804);
xnor UO_1802 (O_1802,N_24855,N_24915);
nor UO_1803 (O_1803,N_24932,N_24945);
nor UO_1804 (O_1804,N_24914,N_24903);
nor UO_1805 (O_1805,N_24823,N_24980);
and UO_1806 (O_1806,N_24928,N_24940);
nand UO_1807 (O_1807,N_24886,N_24824);
and UO_1808 (O_1808,N_24942,N_24993);
xnor UO_1809 (O_1809,N_24953,N_24944);
or UO_1810 (O_1810,N_24834,N_24909);
xnor UO_1811 (O_1811,N_24965,N_24894);
or UO_1812 (O_1812,N_24994,N_24959);
and UO_1813 (O_1813,N_24841,N_24879);
nor UO_1814 (O_1814,N_24832,N_24843);
nand UO_1815 (O_1815,N_24831,N_24943);
or UO_1816 (O_1816,N_24836,N_24830);
nor UO_1817 (O_1817,N_24812,N_24954);
nor UO_1818 (O_1818,N_24909,N_24820);
or UO_1819 (O_1819,N_24815,N_24943);
nand UO_1820 (O_1820,N_24949,N_24864);
and UO_1821 (O_1821,N_24876,N_24883);
nor UO_1822 (O_1822,N_24975,N_24858);
and UO_1823 (O_1823,N_24824,N_24968);
and UO_1824 (O_1824,N_24987,N_24883);
or UO_1825 (O_1825,N_24969,N_24914);
nand UO_1826 (O_1826,N_24982,N_24926);
or UO_1827 (O_1827,N_24886,N_24861);
nand UO_1828 (O_1828,N_24918,N_24827);
xnor UO_1829 (O_1829,N_24970,N_24815);
xnor UO_1830 (O_1830,N_24874,N_24905);
and UO_1831 (O_1831,N_24980,N_24998);
nor UO_1832 (O_1832,N_24893,N_24904);
and UO_1833 (O_1833,N_24895,N_24984);
and UO_1834 (O_1834,N_24974,N_24858);
xnor UO_1835 (O_1835,N_24892,N_24813);
xnor UO_1836 (O_1836,N_24803,N_24836);
nand UO_1837 (O_1837,N_24968,N_24996);
nor UO_1838 (O_1838,N_24970,N_24922);
nor UO_1839 (O_1839,N_24831,N_24856);
nand UO_1840 (O_1840,N_24801,N_24987);
and UO_1841 (O_1841,N_24994,N_24887);
nor UO_1842 (O_1842,N_24960,N_24916);
nand UO_1843 (O_1843,N_24979,N_24875);
and UO_1844 (O_1844,N_24998,N_24917);
or UO_1845 (O_1845,N_24899,N_24920);
or UO_1846 (O_1846,N_24947,N_24990);
and UO_1847 (O_1847,N_24918,N_24955);
or UO_1848 (O_1848,N_24981,N_24925);
nor UO_1849 (O_1849,N_24983,N_24837);
nor UO_1850 (O_1850,N_24975,N_24875);
or UO_1851 (O_1851,N_24829,N_24976);
nor UO_1852 (O_1852,N_24958,N_24811);
xor UO_1853 (O_1853,N_24972,N_24814);
xnor UO_1854 (O_1854,N_24909,N_24887);
nor UO_1855 (O_1855,N_24809,N_24912);
or UO_1856 (O_1856,N_24885,N_24881);
or UO_1857 (O_1857,N_24993,N_24963);
nand UO_1858 (O_1858,N_24813,N_24832);
nand UO_1859 (O_1859,N_24950,N_24946);
nor UO_1860 (O_1860,N_24986,N_24951);
nor UO_1861 (O_1861,N_24934,N_24892);
nand UO_1862 (O_1862,N_24915,N_24804);
nor UO_1863 (O_1863,N_24819,N_24834);
nor UO_1864 (O_1864,N_24919,N_24880);
xnor UO_1865 (O_1865,N_24827,N_24984);
nand UO_1866 (O_1866,N_24890,N_24831);
xor UO_1867 (O_1867,N_24960,N_24846);
nand UO_1868 (O_1868,N_24848,N_24949);
or UO_1869 (O_1869,N_24895,N_24828);
xnor UO_1870 (O_1870,N_24848,N_24965);
or UO_1871 (O_1871,N_24930,N_24898);
or UO_1872 (O_1872,N_24821,N_24809);
or UO_1873 (O_1873,N_24838,N_24943);
or UO_1874 (O_1874,N_24813,N_24979);
and UO_1875 (O_1875,N_24943,N_24932);
and UO_1876 (O_1876,N_24814,N_24848);
nand UO_1877 (O_1877,N_24956,N_24947);
xor UO_1878 (O_1878,N_24984,N_24942);
and UO_1879 (O_1879,N_24907,N_24866);
xor UO_1880 (O_1880,N_24862,N_24929);
and UO_1881 (O_1881,N_24947,N_24934);
and UO_1882 (O_1882,N_24937,N_24960);
and UO_1883 (O_1883,N_24941,N_24835);
and UO_1884 (O_1884,N_24920,N_24941);
nand UO_1885 (O_1885,N_24871,N_24828);
nor UO_1886 (O_1886,N_24904,N_24807);
nor UO_1887 (O_1887,N_24862,N_24950);
or UO_1888 (O_1888,N_24880,N_24962);
xnor UO_1889 (O_1889,N_24970,N_24847);
xnor UO_1890 (O_1890,N_24899,N_24859);
and UO_1891 (O_1891,N_24884,N_24806);
nand UO_1892 (O_1892,N_24932,N_24883);
nor UO_1893 (O_1893,N_24922,N_24956);
or UO_1894 (O_1894,N_24809,N_24999);
nor UO_1895 (O_1895,N_24983,N_24868);
nand UO_1896 (O_1896,N_24839,N_24964);
and UO_1897 (O_1897,N_24813,N_24826);
nand UO_1898 (O_1898,N_24978,N_24809);
nand UO_1899 (O_1899,N_24870,N_24813);
xor UO_1900 (O_1900,N_24952,N_24976);
nor UO_1901 (O_1901,N_24845,N_24801);
nand UO_1902 (O_1902,N_24869,N_24893);
nor UO_1903 (O_1903,N_24942,N_24979);
nand UO_1904 (O_1904,N_24944,N_24806);
nand UO_1905 (O_1905,N_24938,N_24891);
and UO_1906 (O_1906,N_24964,N_24807);
or UO_1907 (O_1907,N_24964,N_24877);
xor UO_1908 (O_1908,N_24873,N_24954);
nand UO_1909 (O_1909,N_24930,N_24905);
nand UO_1910 (O_1910,N_24846,N_24837);
nor UO_1911 (O_1911,N_24906,N_24903);
nor UO_1912 (O_1912,N_24843,N_24873);
or UO_1913 (O_1913,N_24956,N_24853);
nor UO_1914 (O_1914,N_24901,N_24988);
or UO_1915 (O_1915,N_24851,N_24919);
xor UO_1916 (O_1916,N_24859,N_24947);
nand UO_1917 (O_1917,N_24878,N_24939);
nor UO_1918 (O_1918,N_24898,N_24926);
or UO_1919 (O_1919,N_24992,N_24916);
and UO_1920 (O_1920,N_24910,N_24966);
and UO_1921 (O_1921,N_24922,N_24841);
or UO_1922 (O_1922,N_24963,N_24911);
or UO_1923 (O_1923,N_24808,N_24949);
or UO_1924 (O_1924,N_24800,N_24950);
xnor UO_1925 (O_1925,N_24933,N_24908);
nor UO_1926 (O_1926,N_24823,N_24916);
nand UO_1927 (O_1927,N_24820,N_24822);
and UO_1928 (O_1928,N_24910,N_24912);
and UO_1929 (O_1929,N_24956,N_24863);
or UO_1930 (O_1930,N_24945,N_24863);
and UO_1931 (O_1931,N_24970,N_24876);
xnor UO_1932 (O_1932,N_24923,N_24903);
nor UO_1933 (O_1933,N_24982,N_24950);
xor UO_1934 (O_1934,N_24951,N_24993);
nor UO_1935 (O_1935,N_24954,N_24947);
xor UO_1936 (O_1936,N_24910,N_24839);
and UO_1937 (O_1937,N_24849,N_24854);
nand UO_1938 (O_1938,N_24996,N_24884);
nand UO_1939 (O_1939,N_24969,N_24958);
and UO_1940 (O_1940,N_24866,N_24844);
and UO_1941 (O_1941,N_24871,N_24802);
nand UO_1942 (O_1942,N_24948,N_24979);
or UO_1943 (O_1943,N_24817,N_24946);
and UO_1944 (O_1944,N_24923,N_24872);
or UO_1945 (O_1945,N_24829,N_24906);
xnor UO_1946 (O_1946,N_24805,N_24857);
xor UO_1947 (O_1947,N_24809,N_24947);
nand UO_1948 (O_1948,N_24836,N_24809);
and UO_1949 (O_1949,N_24905,N_24812);
nor UO_1950 (O_1950,N_24981,N_24813);
or UO_1951 (O_1951,N_24927,N_24820);
and UO_1952 (O_1952,N_24915,N_24956);
xnor UO_1953 (O_1953,N_24983,N_24856);
nor UO_1954 (O_1954,N_24986,N_24867);
nor UO_1955 (O_1955,N_24900,N_24860);
or UO_1956 (O_1956,N_24985,N_24917);
or UO_1957 (O_1957,N_24995,N_24941);
nand UO_1958 (O_1958,N_24915,N_24913);
or UO_1959 (O_1959,N_24950,N_24881);
nand UO_1960 (O_1960,N_24987,N_24900);
xor UO_1961 (O_1961,N_24879,N_24917);
nand UO_1962 (O_1962,N_24982,N_24981);
or UO_1963 (O_1963,N_24850,N_24832);
nor UO_1964 (O_1964,N_24996,N_24936);
or UO_1965 (O_1965,N_24837,N_24942);
or UO_1966 (O_1966,N_24969,N_24902);
nor UO_1967 (O_1967,N_24889,N_24861);
xor UO_1968 (O_1968,N_24925,N_24814);
or UO_1969 (O_1969,N_24807,N_24934);
nand UO_1970 (O_1970,N_24826,N_24966);
or UO_1971 (O_1971,N_24986,N_24965);
or UO_1972 (O_1972,N_24890,N_24969);
xor UO_1973 (O_1973,N_24917,N_24878);
and UO_1974 (O_1974,N_24815,N_24891);
nand UO_1975 (O_1975,N_24893,N_24940);
nand UO_1976 (O_1976,N_24856,N_24915);
and UO_1977 (O_1977,N_24976,N_24888);
nor UO_1978 (O_1978,N_24956,N_24944);
and UO_1979 (O_1979,N_24882,N_24949);
nor UO_1980 (O_1980,N_24855,N_24972);
and UO_1981 (O_1981,N_24904,N_24927);
or UO_1982 (O_1982,N_24819,N_24934);
or UO_1983 (O_1983,N_24843,N_24937);
or UO_1984 (O_1984,N_24991,N_24810);
and UO_1985 (O_1985,N_24970,N_24916);
or UO_1986 (O_1986,N_24807,N_24811);
nor UO_1987 (O_1987,N_24854,N_24963);
or UO_1988 (O_1988,N_24976,N_24960);
nand UO_1989 (O_1989,N_24953,N_24814);
nor UO_1990 (O_1990,N_24964,N_24892);
nand UO_1991 (O_1991,N_24892,N_24985);
nor UO_1992 (O_1992,N_24945,N_24872);
or UO_1993 (O_1993,N_24907,N_24962);
xnor UO_1994 (O_1994,N_24904,N_24958);
and UO_1995 (O_1995,N_24876,N_24986);
nand UO_1996 (O_1996,N_24938,N_24822);
and UO_1997 (O_1997,N_24919,N_24805);
and UO_1998 (O_1998,N_24878,N_24823);
nor UO_1999 (O_1999,N_24992,N_24959);
and UO_2000 (O_2000,N_24826,N_24809);
nor UO_2001 (O_2001,N_24902,N_24947);
nand UO_2002 (O_2002,N_24877,N_24905);
nor UO_2003 (O_2003,N_24980,N_24820);
and UO_2004 (O_2004,N_24935,N_24936);
xnor UO_2005 (O_2005,N_24933,N_24833);
nand UO_2006 (O_2006,N_24996,N_24880);
xnor UO_2007 (O_2007,N_24894,N_24827);
nand UO_2008 (O_2008,N_24903,N_24984);
nor UO_2009 (O_2009,N_24913,N_24952);
or UO_2010 (O_2010,N_24873,N_24931);
nor UO_2011 (O_2011,N_24946,N_24802);
or UO_2012 (O_2012,N_24983,N_24921);
nor UO_2013 (O_2013,N_24861,N_24821);
or UO_2014 (O_2014,N_24974,N_24870);
or UO_2015 (O_2015,N_24839,N_24940);
xor UO_2016 (O_2016,N_24812,N_24834);
nor UO_2017 (O_2017,N_24803,N_24920);
nor UO_2018 (O_2018,N_24951,N_24989);
nand UO_2019 (O_2019,N_24925,N_24812);
nand UO_2020 (O_2020,N_24863,N_24868);
nand UO_2021 (O_2021,N_24964,N_24987);
nand UO_2022 (O_2022,N_24805,N_24985);
nand UO_2023 (O_2023,N_24930,N_24934);
or UO_2024 (O_2024,N_24816,N_24932);
nor UO_2025 (O_2025,N_24816,N_24827);
xor UO_2026 (O_2026,N_24824,N_24991);
or UO_2027 (O_2027,N_24973,N_24910);
xor UO_2028 (O_2028,N_24819,N_24937);
or UO_2029 (O_2029,N_24921,N_24959);
nor UO_2030 (O_2030,N_24828,N_24818);
xnor UO_2031 (O_2031,N_24966,N_24902);
and UO_2032 (O_2032,N_24959,N_24942);
xor UO_2033 (O_2033,N_24856,N_24910);
nor UO_2034 (O_2034,N_24996,N_24975);
or UO_2035 (O_2035,N_24800,N_24818);
xor UO_2036 (O_2036,N_24861,N_24843);
nand UO_2037 (O_2037,N_24955,N_24952);
or UO_2038 (O_2038,N_24921,N_24968);
nand UO_2039 (O_2039,N_24809,N_24838);
nor UO_2040 (O_2040,N_24899,N_24982);
and UO_2041 (O_2041,N_24914,N_24821);
xor UO_2042 (O_2042,N_24977,N_24822);
nand UO_2043 (O_2043,N_24832,N_24863);
and UO_2044 (O_2044,N_24947,N_24915);
xnor UO_2045 (O_2045,N_24937,N_24814);
nor UO_2046 (O_2046,N_24811,N_24884);
xnor UO_2047 (O_2047,N_24917,N_24997);
nand UO_2048 (O_2048,N_24838,N_24984);
and UO_2049 (O_2049,N_24909,N_24973);
and UO_2050 (O_2050,N_24995,N_24973);
and UO_2051 (O_2051,N_24872,N_24830);
and UO_2052 (O_2052,N_24877,N_24821);
nand UO_2053 (O_2053,N_24926,N_24950);
nand UO_2054 (O_2054,N_24850,N_24836);
or UO_2055 (O_2055,N_24899,N_24850);
xnor UO_2056 (O_2056,N_24947,N_24840);
or UO_2057 (O_2057,N_24917,N_24993);
or UO_2058 (O_2058,N_24845,N_24944);
or UO_2059 (O_2059,N_24841,N_24852);
nor UO_2060 (O_2060,N_24984,N_24947);
xor UO_2061 (O_2061,N_24915,N_24982);
nand UO_2062 (O_2062,N_24850,N_24984);
or UO_2063 (O_2063,N_24911,N_24931);
xor UO_2064 (O_2064,N_24916,N_24810);
or UO_2065 (O_2065,N_24940,N_24867);
or UO_2066 (O_2066,N_24897,N_24848);
xor UO_2067 (O_2067,N_24993,N_24976);
or UO_2068 (O_2068,N_24946,N_24800);
nand UO_2069 (O_2069,N_24882,N_24886);
nand UO_2070 (O_2070,N_24831,N_24932);
or UO_2071 (O_2071,N_24923,N_24915);
xor UO_2072 (O_2072,N_24965,N_24957);
nand UO_2073 (O_2073,N_24942,N_24982);
nand UO_2074 (O_2074,N_24857,N_24853);
nand UO_2075 (O_2075,N_24815,N_24948);
xor UO_2076 (O_2076,N_24949,N_24846);
nor UO_2077 (O_2077,N_24883,N_24897);
or UO_2078 (O_2078,N_24951,N_24803);
nand UO_2079 (O_2079,N_24826,N_24886);
xnor UO_2080 (O_2080,N_24817,N_24912);
nor UO_2081 (O_2081,N_24983,N_24902);
nor UO_2082 (O_2082,N_24898,N_24835);
or UO_2083 (O_2083,N_24853,N_24947);
nand UO_2084 (O_2084,N_24939,N_24813);
nand UO_2085 (O_2085,N_24971,N_24926);
and UO_2086 (O_2086,N_24982,N_24837);
nand UO_2087 (O_2087,N_24941,N_24927);
xnor UO_2088 (O_2088,N_24852,N_24800);
nor UO_2089 (O_2089,N_24845,N_24866);
xor UO_2090 (O_2090,N_24974,N_24802);
nor UO_2091 (O_2091,N_24955,N_24807);
nand UO_2092 (O_2092,N_24875,N_24807);
and UO_2093 (O_2093,N_24835,N_24993);
nor UO_2094 (O_2094,N_24830,N_24833);
xor UO_2095 (O_2095,N_24898,N_24839);
or UO_2096 (O_2096,N_24897,N_24924);
nor UO_2097 (O_2097,N_24837,N_24937);
xor UO_2098 (O_2098,N_24921,N_24818);
xor UO_2099 (O_2099,N_24835,N_24970);
nand UO_2100 (O_2100,N_24895,N_24887);
nor UO_2101 (O_2101,N_24824,N_24839);
or UO_2102 (O_2102,N_24919,N_24903);
and UO_2103 (O_2103,N_24861,N_24941);
nand UO_2104 (O_2104,N_24903,N_24913);
nor UO_2105 (O_2105,N_24904,N_24844);
nor UO_2106 (O_2106,N_24824,N_24942);
and UO_2107 (O_2107,N_24866,N_24938);
nor UO_2108 (O_2108,N_24859,N_24854);
nor UO_2109 (O_2109,N_24875,N_24832);
xor UO_2110 (O_2110,N_24931,N_24984);
xnor UO_2111 (O_2111,N_24816,N_24909);
or UO_2112 (O_2112,N_24925,N_24998);
and UO_2113 (O_2113,N_24928,N_24827);
xor UO_2114 (O_2114,N_24938,N_24927);
xnor UO_2115 (O_2115,N_24988,N_24981);
nor UO_2116 (O_2116,N_24949,N_24923);
and UO_2117 (O_2117,N_24950,N_24915);
and UO_2118 (O_2118,N_24972,N_24984);
nor UO_2119 (O_2119,N_24856,N_24836);
nor UO_2120 (O_2120,N_24997,N_24925);
and UO_2121 (O_2121,N_24998,N_24869);
or UO_2122 (O_2122,N_24986,N_24984);
or UO_2123 (O_2123,N_24920,N_24860);
nand UO_2124 (O_2124,N_24953,N_24883);
xor UO_2125 (O_2125,N_24997,N_24932);
and UO_2126 (O_2126,N_24952,N_24885);
xor UO_2127 (O_2127,N_24950,N_24899);
or UO_2128 (O_2128,N_24922,N_24927);
nor UO_2129 (O_2129,N_24942,N_24815);
nor UO_2130 (O_2130,N_24909,N_24991);
nor UO_2131 (O_2131,N_24894,N_24806);
and UO_2132 (O_2132,N_24921,N_24833);
xor UO_2133 (O_2133,N_24938,N_24908);
and UO_2134 (O_2134,N_24879,N_24844);
xnor UO_2135 (O_2135,N_24827,N_24973);
xnor UO_2136 (O_2136,N_24901,N_24909);
nand UO_2137 (O_2137,N_24963,N_24998);
nor UO_2138 (O_2138,N_24831,N_24892);
nor UO_2139 (O_2139,N_24906,N_24832);
xor UO_2140 (O_2140,N_24825,N_24863);
nand UO_2141 (O_2141,N_24853,N_24927);
xnor UO_2142 (O_2142,N_24902,N_24815);
or UO_2143 (O_2143,N_24969,N_24896);
or UO_2144 (O_2144,N_24959,N_24922);
or UO_2145 (O_2145,N_24991,N_24891);
nand UO_2146 (O_2146,N_24823,N_24892);
xor UO_2147 (O_2147,N_24876,N_24806);
nor UO_2148 (O_2148,N_24966,N_24978);
nor UO_2149 (O_2149,N_24928,N_24987);
or UO_2150 (O_2150,N_24979,N_24914);
nand UO_2151 (O_2151,N_24815,N_24859);
nand UO_2152 (O_2152,N_24995,N_24990);
and UO_2153 (O_2153,N_24882,N_24811);
nand UO_2154 (O_2154,N_24910,N_24808);
nor UO_2155 (O_2155,N_24998,N_24929);
and UO_2156 (O_2156,N_24858,N_24990);
or UO_2157 (O_2157,N_24935,N_24985);
nor UO_2158 (O_2158,N_24886,N_24869);
xnor UO_2159 (O_2159,N_24920,N_24856);
and UO_2160 (O_2160,N_24962,N_24929);
nand UO_2161 (O_2161,N_24895,N_24876);
and UO_2162 (O_2162,N_24912,N_24995);
or UO_2163 (O_2163,N_24829,N_24889);
nand UO_2164 (O_2164,N_24801,N_24892);
and UO_2165 (O_2165,N_24864,N_24879);
and UO_2166 (O_2166,N_24887,N_24874);
nand UO_2167 (O_2167,N_24848,N_24920);
nand UO_2168 (O_2168,N_24917,N_24966);
xor UO_2169 (O_2169,N_24908,N_24972);
nand UO_2170 (O_2170,N_24854,N_24916);
nor UO_2171 (O_2171,N_24902,N_24992);
nand UO_2172 (O_2172,N_24908,N_24814);
nand UO_2173 (O_2173,N_24820,N_24970);
or UO_2174 (O_2174,N_24970,N_24827);
nand UO_2175 (O_2175,N_24886,N_24892);
and UO_2176 (O_2176,N_24870,N_24877);
and UO_2177 (O_2177,N_24939,N_24943);
nor UO_2178 (O_2178,N_24967,N_24981);
or UO_2179 (O_2179,N_24952,N_24908);
xor UO_2180 (O_2180,N_24832,N_24866);
nor UO_2181 (O_2181,N_24826,N_24834);
nand UO_2182 (O_2182,N_24902,N_24940);
nor UO_2183 (O_2183,N_24977,N_24872);
and UO_2184 (O_2184,N_24909,N_24961);
or UO_2185 (O_2185,N_24836,N_24975);
nand UO_2186 (O_2186,N_24844,N_24978);
xor UO_2187 (O_2187,N_24818,N_24822);
and UO_2188 (O_2188,N_24855,N_24964);
nand UO_2189 (O_2189,N_24923,N_24808);
nand UO_2190 (O_2190,N_24845,N_24942);
and UO_2191 (O_2191,N_24821,N_24968);
and UO_2192 (O_2192,N_24959,N_24862);
or UO_2193 (O_2193,N_24887,N_24976);
nand UO_2194 (O_2194,N_24950,N_24907);
xor UO_2195 (O_2195,N_24994,N_24833);
and UO_2196 (O_2196,N_24899,N_24918);
and UO_2197 (O_2197,N_24965,N_24862);
xor UO_2198 (O_2198,N_24906,N_24834);
nand UO_2199 (O_2199,N_24966,N_24968);
xor UO_2200 (O_2200,N_24880,N_24805);
xor UO_2201 (O_2201,N_24870,N_24803);
or UO_2202 (O_2202,N_24990,N_24856);
nor UO_2203 (O_2203,N_24979,N_24866);
xnor UO_2204 (O_2204,N_24996,N_24985);
and UO_2205 (O_2205,N_24891,N_24893);
or UO_2206 (O_2206,N_24859,N_24971);
nor UO_2207 (O_2207,N_24814,N_24891);
nand UO_2208 (O_2208,N_24840,N_24942);
or UO_2209 (O_2209,N_24816,N_24965);
xor UO_2210 (O_2210,N_24945,N_24860);
nand UO_2211 (O_2211,N_24836,N_24852);
nor UO_2212 (O_2212,N_24829,N_24851);
or UO_2213 (O_2213,N_24829,N_24982);
or UO_2214 (O_2214,N_24890,N_24817);
nor UO_2215 (O_2215,N_24819,N_24875);
nor UO_2216 (O_2216,N_24858,N_24852);
xor UO_2217 (O_2217,N_24839,N_24970);
and UO_2218 (O_2218,N_24994,N_24912);
nor UO_2219 (O_2219,N_24961,N_24855);
nand UO_2220 (O_2220,N_24862,N_24891);
xor UO_2221 (O_2221,N_24800,N_24998);
nand UO_2222 (O_2222,N_24853,N_24919);
and UO_2223 (O_2223,N_24989,N_24919);
and UO_2224 (O_2224,N_24821,N_24965);
nor UO_2225 (O_2225,N_24864,N_24876);
nor UO_2226 (O_2226,N_24817,N_24893);
and UO_2227 (O_2227,N_24914,N_24880);
nor UO_2228 (O_2228,N_24964,N_24802);
or UO_2229 (O_2229,N_24972,N_24993);
nand UO_2230 (O_2230,N_24884,N_24933);
and UO_2231 (O_2231,N_24976,N_24925);
and UO_2232 (O_2232,N_24905,N_24979);
nor UO_2233 (O_2233,N_24856,N_24941);
and UO_2234 (O_2234,N_24889,N_24972);
and UO_2235 (O_2235,N_24821,N_24921);
nand UO_2236 (O_2236,N_24934,N_24843);
and UO_2237 (O_2237,N_24907,N_24905);
nand UO_2238 (O_2238,N_24918,N_24823);
and UO_2239 (O_2239,N_24852,N_24905);
xnor UO_2240 (O_2240,N_24897,N_24996);
and UO_2241 (O_2241,N_24877,N_24911);
nor UO_2242 (O_2242,N_24888,N_24851);
xnor UO_2243 (O_2243,N_24966,N_24961);
xor UO_2244 (O_2244,N_24835,N_24968);
nor UO_2245 (O_2245,N_24828,N_24869);
nand UO_2246 (O_2246,N_24944,N_24850);
xnor UO_2247 (O_2247,N_24814,N_24831);
xnor UO_2248 (O_2248,N_24910,N_24899);
and UO_2249 (O_2249,N_24821,N_24970);
or UO_2250 (O_2250,N_24808,N_24972);
xor UO_2251 (O_2251,N_24888,N_24837);
or UO_2252 (O_2252,N_24845,N_24951);
and UO_2253 (O_2253,N_24886,N_24947);
or UO_2254 (O_2254,N_24839,N_24991);
xnor UO_2255 (O_2255,N_24966,N_24829);
and UO_2256 (O_2256,N_24993,N_24824);
nand UO_2257 (O_2257,N_24994,N_24850);
nand UO_2258 (O_2258,N_24953,N_24823);
nor UO_2259 (O_2259,N_24919,N_24971);
xnor UO_2260 (O_2260,N_24912,N_24999);
or UO_2261 (O_2261,N_24997,N_24883);
nand UO_2262 (O_2262,N_24920,N_24877);
xnor UO_2263 (O_2263,N_24866,N_24936);
nor UO_2264 (O_2264,N_24831,N_24939);
xnor UO_2265 (O_2265,N_24918,N_24942);
and UO_2266 (O_2266,N_24994,N_24888);
and UO_2267 (O_2267,N_24884,N_24962);
or UO_2268 (O_2268,N_24807,N_24833);
nor UO_2269 (O_2269,N_24826,N_24932);
or UO_2270 (O_2270,N_24956,N_24871);
nor UO_2271 (O_2271,N_24959,N_24909);
nand UO_2272 (O_2272,N_24957,N_24948);
nor UO_2273 (O_2273,N_24913,N_24919);
and UO_2274 (O_2274,N_24893,N_24915);
nor UO_2275 (O_2275,N_24814,N_24918);
nand UO_2276 (O_2276,N_24922,N_24913);
xnor UO_2277 (O_2277,N_24958,N_24941);
or UO_2278 (O_2278,N_24971,N_24838);
and UO_2279 (O_2279,N_24928,N_24948);
nor UO_2280 (O_2280,N_24953,N_24875);
and UO_2281 (O_2281,N_24934,N_24949);
nand UO_2282 (O_2282,N_24958,N_24999);
or UO_2283 (O_2283,N_24910,N_24999);
nand UO_2284 (O_2284,N_24812,N_24853);
or UO_2285 (O_2285,N_24830,N_24822);
nor UO_2286 (O_2286,N_24867,N_24990);
xnor UO_2287 (O_2287,N_24955,N_24824);
nand UO_2288 (O_2288,N_24833,N_24967);
and UO_2289 (O_2289,N_24972,N_24887);
nor UO_2290 (O_2290,N_24953,N_24971);
or UO_2291 (O_2291,N_24816,N_24850);
and UO_2292 (O_2292,N_24928,N_24807);
nand UO_2293 (O_2293,N_24938,N_24893);
nand UO_2294 (O_2294,N_24808,N_24922);
nand UO_2295 (O_2295,N_24899,N_24836);
or UO_2296 (O_2296,N_24821,N_24995);
nand UO_2297 (O_2297,N_24827,N_24980);
nand UO_2298 (O_2298,N_24880,N_24955);
nand UO_2299 (O_2299,N_24920,N_24981);
or UO_2300 (O_2300,N_24847,N_24912);
nand UO_2301 (O_2301,N_24931,N_24987);
xnor UO_2302 (O_2302,N_24932,N_24890);
nor UO_2303 (O_2303,N_24854,N_24947);
xnor UO_2304 (O_2304,N_24897,N_24825);
and UO_2305 (O_2305,N_24882,N_24867);
nor UO_2306 (O_2306,N_24963,N_24957);
nor UO_2307 (O_2307,N_24838,N_24886);
or UO_2308 (O_2308,N_24935,N_24926);
and UO_2309 (O_2309,N_24859,N_24999);
nand UO_2310 (O_2310,N_24829,N_24916);
xnor UO_2311 (O_2311,N_24983,N_24881);
or UO_2312 (O_2312,N_24843,N_24994);
nor UO_2313 (O_2313,N_24961,N_24883);
xnor UO_2314 (O_2314,N_24860,N_24803);
and UO_2315 (O_2315,N_24921,N_24909);
nor UO_2316 (O_2316,N_24856,N_24960);
xor UO_2317 (O_2317,N_24851,N_24979);
nand UO_2318 (O_2318,N_24952,N_24984);
nand UO_2319 (O_2319,N_24945,N_24838);
nand UO_2320 (O_2320,N_24950,N_24891);
and UO_2321 (O_2321,N_24974,N_24896);
and UO_2322 (O_2322,N_24804,N_24875);
or UO_2323 (O_2323,N_24938,N_24900);
nand UO_2324 (O_2324,N_24921,N_24939);
xnor UO_2325 (O_2325,N_24825,N_24859);
nand UO_2326 (O_2326,N_24881,N_24951);
nand UO_2327 (O_2327,N_24955,N_24910);
and UO_2328 (O_2328,N_24872,N_24846);
or UO_2329 (O_2329,N_24991,N_24946);
nor UO_2330 (O_2330,N_24966,N_24901);
nand UO_2331 (O_2331,N_24919,N_24856);
or UO_2332 (O_2332,N_24896,N_24942);
nand UO_2333 (O_2333,N_24934,N_24933);
or UO_2334 (O_2334,N_24840,N_24957);
or UO_2335 (O_2335,N_24877,N_24894);
nand UO_2336 (O_2336,N_24876,N_24935);
or UO_2337 (O_2337,N_24814,N_24872);
nand UO_2338 (O_2338,N_24866,N_24872);
nor UO_2339 (O_2339,N_24901,N_24942);
or UO_2340 (O_2340,N_24967,N_24864);
nand UO_2341 (O_2341,N_24800,N_24925);
and UO_2342 (O_2342,N_24908,N_24860);
nand UO_2343 (O_2343,N_24964,N_24951);
xor UO_2344 (O_2344,N_24854,N_24863);
or UO_2345 (O_2345,N_24886,N_24809);
or UO_2346 (O_2346,N_24826,N_24838);
nand UO_2347 (O_2347,N_24935,N_24956);
and UO_2348 (O_2348,N_24826,N_24832);
nor UO_2349 (O_2349,N_24830,N_24846);
nand UO_2350 (O_2350,N_24866,N_24934);
and UO_2351 (O_2351,N_24839,N_24810);
nor UO_2352 (O_2352,N_24969,N_24909);
and UO_2353 (O_2353,N_24978,N_24942);
or UO_2354 (O_2354,N_24832,N_24897);
or UO_2355 (O_2355,N_24966,N_24870);
and UO_2356 (O_2356,N_24862,N_24814);
nor UO_2357 (O_2357,N_24989,N_24948);
and UO_2358 (O_2358,N_24994,N_24861);
xnor UO_2359 (O_2359,N_24966,N_24963);
nor UO_2360 (O_2360,N_24920,N_24833);
or UO_2361 (O_2361,N_24878,N_24843);
and UO_2362 (O_2362,N_24804,N_24906);
or UO_2363 (O_2363,N_24899,N_24984);
and UO_2364 (O_2364,N_24968,N_24950);
and UO_2365 (O_2365,N_24883,N_24853);
or UO_2366 (O_2366,N_24912,N_24976);
nand UO_2367 (O_2367,N_24999,N_24802);
nand UO_2368 (O_2368,N_24857,N_24802);
and UO_2369 (O_2369,N_24884,N_24819);
nand UO_2370 (O_2370,N_24879,N_24982);
and UO_2371 (O_2371,N_24821,N_24854);
or UO_2372 (O_2372,N_24991,N_24937);
xnor UO_2373 (O_2373,N_24865,N_24857);
or UO_2374 (O_2374,N_24880,N_24961);
or UO_2375 (O_2375,N_24957,N_24841);
nand UO_2376 (O_2376,N_24956,N_24864);
or UO_2377 (O_2377,N_24802,N_24976);
or UO_2378 (O_2378,N_24854,N_24901);
xnor UO_2379 (O_2379,N_24884,N_24967);
or UO_2380 (O_2380,N_24835,N_24928);
nor UO_2381 (O_2381,N_24887,N_24859);
nand UO_2382 (O_2382,N_24915,N_24903);
and UO_2383 (O_2383,N_24935,N_24860);
and UO_2384 (O_2384,N_24979,N_24982);
or UO_2385 (O_2385,N_24928,N_24874);
xor UO_2386 (O_2386,N_24928,N_24927);
or UO_2387 (O_2387,N_24825,N_24883);
xor UO_2388 (O_2388,N_24978,N_24803);
nand UO_2389 (O_2389,N_24963,N_24812);
nor UO_2390 (O_2390,N_24888,N_24959);
nor UO_2391 (O_2391,N_24803,N_24805);
nand UO_2392 (O_2392,N_24882,N_24942);
or UO_2393 (O_2393,N_24833,N_24944);
xor UO_2394 (O_2394,N_24850,N_24875);
or UO_2395 (O_2395,N_24952,N_24875);
or UO_2396 (O_2396,N_24869,N_24988);
nor UO_2397 (O_2397,N_24938,N_24959);
or UO_2398 (O_2398,N_24932,N_24844);
and UO_2399 (O_2399,N_24861,N_24931);
nand UO_2400 (O_2400,N_24827,N_24968);
xor UO_2401 (O_2401,N_24924,N_24837);
nor UO_2402 (O_2402,N_24817,N_24862);
nor UO_2403 (O_2403,N_24884,N_24944);
nor UO_2404 (O_2404,N_24937,N_24979);
nor UO_2405 (O_2405,N_24828,N_24939);
and UO_2406 (O_2406,N_24834,N_24969);
nor UO_2407 (O_2407,N_24845,N_24991);
xnor UO_2408 (O_2408,N_24881,N_24882);
nor UO_2409 (O_2409,N_24929,N_24835);
and UO_2410 (O_2410,N_24825,N_24980);
or UO_2411 (O_2411,N_24896,N_24872);
xor UO_2412 (O_2412,N_24973,N_24803);
xor UO_2413 (O_2413,N_24945,N_24949);
or UO_2414 (O_2414,N_24813,N_24881);
nor UO_2415 (O_2415,N_24958,N_24901);
xnor UO_2416 (O_2416,N_24858,N_24957);
nor UO_2417 (O_2417,N_24855,N_24917);
xnor UO_2418 (O_2418,N_24948,N_24877);
xnor UO_2419 (O_2419,N_24906,N_24830);
xor UO_2420 (O_2420,N_24934,N_24859);
xor UO_2421 (O_2421,N_24814,N_24822);
nor UO_2422 (O_2422,N_24809,N_24881);
or UO_2423 (O_2423,N_24903,N_24807);
nor UO_2424 (O_2424,N_24966,N_24884);
and UO_2425 (O_2425,N_24953,N_24992);
nand UO_2426 (O_2426,N_24905,N_24935);
nand UO_2427 (O_2427,N_24811,N_24909);
or UO_2428 (O_2428,N_24875,N_24816);
nor UO_2429 (O_2429,N_24811,N_24995);
or UO_2430 (O_2430,N_24983,N_24855);
nor UO_2431 (O_2431,N_24811,N_24888);
nor UO_2432 (O_2432,N_24952,N_24879);
xor UO_2433 (O_2433,N_24886,N_24911);
or UO_2434 (O_2434,N_24953,N_24821);
or UO_2435 (O_2435,N_24991,N_24855);
xor UO_2436 (O_2436,N_24908,N_24807);
nor UO_2437 (O_2437,N_24899,N_24938);
and UO_2438 (O_2438,N_24824,N_24876);
and UO_2439 (O_2439,N_24991,N_24822);
and UO_2440 (O_2440,N_24810,N_24849);
nand UO_2441 (O_2441,N_24953,N_24942);
and UO_2442 (O_2442,N_24888,N_24895);
or UO_2443 (O_2443,N_24953,N_24884);
nand UO_2444 (O_2444,N_24986,N_24871);
nand UO_2445 (O_2445,N_24856,N_24970);
and UO_2446 (O_2446,N_24859,N_24970);
or UO_2447 (O_2447,N_24875,N_24857);
or UO_2448 (O_2448,N_24897,N_24892);
xnor UO_2449 (O_2449,N_24864,N_24863);
xnor UO_2450 (O_2450,N_24980,N_24871);
nand UO_2451 (O_2451,N_24986,N_24832);
or UO_2452 (O_2452,N_24804,N_24907);
nor UO_2453 (O_2453,N_24971,N_24831);
or UO_2454 (O_2454,N_24826,N_24862);
xor UO_2455 (O_2455,N_24962,N_24865);
nor UO_2456 (O_2456,N_24938,N_24918);
nand UO_2457 (O_2457,N_24974,N_24903);
xor UO_2458 (O_2458,N_24994,N_24817);
xnor UO_2459 (O_2459,N_24847,N_24958);
xor UO_2460 (O_2460,N_24948,N_24899);
and UO_2461 (O_2461,N_24996,N_24926);
nor UO_2462 (O_2462,N_24867,N_24885);
and UO_2463 (O_2463,N_24932,N_24882);
xor UO_2464 (O_2464,N_24841,N_24838);
and UO_2465 (O_2465,N_24919,N_24965);
nor UO_2466 (O_2466,N_24906,N_24860);
nor UO_2467 (O_2467,N_24922,N_24965);
and UO_2468 (O_2468,N_24909,N_24978);
and UO_2469 (O_2469,N_24962,N_24981);
nor UO_2470 (O_2470,N_24834,N_24940);
or UO_2471 (O_2471,N_24951,N_24806);
nor UO_2472 (O_2472,N_24957,N_24896);
xnor UO_2473 (O_2473,N_24993,N_24929);
or UO_2474 (O_2474,N_24909,N_24806);
and UO_2475 (O_2475,N_24861,N_24928);
xor UO_2476 (O_2476,N_24801,N_24942);
nor UO_2477 (O_2477,N_24919,N_24872);
nand UO_2478 (O_2478,N_24917,N_24899);
or UO_2479 (O_2479,N_24897,N_24923);
xor UO_2480 (O_2480,N_24869,N_24980);
nand UO_2481 (O_2481,N_24852,N_24902);
and UO_2482 (O_2482,N_24809,N_24871);
xnor UO_2483 (O_2483,N_24943,N_24930);
xnor UO_2484 (O_2484,N_24922,N_24850);
and UO_2485 (O_2485,N_24855,N_24817);
nor UO_2486 (O_2486,N_24909,N_24985);
nand UO_2487 (O_2487,N_24832,N_24980);
nor UO_2488 (O_2488,N_24907,N_24951);
or UO_2489 (O_2489,N_24985,N_24997);
nor UO_2490 (O_2490,N_24911,N_24821);
or UO_2491 (O_2491,N_24812,N_24813);
and UO_2492 (O_2492,N_24966,N_24948);
nor UO_2493 (O_2493,N_24801,N_24886);
xor UO_2494 (O_2494,N_24915,N_24829);
or UO_2495 (O_2495,N_24900,N_24916);
nand UO_2496 (O_2496,N_24856,N_24976);
and UO_2497 (O_2497,N_24904,N_24918);
nand UO_2498 (O_2498,N_24991,N_24971);
xor UO_2499 (O_2499,N_24831,N_24850);
xnor UO_2500 (O_2500,N_24878,N_24982);
and UO_2501 (O_2501,N_24880,N_24945);
or UO_2502 (O_2502,N_24946,N_24828);
nor UO_2503 (O_2503,N_24894,N_24900);
nor UO_2504 (O_2504,N_24850,N_24975);
nor UO_2505 (O_2505,N_24996,N_24895);
nor UO_2506 (O_2506,N_24879,N_24896);
and UO_2507 (O_2507,N_24928,N_24908);
xor UO_2508 (O_2508,N_24848,N_24898);
nor UO_2509 (O_2509,N_24968,N_24818);
and UO_2510 (O_2510,N_24972,N_24964);
and UO_2511 (O_2511,N_24806,N_24851);
and UO_2512 (O_2512,N_24951,N_24933);
xor UO_2513 (O_2513,N_24832,N_24817);
xnor UO_2514 (O_2514,N_24862,N_24910);
nor UO_2515 (O_2515,N_24988,N_24846);
or UO_2516 (O_2516,N_24867,N_24914);
and UO_2517 (O_2517,N_24825,N_24828);
or UO_2518 (O_2518,N_24925,N_24996);
and UO_2519 (O_2519,N_24888,N_24819);
and UO_2520 (O_2520,N_24951,N_24996);
xnor UO_2521 (O_2521,N_24879,N_24882);
and UO_2522 (O_2522,N_24841,N_24807);
nor UO_2523 (O_2523,N_24821,N_24918);
nand UO_2524 (O_2524,N_24928,N_24822);
and UO_2525 (O_2525,N_24816,N_24934);
nand UO_2526 (O_2526,N_24836,N_24925);
nand UO_2527 (O_2527,N_24968,N_24900);
nor UO_2528 (O_2528,N_24988,N_24957);
or UO_2529 (O_2529,N_24978,N_24846);
or UO_2530 (O_2530,N_24933,N_24969);
and UO_2531 (O_2531,N_24840,N_24907);
and UO_2532 (O_2532,N_24923,N_24909);
nor UO_2533 (O_2533,N_24909,N_24933);
or UO_2534 (O_2534,N_24808,N_24916);
or UO_2535 (O_2535,N_24894,N_24961);
or UO_2536 (O_2536,N_24993,N_24898);
nor UO_2537 (O_2537,N_24978,N_24811);
nor UO_2538 (O_2538,N_24826,N_24992);
xnor UO_2539 (O_2539,N_24901,N_24829);
xor UO_2540 (O_2540,N_24835,N_24975);
and UO_2541 (O_2541,N_24864,N_24908);
nand UO_2542 (O_2542,N_24892,N_24926);
xor UO_2543 (O_2543,N_24971,N_24872);
nand UO_2544 (O_2544,N_24989,N_24996);
nor UO_2545 (O_2545,N_24955,N_24948);
and UO_2546 (O_2546,N_24926,N_24851);
and UO_2547 (O_2547,N_24809,N_24825);
or UO_2548 (O_2548,N_24815,N_24836);
or UO_2549 (O_2549,N_24847,N_24890);
nand UO_2550 (O_2550,N_24979,N_24940);
and UO_2551 (O_2551,N_24858,N_24885);
nor UO_2552 (O_2552,N_24958,N_24823);
nor UO_2553 (O_2553,N_24968,N_24960);
xnor UO_2554 (O_2554,N_24903,N_24977);
xnor UO_2555 (O_2555,N_24899,N_24831);
and UO_2556 (O_2556,N_24860,N_24857);
xor UO_2557 (O_2557,N_24890,N_24881);
nand UO_2558 (O_2558,N_24893,N_24847);
or UO_2559 (O_2559,N_24968,N_24884);
or UO_2560 (O_2560,N_24939,N_24936);
nand UO_2561 (O_2561,N_24948,N_24960);
nand UO_2562 (O_2562,N_24818,N_24809);
and UO_2563 (O_2563,N_24993,N_24870);
nand UO_2564 (O_2564,N_24833,N_24861);
or UO_2565 (O_2565,N_24974,N_24914);
nor UO_2566 (O_2566,N_24938,N_24802);
nor UO_2567 (O_2567,N_24845,N_24837);
or UO_2568 (O_2568,N_24940,N_24859);
or UO_2569 (O_2569,N_24923,N_24861);
or UO_2570 (O_2570,N_24948,N_24975);
nand UO_2571 (O_2571,N_24907,N_24847);
or UO_2572 (O_2572,N_24929,N_24996);
nor UO_2573 (O_2573,N_24890,N_24940);
or UO_2574 (O_2574,N_24849,N_24858);
nor UO_2575 (O_2575,N_24865,N_24935);
and UO_2576 (O_2576,N_24800,N_24817);
nand UO_2577 (O_2577,N_24825,N_24896);
xor UO_2578 (O_2578,N_24827,N_24982);
nor UO_2579 (O_2579,N_24985,N_24896);
or UO_2580 (O_2580,N_24928,N_24882);
xnor UO_2581 (O_2581,N_24822,N_24915);
or UO_2582 (O_2582,N_24984,N_24858);
nor UO_2583 (O_2583,N_24929,N_24815);
xor UO_2584 (O_2584,N_24832,N_24915);
nor UO_2585 (O_2585,N_24976,N_24936);
and UO_2586 (O_2586,N_24904,N_24930);
or UO_2587 (O_2587,N_24862,N_24828);
nor UO_2588 (O_2588,N_24976,N_24988);
nor UO_2589 (O_2589,N_24806,N_24871);
xor UO_2590 (O_2590,N_24980,N_24942);
or UO_2591 (O_2591,N_24873,N_24897);
or UO_2592 (O_2592,N_24867,N_24804);
nor UO_2593 (O_2593,N_24812,N_24923);
nand UO_2594 (O_2594,N_24950,N_24980);
nor UO_2595 (O_2595,N_24865,N_24815);
nand UO_2596 (O_2596,N_24891,N_24916);
and UO_2597 (O_2597,N_24990,N_24828);
and UO_2598 (O_2598,N_24992,N_24803);
or UO_2599 (O_2599,N_24933,N_24840);
or UO_2600 (O_2600,N_24966,N_24821);
nand UO_2601 (O_2601,N_24802,N_24817);
nand UO_2602 (O_2602,N_24869,N_24963);
nand UO_2603 (O_2603,N_24897,N_24859);
xnor UO_2604 (O_2604,N_24913,N_24821);
or UO_2605 (O_2605,N_24871,N_24821);
nand UO_2606 (O_2606,N_24883,N_24995);
or UO_2607 (O_2607,N_24842,N_24936);
nand UO_2608 (O_2608,N_24861,N_24855);
nand UO_2609 (O_2609,N_24859,N_24984);
and UO_2610 (O_2610,N_24955,N_24814);
nor UO_2611 (O_2611,N_24915,N_24824);
or UO_2612 (O_2612,N_24847,N_24881);
nor UO_2613 (O_2613,N_24997,N_24980);
nor UO_2614 (O_2614,N_24838,N_24997);
xnor UO_2615 (O_2615,N_24990,N_24809);
xor UO_2616 (O_2616,N_24922,N_24962);
nand UO_2617 (O_2617,N_24842,N_24879);
nand UO_2618 (O_2618,N_24841,N_24905);
and UO_2619 (O_2619,N_24931,N_24879);
xnor UO_2620 (O_2620,N_24924,N_24894);
or UO_2621 (O_2621,N_24897,N_24915);
nand UO_2622 (O_2622,N_24906,N_24896);
nor UO_2623 (O_2623,N_24962,N_24996);
nor UO_2624 (O_2624,N_24861,N_24806);
nor UO_2625 (O_2625,N_24844,N_24829);
nor UO_2626 (O_2626,N_24903,N_24889);
or UO_2627 (O_2627,N_24997,N_24882);
nor UO_2628 (O_2628,N_24898,N_24850);
xor UO_2629 (O_2629,N_24955,N_24959);
and UO_2630 (O_2630,N_24978,N_24810);
nand UO_2631 (O_2631,N_24869,N_24854);
nor UO_2632 (O_2632,N_24853,N_24828);
nand UO_2633 (O_2633,N_24905,N_24916);
and UO_2634 (O_2634,N_24836,N_24839);
or UO_2635 (O_2635,N_24871,N_24848);
nor UO_2636 (O_2636,N_24928,N_24974);
and UO_2637 (O_2637,N_24897,N_24916);
nor UO_2638 (O_2638,N_24836,N_24917);
nor UO_2639 (O_2639,N_24837,N_24824);
nor UO_2640 (O_2640,N_24801,N_24867);
nand UO_2641 (O_2641,N_24988,N_24903);
or UO_2642 (O_2642,N_24880,N_24848);
xnor UO_2643 (O_2643,N_24921,N_24955);
or UO_2644 (O_2644,N_24826,N_24915);
and UO_2645 (O_2645,N_24912,N_24920);
xnor UO_2646 (O_2646,N_24997,N_24835);
xor UO_2647 (O_2647,N_24954,N_24916);
or UO_2648 (O_2648,N_24942,N_24926);
xnor UO_2649 (O_2649,N_24930,N_24907);
or UO_2650 (O_2650,N_24852,N_24811);
nand UO_2651 (O_2651,N_24943,N_24846);
and UO_2652 (O_2652,N_24885,N_24976);
or UO_2653 (O_2653,N_24884,N_24802);
xnor UO_2654 (O_2654,N_24985,N_24974);
nor UO_2655 (O_2655,N_24800,N_24842);
nor UO_2656 (O_2656,N_24906,N_24974);
xor UO_2657 (O_2657,N_24903,N_24861);
xnor UO_2658 (O_2658,N_24821,N_24872);
or UO_2659 (O_2659,N_24933,N_24881);
and UO_2660 (O_2660,N_24817,N_24882);
or UO_2661 (O_2661,N_24927,N_24874);
nand UO_2662 (O_2662,N_24825,N_24972);
nor UO_2663 (O_2663,N_24955,N_24913);
nand UO_2664 (O_2664,N_24986,N_24829);
and UO_2665 (O_2665,N_24811,N_24887);
nand UO_2666 (O_2666,N_24937,N_24901);
nand UO_2667 (O_2667,N_24939,N_24855);
and UO_2668 (O_2668,N_24837,N_24989);
and UO_2669 (O_2669,N_24963,N_24991);
xor UO_2670 (O_2670,N_24822,N_24887);
or UO_2671 (O_2671,N_24823,N_24982);
and UO_2672 (O_2672,N_24910,N_24892);
nor UO_2673 (O_2673,N_24902,N_24949);
or UO_2674 (O_2674,N_24954,N_24848);
and UO_2675 (O_2675,N_24900,N_24829);
xor UO_2676 (O_2676,N_24971,N_24886);
or UO_2677 (O_2677,N_24829,N_24814);
and UO_2678 (O_2678,N_24844,N_24867);
nand UO_2679 (O_2679,N_24908,N_24879);
nor UO_2680 (O_2680,N_24820,N_24974);
xor UO_2681 (O_2681,N_24879,N_24977);
xor UO_2682 (O_2682,N_24922,N_24972);
or UO_2683 (O_2683,N_24851,N_24935);
and UO_2684 (O_2684,N_24888,N_24988);
nand UO_2685 (O_2685,N_24954,N_24925);
nor UO_2686 (O_2686,N_24810,N_24982);
or UO_2687 (O_2687,N_24811,N_24982);
nor UO_2688 (O_2688,N_24869,N_24850);
xnor UO_2689 (O_2689,N_24988,N_24854);
or UO_2690 (O_2690,N_24822,N_24911);
nor UO_2691 (O_2691,N_24965,N_24880);
nand UO_2692 (O_2692,N_24954,N_24857);
xor UO_2693 (O_2693,N_24888,N_24929);
nor UO_2694 (O_2694,N_24917,N_24988);
nand UO_2695 (O_2695,N_24928,N_24812);
and UO_2696 (O_2696,N_24919,N_24964);
nor UO_2697 (O_2697,N_24814,N_24986);
or UO_2698 (O_2698,N_24807,N_24899);
and UO_2699 (O_2699,N_24842,N_24929);
nor UO_2700 (O_2700,N_24913,N_24884);
or UO_2701 (O_2701,N_24948,N_24962);
nor UO_2702 (O_2702,N_24824,N_24934);
nor UO_2703 (O_2703,N_24898,N_24893);
nand UO_2704 (O_2704,N_24840,N_24985);
nor UO_2705 (O_2705,N_24861,N_24881);
xnor UO_2706 (O_2706,N_24839,N_24998);
nand UO_2707 (O_2707,N_24847,N_24834);
and UO_2708 (O_2708,N_24969,N_24971);
nand UO_2709 (O_2709,N_24828,N_24902);
nand UO_2710 (O_2710,N_24947,N_24825);
xnor UO_2711 (O_2711,N_24923,N_24980);
or UO_2712 (O_2712,N_24990,N_24864);
nor UO_2713 (O_2713,N_24849,N_24838);
nor UO_2714 (O_2714,N_24995,N_24807);
nand UO_2715 (O_2715,N_24889,N_24850);
or UO_2716 (O_2716,N_24800,N_24885);
and UO_2717 (O_2717,N_24926,N_24934);
nand UO_2718 (O_2718,N_24967,N_24893);
xnor UO_2719 (O_2719,N_24958,N_24800);
or UO_2720 (O_2720,N_24919,N_24981);
nand UO_2721 (O_2721,N_24858,N_24960);
xnor UO_2722 (O_2722,N_24818,N_24918);
or UO_2723 (O_2723,N_24864,N_24855);
or UO_2724 (O_2724,N_24836,N_24843);
nor UO_2725 (O_2725,N_24832,N_24964);
or UO_2726 (O_2726,N_24834,N_24870);
nand UO_2727 (O_2727,N_24811,N_24951);
xnor UO_2728 (O_2728,N_24825,N_24827);
and UO_2729 (O_2729,N_24867,N_24977);
nor UO_2730 (O_2730,N_24884,N_24925);
nand UO_2731 (O_2731,N_24972,N_24859);
or UO_2732 (O_2732,N_24974,N_24817);
nor UO_2733 (O_2733,N_24917,N_24957);
nand UO_2734 (O_2734,N_24845,N_24914);
xor UO_2735 (O_2735,N_24900,N_24858);
and UO_2736 (O_2736,N_24969,N_24862);
or UO_2737 (O_2737,N_24895,N_24966);
xor UO_2738 (O_2738,N_24981,N_24976);
xor UO_2739 (O_2739,N_24874,N_24960);
xnor UO_2740 (O_2740,N_24985,N_24852);
xnor UO_2741 (O_2741,N_24865,N_24964);
xnor UO_2742 (O_2742,N_24970,N_24935);
nand UO_2743 (O_2743,N_24971,N_24973);
and UO_2744 (O_2744,N_24904,N_24951);
xnor UO_2745 (O_2745,N_24800,N_24917);
xor UO_2746 (O_2746,N_24801,N_24814);
and UO_2747 (O_2747,N_24906,N_24861);
nor UO_2748 (O_2748,N_24847,N_24841);
xnor UO_2749 (O_2749,N_24906,N_24927);
nor UO_2750 (O_2750,N_24999,N_24939);
or UO_2751 (O_2751,N_24888,N_24946);
nor UO_2752 (O_2752,N_24845,N_24938);
nor UO_2753 (O_2753,N_24946,N_24885);
xor UO_2754 (O_2754,N_24809,N_24844);
and UO_2755 (O_2755,N_24925,N_24879);
or UO_2756 (O_2756,N_24901,N_24944);
xnor UO_2757 (O_2757,N_24990,N_24832);
nor UO_2758 (O_2758,N_24823,N_24899);
xor UO_2759 (O_2759,N_24851,N_24856);
nand UO_2760 (O_2760,N_24853,N_24966);
nand UO_2761 (O_2761,N_24881,N_24874);
nor UO_2762 (O_2762,N_24857,N_24984);
nand UO_2763 (O_2763,N_24971,N_24880);
nand UO_2764 (O_2764,N_24891,N_24952);
or UO_2765 (O_2765,N_24805,N_24837);
and UO_2766 (O_2766,N_24918,N_24895);
nand UO_2767 (O_2767,N_24914,N_24853);
nand UO_2768 (O_2768,N_24885,N_24843);
nor UO_2769 (O_2769,N_24895,N_24885);
or UO_2770 (O_2770,N_24811,N_24956);
nand UO_2771 (O_2771,N_24957,N_24933);
or UO_2772 (O_2772,N_24817,N_24991);
nor UO_2773 (O_2773,N_24964,N_24967);
and UO_2774 (O_2774,N_24953,N_24998);
nor UO_2775 (O_2775,N_24808,N_24935);
or UO_2776 (O_2776,N_24868,N_24827);
or UO_2777 (O_2777,N_24834,N_24825);
or UO_2778 (O_2778,N_24886,N_24988);
xor UO_2779 (O_2779,N_24836,N_24864);
nor UO_2780 (O_2780,N_24997,N_24843);
nand UO_2781 (O_2781,N_24863,N_24874);
xor UO_2782 (O_2782,N_24939,N_24927);
nor UO_2783 (O_2783,N_24814,N_24965);
xnor UO_2784 (O_2784,N_24952,N_24973);
or UO_2785 (O_2785,N_24825,N_24904);
or UO_2786 (O_2786,N_24985,N_24847);
or UO_2787 (O_2787,N_24854,N_24907);
nand UO_2788 (O_2788,N_24976,N_24844);
or UO_2789 (O_2789,N_24801,N_24828);
nand UO_2790 (O_2790,N_24915,N_24924);
xnor UO_2791 (O_2791,N_24826,N_24819);
xor UO_2792 (O_2792,N_24882,N_24938);
or UO_2793 (O_2793,N_24929,N_24851);
xnor UO_2794 (O_2794,N_24862,N_24856);
nand UO_2795 (O_2795,N_24823,N_24912);
or UO_2796 (O_2796,N_24833,N_24852);
nand UO_2797 (O_2797,N_24939,N_24947);
and UO_2798 (O_2798,N_24918,N_24839);
nor UO_2799 (O_2799,N_24916,N_24936);
and UO_2800 (O_2800,N_24877,N_24924);
and UO_2801 (O_2801,N_24804,N_24865);
or UO_2802 (O_2802,N_24849,N_24992);
xnor UO_2803 (O_2803,N_24814,N_24881);
and UO_2804 (O_2804,N_24806,N_24811);
or UO_2805 (O_2805,N_24982,N_24928);
xnor UO_2806 (O_2806,N_24890,N_24935);
and UO_2807 (O_2807,N_24868,N_24935);
or UO_2808 (O_2808,N_24991,N_24907);
xor UO_2809 (O_2809,N_24951,N_24973);
nand UO_2810 (O_2810,N_24928,N_24970);
or UO_2811 (O_2811,N_24957,N_24863);
nand UO_2812 (O_2812,N_24998,N_24830);
and UO_2813 (O_2813,N_24945,N_24974);
nor UO_2814 (O_2814,N_24847,N_24926);
or UO_2815 (O_2815,N_24937,N_24802);
nand UO_2816 (O_2816,N_24836,N_24878);
and UO_2817 (O_2817,N_24891,N_24861);
nand UO_2818 (O_2818,N_24956,N_24845);
or UO_2819 (O_2819,N_24886,N_24934);
and UO_2820 (O_2820,N_24871,N_24920);
or UO_2821 (O_2821,N_24970,N_24920);
and UO_2822 (O_2822,N_24806,N_24935);
or UO_2823 (O_2823,N_24897,N_24861);
and UO_2824 (O_2824,N_24847,N_24951);
or UO_2825 (O_2825,N_24894,N_24913);
and UO_2826 (O_2826,N_24997,N_24839);
nor UO_2827 (O_2827,N_24878,N_24927);
nand UO_2828 (O_2828,N_24961,N_24913);
nor UO_2829 (O_2829,N_24801,N_24907);
and UO_2830 (O_2830,N_24929,N_24984);
xor UO_2831 (O_2831,N_24911,N_24815);
and UO_2832 (O_2832,N_24849,N_24875);
nor UO_2833 (O_2833,N_24905,N_24857);
or UO_2834 (O_2834,N_24946,N_24927);
xor UO_2835 (O_2835,N_24986,N_24933);
or UO_2836 (O_2836,N_24826,N_24957);
xnor UO_2837 (O_2837,N_24959,N_24880);
nor UO_2838 (O_2838,N_24907,N_24952);
or UO_2839 (O_2839,N_24867,N_24928);
nand UO_2840 (O_2840,N_24968,N_24926);
or UO_2841 (O_2841,N_24870,N_24895);
and UO_2842 (O_2842,N_24938,N_24992);
nor UO_2843 (O_2843,N_24990,N_24884);
xnor UO_2844 (O_2844,N_24834,N_24902);
nor UO_2845 (O_2845,N_24819,N_24843);
or UO_2846 (O_2846,N_24940,N_24842);
and UO_2847 (O_2847,N_24982,N_24952);
or UO_2848 (O_2848,N_24896,N_24990);
nor UO_2849 (O_2849,N_24891,N_24841);
or UO_2850 (O_2850,N_24811,N_24974);
xnor UO_2851 (O_2851,N_24800,N_24882);
nor UO_2852 (O_2852,N_24837,N_24904);
nand UO_2853 (O_2853,N_24933,N_24931);
nand UO_2854 (O_2854,N_24852,N_24819);
and UO_2855 (O_2855,N_24891,N_24984);
and UO_2856 (O_2856,N_24898,N_24846);
xnor UO_2857 (O_2857,N_24981,N_24825);
and UO_2858 (O_2858,N_24856,N_24900);
or UO_2859 (O_2859,N_24929,N_24810);
nor UO_2860 (O_2860,N_24915,N_24962);
xnor UO_2861 (O_2861,N_24848,N_24824);
xor UO_2862 (O_2862,N_24997,N_24803);
nand UO_2863 (O_2863,N_24900,N_24878);
and UO_2864 (O_2864,N_24851,N_24901);
or UO_2865 (O_2865,N_24833,N_24801);
nor UO_2866 (O_2866,N_24954,N_24880);
xor UO_2867 (O_2867,N_24835,N_24865);
nor UO_2868 (O_2868,N_24938,N_24800);
nor UO_2869 (O_2869,N_24976,N_24894);
and UO_2870 (O_2870,N_24907,N_24908);
or UO_2871 (O_2871,N_24975,N_24987);
and UO_2872 (O_2872,N_24837,N_24918);
nor UO_2873 (O_2873,N_24867,N_24830);
xnor UO_2874 (O_2874,N_24930,N_24867);
nand UO_2875 (O_2875,N_24811,N_24843);
nand UO_2876 (O_2876,N_24852,N_24821);
nand UO_2877 (O_2877,N_24953,N_24974);
nand UO_2878 (O_2878,N_24914,N_24834);
nand UO_2879 (O_2879,N_24983,N_24942);
or UO_2880 (O_2880,N_24874,N_24976);
nor UO_2881 (O_2881,N_24835,N_24868);
or UO_2882 (O_2882,N_24960,N_24870);
xnor UO_2883 (O_2883,N_24962,N_24875);
or UO_2884 (O_2884,N_24926,N_24864);
xnor UO_2885 (O_2885,N_24892,N_24958);
nor UO_2886 (O_2886,N_24852,N_24883);
and UO_2887 (O_2887,N_24844,N_24875);
or UO_2888 (O_2888,N_24887,N_24817);
nand UO_2889 (O_2889,N_24964,N_24836);
or UO_2890 (O_2890,N_24954,N_24871);
nor UO_2891 (O_2891,N_24973,N_24978);
nor UO_2892 (O_2892,N_24983,N_24988);
nor UO_2893 (O_2893,N_24948,N_24892);
xnor UO_2894 (O_2894,N_24979,N_24991);
xor UO_2895 (O_2895,N_24880,N_24964);
xor UO_2896 (O_2896,N_24969,N_24836);
or UO_2897 (O_2897,N_24812,N_24988);
or UO_2898 (O_2898,N_24966,N_24809);
or UO_2899 (O_2899,N_24907,N_24815);
nand UO_2900 (O_2900,N_24989,N_24825);
or UO_2901 (O_2901,N_24817,N_24834);
nand UO_2902 (O_2902,N_24926,N_24972);
nand UO_2903 (O_2903,N_24865,N_24819);
or UO_2904 (O_2904,N_24864,N_24853);
and UO_2905 (O_2905,N_24864,N_24914);
xnor UO_2906 (O_2906,N_24909,N_24815);
nand UO_2907 (O_2907,N_24931,N_24961);
and UO_2908 (O_2908,N_24913,N_24904);
xor UO_2909 (O_2909,N_24909,N_24838);
or UO_2910 (O_2910,N_24922,N_24868);
nand UO_2911 (O_2911,N_24857,N_24913);
and UO_2912 (O_2912,N_24807,N_24926);
nor UO_2913 (O_2913,N_24822,N_24942);
nor UO_2914 (O_2914,N_24994,N_24893);
xor UO_2915 (O_2915,N_24871,N_24856);
xor UO_2916 (O_2916,N_24925,N_24861);
and UO_2917 (O_2917,N_24842,N_24943);
or UO_2918 (O_2918,N_24982,N_24939);
and UO_2919 (O_2919,N_24919,N_24891);
nand UO_2920 (O_2920,N_24892,N_24890);
xnor UO_2921 (O_2921,N_24874,N_24896);
xnor UO_2922 (O_2922,N_24851,N_24896);
xor UO_2923 (O_2923,N_24906,N_24852);
xor UO_2924 (O_2924,N_24903,N_24838);
and UO_2925 (O_2925,N_24963,N_24986);
nand UO_2926 (O_2926,N_24991,N_24985);
and UO_2927 (O_2927,N_24831,N_24944);
or UO_2928 (O_2928,N_24857,N_24863);
or UO_2929 (O_2929,N_24804,N_24944);
and UO_2930 (O_2930,N_24844,N_24949);
xor UO_2931 (O_2931,N_24880,N_24907);
nand UO_2932 (O_2932,N_24800,N_24987);
nand UO_2933 (O_2933,N_24918,N_24908);
nand UO_2934 (O_2934,N_24945,N_24806);
or UO_2935 (O_2935,N_24996,N_24886);
xor UO_2936 (O_2936,N_24848,N_24958);
and UO_2937 (O_2937,N_24927,N_24979);
xor UO_2938 (O_2938,N_24881,N_24963);
xnor UO_2939 (O_2939,N_24815,N_24955);
xor UO_2940 (O_2940,N_24861,N_24913);
xnor UO_2941 (O_2941,N_24873,N_24968);
nand UO_2942 (O_2942,N_24992,N_24998);
nor UO_2943 (O_2943,N_24953,N_24917);
xor UO_2944 (O_2944,N_24849,N_24971);
nor UO_2945 (O_2945,N_24810,N_24873);
nand UO_2946 (O_2946,N_24865,N_24843);
xor UO_2947 (O_2947,N_24862,N_24880);
xor UO_2948 (O_2948,N_24875,N_24980);
and UO_2949 (O_2949,N_24960,N_24859);
nand UO_2950 (O_2950,N_24985,N_24975);
or UO_2951 (O_2951,N_24864,N_24828);
nor UO_2952 (O_2952,N_24917,N_24946);
and UO_2953 (O_2953,N_24984,N_24854);
or UO_2954 (O_2954,N_24919,N_24916);
nor UO_2955 (O_2955,N_24994,N_24998);
or UO_2956 (O_2956,N_24874,N_24977);
nand UO_2957 (O_2957,N_24928,N_24907);
nand UO_2958 (O_2958,N_24921,N_24994);
xor UO_2959 (O_2959,N_24882,N_24860);
xnor UO_2960 (O_2960,N_24803,N_24875);
nand UO_2961 (O_2961,N_24857,N_24890);
or UO_2962 (O_2962,N_24996,N_24921);
or UO_2963 (O_2963,N_24991,N_24899);
or UO_2964 (O_2964,N_24859,N_24954);
and UO_2965 (O_2965,N_24831,N_24937);
nor UO_2966 (O_2966,N_24922,N_24849);
nand UO_2967 (O_2967,N_24921,N_24928);
or UO_2968 (O_2968,N_24854,N_24940);
and UO_2969 (O_2969,N_24945,N_24891);
and UO_2970 (O_2970,N_24820,N_24870);
nand UO_2971 (O_2971,N_24958,N_24895);
or UO_2972 (O_2972,N_24801,N_24972);
and UO_2973 (O_2973,N_24924,N_24984);
or UO_2974 (O_2974,N_24946,N_24992);
and UO_2975 (O_2975,N_24813,N_24955);
xor UO_2976 (O_2976,N_24985,N_24926);
and UO_2977 (O_2977,N_24965,N_24882);
nor UO_2978 (O_2978,N_24918,N_24931);
or UO_2979 (O_2979,N_24829,N_24859);
or UO_2980 (O_2980,N_24954,N_24824);
nand UO_2981 (O_2981,N_24811,N_24985);
nand UO_2982 (O_2982,N_24800,N_24833);
and UO_2983 (O_2983,N_24916,N_24853);
and UO_2984 (O_2984,N_24963,N_24904);
xor UO_2985 (O_2985,N_24869,N_24924);
nand UO_2986 (O_2986,N_24904,N_24827);
xor UO_2987 (O_2987,N_24892,N_24818);
nor UO_2988 (O_2988,N_24979,N_24999);
and UO_2989 (O_2989,N_24916,N_24895);
xnor UO_2990 (O_2990,N_24973,N_24914);
nand UO_2991 (O_2991,N_24991,N_24944);
nor UO_2992 (O_2992,N_24884,N_24987);
and UO_2993 (O_2993,N_24908,N_24977);
nor UO_2994 (O_2994,N_24965,N_24841);
nand UO_2995 (O_2995,N_24996,N_24923);
or UO_2996 (O_2996,N_24968,N_24811);
and UO_2997 (O_2997,N_24878,N_24943);
nand UO_2998 (O_2998,N_24919,N_24878);
and UO_2999 (O_2999,N_24902,N_24967);
endmodule