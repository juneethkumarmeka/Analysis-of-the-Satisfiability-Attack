module basic_750_5000_1000_10_levels_10xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
nor U0 (N_0,In_22,In_151);
nand U1 (N_1,In_442,In_309);
nand U2 (N_2,In_488,In_297);
or U3 (N_3,In_667,In_703);
or U4 (N_4,In_135,In_199);
nor U5 (N_5,In_456,In_547);
xnor U6 (N_6,In_458,In_330);
nor U7 (N_7,In_450,In_7);
xnor U8 (N_8,In_413,In_747);
or U9 (N_9,In_497,In_108);
xnor U10 (N_10,In_736,In_167);
nand U11 (N_11,In_666,In_709);
nand U12 (N_12,In_604,In_229);
or U13 (N_13,In_144,In_624);
nor U14 (N_14,In_725,In_274);
nand U15 (N_15,In_618,In_18);
or U16 (N_16,In_341,In_622);
nand U17 (N_17,In_401,In_690);
nor U18 (N_18,In_556,In_188);
xor U19 (N_19,In_222,In_143);
xnor U20 (N_20,In_524,In_6);
nand U21 (N_21,In_223,In_14);
or U22 (N_22,In_713,In_501);
or U23 (N_23,In_321,In_688);
or U24 (N_24,In_452,In_418);
nand U25 (N_25,In_294,In_338);
xor U26 (N_26,In_724,In_68);
xnor U27 (N_27,In_555,In_179);
nand U28 (N_28,In_308,In_138);
nor U29 (N_29,In_689,In_708);
xor U30 (N_30,In_592,In_542);
and U31 (N_31,In_496,In_665);
and U32 (N_32,In_124,In_640);
xor U33 (N_33,In_739,In_517);
xor U34 (N_34,In_216,In_370);
xor U35 (N_35,In_516,In_212);
or U36 (N_36,In_293,In_434);
nand U37 (N_37,In_148,In_656);
and U38 (N_38,In_535,In_530);
nor U39 (N_39,In_463,In_11);
and U40 (N_40,In_489,In_61);
xor U41 (N_41,In_340,In_186);
and U42 (N_42,In_596,In_625);
xnor U43 (N_43,In_176,In_173);
or U44 (N_44,In_66,In_242);
or U45 (N_45,In_393,In_718);
nand U46 (N_46,In_500,In_270);
or U47 (N_47,In_553,In_634);
nand U48 (N_48,In_78,In_268);
nand U49 (N_49,In_165,In_443);
xor U50 (N_50,In_280,In_379);
nand U51 (N_51,In_470,In_531);
and U52 (N_52,In_390,In_536);
and U53 (N_53,In_244,In_64);
nand U54 (N_54,In_552,In_210);
xor U55 (N_55,In_478,In_17);
or U56 (N_56,In_55,In_142);
nand U57 (N_57,In_544,In_363);
or U58 (N_58,In_183,In_473);
nand U59 (N_59,In_355,In_594);
nand U60 (N_60,In_91,In_70);
or U61 (N_61,In_372,In_217);
xnor U62 (N_62,In_324,In_349);
nor U63 (N_63,In_354,In_570);
nor U64 (N_64,In_737,In_661);
and U65 (N_65,In_684,In_482);
nor U66 (N_66,In_265,In_518);
or U67 (N_67,In_284,In_331);
nand U68 (N_68,In_520,In_56);
xnor U69 (N_69,In_360,In_662);
xor U70 (N_70,In_352,In_735);
or U71 (N_71,In_484,In_712);
xor U72 (N_72,In_146,In_700);
nand U73 (N_73,In_749,In_566);
nand U74 (N_74,In_261,In_203);
nor U75 (N_75,In_691,In_441);
nand U76 (N_76,In_638,In_546);
and U77 (N_77,In_136,In_494);
or U78 (N_78,In_333,In_527);
nor U79 (N_79,In_499,In_278);
nand U80 (N_80,In_522,In_586);
xnor U81 (N_81,In_112,In_342);
or U82 (N_82,In_400,In_502);
nand U83 (N_83,In_741,In_402);
nand U84 (N_84,In_600,In_587);
and U85 (N_85,In_632,In_164);
xor U86 (N_86,In_163,In_271);
nand U87 (N_87,In_433,In_562);
xnor U88 (N_88,In_62,In_15);
or U89 (N_89,In_475,In_710);
xor U90 (N_90,In_436,In_344);
nand U91 (N_91,In_234,In_351);
xnor U92 (N_92,In_246,In_481);
or U93 (N_93,In_579,In_512);
nor U94 (N_94,In_446,In_157);
nand U95 (N_95,In_744,In_235);
or U96 (N_96,In_748,In_40);
nand U97 (N_97,In_541,In_154);
or U98 (N_98,In_384,In_394);
or U99 (N_99,In_30,In_564);
and U100 (N_100,In_723,In_162);
nand U101 (N_101,In_629,In_707);
xnor U102 (N_102,In_730,In_651);
or U103 (N_103,In_514,In_362);
or U104 (N_104,In_83,In_699);
nor U105 (N_105,In_540,In_715);
xor U106 (N_106,In_606,In_399);
nand U107 (N_107,In_589,In_13);
xnor U108 (N_108,In_187,In_539);
nor U109 (N_109,In_155,In_357);
nor U110 (N_110,In_51,In_609);
or U111 (N_111,In_576,In_490);
and U112 (N_112,In_75,In_716);
and U113 (N_113,In_406,In_134);
nand U114 (N_114,In_277,In_122);
and U115 (N_115,In_693,In_27);
nor U116 (N_116,In_103,In_407);
or U117 (N_117,In_664,In_746);
nor U118 (N_118,In_578,In_272);
nand U119 (N_119,In_291,In_358);
xor U120 (N_120,In_639,In_137);
nand U121 (N_121,In_161,In_171);
nand U122 (N_122,In_314,In_230);
xnor U123 (N_123,In_595,In_461);
nand U124 (N_124,In_419,In_53);
nand U125 (N_125,In_695,In_100);
nor U126 (N_126,In_237,In_104);
nand U127 (N_127,In_559,In_109);
nor U128 (N_128,In_87,In_0);
nand U129 (N_129,In_335,In_300);
and U130 (N_130,In_416,In_410);
and U131 (N_131,In_571,In_114);
nor U132 (N_132,In_677,In_367);
and U133 (N_133,In_431,In_37);
nor U134 (N_134,In_649,In_282);
xnor U135 (N_135,In_254,In_637);
nor U136 (N_136,In_125,In_660);
and U137 (N_137,In_567,In_249);
or U138 (N_138,In_510,In_126);
nand U139 (N_139,In_616,In_474);
and U140 (N_140,In_86,In_425);
and U141 (N_141,In_185,In_224);
and U142 (N_142,In_213,In_597);
or U143 (N_143,In_658,In_46);
and U144 (N_144,In_580,In_591);
xnor U145 (N_145,In_375,In_380);
xor U146 (N_146,In_529,In_371);
xnor U147 (N_147,In_285,In_159);
nand U148 (N_148,In_655,In_459);
nor U149 (N_149,In_287,In_593);
nand U150 (N_150,In_356,In_194);
and U151 (N_151,In_275,In_376);
nand U152 (N_152,In_449,In_267);
xnor U153 (N_153,In_334,In_117);
and U154 (N_154,In_192,In_728);
nor U155 (N_155,In_588,In_545);
xnor U156 (N_156,In_263,In_603);
nand U157 (N_157,In_727,In_428);
or U158 (N_158,In_430,In_264);
xnor U159 (N_159,In_647,In_534);
and U160 (N_160,In_209,In_694);
or U161 (N_161,In_153,In_605);
and U162 (N_162,In_184,In_558);
and U163 (N_163,In_628,In_472);
and U164 (N_164,In_92,In_692);
nand U165 (N_165,In_311,In_361);
xnor U166 (N_166,In_438,In_110);
xor U167 (N_167,In_644,In_627);
or U168 (N_168,In_598,In_633);
nand U169 (N_169,In_160,In_641);
and U170 (N_170,In_49,In_455);
nor U171 (N_171,In_601,In_615);
or U172 (N_172,In_387,In_9);
and U173 (N_173,In_674,In_672);
nor U174 (N_174,In_421,In_584);
and U175 (N_175,In_181,In_320);
and U176 (N_176,In_528,In_717);
nor U177 (N_177,In_635,In_123);
xor U178 (N_178,In_396,In_328);
and U179 (N_179,In_670,In_317);
and U180 (N_180,In_140,In_424);
or U181 (N_181,In_669,In_479);
nand U182 (N_182,In_648,In_326);
nor U183 (N_183,In_548,In_602);
nor U184 (N_184,In_156,In_610);
and U185 (N_185,In_2,In_706);
and U186 (N_186,In_65,In_303);
nor U187 (N_187,In_130,In_630);
nand U188 (N_188,In_74,In_513);
xor U189 (N_189,In_292,In_733);
or U190 (N_190,In_286,In_28);
nor U191 (N_191,In_585,In_169);
xor U192 (N_192,In_437,In_107);
nand U193 (N_193,In_671,In_683);
and U194 (N_194,In_581,In_197);
nor U195 (N_195,In_368,In_133);
nor U196 (N_196,In_57,In_582);
nor U197 (N_197,In_705,In_668);
and U198 (N_198,In_118,In_139);
nor U199 (N_199,In_503,In_734);
nor U200 (N_200,In_205,In_221);
xor U201 (N_201,In_69,In_636);
nand U202 (N_202,In_247,In_374);
nand U203 (N_203,In_127,In_623);
and U204 (N_204,In_20,In_557);
xnor U205 (N_205,In_397,In_200);
nor U206 (N_206,In_572,In_283);
and U207 (N_207,In_208,In_8);
or U208 (N_208,In_532,In_432);
or U209 (N_209,In_676,In_238);
or U210 (N_210,In_266,In_462);
xor U211 (N_211,In_621,In_190);
xnor U212 (N_212,In_526,In_533);
xnor U213 (N_213,In_31,In_332);
nand U214 (N_214,In_289,In_339);
nor U215 (N_215,In_619,In_345);
or U216 (N_216,In_177,In_93);
nor U217 (N_217,In_697,In_422);
or U218 (N_218,In_214,In_701);
nor U219 (N_219,In_369,In_409);
nand U220 (N_220,In_465,In_231);
nor U221 (N_221,In_98,In_131);
or U222 (N_222,In_411,In_395);
and U223 (N_223,In_732,In_505);
xor U224 (N_224,In_236,In_611);
or U225 (N_225,In_454,In_195);
xnor U226 (N_226,In_714,In_202);
nor U227 (N_227,In_679,In_304);
nand U228 (N_228,In_85,In_113);
xnor U229 (N_229,In_152,In_412);
or U230 (N_230,In_43,In_141);
xor U231 (N_231,In_25,In_511);
or U232 (N_232,In_302,In_73);
nor U233 (N_233,In_486,In_175);
and U234 (N_234,In_464,In_1);
or U235 (N_235,In_241,In_48);
nand U236 (N_236,In_523,In_81);
xor U237 (N_237,In_239,In_329);
xor U238 (N_238,In_573,In_269);
nor U239 (N_239,In_398,In_240);
or U240 (N_240,In_495,In_39);
nand U241 (N_241,In_740,In_702);
nor U242 (N_242,In_569,In_415);
nand U243 (N_243,In_742,In_346);
nand U244 (N_244,In_71,In_719);
and U245 (N_245,In_276,In_642);
nor U246 (N_246,In_687,In_226);
xnor U247 (N_247,In_408,In_206);
nor U248 (N_248,In_453,In_439);
or U249 (N_249,In_312,In_467);
and U250 (N_250,In_696,In_307);
or U251 (N_251,In_211,In_166);
nor U252 (N_252,In_391,In_720);
and U253 (N_253,In_299,In_5);
and U254 (N_254,In_279,In_215);
and U255 (N_255,In_132,In_322);
xnor U256 (N_256,In_353,In_575);
nor U257 (N_257,In_417,In_233);
or U258 (N_258,In_172,In_493);
nand U259 (N_259,In_426,In_451);
nor U260 (N_260,In_498,In_617);
nand U261 (N_261,In_568,In_471);
xnor U262 (N_262,In_201,In_77);
and U263 (N_263,In_318,In_32);
nand U264 (N_264,In_225,In_631);
and U265 (N_265,In_469,In_301);
nand U266 (N_266,In_207,In_52);
xnor U267 (N_267,In_743,In_180);
xor U268 (N_268,In_613,In_305);
xnor U269 (N_269,In_577,In_158);
nor U270 (N_270,In_256,In_681);
xor U271 (N_271,In_366,In_21);
or U272 (N_272,In_650,In_435);
or U273 (N_273,In_405,In_698);
xor U274 (N_274,In_41,In_348);
and U275 (N_275,In_248,In_359);
or U276 (N_276,In_738,In_383);
nand U277 (N_277,In_128,In_504);
or U278 (N_278,In_258,In_457);
or U279 (N_279,In_445,In_54);
and U280 (N_280,In_614,In_508);
xor U281 (N_281,In_47,In_96);
nor U282 (N_282,In_89,In_336);
xnor U283 (N_283,In_227,In_364);
nor U284 (N_284,In_4,In_659);
and U285 (N_285,In_560,In_382);
xnor U286 (N_286,In_440,In_319);
nand U287 (N_287,In_347,In_33);
nand U288 (N_288,In_704,In_88);
xnor U289 (N_289,In_257,In_24);
nor U290 (N_290,In_76,In_444);
and U291 (N_291,In_466,In_515);
nor U292 (N_292,In_731,In_29);
and U293 (N_293,In_67,In_476);
nor U294 (N_294,In_63,In_590);
nor U295 (N_295,In_643,In_491);
nand U296 (N_296,In_178,In_682);
nand U297 (N_297,In_663,In_626);
or U298 (N_298,In_50,In_145);
xor U299 (N_299,In_19,In_228);
or U300 (N_300,In_509,In_129);
and U301 (N_301,In_306,In_599);
nand U302 (N_302,In_106,In_281);
nand U303 (N_303,In_745,In_608);
nand U304 (N_304,In_182,In_350);
nand U305 (N_305,In_115,In_259);
nand U306 (N_306,In_12,In_549);
nand U307 (N_307,In_251,In_685);
xnor U308 (N_308,In_253,In_388);
or U309 (N_309,In_377,In_492);
nor U310 (N_310,In_551,In_480);
nand U311 (N_311,In_607,In_262);
xnor U312 (N_312,In_654,In_543);
xor U313 (N_313,In_565,In_373);
nor U314 (N_314,In_290,In_561);
xor U315 (N_315,In_44,In_3);
nor U316 (N_316,In_386,In_711);
and U317 (N_317,In_34,In_507);
or U318 (N_318,In_645,In_427);
nor U319 (N_319,In_298,In_150);
or U320 (N_320,In_538,In_487);
nor U321 (N_321,In_554,In_477);
xnor U322 (N_322,In_260,In_219);
nor U323 (N_323,In_722,In_250);
or U324 (N_324,In_612,In_245);
nor U325 (N_325,In_174,In_147);
and U326 (N_326,In_483,In_726);
and U327 (N_327,In_26,In_119);
nand U328 (N_328,In_310,In_90);
xnor U329 (N_329,In_657,In_678);
nand U330 (N_330,In_337,In_447);
xnor U331 (N_331,In_84,In_97);
xnor U332 (N_332,In_563,In_385);
nor U333 (N_333,In_36,In_403);
and U334 (N_334,In_519,In_220);
or U335 (N_335,In_80,In_196);
xnor U336 (N_336,In_116,In_82);
or U337 (N_337,In_243,In_325);
nand U338 (N_338,In_414,In_404);
nand U339 (N_339,In_60,In_101);
xor U340 (N_340,In_381,In_232);
or U341 (N_341,In_525,In_423);
nand U342 (N_342,In_506,In_537);
nor U343 (N_343,In_323,In_273);
nand U344 (N_344,In_99,In_204);
nand U345 (N_345,In_59,In_392);
nor U346 (N_346,In_468,In_313);
or U347 (N_347,In_16,In_420);
xnor U348 (N_348,In_10,In_111);
xnor U349 (N_349,In_652,In_102);
or U350 (N_350,In_721,In_198);
nor U351 (N_351,In_45,In_23);
or U352 (N_352,In_620,In_343);
or U353 (N_353,In_315,In_583);
nor U354 (N_354,In_327,In_121);
and U355 (N_355,In_42,In_170);
or U356 (N_356,In_38,In_673);
xor U357 (N_357,In_378,In_485);
or U358 (N_358,In_149,In_218);
or U359 (N_359,In_295,In_574);
nand U360 (N_360,In_288,In_79);
nor U361 (N_361,In_94,In_389);
and U362 (N_362,In_429,In_686);
nand U363 (N_363,In_72,In_120);
nor U364 (N_364,In_95,In_729);
nand U365 (N_365,In_675,In_168);
xnor U366 (N_366,In_255,In_365);
nor U367 (N_367,In_193,In_296);
or U368 (N_368,In_105,In_448);
nand U369 (N_369,In_653,In_550);
xnor U370 (N_370,In_35,In_189);
xnor U371 (N_371,In_191,In_316);
or U372 (N_372,In_646,In_521);
xnor U373 (N_373,In_680,In_460);
or U374 (N_374,In_252,In_58);
or U375 (N_375,In_378,In_544);
or U376 (N_376,In_561,In_585);
nand U377 (N_377,In_538,In_183);
or U378 (N_378,In_317,In_198);
xnor U379 (N_379,In_593,In_284);
xnor U380 (N_380,In_207,In_518);
or U381 (N_381,In_88,In_541);
and U382 (N_382,In_645,In_98);
and U383 (N_383,In_692,In_127);
and U384 (N_384,In_512,In_473);
xor U385 (N_385,In_662,In_430);
nor U386 (N_386,In_466,In_132);
or U387 (N_387,In_574,In_531);
or U388 (N_388,In_698,In_170);
and U389 (N_389,In_379,In_121);
nor U390 (N_390,In_235,In_284);
or U391 (N_391,In_598,In_247);
nand U392 (N_392,In_492,In_496);
xnor U393 (N_393,In_138,In_266);
xor U394 (N_394,In_350,In_706);
or U395 (N_395,In_662,In_667);
or U396 (N_396,In_694,In_745);
xor U397 (N_397,In_38,In_281);
and U398 (N_398,In_373,In_313);
nand U399 (N_399,In_196,In_386);
nand U400 (N_400,In_214,In_13);
or U401 (N_401,In_334,In_61);
and U402 (N_402,In_578,In_37);
nand U403 (N_403,In_442,In_213);
xnor U404 (N_404,In_398,In_231);
xor U405 (N_405,In_653,In_160);
or U406 (N_406,In_302,In_304);
and U407 (N_407,In_121,In_365);
nor U408 (N_408,In_467,In_183);
and U409 (N_409,In_412,In_150);
nor U410 (N_410,In_661,In_189);
xor U411 (N_411,In_112,In_617);
nor U412 (N_412,In_695,In_573);
xor U413 (N_413,In_225,In_283);
or U414 (N_414,In_582,In_22);
or U415 (N_415,In_554,In_715);
nor U416 (N_416,In_314,In_205);
nand U417 (N_417,In_259,In_385);
nor U418 (N_418,In_72,In_266);
xor U419 (N_419,In_654,In_314);
and U420 (N_420,In_491,In_285);
nand U421 (N_421,In_121,In_295);
and U422 (N_422,In_664,In_514);
nand U423 (N_423,In_6,In_139);
xnor U424 (N_424,In_88,In_537);
or U425 (N_425,In_356,In_343);
and U426 (N_426,In_308,In_508);
and U427 (N_427,In_23,In_30);
and U428 (N_428,In_67,In_136);
or U429 (N_429,In_306,In_635);
or U430 (N_430,In_73,In_573);
or U431 (N_431,In_397,In_235);
xnor U432 (N_432,In_132,In_370);
xor U433 (N_433,In_546,In_520);
or U434 (N_434,In_349,In_544);
or U435 (N_435,In_741,In_283);
nor U436 (N_436,In_34,In_212);
xor U437 (N_437,In_308,In_61);
and U438 (N_438,In_470,In_257);
nand U439 (N_439,In_410,In_261);
xnor U440 (N_440,In_709,In_193);
or U441 (N_441,In_138,In_724);
and U442 (N_442,In_466,In_159);
xor U443 (N_443,In_66,In_363);
and U444 (N_444,In_461,In_528);
nand U445 (N_445,In_439,In_523);
nand U446 (N_446,In_677,In_320);
or U447 (N_447,In_104,In_419);
nand U448 (N_448,In_284,In_392);
nor U449 (N_449,In_581,In_145);
and U450 (N_450,In_166,In_82);
nor U451 (N_451,In_297,In_125);
or U452 (N_452,In_166,In_66);
and U453 (N_453,In_654,In_144);
or U454 (N_454,In_284,In_704);
nor U455 (N_455,In_621,In_565);
nand U456 (N_456,In_260,In_246);
nand U457 (N_457,In_297,In_692);
nor U458 (N_458,In_24,In_29);
and U459 (N_459,In_10,In_663);
and U460 (N_460,In_508,In_53);
nand U461 (N_461,In_580,In_23);
nand U462 (N_462,In_253,In_3);
and U463 (N_463,In_497,In_312);
nand U464 (N_464,In_61,In_523);
nand U465 (N_465,In_713,In_247);
nor U466 (N_466,In_121,In_112);
nand U467 (N_467,In_719,In_125);
nor U468 (N_468,In_63,In_402);
xnor U469 (N_469,In_509,In_738);
xor U470 (N_470,In_157,In_119);
nor U471 (N_471,In_666,In_502);
xor U472 (N_472,In_452,In_276);
xnor U473 (N_473,In_58,In_572);
nand U474 (N_474,In_246,In_692);
xnor U475 (N_475,In_69,In_178);
or U476 (N_476,In_114,In_439);
xnor U477 (N_477,In_621,In_638);
xor U478 (N_478,In_718,In_732);
nor U479 (N_479,In_649,In_5);
or U480 (N_480,In_37,In_342);
nand U481 (N_481,In_215,In_723);
xor U482 (N_482,In_90,In_268);
nand U483 (N_483,In_129,In_65);
nor U484 (N_484,In_76,In_141);
or U485 (N_485,In_142,In_335);
nor U486 (N_486,In_120,In_81);
and U487 (N_487,In_489,In_348);
nor U488 (N_488,In_90,In_710);
and U489 (N_489,In_36,In_601);
and U490 (N_490,In_145,In_667);
xor U491 (N_491,In_670,In_550);
xor U492 (N_492,In_145,In_124);
nor U493 (N_493,In_414,In_317);
nor U494 (N_494,In_134,In_208);
and U495 (N_495,In_411,In_190);
or U496 (N_496,In_544,In_494);
and U497 (N_497,In_374,In_146);
nand U498 (N_498,In_485,In_715);
xnor U499 (N_499,In_312,In_177);
nand U500 (N_500,N_122,N_70);
xnor U501 (N_501,N_236,N_223);
nor U502 (N_502,N_422,N_437);
nor U503 (N_503,N_20,N_23);
nor U504 (N_504,N_435,N_163);
nor U505 (N_505,N_349,N_282);
nand U506 (N_506,N_81,N_446);
or U507 (N_507,N_108,N_451);
nor U508 (N_508,N_232,N_487);
nor U509 (N_509,N_174,N_88);
xor U510 (N_510,N_477,N_116);
or U511 (N_511,N_140,N_271);
nor U512 (N_512,N_469,N_227);
and U513 (N_513,N_332,N_95);
and U514 (N_514,N_14,N_331);
xor U515 (N_515,N_294,N_45);
and U516 (N_516,N_52,N_409);
xor U517 (N_517,N_71,N_53);
xnor U518 (N_518,N_27,N_342);
nor U519 (N_519,N_335,N_36);
nand U520 (N_520,N_492,N_19);
xnor U521 (N_521,N_378,N_136);
nor U522 (N_522,N_22,N_86);
xor U523 (N_523,N_65,N_486);
xnor U524 (N_524,N_191,N_348);
xnor U525 (N_525,N_113,N_44);
xnor U526 (N_526,N_181,N_319);
xnor U527 (N_527,N_382,N_473);
or U528 (N_528,N_215,N_419);
nor U529 (N_529,N_10,N_48);
and U530 (N_530,N_220,N_428);
nor U531 (N_531,N_147,N_260);
or U532 (N_532,N_499,N_31);
xor U533 (N_533,N_457,N_33);
xnor U534 (N_534,N_133,N_393);
nor U535 (N_535,N_103,N_56);
or U536 (N_536,N_196,N_447);
and U537 (N_537,N_148,N_443);
or U538 (N_538,N_173,N_289);
nor U539 (N_539,N_194,N_471);
nand U540 (N_540,N_154,N_302);
nor U541 (N_541,N_412,N_263);
xor U542 (N_542,N_169,N_198);
and U543 (N_543,N_50,N_366);
nor U544 (N_544,N_61,N_89);
nand U545 (N_545,N_273,N_197);
or U546 (N_546,N_75,N_281);
and U547 (N_547,N_436,N_94);
xnor U548 (N_548,N_41,N_221);
xnor U549 (N_549,N_24,N_401);
nor U550 (N_550,N_129,N_93);
and U551 (N_551,N_455,N_30);
nor U552 (N_552,N_286,N_309);
nand U553 (N_553,N_107,N_190);
xnor U554 (N_554,N_311,N_363);
nand U555 (N_555,N_85,N_139);
or U556 (N_556,N_167,N_255);
nor U557 (N_557,N_429,N_79);
nand U558 (N_558,N_327,N_396);
xnor U559 (N_559,N_465,N_365);
nor U560 (N_560,N_249,N_397);
xor U561 (N_561,N_143,N_308);
or U562 (N_562,N_46,N_270);
xnor U563 (N_563,N_150,N_49);
or U564 (N_564,N_151,N_464);
nor U565 (N_565,N_267,N_4);
nor U566 (N_566,N_180,N_411);
or U567 (N_567,N_445,N_418);
or U568 (N_568,N_149,N_239);
or U569 (N_569,N_256,N_385);
nand U570 (N_570,N_185,N_277);
nor U571 (N_571,N_182,N_470);
and U572 (N_572,N_171,N_230);
or U573 (N_573,N_164,N_64);
xor U574 (N_574,N_26,N_117);
or U575 (N_575,N_293,N_497);
and U576 (N_576,N_138,N_121);
nor U577 (N_577,N_152,N_246);
nor U578 (N_578,N_417,N_11);
nor U579 (N_579,N_390,N_224);
xnor U580 (N_580,N_102,N_105);
nor U581 (N_581,N_7,N_355);
and U582 (N_582,N_427,N_214);
nand U583 (N_583,N_141,N_384);
nor U584 (N_584,N_414,N_120);
or U585 (N_585,N_391,N_388);
nor U586 (N_586,N_91,N_405);
or U587 (N_587,N_200,N_254);
and U588 (N_588,N_132,N_114);
and U589 (N_589,N_233,N_336);
xnor U590 (N_590,N_125,N_186);
and U591 (N_591,N_279,N_431);
and U592 (N_592,N_28,N_369);
nor U593 (N_593,N_361,N_63);
nand U594 (N_594,N_290,N_299);
or U595 (N_595,N_127,N_442);
or U596 (N_596,N_12,N_156);
nand U597 (N_597,N_234,N_145);
and U598 (N_598,N_344,N_439);
xnor U599 (N_599,N_195,N_179);
or U600 (N_600,N_280,N_124);
and U601 (N_601,N_206,N_13);
or U602 (N_602,N_134,N_312);
nand U603 (N_603,N_298,N_212);
nand U604 (N_604,N_57,N_72);
nor U605 (N_605,N_493,N_496);
nand U606 (N_606,N_216,N_83);
nand U607 (N_607,N_1,N_479);
nand U608 (N_608,N_137,N_118);
xnor U609 (N_609,N_39,N_187);
and U610 (N_610,N_490,N_373);
nand U611 (N_611,N_482,N_315);
xor U612 (N_612,N_372,N_456);
xnor U613 (N_613,N_370,N_351);
and U614 (N_614,N_303,N_322);
nor U615 (N_615,N_168,N_358);
and U616 (N_616,N_381,N_306);
nor U617 (N_617,N_288,N_326);
or U618 (N_618,N_475,N_37);
or U619 (N_619,N_172,N_183);
nand U620 (N_620,N_426,N_489);
nor U621 (N_621,N_440,N_450);
nand U622 (N_622,N_38,N_146);
xor U623 (N_623,N_467,N_448);
and U624 (N_624,N_98,N_217);
nor U625 (N_625,N_374,N_462);
xnor U626 (N_626,N_258,N_15);
nand U627 (N_627,N_420,N_276);
nor U628 (N_628,N_259,N_421);
xnor U629 (N_629,N_380,N_35);
and U630 (N_630,N_398,N_416);
nor U631 (N_631,N_43,N_399);
xor U632 (N_632,N_444,N_481);
xnor U633 (N_633,N_55,N_343);
and U634 (N_634,N_205,N_74);
nand U635 (N_635,N_438,N_250);
and U636 (N_636,N_352,N_34);
nand U637 (N_637,N_203,N_245);
and U638 (N_638,N_345,N_0);
and U639 (N_639,N_192,N_222);
nor U640 (N_640,N_51,N_123);
or U641 (N_641,N_243,N_131);
nor U642 (N_642,N_459,N_310);
or U643 (N_643,N_175,N_92);
or U644 (N_644,N_235,N_58);
nand U645 (N_645,N_106,N_339);
or U646 (N_646,N_283,N_297);
nand U647 (N_647,N_211,N_408);
nand U648 (N_648,N_84,N_265);
nor U649 (N_649,N_354,N_313);
nand U650 (N_650,N_119,N_248);
or U651 (N_651,N_295,N_47);
xnor U652 (N_652,N_60,N_458);
xor U653 (N_653,N_353,N_157);
and U654 (N_654,N_62,N_321);
nand U655 (N_655,N_434,N_40);
or U656 (N_656,N_219,N_252);
and U657 (N_657,N_153,N_472);
nand U658 (N_658,N_87,N_485);
nand U659 (N_659,N_32,N_350);
and U660 (N_660,N_320,N_231);
and U661 (N_661,N_269,N_424);
or U662 (N_662,N_314,N_257);
nand U663 (N_663,N_17,N_226);
nand U664 (N_664,N_386,N_359);
nand U665 (N_665,N_76,N_430);
xor U666 (N_666,N_453,N_142);
nand U667 (N_667,N_253,N_425);
or U668 (N_668,N_213,N_18);
nor U669 (N_669,N_460,N_347);
xor U670 (N_670,N_160,N_155);
nand U671 (N_671,N_466,N_251);
nand U672 (N_672,N_484,N_42);
or U673 (N_673,N_376,N_6);
nor U674 (N_674,N_68,N_199);
xnor U675 (N_675,N_407,N_104);
nand U676 (N_676,N_452,N_90);
or U677 (N_677,N_158,N_228);
nand U678 (N_678,N_135,N_97);
nor U679 (N_679,N_225,N_483);
nor U680 (N_680,N_375,N_238);
and U681 (N_681,N_274,N_406);
nand U682 (N_682,N_126,N_480);
nand U683 (N_683,N_304,N_337);
nor U684 (N_684,N_284,N_449);
nor U685 (N_685,N_291,N_461);
and U686 (N_686,N_413,N_77);
nand U687 (N_687,N_262,N_368);
nor U688 (N_688,N_59,N_491);
nand U689 (N_689,N_66,N_82);
and U690 (N_690,N_423,N_162);
and U691 (N_691,N_275,N_329);
and U692 (N_692,N_29,N_202);
xnor U693 (N_693,N_189,N_325);
nand U694 (N_694,N_242,N_341);
or U695 (N_695,N_360,N_296);
nand U696 (N_696,N_111,N_159);
xor U697 (N_697,N_69,N_395);
and U698 (N_698,N_316,N_161);
or U699 (N_699,N_96,N_218);
nand U700 (N_700,N_237,N_264);
or U701 (N_701,N_184,N_498);
nand U702 (N_702,N_99,N_494);
or U703 (N_703,N_287,N_402);
and U704 (N_704,N_371,N_305);
xnor U705 (N_705,N_3,N_144);
xnor U706 (N_706,N_244,N_101);
xor U707 (N_707,N_410,N_338);
xor U708 (N_708,N_403,N_478);
nand U709 (N_709,N_387,N_463);
nand U710 (N_710,N_474,N_404);
or U711 (N_711,N_323,N_112);
nand U712 (N_712,N_165,N_333);
nor U713 (N_713,N_109,N_324);
nor U714 (N_714,N_300,N_488);
and U715 (N_715,N_170,N_301);
and U716 (N_716,N_364,N_229);
nor U717 (N_717,N_383,N_130);
nor U718 (N_718,N_110,N_272);
and U719 (N_719,N_8,N_177);
and U720 (N_720,N_5,N_261);
nor U721 (N_721,N_356,N_379);
xor U722 (N_722,N_468,N_2);
nor U723 (N_723,N_415,N_318);
and U724 (N_724,N_377,N_115);
and U725 (N_725,N_16,N_292);
and U726 (N_726,N_178,N_241);
nand U727 (N_727,N_73,N_166);
and U728 (N_728,N_476,N_208);
or U729 (N_729,N_67,N_400);
or U730 (N_730,N_176,N_100);
xnor U731 (N_731,N_334,N_9);
or U732 (N_732,N_193,N_340);
nor U733 (N_733,N_330,N_346);
or U734 (N_734,N_394,N_392);
nand U735 (N_735,N_204,N_268);
xnor U736 (N_736,N_247,N_495);
nor U737 (N_737,N_201,N_357);
nand U738 (N_738,N_389,N_278);
and U739 (N_739,N_128,N_454);
or U740 (N_740,N_188,N_25);
nor U741 (N_741,N_307,N_285);
nand U742 (N_742,N_266,N_328);
and U743 (N_743,N_240,N_441);
nand U744 (N_744,N_367,N_362);
and U745 (N_745,N_78,N_433);
xnor U746 (N_746,N_432,N_21);
or U747 (N_747,N_207,N_210);
nor U748 (N_748,N_80,N_317);
nand U749 (N_749,N_54,N_209);
nor U750 (N_750,N_342,N_433);
nand U751 (N_751,N_355,N_487);
nand U752 (N_752,N_331,N_111);
nor U753 (N_753,N_373,N_128);
nand U754 (N_754,N_318,N_386);
and U755 (N_755,N_334,N_255);
or U756 (N_756,N_237,N_57);
and U757 (N_757,N_436,N_430);
or U758 (N_758,N_18,N_228);
nor U759 (N_759,N_105,N_81);
or U760 (N_760,N_402,N_227);
or U761 (N_761,N_249,N_193);
or U762 (N_762,N_198,N_486);
xnor U763 (N_763,N_316,N_232);
xor U764 (N_764,N_295,N_160);
or U765 (N_765,N_247,N_380);
xor U766 (N_766,N_172,N_373);
nor U767 (N_767,N_244,N_324);
nor U768 (N_768,N_166,N_332);
or U769 (N_769,N_351,N_393);
nand U770 (N_770,N_82,N_61);
and U771 (N_771,N_496,N_246);
xnor U772 (N_772,N_290,N_498);
and U773 (N_773,N_380,N_412);
or U774 (N_774,N_275,N_313);
xor U775 (N_775,N_467,N_483);
xnor U776 (N_776,N_184,N_215);
nor U777 (N_777,N_254,N_143);
and U778 (N_778,N_119,N_101);
nor U779 (N_779,N_310,N_440);
and U780 (N_780,N_5,N_362);
xor U781 (N_781,N_169,N_185);
nand U782 (N_782,N_102,N_49);
and U783 (N_783,N_48,N_207);
nand U784 (N_784,N_315,N_486);
nor U785 (N_785,N_121,N_169);
nand U786 (N_786,N_298,N_445);
xnor U787 (N_787,N_305,N_470);
nor U788 (N_788,N_91,N_363);
and U789 (N_789,N_177,N_486);
nor U790 (N_790,N_495,N_226);
nand U791 (N_791,N_67,N_94);
or U792 (N_792,N_30,N_11);
or U793 (N_793,N_345,N_166);
nor U794 (N_794,N_100,N_71);
xnor U795 (N_795,N_150,N_187);
xor U796 (N_796,N_416,N_265);
nand U797 (N_797,N_148,N_120);
xor U798 (N_798,N_227,N_421);
and U799 (N_799,N_67,N_54);
or U800 (N_800,N_440,N_146);
nand U801 (N_801,N_265,N_333);
nand U802 (N_802,N_475,N_187);
and U803 (N_803,N_114,N_483);
xnor U804 (N_804,N_321,N_286);
nand U805 (N_805,N_103,N_499);
xnor U806 (N_806,N_54,N_256);
xor U807 (N_807,N_241,N_286);
xnor U808 (N_808,N_450,N_388);
xor U809 (N_809,N_148,N_386);
or U810 (N_810,N_155,N_346);
and U811 (N_811,N_140,N_204);
nor U812 (N_812,N_110,N_131);
nand U813 (N_813,N_293,N_96);
nor U814 (N_814,N_100,N_167);
and U815 (N_815,N_155,N_436);
nand U816 (N_816,N_153,N_84);
nor U817 (N_817,N_99,N_339);
or U818 (N_818,N_330,N_119);
or U819 (N_819,N_337,N_178);
nor U820 (N_820,N_324,N_330);
nand U821 (N_821,N_258,N_247);
or U822 (N_822,N_183,N_112);
and U823 (N_823,N_415,N_181);
nor U824 (N_824,N_38,N_71);
nand U825 (N_825,N_345,N_255);
or U826 (N_826,N_59,N_485);
xnor U827 (N_827,N_27,N_496);
xor U828 (N_828,N_219,N_274);
xor U829 (N_829,N_95,N_116);
or U830 (N_830,N_375,N_478);
nand U831 (N_831,N_18,N_280);
or U832 (N_832,N_179,N_380);
nor U833 (N_833,N_124,N_470);
and U834 (N_834,N_27,N_488);
xnor U835 (N_835,N_132,N_285);
and U836 (N_836,N_441,N_90);
nor U837 (N_837,N_169,N_8);
nor U838 (N_838,N_31,N_70);
or U839 (N_839,N_249,N_175);
xor U840 (N_840,N_442,N_346);
xor U841 (N_841,N_399,N_240);
and U842 (N_842,N_292,N_406);
nand U843 (N_843,N_118,N_272);
and U844 (N_844,N_412,N_206);
or U845 (N_845,N_263,N_23);
xnor U846 (N_846,N_380,N_469);
or U847 (N_847,N_231,N_101);
or U848 (N_848,N_474,N_305);
nand U849 (N_849,N_232,N_418);
or U850 (N_850,N_419,N_360);
nor U851 (N_851,N_358,N_131);
xor U852 (N_852,N_22,N_77);
xnor U853 (N_853,N_92,N_224);
xnor U854 (N_854,N_20,N_410);
xor U855 (N_855,N_66,N_154);
xnor U856 (N_856,N_491,N_147);
and U857 (N_857,N_472,N_110);
xor U858 (N_858,N_0,N_290);
xor U859 (N_859,N_490,N_287);
or U860 (N_860,N_125,N_216);
nor U861 (N_861,N_199,N_189);
xor U862 (N_862,N_352,N_50);
nand U863 (N_863,N_415,N_440);
and U864 (N_864,N_5,N_386);
or U865 (N_865,N_145,N_275);
nor U866 (N_866,N_161,N_212);
nand U867 (N_867,N_189,N_235);
and U868 (N_868,N_292,N_83);
or U869 (N_869,N_386,N_486);
nand U870 (N_870,N_411,N_284);
and U871 (N_871,N_147,N_127);
and U872 (N_872,N_275,N_240);
or U873 (N_873,N_133,N_67);
nand U874 (N_874,N_123,N_414);
or U875 (N_875,N_263,N_196);
or U876 (N_876,N_307,N_372);
and U877 (N_877,N_112,N_304);
xor U878 (N_878,N_308,N_31);
nor U879 (N_879,N_42,N_304);
xor U880 (N_880,N_176,N_477);
and U881 (N_881,N_199,N_334);
nand U882 (N_882,N_392,N_123);
xor U883 (N_883,N_190,N_91);
or U884 (N_884,N_402,N_278);
or U885 (N_885,N_103,N_473);
xor U886 (N_886,N_466,N_397);
nor U887 (N_887,N_496,N_456);
and U888 (N_888,N_156,N_135);
xor U889 (N_889,N_336,N_323);
xnor U890 (N_890,N_257,N_477);
xnor U891 (N_891,N_51,N_194);
nand U892 (N_892,N_269,N_432);
nand U893 (N_893,N_82,N_381);
nor U894 (N_894,N_313,N_394);
nor U895 (N_895,N_215,N_395);
nand U896 (N_896,N_417,N_475);
nor U897 (N_897,N_362,N_251);
and U898 (N_898,N_215,N_368);
and U899 (N_899,N_362,N_204);
and U900 (N_900,N_19,N_355);
xor U901 (N_901,N_220,N_336);
nor U902 (N_902,N_77,N_283);
and U903 (N_903,N_124,N_18);
and U904 (N_904,N_114,N_156);
or U905 (N_905,N_360,N_195);
nand U906 (N_906,N_212,N_451);
nor U907 (N_907,N_157,N_346);
nor U908 (N_908,N_477,N_155);
or U909 (N_909,N_323,N_107);
and U910 (N_910,N_337,N_447);
nor U911 (N_911,N_286,N_24);
nor U912 (N_912,N_141,N_428);
and U913 (N_913,N_387,N_296);
xor U914 (N_914,N_216,N_10);
xnor U915 (N_915,N_450,N_102);
nor U916 (N_916,N_477,N_48);
and U917 (N_917,N_394,N_39);
and U918 (N_918,N_319,N_453);
and U919 (N_919,N_217,N_115);
or U920 (N_920,N_142,N_151);
nor U921 (N_921,N_40,N_386);
or U922 (N_922,N_90,N_499);
nor U923 (N_923,N_233,N_469);
and U924 (N_924,N_353,N_115);
nor U925 (N_925,N_308,N_283);
or U926 (N_926,N_331,N_124);
xnor U927 (N_927,N_130,N_390);
xor U928 (N_928,N_392,N_151);
xor U929 (N_929,N_484,N_391);
nand U930 (N_930,N_390,N_258);
or U931 (N_931,N_179,N_264);
and U932 (N_932,N_486,N_156);
nor U933 (N_933,N_130,N_264);
or U934 (N_934,N_293,N_215);
nand U935 (N_935,N_96,N_130);
nand U936 (N_936,N_289,N_322);
or U937 (N_937,N_142,N_444);
and U938 (N_938,N_143,N_369);
nand U939 (N_939,N_329,N_32);
nor U940 (N_940,N_12,N_315);
nand U941 (N_941,N_98,N_51);
or U942 (N_942,N_485,N_172);
nor U943 (N_943,N_242,N_312);
nor U944 (N_944,N_224,N_37);
nand U945 (N_945,N_376,N_64);
and U946 (N_946,N_326,N_248);
xor U947 (N_947,N_91,N_192);
nand U948 (N_948,N_362,N_135);
xor U949 (N_949,N_222,N_364);
xnor U950 (N_950,N_385,N_5);
xnor U951 (N_951,N_456,N_264);
and U952 (N_952,N_302,N_27);
nor U953 (N_953,N_148,N_176);
nor U954 (N_954,N_49,N_489);
nand U955 (N_955,N_205,N_222);
nor U956 (N_956,N_243,N_454);
nand U957 (N_957,N_277,N_485);
nor U958 (N_958,N_433,N_356);
and U959 (N_959,N_143,N_348);
xor U960 (N_960,N_276,N_343);
nand U961 (N_961,N_445,N_419);
xor U962 (N_962,N_226,N_267);
or U963 (N_963,N_198,N_222);
nor U964 (N_964,N_180,N_56);
or U965 (N_965,N_216,N_20);
and U966 (N_966,N_144,N_281);
nor U967 (N_967,N_399,N_291);
and U968 (N_968,N_317,N_230);
and U969 (N_969,N_289,N_151);
or U970 (N_970,N_184,N_440);
and U971 (N_971,N_393,N_245);
and U972 (N_972,N_210,N_206);
nor U973 (N_973,N_427,N_101);
and U974 (N_974,N_194,N_282);
and U975 (N_975,N_225,N_457);
nor U976 (N_976,N_10,N_146);
xnor U977 (N_977,N_134,N_283);
and U978 (N_978,N_426,N_263);
and U979 (N_979,N_31,N_256);
and U980 (N_980,N_420,N_157);
nor U981 (N_981,N_384,N_160);
or U982 (N_982,N_289,N_443);
and U983 (N_983,N_279,N_159);
or U984 (N_984,N_224,N_165);
xnor U985 (N_985,N_165,N_299);
or U986 (N_986,N_462,N_97);
xnor U987 (N_987,N_29,N_343);
nor U988 (N_988,N_322,N_151);
and U989 (N_989,N_153,N_461);
nand U990 (N_990,N_436,N_183);
xor U991 (N_991,N_236,N_74);
and U992 (N_992,N_173,N_409);
xor U993 (N_993,N_74,N_298);
or U994 (N_994,N_218,N_248);
and U995 (N_995,N_185,N_68);
nor U996 (N_996,N_17,N_108);
or U997 (N_997,N_309,N_68);
and U998 (N_998,N_324,N_426);
xor U999 (N_999,N_290,N_382);
nor U1000 (N_1000,N_819,N_759);
nor U1001 (N_1001,N_864,N_991);
nor U1002 (N_1002,N_731,N_815);
nor U1003 (N_1003,N_609,N_556);
xnor U1004 (N_1004,N_530,N_717);
nand U1005 (N_1005,N_937,N_936);
nor U1006 (N_1006,N_694,N_649);
nand U1007 (N_1007,N_776,N_661);
or U1008 (N_1008,N_598,N_899);
or U1009 (N_1009,N_977,N_749);
nor U1010 (N_1010,N_935,N_519);
nand U1011 (N_1011,N_761,N_600);
xnor U1012 (N_1012,N_954,N_697);
or U1013 (N_1013,N_788,N_763);
nor U1014 (N_1014,N_770,N_754);
nand U1015 (N_1015,N_608,N_507);
nand U1016 (N_1016,N_943,N_523);
nand U1017 (N_1017,N_982,N_769);
nor U1018 (N_1018,N_590,N_660);
and U1019 (N_1019,N_879,N_520);
xor U1020 (N_1020,N_980,N_675);
xnor U1021 (N_1021,N_545,N_571);
xnor U1022 (N_1022,N_536,N_566);
nand U1023 (N_1023,N_895,N_939);
xnor U1024 (N_1024,N_730,N_510);
or U1025 (N_1025,N_656,N_782);
nor U1026 (N_1026,N_626,N_881);
xor U1027 (N_1027,N_984,N_762);
xor U1028 (N_1028,N_647,N_906);
nor U1029 (N_1029,N_527,N_544);
nor U1030 (N_1030,N_687,N_959);
nor U1031 (N_1031,N_996,N_718);
or U1032 (N_1032,N_871,N_514);
xor U1033 (N_1033,N_888,N_669);
and U1034 (N_1034,N_909,N_990);
and U1035 (N_1035,N_757,N_809);
nor U1036 (N_1036,N_646,N_911);
nor U1037 (N_1037,N_618,N_604);
xor U1038 (N_1038,N_720,N_534);
xor U1039 (N_1039,N_812,N_563);
nor U1040 (N_1040,N_639,N_829);
nand U1041 (N_1041,N_612,N_630);
nand U1042 (N_1042,N_771,N_575);
or U1043 (N_1043,N_845,N_508);
xor U1044 (N_1044,N_746,N_512);
xnor U1045 (N_1045,N_709,N_693);
and U1046 (N_1046,N_617,N_968);
nor U1047 (N_1047,N_650,N_930);
and U1048 (N_1048,N_925,N_821);
and U1049 (N_1049,N_831,N_651);
nand U1050 (N_1050,N_503,N_594);
nand U1051 (N_1051,N_840,N_802);
nor U1052 (N_1052,N_572,N_973);
nor U1053 (N_1053,N_706,N_509);
or U1054 (N_1054,N_934,N_768);
and U1055 (N_1055,N_637,N_532);
nor U1056 (N_1056,N_521,N_997);
or U1057 (N_1057,N_711,N_978);
or U1058 (N_1058,N_903,N_995);
nor U1059 (N_1059,N_565,N_953);
xor U1060 (N_1060,N_505,N_947);
and U1061 (N_1061,N_601,N_862);
or U1062 (N_1062,N_538,N_867);
nor U1063 (N_1063,N_698,N_874);
nand U1064 (N_1064,N_950,N_500);
xor U1065 (N_1065,N_961,N_781);
xnor U1066 (N_1066,N_549,N_832);
nand U1067 (N_1067,N_570,N_584);
or U1068 (N_1068,N_680,N_872);
and U1069 (N_1069,N_506,N_644);
and U1070 (N_1070,N_585,N_922);
or U1071 (N_1071,N_932,N_504);
nand U1072 (N_1072,N_736,N_791);
nor U1073 (N_1073,N_855,N_919);
xor U1074 (N_1074,N_869,N_582);
nand U1075 (N_1075,N_779,N_786);
xnor U1076 (N_1076,N_688,N_743);
nor U1077 (N_1077,N_798,N_852);
and U1078 (N_1078,N_865,N_866);
nor U1079 (N_1079,N_785,N_702);
xor U1080 (N_1080,N_800,N_628);
nor U1081 (N_1081,N_884,N_989);
nor U1082 (N_1082,N_857,N_648);
or U1083 (N_1083,N_684,N_654);
or U1084 (N_1084,N_524,N_823);
or U1085 (N_1085,N_926,N_976);
nor U1086 (N_1086,N_540,N_963);
nor U1087 (N_1087,N_933,N_913);
and U1088 (N_1088,N_817,N_778);
and U1089 (N_1089,N_877,N_971);
or U1090 (N_1090,N_795,N_547);
and U1091 (N_1091,N_655,N_940);
and U1092 (N_1092,N_671,N_880);
and U1093 (N_1093,N_994,N_610);
nand U1094 (N_1094,N_576,N_780);
and U1095 (N_1095,N_797,N_905);
nor U1096 (N_1096,N_573,N_870);
nor U1097 (N_1097,N_517,N_772);
nand U1098 (N_1098,N_587,N_535);
xor U1099 (N_1099,N_957,N_787);
xor U1100 (N_1100,N_712,N_674);
nand U1101 (N_1101,N_657,N_659);
nor U1102 (N_1102,N_635,N_955);
nor U1103 (N_1103,N_685,N_902);
nor U1104 (N_1104,N_607,N_901);
or U1105 (N_1105,N_511,N_945);
nand U1106 (N_1106,N_613,N_828);
and U1107 (N_1107,N_890,N_752);
nor U1108 (N_1108,N_733,N_526);
and U1109 (N_1109,N_992,N_773);
xor U1110 (N_1110,N_673,N_859);
or U1111 (N_1111,N_632,N_960);
xnor U1112 (N_1112,N_695,N_689);
nand U1113 (N_1113,N_701,N_597);
nor U1114 (N_1114,N_836,N_846);
or U1115 (N_1115,N_723,N_696);
xnor U1116 (N_1116,N_889,N_665);
and U1117 (N_1117,N_741,N_917);
nand U1118 (N_1118,N_558,N_924);
xor U1119 (N_1119,N_588,N_814);
or U1120 (N_1120,N_948,N_686);
nor U1121 (N_1121,N_619,N_750);
nor U1122 (N_1122,N_586,N_589);
and U1123 (N_1123,N_988,N_850);
xnor U1124 (N_1124,N_887,N_860);
xor U1125 (N_1125,N_810,N_580);
nor U1126 (N_1126,N_708,N_550);
nand U1127 (N_1127,N_897,N_986);
nand U1128 (N_1128,N_966,N_638);
nand U1129 (N_1129,N_987,N_641);
nor U1130 (N_1130,N_863,N_942);
or U1131 (N_1131,N_502,N_921);
and U1132 (N_1132,N_541,N_513);
nor U1133 (N_1133,N_844,N_858);
nand U1134 (N_1134,N_783,N_679);
and U1135 (N_1135,N_652,N_908);
and U1136 (N_1136,N_719,N_611);
nand U1137 (N_1137,N_807,N_923);
nor U1138 (N_1138,N_816,N_559);
xor U1139 (N_1139,N_525,N_591);
nor U1140 (N_1140,N_876,N_891);
nor U1141 (N_1141,N_985,N_835);
xnor U1142 (N_1142,N_636,N_803);
xor U1143 (N_1143,N_843,N_699);
xnor U1144 (N_1144,N_837,N_965);
and U1145 (N_1145,N_554,N_929);
nand U1146 (N_1146,N_537,N_581);
or U1147 (N_1147,N_893,N_668);
nand U1148 (N_1148,N_931,N_678);
or U1149 (N_1149,N_725,N_755);
nand U1150 (N_1150,N_993,N_561);
and U1151 (N_1151,N_777,N_842);
xor U1152 (N_1152,N_516,N_818);
xor U1153 (N_1153,N_753,N_599);
or U1154 (N_1154,N_744,N_577);
xor U1155 (N_1155,N_643,N_910);
nand U1156 (N_1156,N_907,N_670);
xnor U1157 (N_1157,N_622,N_546);
and U1158 (N_1158,N_751,N_894);
xnor U1159 (N_1159,N_825,N_605);
or U1160 (N_1160,N_642,N_898);
and U1161 (N_1161,N_841,N_557);
nand U1162 (N_1162,N_713,N_806);
nor U1163 (N_1163,N_794,N_826);
and U1164 (N_1164,N_515,N_710);
nor U1165 (N_1165,N_574,N_562);
nor U1166 (N_1166,N_813,N_774);
nor U1167 (N_1167,N_822,N_539);
nor U1168 (N_1168,N_981,N_830);
nor U1169 (N_1169,N_951,N_533);
xnor U1170 (N_1170,N_677,N_956);
and U1171 (N_1171,N_676,N_827);
nand U1172 (N_1172,N_705,N_716);
or U1173 (N_1173,N_734,N_567);
nand U1174 (N_1174,N_735,N_592);
and U1175 (N_1175,N_969,N_804);
and U1176 (N_1176,N_707,N_760);
xor U1177 (N_1177,N_729,N_764);
nand U1178 (N_1178,N_972,N_928);
or U1179 (N_1179,N_914,N_727);
nand U1180 (N_1180,N_501,N_805);
xnor U1181 (N_1181,N_682,N_738);
and U1182 (N_1182,N_737,N_811);
xor U1183 (N_1183,N_531,N_944);
nand U1184 (N_1184,N_834,N_756);
and U1185 (N_1185,N_662,N_854);
and U1186 (N_1186,N_724,N_873);
and U1187 (N_1187,N_593,N_904);
xor U1188 (N_1188,N_569,N_915);
or U1189 (N_1189,N_624,N_740);
and U1190 (N_1190,N_667,N_529);
xnor U1191 (N_1191,N_579,N_595);
xor U1192 (N_1192,N_542,N_900);
xor U1193 (N_1193,N_664,N_853);
and U1194 (N_1194,N_583,N_745);
nand U1195 (N_1195,N_875,N_918);
or U1196 (N_1196,N_998,N_789);
nor U1197 (N_1197,N_967,N_615);
and U1198 (N_1198,N_621,N_596);
or U1199 (N_1199,N_927,N_518);
and U1200 (N_1200,N_847,N_726);
xnor U1201 (N_1201,N_946,N_748);
or U1202 (N_1202,N_747,N_883);
nor U1203 (N_1203,N_616,N_640);
nor U1204 (N_1204,N_801,N_672);
or U1205 (N_1205,N_742,N_790);
or U1206 (N_1206,N_663,N_775);
nand U1207 (N_1207,N_633,N_896);
nor U1208 (N_1208,N_808,N_970);
or U1209 (N_1209,N_999,N_949);
xor U1210 (N_1210,N_551,N_728);
and U1211 (N_1211,N_848,N_849);
xnor U1212 (N_1212,N_784,N_938);
nor U1213 (N_1213,N_560,N_627);
xor U1214 (N_1214,N_912,N_962);
nor U1215 (N_1215,N_690,N_552);
and U1216 (N_1216,N_974,N_824);
or U1217 (N_1217,N_623,N_920);
or U1218 (N_1218,N_722,N_653);
nor U1219 (N_1219,N_839,N_838);
xor U1220 (N_1220,N_658,N_861);
xor U1221 (N_1221,N_941,N_692);
nand U1222 (N_1222,N_564,N_631);
nand U1223 (N_1223,N_952,N_614);
and U1224 (N_1224,N_765,N_634);
and U1225 (N_1225,N_758,N_700);
nand U1226 (N_1226,N_666,N_796);
and U1227 (N_1227,N_704,N_766);
xor U1228 (N_1228,N_739,N_792);
xor U1229 (N_1229,N_555,N_645);
xor U1230 (N_1230,N_975,N_721);
xor U1231 (N_1231,N_958,N_820);
xor U1232 (N_1232,N_856,N_578);
xnor U1233 (N_1233,N_767,N_983);
xnor U1234 (N_1234,N_886,N_715);
nor U1235 (N_1235,N_606,N_553);
or U1236 (N_1236,N_892,N_851);
or U1237 (N_1237,N_714,N_979);
or U1238 (N_1238,N_916,N_522);
and U1239 (N_1239,N_603,N_793);
xnor U1240 (N_1240,N_625,N_799);
xor U1241 (N_1241,N_868,N_568);
xnor U1242 (N_1242,N_681,N_548);
nand U1243 (N_1243,N_964,N_833);
or U1244 (N_1244,N_602,N_732);
or U1245 (N_1245,N_885,N_878);
and U1246 (N_1246,N_683,N_543);
or U1247 (N_1247,N_528,N_691);
xnor U1248 (N_1248,N_703,N_629);
nand U1249 (N_1249,N_882,N_620);
nand U1250 (N_1250,N_877,N_920);
xor U1251 (N_1251,N_740,N_718);
or U1252 (N_1252,N_936,N_611);
nand U1253 (N_1253,N_895,N_800);
nand U1254 (N_1254,N_897,N_575);
xnor U1255 (N_1255,N_586,N_554);
or U1256 (N_1256,N_594,N_891);
nor U1257 (N_1257,N_732,N_870);
and U1258 (N_1258,N_984,N_731);
nor U1259 (N_1259,N_889,N_945);
nand U1260 (N_1260,N_777,N_718);
xor U1261 (N_1261,N_543,N_958);
xor U1262 (N_1262,N_627,N_715);
xnor U1263 (N_1263,N_515,N_890);
or U1264 (N_1264,N_891,N_962);
nand U1265 (N_1265,N_840,N_757);
nand U1266 (N_1266,N_556,N_841);
nand U1267 (N_1267,N_916,N_692);
or U1268 (N_1268,N_729,N_507);
nor U1269 (N_1269,N_548,N_600);
or U1270 (N_1270,N_637,N_522);
or U1271 (N_1271,N_551,N_797);
nor U1272 (N_1272,N_574,N_563);
and U1273 (N_1273,N_557,N_894);
nor U1274 (N_1274,N_642,N_730);
nand U1275 (N_1275,N_696,N_633);
nor U1276 (N_1276,N_798,N_853);
nor U1277 (N_1277,N_970,N_916);
nand U1278 (N_1278,N_987,N_549);
and U1279 (N_1279,N_872,N_544);
nand U1280 (N_1280,N_852,N_524);
nand U1281 (N_1281,N_547,N_913);
nor U1282 (N_1282,N_668,N_820);
xnor U1283 (N_1283,N_516,N_609);
nand U1284 (N_1284,N_749,N_912);
nor U1285 (N_1285,N_865,N_851);
xor U1286 (N_1286,N_573,N_864);
nor U1287 (N_1287,N_814,N_895);
nand U1288 (N_1288,N_590,N_702);
xor U1289 (N_1289,N_506,N_795);
nor U1290 (N_1290,N_570,N_563);
nand U1291 (N_1291,N_797,N_866);
nor U1292 (N_1292,N_791,N_896);
or U1293 (N_1293,N_694,N_841);
nand U1294 (N_1294,N_754,N_790);
xor U1295 (N_1295,N_900,N_841);
and U1296 (N_1296,N_523,N_772);
nor U1297 (N_1297,N_660,N_906);
or U1298 (N_1298,N_578,N_912);
nor U1299 (N_1299,N_591,N_665);
nor U1300 (N_1300,N_843,N_630);
nand U1301 (N_1301,N_524,N_982);
or U1302 (N_1302,N_880,N_557);
xor U1303 (N_1303,N_873,N_648);
and U1304 (N_1304,N_625,N_723);
or U1305 (N_1305,N_702,N_818);
nand U1306 (N_1306,N_512,N_714);
nor U1307 (N_1307,N_752,N_760);
nand U1308 (N_1308,N_957,N_921);
nor U1309 (N_1309,N_649,N_596);
or U1310 (N_1310,N_504,N_630);
and U1311 (N_1311,N_783,N_844);
xor U1312 (N_1312,N_932,N_611);
xor U1313 (N_1313,N_874,N_527);
or U1314 (N_1314,N_669,N_816);
nand U1315 (N_1315,N_952,N_759);
or U1316 (N_1316,N_974,N_644);
xnor U1317 (N_1317,N_731,N_834);
xnor U1318 (N_1318,N_929,N_712);
and U1319 (N_1319,N_995,N_715);
or U1320 (N_1320,N_618,N_959);
xor U1321 (N_1321,N_596,N_559);
nor U1322 (N_1322,N_905,N_504);
xor U1323 (N_1323,N_978,N_702);
xor U1324 (N_1324,N_724,N_935);
nand U1325 (N_1325,N_721,N_863);
or U1326 (N_1326,N_968,N_944);
and U1327 (N_1327,N_596,N_537);
nand U1328 (N_1328,N_795,N_504);
nor U1329 (N_1329,N_668,N_523);
and U1330 (N_1330,N_705,N_900);
or U1331 (N_1331,N_516,N_664);
and U1332 (N_1332,N_861,N_715);
nand U1333 (N_1333,N_960,N_900);
or U1334 (N_1334,N_588,N_878);
or U1335 (N_1335,N_586,N_598);
or U1336 (N_1336,N_526,N_667);
nor U1337 (N_1337,N_760,N_932);
nand U1338 (N_1338,N_880,N_938);
and U1339 (N_1339,N_782,N_860);
and U1340 (N_1340,N_766,N_620);
and U1341 (N_1341,N_607,N_889);
xor U1342 (N_1342,N_611,N_749);
and U1343 (N_1343,N_852,N_859);
or U1344 (N_1344,N_993,N_601);
xor U1345 (N_1345,N_569,N_840);
xor U1346 (N_1346,N_668,N_838);
nand U1347 (N_1347,N_764,N_785);
or U1348 (N_1348,N_987,N_893);
xor U1349 (N_1349,N_938,N_995);
xnor U1350 (N_1350,N_785,N_810);
xnor U1351 (N_1351,N_881,N_733);
nor U1352 (N_1352,N_811,N_796);
nor U1353 (N_1353,N_523,N_813);
xnor U1354 (N_1354,N_798,N_731);
xnor U1355 (N_1355,N_784,N_935);
or U1356 (N_1356,N_793,N_789);
or U1357 (N_1357,N_731,N_523);
nor U1358 (N_1358,N_892,N_627);
and U1359 (N_1359,N_791,N_980);
nor U1360 (N_1360,N_910,N_771);
or U1361 (N_1361,N_969,N_814);
xor U1362 (N_1362,N_944,N_511);
or U1363 (N_1363,N_621,N_810);
and U1364 (N_1364,N_823,N_571);
and U1365 (N_1365,N_782,N_924);
xor U1366 (N_1366,N_643,N_973);
and U1367 (N_1367,N_587,N_811);
and U1368 (N_1368,N_620,N_614);
nor U1369 (N_1369,N_924,N_891);
nand U1370 (N_1370,N_953,N_692);
nand U1371 (N_1371,N_993,N_833);
xor U1372 (N_1372,N_502,N_850);
nand U1373 (N_1373,N_596,N_910);
and U1374 (N_1374,N_660,N_523);
nor U1375 (N_1375,N_616,N_685);
nor U1376 (N_1376,N_677,N_870);
or U1377 (N_1377,N_868,N_806);
nand U1378 (N_1378,N_958,N_700);
xnor U1379 (N_1379,N_777,N_983);
nand U1380 (N_1380,N_668,N_975);
nand U1381 (N_1381,N_587,N_863);
and U1382 (N_1382,N_830,N_837);
nor U1383 (N_1383,N_563,N_627);
or U1384 (N_1384,N_957,N_580);
or U1385 (N_1385,N_950,N_649);
nand U1386 (N_1386,N_936,N_546);
or U1387 (N_1387,N_845,N_503);
nor U1388 (N_1388,N_837,N_901);
xnor U1389 (N_1389,N_909,N_628);
nor U1390 (N_1390,N_934,N_523);
and U1391 (N_1391,N_592,N_657);
nor U1392 (N_1392,N_714,N_758);
nand U1393 (N_1393,N_635,N_732);
xnor U1394 (N_1394,N_712,N_989);
or U1395 (N_1395,N_656,N_624);
or U1396 (N_1396,N_972,N_891);
nand U1397 (N_1397,N_929,N_642);
nand U1398 (N_1398,N_675,N_777);
or U1399 (N_1399,N_738,N_861);
and U1400 (N_1400,N_667,N_568);
nor U1401 (N_1401,N_707,N_779);
nor U1402 (N_1402,N_987,N_674);
nand U1403 (N_1403,N_807,N_599);
nand U1404 (N_1404,N_760,N_628);
and U1405 (N_1405,N_658,N_858);
nand U1406 (N_1406,N_811,N_847);
xor U1407 (N_1407,N_614,N_851);
xor U1408 (N_1408,N_988,N_768);
nand U1409 (N_1409,N_655,N_653);
or U1410 (N_1410,N_514,N_712);
xnor U1411 (N_1411,N_791,N_900);
and U1412 (N_1412,N_599,N_658);
or U1413 (N_1413,N_532,N_734);
nand U1414 (N_1414,N_549,N_735);
or U1415 (N_1415,N_996,N_820);
and U1416 (N_1416,N_773,N_525);
nor U1417 (N_1417,N_598,N_675);
nand U1418 (N_1418,N_531,N_670);
nor U1419 (N_1419,N_777,N_609);
and U1420 (N_1420,N_840,N_744);
and U1421 (N_1421,N_508,N_773);
nand U1422 (N_1422,N_557,N_622);
xnor U1423 (N_1423,N_789,N_521);
or U1424 (N_1424,N_980,N_796);
and U1425 (N_1425,N_778,N_998);
and U1426 (N_1426,N_580,N_669);
nand U1427 (N_1427,N_889,N_835);
xnor U1428 (N_1428,N_508,N_877);
nor U1429 (N_1429,N_790,N_845);
or U1430 (N_1430,N_598,N_897);
or U1431 (N_1431,N_592,N_991);
xor U1432 (N_1432,N_658,N_765);
and U1433 (N_1433,N_983,N_580);
or U1434 (N_1434,N_738,N_586);
or U1435 (N_1435,N_534,N_997);
nor U1436 (N_1436,N_944,N_754);
nand U1437 (N_1437,N_951,N_594);
nor U1438 (N_1438,N_542,N_549);
and U1439 (N_1439,N_652,N_728);
and U1440 (N_1440,N_631,N_866);
nand U1441 (N_1441,N_594,N_502);
nor U1442 (N_1442,N_530,N_659);
or U1443 (N_1443,N_617,N_718);
nor U1444 (N_1444,N_833,N_659);
or U1445 (N_1445,N_640,N_808);
and U1446 (N_1446,N_846,N_848);
nand U1447 (N_1447,N_559,N_512);
nand U1448 (N_1448,N_512,N_533);
xnor U1449 (N_1449,N_701,N_922);
or U1450 (N_1450,N_945,N_824);
and U1451 (N_1451,N_956,N_614);
xnor U1452 (N_1452,N_642,N_974);
and U1453 (N_1453,N_612,N_895);
nand U1454 (N_1454,N_712,N_560);
or U1455 (N_1455,N_898,N_938);
xor U1456 (N_1456,N_706,N_918);
or U1457 (N_1457,N_876,N_685);
xnor U1458 (N_1458,N_671,N_966);
and U1459 (N_1459,N_508,N_744);
xnor U1460 (N_1460,N_869,N_755);
and U1461 (N_1461,N_908,N_806);
or U1462 (N_1462,N_785,N_502);
or U1463 (N_1463,N_695,N_831);
xnor U1464 (N_1464,N_792,N_800);
xor U1465 (N_1465,N_707,N_538);
and U1466 (N_1466,N_649,N_677);
nor U1467 (N_1467,N_598,N_739);
nand U1468 (N_1468,N_590,N_500);
nor U1469 (N_1469,N_720,N_838);
nand U1470 (N_1470,N_858,N_784);
or U1471 (N_1471,N_719,N_709);
nand U1472 (N_1472,N_584,N_675);
nor U1473 (N_1473,N_543,N_618);
xor U1474 (N_1474,N_888,N_727);
nand U1475 (N_1475,N_537,N_773);
xnor U1476 (N_1476,N_607,N_587);
nand U1477 (N_1477,N_743,N_521);
xnor U1478 (N_1478,N_874,N_810);
xor U1479 (N_1479,N_850,N_990);
xnor U1480 (N_1480,N_543,N_770);
and U1481 (N_1481,N_557,N_943);
and U1482 (N_1482,N_809,N_631);
nor U1483 (N_1483,N_548,N_610);
nand U1484 (N_1484,N_745,N_667);
or U1485 (N_1485,N_642,N_704);
or U1486 (N_1486,N_745,N_818);
or U1487 (N_1487,N_897,N_519);
nand U1488 (N_1488,N_795,N_773);
xor U1489 (N_1489,N_769,N_853);
or U1490 (N_1490,N_580,N_935);
or U1491 (N_1491,N_617,N_516);
xnor U1492 (N_1492,N_935,N_682);
or U1493 (N_1493,N_588,N_504);
and U1494 (N_1494,N_956,N_778);
or U1495 (N_1495,N_922,N_706);
or U1496 (N_1496,N_675,N_589);
or U1497 (N_1497,N_791,N_779);
xnor U1498 (N_1498,N_701,N_932);
nor U1499 (N_1499,N_889,N_962);
and U1500 (N_1500,N_1036,N_1266);
or U1501 (N_1501,N_1244,N_1462);
xnor U1502 (N_1502,N_1281,N_1476);
or U1503 (N_1503,N_1322,N_1238);
nor U1504 (N_1504,N_1091,N_1202);
nor U1505 (N_1505,N_1320,N_1215);
nand U1506 (N_1506,N_1090,N_1368);
nand U1507 (N_1507,N_1358,N_1373);
or U1508 (N_1508,N_1068,N_1415);
nand U1509 (N_1509,N_1159,N_1121);
xnor U1510 (N_1510,N_1458,N_1242);
nand U1511 (N_1511,N_1118,N_1126);
and U1512 (N_1512,N_1265,N_1097);
xor U1513 (N_1513,N_1285,N_1189);
and U1514 (N_1514,N_1143,N_1085);
or U1515 (N_1515,N_1472,N_1117);
nor U1516 (N_1516,N_1195,N_1457);
and U1517 (N_1517,N_1404,N_1182);
and U1518 (N_1518,N_1475,N_1100);
and U1519 (N_1519,N_1257,N_1443);
and U1520 (N_1520,N_1156,N_1024);
nand U1521 (N_1521,N_1372,N_1310);
or U1522 (N_1522,N_1383,N_1234);
and U1523 (N_1523,N_1104,N_1335);
nor U1524 (N_1524,N_1101,N_1453);
and U1525 (N_1525,N_1173,N_1051);
nand U1526 (N_1526,N_1055,N_1108);
xor U1527 (N_1527,N_1154,N_1141);
xor U1528 (N_1528,N_1066,N_1326);
or U1529 (N_1529,N_1390,N_1021);
nand U1530 (N_1530,N_1218,N_1065);
and U1531 (N_1531,N_1345,N_1003);
or U1532 (N_1532,N_1061,N_1305);
nor U1533 (N_1533,N_1029,N_1431);
nor U1534 (N_1534,N_1371,N_1214);
xnor U1535 (N_1535,N_1325,N_1317);
and U1536 (N_1536,N_1425,N_1471);
xor U1537 (N_1537,N_1445,N_1174);
xnor U1538 (N_1538,N_1172,N_1137);
or U1539 (N_1539,N_1083,N_1221);
nor U1540 (N_1540,N_1228,N_1477);
xor U1541 (N_1541,N_1275,N_1247);
nand U1542 (N_1542,N_1171,N_1451);
or U1543 (N_1543,N_1349,N_1364);
and U1544 (N_1544,N_1348,N_1395);
or U1545 (N_1545,N_1139,N_1303);
nand U1546 (N_1546,N_1329,N_1054);
nand U1547 (N_1547,N_1465,N_1463);
or U1548 (N_1548,N_1336,N_1180);
nand U1549 (N_1549,N_1072,N_1384);
and U1550 (N_1550,N_1352,N_1089);
nor U1551 (N_1551,N_1488,N_1170);
xnor U1552 (N_1552,N_1338,N_1005);
and U1553 (N_1553,N_1304,N_1071);
nand U1554 (N_1554,N_1355,N_1436);
xor U1555 (N_1555,N_1429,N_1125);
xnor U1556 (N_1556,N_1251,N_1119);
nor U1557 (N_1557,N_1194,N_1366);
nor U1558 (N_1558,N_1363,N_1239);
xnor U1559 (N_1559,N_1377,N_1216);
xnor U1560 (N_1560,N_1403,N_1058);
nand U1561 (N_1561,N_1049,N_1205);
nor U1562 (N_1562,N_1070,N_1427);
nor U1563 (N_1563,N_1344,N_1045);
or U1564 (N_1564,N_1290,N_1032);
nor U1565 (N_1565,N_1387,N_1056);
nor U1566 (N_1566,N_1134,N_1080);
xor U1567 (N_1567,N_1292,N_1002);
nand U1568 (N_1568,N_1016,N_1319);
nor U1569 (N_1569,N_1167,N_1391);
and U1570 (N_1570,N_1294,N_1069);
nor U1571 (N_1571,N_1004,N_1213);
or U1572 (N_1572,N_1444,N_1494);
nand U1573 (N_1573,N_1112,N_1008);
and U1574 (N_1574,N_1307,N_1035);
nand U1575 (N_1575,N_1144,N_1411);
nor U1576 (N_1576,N_1313,N_1116);
and U1577 (N_1577,N_1256,N_1211);
and U1578 (N_1578,N_1258,N_1152);
or U1579 (N_1579,N_1284,N_1495);
nor U1580 (N_1580,N_1074,N_1460);
and U1581 (N_1581,N_1375,N_1400);
nor U1582 (N_1582,N_1081,N_1381);
and U1583 (N_1583,N_1276,N_1064);
and U1584 (N_1584,N_1176,N_1379);
xnor U1585 (N_1585,N_1146,N_1328);
or U1586 (N_1586,N_1461,N_1433);
or U1587 (N_1587,N_1014,N_1198);
nand U1588 (N_1588,N_1306,N_1380);
or U1589 (N_1589,N_1127,N_1405);
and U1590 (N_1590,N_1470,N_1434);
or U1591 (N_1591,N_1190,N_1267);
nand U1592 (N_1592,N_1446,N_1374);
nor U1593 (N_1593,N_1034,N_1312);
nand U1594 (N_1594,N_1212,N_1426);
or U1595 (N_1595,N_1455,N_1311);
nand U1596 (N_1596,N_1342,N_1327);
nor U1597 (N_1597,N_1086,N_1210);
xnor U1598 (N_1598,N_1224,N_1177);
and U1599 (N_1599,N_1407,N_1401);
nor U1600 (N_1600,N_1498,N_1353);
or U1601 (N_1601,N_1454,N_1044);
nand U1602 (N_1602,N_1236,N_1011);
nor U1603 (N_1603,N_1145,N_1038);
xnor U1604 (N_1604,N_1408,N_1330);
nor U1605 (N_1605,N_1122,N_1283);
nand U1606 (N_1606,N_1492,N_1356);
or U1607 (N_1607,N_1113,N_1346);
xnor U1608 (N_1608,N_1094,N_1042);
xor U1609 (N_1609,N_1006,N_1023);
nand U1610 (N_1610,N_1447,N_1440);
nor U1611 (N_1611,N_1120,N_1343);
xnor U1612 (N_1612,N_1262,N_1153);
and U1613 (N_1613,N_1333,N_1027);
nand U1614 (N_1614,N_1482,N_1417);
nand U1615 (N_1615,N_1199,N_1208);
xnor U1616 (N_1616,N_1220,N_1332);
or U1617 (N_1617,N_1123,N_1273);
nor U1618 (N_1618,N_1192,N_1219);
xor U1619 (N_1619,N_1413,N_1428);
nor U1620 (N_1620,N_1481,N_1206);
nor U1621 (N_1621,N_1160,N_1185);
or U1622 (N_1622,N_1250,N_1450);
xor U1623 (N_1623,N_1389,N_1225);
xor U1624 (N_1624,N_1394,N_1111);
and U1625 (N_1625,N_1323,N_1217);
nand U1626 (N_1626,N_1102,N_1096);
nand U1627 (N_1627,N_1485,N_1286);
nand U1628 (N_1628,N_1232,N_1186);
and U1629 (N_1629,N_1196,N_1288);
nor U1630 (N_1630,N_1249,N_1017);
nor U1631 (N_1631,N_1204,N_1087);
or U1632 (N_1632,N_1388,N_1253);
or U1633 (N_1633,N_1489,N_1063);
and U1634 (N_1634,N_1382,N_1149);
nor U1635 (N_1635,N_1001,N_1359);
xor U1636 (N_1636,N_1077,N_1438);
nor U1637 (N_1637,N_1106,N_1222);
xor U1638 (N_1638,N_1295,N_1264);
nor U1639 (N_1639,N_1135,N_1420);
nor U1640 (N_1640,N_1050,N_1230);
xor U1641 (N_1641,N_1467,N_1015);
xor U1642 (N_1642,N_1059,N_1132);
or U1643 (N_1643,N_1456,N_1191);
and U1644 (N_1644,N_1103,N_1107);
xnor U1645 (N_1645,N_1184,N_1291);
xor U1646 (N_1646,N_1398,N_1200);
nor U1647 (N_1647,N_1067,N_1164);
or U1648 (N_1648,N_1270,N_1010);
nand U1649 (N_1649,N_1496,N_1115);
nor U1650 (N_1650,N_1020,N_1399);
and U1651 (N_1651,N_1130,N_1142);
nand U1652 (N_1652,N_1110,N_1442);
nand U1653 (N_1653,N_1278,N_1478);
xor U1654 (N_1654,N_1412,N_1047);
or U1655 (N_1655,N_1084,N_1298);
xnor U1656 (N_1656,N_1252,N_1223);
and U1657 (N_1657,N_1423,N_1314);
nand U1658 (N_1658,N_1009,N_1464);
nand U1659 (N_1659,N_1237,N_1088);
nor U1660 (N_1660,N_1316,N_1293);
and U1661 (N_1661,N_1357,N_1497);
nand U1662 (N_1662,N_1486,N_1227);
or U1663 (N_1663,N_1337,N_1255);
nand U1664 (N_1664,N_1057,N_1155);
nand U1665 (N_1665,N_1421,N_1441);
or U1666 (N_1666,N_1432,N_1300);
xor U1667 (N_1667,N_1233,N_1302);
nor U1668 (N_1668,N_1261,N_1490);
and U1669 (N_1669,N_1414,N_1148);
and U1670 (N_1670,N_1028,N_1416);
and U1671 (N_1671,N_1092,N_1370);
xnor U1672 (N_1672,N_1402,N_1385);
xnor U1673 (N_1673,N_1183,N_1289);
nor U1674 (N_1674,N_1165,N_1272);
nand U1675 (N_1675,N_1138,N_1282);
nand U1676 (N_1676,N_1422,N_1297);
nand U1677 (N_1677,N_1339,N_1157);
nand U1678 (N_1678,N_1109,N_1140);
or U1679 (N_1679,N_1075,N_1324);
or U1680 (N_1680,N_1240,N_1062);
xnor U1681 (N_1681,N_1418,N_1361);
nand U1682 (N_1682,N_1147,N_1365);
and U1683 (N_1683,N_1133,N_1287);
or U1684 (N_1684,N_1318,N_1207);
and U1685 (N_1685,N_1340,N_1007);
nand U1686 (N_1686,N_1060,N_1301);
or U1687 (N_1687,N_1452,N_1019);
and U1688 (N_1688,N_1468,N_1277);
or U1689 (N_1689,N_1181,N_1201);
or U1690 (N_1690,N_1248,N_1095);
nand U1691 (N_1691,N_1169,N_1082);
or U1692 (N_1692,N_1309,N_1025);
nand U1693 (N_1693,N_1410,N_1166);
nor U1694 (N_1694,N_1033,N_1136);
and U1695 (N_1695,N_1269,N_1271);
xor U1696 (N_1696,N_1026,N_1168);
nand U1697 (N_1697,N_1376,N_1052);
nand U1698 (N_1698,N_1079,N_1369);
xnor U1699 (N_1699,N_1430,N_1041);
xor U1700 (N_1700,N_1012,N_1279);
xor U1701 (N_1701,N_1483,N_1437);
nor U1702 (N_1702,N_1243,N_1193);
xnor U1703 (N_1703,N_1474,N_1098);
xnor U1704 (N_1704,N_1076,N_1209);
and U1705 (N_1705,N_1179,N_1484);
and U1706 (N_1706,N_1048,N_1254);
xnor U1707 (N_1707,N_1280,N_1000);
nor U1708 (N_1708,N_1499,N_1334);
nor U1709 (N_1709,N_1386,N_1274);
or U1710 (N_1710,N_1321,N_1073);
or U1711 (N_1711,N_1187,N_1362);
xor U1712 (N_1712,N_1435,N_1131);
xor U1713 (N_1713,N_1093,N_1259);
and U1714 (N_1714,N_1392,N_1473);
and U1715 (N_1715,N_1053,N_1161);
xor U1716 (N_1716,N_1409,N_1491);
xor U1717 (N_1717,N_1203,N_1449);
nand U1718 (N_1718,N_1018,N_1099);
xor U1719 (N_1719,N_1378,N_1393);
nand U1720 (N_1720,N_1396,N_1299);
xnor U1721 (N_1721,N_1162,N_1235);
and U1722 (N_1722,N_1479,N_1163);
xor U1723 (N_1723,N_1241,N_1448);
or U1724 (N_1724,N_1040,N_1360);
nand U1725 (N_1725,N_1022,N_1188);
nor U1726 (N_1726,N_1459,N_1078);
nor U1727 (N_1727,N_1031,N_1397);
or U1728 (N_1728,N_1175,N_1331);
or U1729 (N_1729,N_1341,N_1351);
xor U1730 (N_1730,N_1487,N_1150);
or U1731 (N_1731,N_1229,N_1129);
nand U1732 (N_1732,N_1354,N_1114);
and U1733 (N_1733,N_1367,N_1406);
nand U1734 (N_1734,N_1151,N_1480);
or U1735 (N_1735,N_1124,N_1037);
or U1736 (N_1736,N_1493,N_1296);
xor U1737 (N_1737,N_1043,N_1030);
nor U1738 (N_1738,N_1231,N_1245);
and U1739 (N_1739,N_1246,N_1347);
xnor U1740 (N_1740,N_1178,N_1197);
nand U1741 (N_1741,N_1424,N_1350);
nor U1742 (N_1742,N_1039,N_1013);
nor U1743 (N_1743,N_1466,N_1308);
and U1744 (N_1744,N_1128,N_1315);
xor U1745 (N_1745,N_1268,N_1226);
or U1746 (N_1746,N_1439,N_1105);
or U1747 (N_1747,N_1419,N_1263);
nand U1748 (N_1748,N_1469,N_1158);
or U1749 (N_1749,N_1046,N_1260);
and U1750 (N_1750,N_1195,N_1199);
nor U1751 (N_1751,N_1318,N_1179);
xor U1752 (N_1752,N_1371,N_1370);
xnor U1753 (N_1753,N_1302,N_1305);
or U1754 (N_1754,N_1383,N_1041);
xor U1755 (N_1755,N_1314,N_1190);
or U1756 (N_1756,N_1093,N_1304);
xor U1757 (N_1757,N_1126,N_1260);
nor U1758 (N_1758,N_1144,N_1431);
xnor U1759 (N_1759,N_1076,N_1037);
and U1760 (N_1760,N_1107,N_1203);
nand U1761 (N_1761,N_1217,N_1236);
xor U1762 (N_1762,N_1310,N_1138);
or U1763 (N_1763,N_1419,N_1255);
or U1764 (N_1764,N_1480,N_1234);
or U1765 (N_1765,N_1133,N_1466);
nand U1766 (N_1766,N_1230,N_1034);
and U1767 (N_1767,N_1134,N_1160);
xnor U1768 (N_1768,N_1121,N_1313);
nor U1769 (N_1769,N_1056,N_1475);
and U1770 (N_1770,N_1300,N_1028);
and U1771 (N_1771,N_1161,N_1042);
and U1772 (N_1772,N_1270,N_1415);
xor U1773 (N_1773,N_1212,N_1187);
xnor U1774 (N_1774,N_1255,N_1119);
xor U1775 (N_1775,N_1410,N_1446);
or U1776 (N_1776,N_1323,N_1335);
and U1777 (N_1777,N_1462,N_1204);
nor U1778 (N_1778,N_1210,N_1221);
or U1779 (N_1779,N_1339,N_1483);
nor U1780 (N_1780,N_1206,N_1182);
nand U1781 (N_1781,N_1321,N_1464);
nor U1782 (N_1782,N_1379,N_1237);
xnor U1783 (N_1783,N_1383,N_1084);
nor U1784 (N_1784,N_1242,N_1219);
nand U1785 (N_1785,N_1384,N_1185);
or U1786 (N_1786,N_1492,N_1363);
and U1787 (N_1787,N_1406,N_1114);
nor U1788 (N_1788,N_1216,N_1410);
or U1789 (N_1789,N_1356,N_1144);
xnor U1790 (N_1790,N_1325,N_1132);
or U1791 (N_1791,N_1177,N_1084);
nor U1792 (N_1792,N_1159,N_1180);
and U1793 (N_1793,N_1077,N_1295);
nand U1794 (N_1794,N_1253,N_1000);
and U1795 (N_1795,N_1168,N_1084);
or U1796 (N_1796,N_1288,N_1383);
nand U1797 (N_1797,N_1489,N_1183);
or U1798 (N_1798,N_1412,N_1499);
and U1799 (N_1799,N_1234,N_1349);
or U1800 (N_1800,N_1376,N_1455);
nand U1801 (N_1801,N_1306,N_1447);
xor U1802 (N_1802,N_1441,N_1037);
xnor U1803 (N_1803,N_1061,N_1082);
and U1804 (N_1804,N_1372,N_1365);
nand U1805 (N_1805,N_1015,N_1390);
nor U1806 (N_1806,N_1077,N_1366);
nor U1807 (N_1807,N_1264,N_1066);
and U1808 (N_1808,N_1020,N_1496);
nor U1809 (N_1809,N_1164,N_1269);
nor U1810 (N_1810,N_1115,N_1374);
nor U1811 (N_1811,N_1048,N_1059);
or U1812 (N_1812,N_1066,N_1078);
xor U1813 (N_1813,N_1260,N_1433);
nor U1814 (N_1814,N_1267,N_1227);
and U1815 (N_1815,N_1217,N_1290);
or U1816 (N_1816,N_1381,N_1045);
and U1817 (N_1817,N_1436,N_1267);
and U1818 (N_1818,N_1381,N_1040);
nand U1819 (N_1819,N_1098,N_1273);
or U1820 (N_1820,N_1478,N_1030);
and U1821 (N_1821,N_1296,N_1344);
and U1822 (N_1822,N_1236,N_1021);
nor U1823 (N_1823,N_1271,N_1305);
nor U1824 (N_1824,N_1448,N_1267);
xor U1825 (N_1825,N_1487,N_1271);
and U1826 (N_1826,N_1026,N_1377);
nand U1827 (N_1827,N_1033,N_1060);
nand U1828 (N_1828,N_1384,N_1281);
and U1829 (N_1829,N_1335,N_1424);
and U1830 (N_1830,N_1092,N_1234);
nor U1831 (N_1831,N_1141,N_1348);
nor U1832 (N_1832,N_1086,N_1327);
nand U1833 (N_1833,N_1364,N_1130);
xor U1834 (N_1834,N_1465,N_1333);
or U1835 (N_1835,N_1204,N_1088);
and U1836 (N_1836,N_1215,N_1345);
and U1837 (N_1837,N_1035,N_1433);
nor U1838 (N_1838,N_1209,N_1486);
or U1839 (N_1839,N_1191,N_1148);
and U1840 (N_1840,N_1429,N_1188);
and U1841 (N_1841,N_1427,N_1140);
nand U1842 (N_1842,N_1432,N_1178);
nand U1843 (N_1843,N_1155,N_1494);
or U1844 (N_1844,N_1215,N_1458);
nand U1845 (N_1845,N_1047,N_1291);
xnor U1846 (N_1846,N_1333,N_1249);
nand U1847 (N_1847,N_1282,N_1210);
and U1848 (N_1848,N_1071,N_1350);
nor U1849 (N_1849,N_1457,N_1283);
or U1850 (N_1850,N_1164,N_1185);
xnor U1851 (N_1851,N_1326,N_1152);
or U1852 (N_1852,N_1296,N_1314);
nor U1853 (N_1853,N_1122,N_1323);
nor U1854 (N_1854,N_1456,N_1355);
and U1855 (N_1855,N_1138,N_1055);
nand U1856 (N_1856,N_1240,N_1013);
nand U1857 (N_1857,N_1452,N_1426);
or U1858 (N_1858,N_1137,N_1428);
and U1859 (N_1859,N_1104,N_1271);
xor U1860 (N_1860,N_1065,N_1354);
or U1861 (N_1861,N_1027,N_1324);
and U1862 (N_1862,N_1497,N_1150);
nand U1863 (N_1863,N_1099,N_1063);
and U1864 (N_1864,N_1179,N_1449);
and U1865 (N_1865,N_1092,N_1240);
xnor U1866 (N_1866,N_1008,N_1044);
or U1867 (N_1867,N_1329,N_1200);
xor U1868 (N_1868,N_1234,N_1239);
nand U1869 (N_1869,N_1111,N_1372);
and U1870 (N_1870,N_1244,N_1461);
nand U1871 (N_1871,N_1124,N_1287);
or U1872 (N_1872,N_1468,N_1306);
or U1873 (N_1873,N_1027,N_1371);
xnor U1874 (N_1874,N_1189,N_1323);
nor U1875 (N_1875,N_1498,N_1010);
and U1876 (N_1876,N_1459,N_1021);
xnor U1877 (N_1877,N_1382,N_1081);
or U1878 (N_1878,N_1407,N_1249);
and U1879 (N_1879,N_1293,N_1425);
or U1880 (N_1880,N_1196,N_1323);
xnor U1881 (N_1881,N_1042,N_1123);
or U1882 (N_1882,N_1160,N_1279);
nand U1883 (N_1883,N_1417,N_1065);
nand U1884 (N_1884,N_1050,N_1156);
and U1885 (N_1885,N_1004,N_1104);
and U1886 (N_1886,N_1138,N_1359);
or U1887 (N_1887,N_1459,N_1139);
nand U1888 (N_1888,N_1400,N_1270);
or U1889 (N_1889,N_1201,N_1117);
xor U1890 (N_1890,N_1341,N_1011);
and U1891 (N_1891,N_1233,N_1184);
xor U1892 (N_1892,N_1032,N_1168);
nand U1893 (N_1893,N_1219,N_1479);
nand U1894 (N_1894,N_1077,N_1495);
or U1895 (N_1895,N_1331,N_1248);
and U1896 (N_1896,N_1492,N_1493);
xor U1897 (N_1897,N_1327,N_1077);
and U1898 (N_1898,N_1318,N_1157);
nand U1899 (N_1899,N_1096,N_1339);
or U1900 (N_1900,N_1182,N_1057);
and U1901 (N_1901,N_1247,N_1484);
nor U1902 (N_1902,N_1256,N_1411);
or U1903 (N_1903,N_1203,N_1087);
and U1904 (N_1904,N_1362,N_1057);
and U1905 (N_1905,N_1471,N_1163);
nor U1906 (N_1906,N_1417,N_1268);
or U1907 (N_1907,N_1270,N_1022);
nor U1908 (N_1908,N_1004,N_1324);
xor U1909 (N_1909,N_1115,N_1381);
or U1910 (N_1910,N_1471,N_1279);
nand U1911 (N_1911,N_1456,N_1468);
and U1912 (N_1912,N_1364,N_1206);
nor U1913 (N_1913,N_1302,N_1091);
nor U1914 (N_1914,N_1038,N_1162);
or U1915 (N_1915,N_1016,N_1054);
xnor U1916 (N_1916,N_1286,N_1021);
nand U1917 (N_1917,N_1238,N_1282);
nor U1918 (N_1918,N_1291,N_1163);
nand U1919 (N_1919,N_1191,N_1105);
or U1920 (N_1920,N_1472,N_1257);
and U1921 (N_1921,N_1269,N_1275);
nor U1922 (N_1922,N_1301,N_1377);
nand U1923 (N_1923,N_1006,N_1005);
nor U1924 (N_1924,N_1095,N_1429);
xnor U1925 (N_1925,N_1155,N_1224);
and U1926 (N_1926,N_1352,N_1255);
xor U1927 (N_1927,N_1489,N_1497);
nor U1928 (N_1928,N_1490,N_1472);
or U1929 (N_1929,N_1149,N_1165);
nor U1930 (N_1930,N_1265,N_1412);
nor U1931 (N_1931,N_1239,N_1175);
or U1932 (N_1932,N_1120,N_1084);
or U1933 (N_1933,N_1460,N_1145);
and U1934 (N_1934,N_1389,N_1332);
nor U1935 (N_1935,N_1350,N_1042);
nand U1936 (N_1936,N_1252,N_1255);
and U1937 (N_1937,N_1306,N_1079);
nor U1938 (N_1938,N_1174,N_1074);
nand U1939 (N_1939,N_1411,N_1038);
and U1940 (N_1940,N_1200,N_1063);
and U1941 (N_1941,N_1206,N_1025);
nand U1942 (N_1942,N_1083,N_1293);
xnor U1943 (N_1943,N_1304,N_1020);
nor U1944 (N_1944,N_1172,N_1216);
nand U1945 (N_1945,N_1246,N_1013);
nor U1946 (N_1946,N_1035,N_1334);
xnor U1947 (N_1947,N_1290,N_1136);
xor U1948 (N_1948,N_1217,N_1477);
xor U1949 (N_1949,N_1294,N_1362);
or U1950 (N_1950,N_1490,N_1306);
and U1951 (N_1951,N_1394,N_1441);
nor U1952 (N_1952,N_1238,N_1296);
nand U1953 (N_1953,N_1361,N_1409);
or U1954 (N_1954,N_1480,N_1073);
or U1955 (N_1955,N_1389,N_1254);
and U1956 (N_1956,N_1129,N_1362);
and U1957 (N_1957,N_1115,N_1101);
nor U1958 (N_1958,N_1400,N_1319);
nand U1959 (N_1959,N_1156,N_1040);
or U1960 (N_1960,N_1411,N_1145);
and U1961 (N_1961,N_1263,N_1359);
and U1962 (N_1962,N_1290,N_1078);
xor U1963 (N_1963,N_1468,N_1385);
and U1964 (N_1964,N_1327,N_1223);
or U1965 (N_1965,N_1188,N_1450);
xnor U1966 (N_1966,N_1426,N_1477);
xnor U1967 (N_1967,N_1246,N_1049);
or U1968 (N_1968,N_1085,N_1431);
nor U1969 (N_1969,N_1352,N_1380);
nand U1970 (N_1970,N_1016,N_1071);
nand U1971 (N_1971,N_1260,N_1421);
nand U1972 (N_1972,N_1469,N_1421);
xor U1973 (N_1973,N_1099,N_1219);
nor U1974 (N_1974,N_1212,N_1018);
or U1975 (N_1975,N_1367,N_1412);
and U1976 (N_1976,N_1187,N_1301);
or U1977 (N_1977,N_1403,N_1492);
and U1978 (N_1978,N_1240,N_1449);
nand U1979 (N_1979,N_1247,N_1161);
nand U1980 (N_1980,N_1364,N_1272);
and U1981 (N_1981,N_1486,N_1472);
or U1982 (N_1982,N_1185,N_1007);
nand U1983 (N_1983,N_1113,N_1473);
xor U1984 (N_1984,N_1206,N_1411);
nand U1985 (N_1985,N_1061,N_1410);
and U1986 (N_1986,N_1001,N_1387);
nor U1987 (N_1987,N_1285,N_1340);
or U1988 (N_1988,N_1022,N_1350);
nor U1989 (N_1989,N_1273,N_1375);
nor U1990 (N_1990,N_1095,N_1259);
and U1991 (N_1991,N_1142,N_1297);
and U1992 (N_1992,N_1179,N_1386);
or U1993 (N_1993,N_1050,N_1082);
and U1994 (N_1994,N_1148,N_1327);
nor U1995 (N_1995,N_1139,N_1105);
nand U1996 (N_1996,N_1191,N_1131);
or U1997 (N_1997,N_1079,N_1284);
xnor U1998 (N_1998,N_1369,N_1312);
or U1999 (N_1999,N_1226,N_1316);
and U2000 (N_2000,N_1811,N_1921);
nor U2001 (N_2001,N_1567,N_1850);
xnor U2002 (N_2002,N_1572,N_1605);
xnor U2003 (N_2003,N_1949,N_1543);
or U2004 (N_2004,N_1564,N_1535);
xor U2005 (N_2005,N_1731,N_1941);
xnor U2006 (N_2006,N_1808,N_1822);
xor U2007 (N_2007,N_1976,N_1788);
nor U2008 (N_2008,N_1696,N_1719);
or U2009 (N_2009,N_1958,N_1702);
nand U2010 (N_2010,N_1926,N_1757);
nor U2011 (N_2011,N_1574,N_1721);
xnor U2012 (N_2012,N_1910,N_1549);
and U2013 (N_2013,N_1909,N_1751);
nand U2014 (N_2014,N_1943,N_1935);
nand U2015 (N_2015,N_1982,N_1857);
and U2016 (N_2016,N_1652,N_1948);
or U2017 (N_2017,N_1946,N_1749);
or U2018 (N_2018,N_1710,N_1825);
nor U2019 (N_2019,N_1806,N_1783);
nand U2020 (N_2020,N_1858,N_1810);
or U2021 (N_2021,N_1873,N_1699);
and U2022 (N_2022,N_1888,N_1595);
nand U2023 (N_2023,N_1774,N_1604);
and U2024 (N_2024,N_1724,N_1578);
xor U2025 (N_2025,N_1905,N_1688);
or U2026 (N_2026,N_1633,N_1695);
and U2027 (N_2027,N_1869,N_1678);
nand U2028 (N_2028,N_1720,N_1996);
or U2029 (N_2029,N_1944,N_1534);
nand U2030 (N_2030,N_1738,N_1583);
xor U2031 (N_2031,N_1906,N_1883);
and U2032 (N_2032,N_1853,N_1815);
or U2033 (N_2033,N_1507,N_1927);
and U2034 (N_2034,N_1668,N_1548);
or U2035 (N_2035,N_1618,N_1840);
nand U2036 (N_2036,N_1653,N_1615);
and U2037 (N_2037,N_1860,N_1947);
nand U2038 (N_2038,N_1940,N_1813);
nand U2039 (N_2039,N_1717,N_1861);
or U2040 (N_2040,N_1977,N_1991);
or U2041 (N_2041,N_1586,N_1866);
nand U2042 (N_2042,N_1638,N_1966);
and U2043 (N_2043,N_1832,N_1989);
and U2044 (N_2044,N_1786,N_1896);
xnor U2045 (N_2045,N_1609,N_1684);
and U2046 (N_2046,N_1865,N_1831);
xnor U2047 (N_2047,N_1995,N_1864);
or U2048 (N_2048,N_1672,N_1826);
and U2049 (N_2049,N_1558,N_1670);
or U2050 (N_2050,N_1990,N_1796);
and U2051 (N_2051,N_1552,N_1897);
nor U2052 (N_2052,N_1907,N_1664);
xor U2053 (N_2053,N_1568,N_1761);
nand U2054 (N_2054,N_1758,N_1984);
nor U2055 (N_2055,N_1703,N_1630);
nor U2056 (N_2056,N_1973,N_1562);
and U2057 (N_2057,N_1818,N_1854);
or U2058 (N_2058,N_1537,N_1592);
and U2059 (N_2059,N_1878,N_1817);
xor U2060 (N_2060,N_1621,N_1685);
xnor U2061 (N_2061,N_1521,N_1506);
or U2062 (N_2062,N_1950,N_1980);
or U2063 (N_2063,N_1975,N_1573);
nor U2064 (N_2064,N_1561,N_1901);
nand U2065 (N_2065,N_1848,N_1969);
xor U2066 (N_2066,N_1974,N_1683);
nand U2067 (N_2067,N_1563,N_1928);
nor U2068 (N_2068,N_1547,N_1899);
xnor U2069 (N_2069,N_1747,N_1934);
nand U2070 (N_2070,N_1556,N_1530);
nor U2071 (N_2071,N_1663,N_1654);
and U2072 (N_2072,N_1734,N_1765);
nor U2073 (N_2073,N_1676,N_1797);
nand U2074 (N_2074,N_1518,N_1776);
and U2075 (N_2075,N_1784,N_1704);
or U2076 (N_2076,N_1687,N_1740);
or U2077 (N_2077,N_1876,N_1802);
nand U2078 (N_2078,N_1525,N_1744);
nor U2079 (N_2079,N_1642,N_1753);
or U2080 (N_2080,N_1680,N_1903);
or U2081 (N_2081,N_1904,N_1780);
or U2082 (N_2082,N_1644,N_1871);
or U2083 (N_2083,N_1646,N_1951);
and U2084 (N_2084,N_1924,N_1981);
xnor U2085 (N_2085,N_1994,N_1536);
xor U2086 (N_2086,N_1681,N_1546);
and U2087 (N_2087,N_1775,N_1824);
or U2088 (N_2088,N_1849,N_1730);
nand U2089 (N_2089,N_1637,N_1691);
or U2090 (N_2090,N_1819,N_1656);
or U2091 (N_2091,N_1659,N_1891);
nor U2092 (N_2092,N_1533,N_1713);
xnor U2093 (N_2093,N_1885,N_1725);
and U2094 (N_2094,N_1660,N_1877);
xor U2095 (N_2095,N_1698,N_1580);
nand U2096 (N_2096,N_1922,N_1923);
or U2097 (N_2097,N_1560,N_1636);
xor U2098 (N_2098,N_1581,N_1576);
xor U2099 (N_2099,N_1998,N_1961);
and U2100 (N_2100,N_1963,N_1945);
nor U2101 (N_2101,N_1647,N_1508);
and U2102 (N_2102,N_1942,N_1582);
or U2103 (N_2103,N_1515,N_1862);
nand U2104 (N_2104,N_1985,N_1787);
xor U2105 (N_2105,N_1502,N_1575);
xnor U2106 (N_2106,N_1657,N_1809);
nand U2107 (N_2107,N_1778,N_1844);
xnor U2108 (N_2108,N_1953,N_1614);
xnor U2109 (N_2109,N_1514,N_1645);
nand U2110 (N_2110,N_1754,N_1523);
or U2111 (N_2111,N_1544,N_1936);
xor U2112 (N_2112,N_1594,N_1920);
or U2113 (N_2113,N_1629,N_1735);
and U2114 (N_2114,N_1919,N_1870);
nand U2115 (N_2115,N_1500,N_1895);
nor U2116 (N_2116,N_1624,N_1827);
nand U2117 (N_2117,N_1643,N_1954);
and U2118 (N_2118,N_1671,N_1874);
nand U2119 (N_2119,N_1501,N_1690);
or U2120 (N_2120,N_1988,N_1913);
and U2121 (N_2121,N_1992,N_1833);
and U2122 (N_2122,N_1750,N_1851);
or U2123 (N_2123,N_1807,N_1520);
or U2124 (N_2124,N_1596,N_1569);
nor U2125 (N_2125,N_1606,N_1872);
or U2126 (N_2126,N_1648,N_1804);
nand U2127 (N_2127,N_1587,N_1829);
nand U2128 (N_2128,N_1799,N_1839);
xnor U2129 (N_2129,N_1894,N_1939);
or U2130 (N_2130,N_1540,N_1759);
and U2131 (N_2131,N_1612,N_1771);
nand U2132 (N_2132,N_1768,N_1639);
and U2133 (N_2133,N_1728,N_1798);
xor U2134 (N_2134,N_1886,N_1686);
xor U2135 (N_2135,N_1957,N_1741);
xor U2136 (N_2136,N_1952,N_1979);
nor U2137 (N_2137,N_1841,N_1938);
and U2138 (N_2138,N_1760,N_1709);
nand U2139 (N_2139,N_1529,N_1599);
or U2140 (N_2140,N_1673,N_1541);
and U2141 (N_2141,N_1522,N_1694);
or U2142 (N_2142,N_1800,N_1737);
xnor U2143 (N_2143,N_1627,N_1843);
xor U2144 (N_2144,N_1640,N_1579);
xnor U2145 (N_2145,N_1565,N_1880);
or U2146 (N_2146,N_1661,N_1527);
xor U2147 (N_2147,N_1727,N_1812);
or U2148 (N_2148,N_1912,N_1613);
and U2149 (N_2149,N_1603,N_1908);
and U2150 (N_2150,N_1968,N_1859);
xnor U2151 (N_2151,N_1511,N_1987);
and U2152 (N_2152,N_1707,N_1902);
or U2153 (N_2153,N_1742,N_1675);
nand U2154 (N_2154,N_1632,N_1836);
or U2155 (N_2155,N_1539,N_1714);
nand U2156 (N_2156,N_1504,N_1589);
xnor U2157 (N_2157,N_1887,N_1916);
and U2158 (N_2158,N_1597,N_1925);
or U2159 (N_2159,N_1962,N_1693);
nor U2160 (N_2160,N_1538,N_1611);
xnor U2161 (N_2161,N_1689,N_1965);
nand U2162 (N_2162,N_1879,N_1900);
nor U2163 (N_2163,N_1513,N_1723);
and U2164 (N_2164,N_1762,N_1649);
xor U2165 (N_2165,N_1960,N_1845);
and U2166 (N_2166,N_1557,N_1666);
nand U2167 (N_2167,N_1566,N_1732);
or U2168 (N_2168,N_1739,N_1718);
and U2169 (N_2169,N_1830,N_1634);
xor U2170 (N_2170,N_1662,N_1610);
nor U2171 (N_2171,N_1838,N_1677);
xnor U2172 (N_2172,N_1855,N_1708);
and U2173 (N_2173,N_1816,N_1593);
nand U2174 (N_2174,N_1545,N_1598);
nand U2175 (N_2175,N_1970,N_1600);
xor U2176 (N_2176,N_1999,N_1674);
nand U2177 (N_2177,N_1914,N_1641);
xnor U2178 (N_2178,N_1553,N_1716);
xnor U2179 (N_2179,N_1650,N_1867);
xor U2180 (N_2180,N_1803,N_1616);
nor U2181 (N_2181,N_1875,N_1591);
xnor U2182 (N_2182,N_1510,N_1978);
and U2183 (N_2183,N_1651,N_1628);
or U2184 (N_2184,N_1555,N_1526);
or U2185 (N_2185,N_1917,N_1584);
nand U2186 (N_2186,N_1889,N_1517);
nor U2187 (N_2187,N_1752,N_1745);
nor U2188 (N_2188,N_1590,N_1617);
nor U2189 (N_2189,N_1625,N_1692);
and U2190 (N_2190,N_1789,N_1834);
nor U2191 (N_2191,N_1781,N_1588);
xnor U2192 (N_2192,N_1554,N_1531);
or U2193 (N_2193,N_1931,N_1868);
nand U2194 (N_2194,N_1509,N_1697);
and U2195 (N_2195,N_1626,N_1821);
and U2196 (N_2196,N_1505,N_1842);
xnor U2197 (N_2197,N_1790,N_1884);
and U2198 (N_2198,N_1837,N_1542);
nand U2199 (N_2199,N_1551,N_1779);
or U2200 (N_2200,N_1736,N_1519);
xor U2201 (N_2201,N_1930,N_1550);
xor U2202 (N_2202,N_1795,N_1986);
or U2203 (N_2203,N_1892,N_1955);
xnor U2204 (N_2204,N_1571,N_1814);
and U2205 (N_2205,N_1846,N_1601);
nand U2206 (N_2206,N_1715,N_1655);
or U2207 (N_2207,N_1997,N_1722);
nor U2208 (N_2208,N_1679,N_1512);
or U2209 (N_2209,N_1772,N_1918);
nor U2210 (N_2210,N_1915,N_1937);
nor U2211 (N_2211,N_1828,N_1964);
xor U2212 (N_2212,N_1712,N_1748);
and U2213 (N_2213,N_1711,N_1770);
or U2214 (N_2214,N_1623,N_1619);
xnor U2215 (N_2215,N_1524,N_1516);
and U2216 (N_2216,N_1766,N_1893);
or U2217 (N_2217,N_1532,N_1729);
nand U2218 (N_2218,N_1794,N_1763);
or U2219 (N_2219,N_1706,N_1726);
and U2220 (N_2220,N_1756,N_1890);
or U2221 (N_2221,N_1585,N_1881);
nor U2222 (N_2222,N_1898,N_1863);
nor U2223 (N_2223,N_1635,N_1767);
nor U2224 (N_2224,N_1503,N_1911);
nand U2225 (N_2225,N_1847,N_1967);
and U2226 (N_2226,N_1620,N_1852);
and U2227 (N_2227,N_1820,N_1801);
xor U2228 (N_2228,N_1733,N_1700);
xnor U2229 (N_2229,N_1559,N_1793);
or U2230 (N_2230,N_1792,N_1805);
nand U2231 (N_2231,N_1959,N_1956);
and U2232 (N_2232,N_1777,N_1983);
nor U2233 (N_2233,N_1667,N_1631);
or U2234 (N_2234,N_1669,N_1701);
and U2235 (N_2235,N_1932,N_1764);
xnor U2236 (N_2236,N_1602,N_1665);
nor U2237 (N_2237,N_1570,N_1769);
or U2238 (N_2238,N_1743,N_1577);
nand U2239 (N_2239,N_1705,N_1993);
nand U2240 (N_2240,N_1607,N_1755);
xor U2241 (N_2241,N_1856,N_1882);
and U2242 (N_2242,N_1782,N_1835);
or U2243 (N_2243,N_1971,N_1791);
nor U2244 (N_2244,N_1528,N_1972);
nor U2245 (N_2245,N_1785,N_1746);
nand U2246 (N_2246,N_1622,N_1608);
or U2247 (N_2247,N_1933,N_1773);
or U2248 (N_2248,N_1658,N_1823);
and U2249 (N_2249,N_1682,N_1929);
or U2250 (N_2250,N_1557,N_1982);
or U2251 (N_2251,N_1735,N_1717);
or U2252 (N_2252,N_1795,N_1728);
xor U2253 (N_2253,N_1781,N_1976);
and U2254 (N_2254,N_1906,N_1694);
nor U2255 (N_2255,N_1532,N_1989);
or U2256 (N_2256,N_1728,N_1700);
xnor U2257 (N_2257,N_1537,N_1786);
or U2258 (N_2258,N_1725,N_1995);
xor U2259 (N_2259,N_1534,N_1972);
or U2260 (N_2260,N_1884,N_1795);
xnor U2261 (N_2261,N_1720,N_1949);
or U2262 (N_2262,N_1504,N_1888);
xor U2263 (N_2263,N_1732,N_1636);
and U2264 (N_2264,N_1947,N_1740);
nand U2265 (N_2265,N_1923,N_1926);
and U2266 (N_2266,N_1622,N_1559);
xor U2267 (N_2267,N_1636,N_1775);
nor U2268 (N_2268,N_1931,N_1772);
or U2269 (N_2269,N_1862,N_1651);
or U2270 (N_2270,N_1924,N_1595);
nand U2271 (N_2271,N_1929,N_1543);
nand U2272 (N_2272,N_1908,N_1571);
nand U2273 (N_2273,N_1517,N_1702);
and U2274 (N_2274,N_1688,N_1825);
xnor U2275 (N_2275,N_1635,N_1905);
nor U2276 (N_2276,N_1852,N_1890);
nand U2277 (N_2277,N_1945,N_1571);
and U2278 (N_2278,N_1950,N_1526);
nand U2279 (N_2279,N_1919,N_1910);
nor U2280 (N_2280,N_1565,N_1769);
xnor U2281 (N_2281,N_1622,N_1609);
nand U2282 (N_2282,N_1833,N_1666);
nand U2283 (N_2283,N_1675,N_1711);
xnor U2284 (N_2284,N_1870,N_1814);
nor U2285 (N_2285,N_1771,N_1955);
nor U2286 (N_2286,N_1552,N_1921);
or U2287 (N_2287,N_1564,N_1891);
xor U2288 (N_2288,N_1622,N_1872);
nor U2289 (N_2289,N_1972,N_1992);
nand U2290 (N_2290,N_1961,N_1561);
and U2291 (N_2291,N_1676,N_1820);
and U2292 (N_2292,N_1886,N_1623);
nand U2293 (N_2293,N_1802,N_1996);
or U2294 (N_2294,N_1956,N_1603);
or U2295 (N_2295,N_1769,N_1991);
or U2296 (N_2296,N_1576,N_1835);
or U2297 (N_2297,N_1625,N_1590);
nor U2298 (N_2298,N_1520,N_1988);
and U2299 (N_2299,N_1715,N_1775);
xor U2300 (N_2300,N_1819,N_1889);
nand U2301 (N_2301,N_1802,N_1742);
nor U2302 (N_2302,N_1727,N_1663);
xnor U2303 (N_2303,N_1921,N_1771);
nor U2304 (N_2304,N_1557,N_1967);
xnor U2305 (N_2305,N_1503,N_1770);
and U2306 (N_2306,N_1716,N_1570);
xor U2307 (N_2307,N_1657,N_1646);
and U2308 (N_2308,N_1919,N_1885);
xor U2309 (N_2309,N_1557,N_1618);
and U2310 (N_2310,N_1820,N_1946);
and U2311 (N_2311,N_1530,N_1674);
or U2312 (N_2312,N_1996,N_1774);
and U2313 (N_2313,N_1834,N_1666);
xor U2314 (N_2314,N_1589,N_1727);
and U2315 (N_2315,N_1503,N_1861);
nand U2316 (N_2316,N_1752,N_1715);
nor U2317 (N_2317,N_1571,N_1610);
or U2318 (N_2318,N_1993,N_1697);
nand U2319 (N_2319,N_1728,N_1725);
nor U2320 (N_2320,N_1610,N_1665);
nor U2321 (N_2321,N_1746,N_1735);
or U2322 (N_2322,N_1549,N_1985);
nand U2323 (N_2323,N_1963,N_1917);
nor U2324 (N_2324,N_1510,N_1740);
and U2325 (N_2325,N_1792,N_1670);
nand U2326 (N_2326,N_1639,N_1523);
and U2327 (N_2327,N_1817,N_1972);
xor U2328 (N_2328,N_1817,N_1937);
nor U2329 (N_2329,N_1926,N_1833);
or U2330 (N_2330,N_1528,N_1760);
or U2331 (N_2331,N_1759,N_1531);
or U2332 (N_2332,N_1870,N_1546);
xnor U2333 (N_2333,N_1763,N_1882);
nor U2334 (N_2334,N_1929,N_1828);
nand U2335 (N_2335,N_1906,N_1679);
and U2336 (N_2336,N_1975,N_1905);
nor U2337 (N_2337,N_1687,N_1929);
nor U2338 (N_2338,N_1740,N_1691);
xnor U2339 (N_2339,N_1752,N_1524);
xor U2340 (N_2340,N_1756,N_1564);
or U2341 (N_2341,N_1862,N_1903);
xnor U2342 (N_2342,N_1670,N_1883);
and U2343 (N_2343,N_1824,N_1929);
xnor U2344 (N_2344,N_1888,N_1883);
nand U2345 (N_2345,N_1656,N_1916);
nor U2346 (N_2346,N_1597,N_1592);
and U2347 (N_2347,N_1526,N_1995);
or U2348 (N_2348,N_1869,N_1786);
xor U2349 (N_2349,N_1693,N_1745);
and U2350 (N_2350,N_1544,N_1908);
and U2351 (N_2351,N_1522,N_1887);
xnor U2352 (N_2352,N_1718,N_1727);
nand U2353 (N_2353,N_1798,N_1625);
or U2354 (N_2354,N_1924,N_1625);
or U2355 (N_2355,N_1914,N_1609);
and U2356 (N_2356,N_1678,N_1526);
and U2357 (N_2357,N_1945,N_1740);
or U2358 (N_2358,N_1505,N_1726);
and U2359 (N_2359,N_1587,N_1750);
xor U2360 (N_2360,N_1586,N_1802);
nor U2361 (N_2361,N_1738,N_1653);
or U2362 (N_2362,N_1671,N_1524);
nand U2363 (N_2363,N_1924,N_1665);
xor U2364 (N_2364,N_1580,N_1508);
or U2365 (N_2365,N_1792,N_1862);
nor U2366 (N_2366,N_1618,N_1525);
xnor U2367 (N_2367,N_1567,N_1798);
or U2368 (N_2368,N_1568,N_1976);
xnor U2369 (N_2369,N_1556,N_1574);
nand U2370 (N_2370,N_1542,N_1602);
nor U2371 (N_2371,N_1820,N_1613);
nor U2372 (N_2372,N_1628,N_1904);
nor U2373 (N_2373,N_1861,N_1696);
nor U2374 (N_2374,N_1698,N_1515);
or U2375 (N_2375,N_1713,N_1633);
and U2376 (N_2376,N_1822,N_1791);
nand U2377 (N_2377,N_1532,N_1543);
nor U2378 (N_2378,N_1522,N_1686);
xor U2379 (N_2379,N_1953,N_1576);
nor U2380 (N_2380,N_1869,N_1920);
nand U2381 (N_2381,N_1856,N_1906);
and U2382 (N_2382,N_1565,N_1698);
xnor U2383 (N_2383,N_1673,N_1942);
nand U2384 (N_2384,N_1581,N_1685);
xnor U2385 (N_2385,N_1611,N_1840);
or U2386 (N_2386,N_1602,N_1897);
and U2387 (N_2387,N_1828,N_1819);
and U2388 (N_2388,N_1734,N_1925);
nand U2389 (N_2389,N_1620,N_1923);
and U2390 (N_2390,N_1646,N_1613);
nor U2391 (N_2391,N_1825,N_1647);
and U2392 (N_2392,N_1601,N_1514);
nand U2393 (N_2393,N_1844,N_1614);
or U2394 (N_2394,N_1847,N_1687);
nand U2395 (N_2395,N_1616,N_1838);
or U2396 (N_2396,N_1943,N_1965);
nand U2397 (N_2397,N_1948,N_1720);
or U2398 (N_2398,N_1776,N_1646);
xnor U2399 (N_2399,N_1623,N_1545);
or U2400 (N_2400,N_1959,N_1954);
or U2401 (N_2401,N_1918,N_1514);
nand U2402 (N_2402,N_1582,N_1931);
nand U2403 (N_2403,N_1650,N_1830);
and U2404 (N_2404,N_1957,N_1746);
and U2405 (N_2405,N_1836,N_1768);
or U2406 (N_2406,N_1769,N_1505);
xnor U2407 (N_2407,N_1979,N_1942);
nand U2408 (N_2408,N_1644,N_1847);
and U2409 (N_2409,N_1732,N_1609);
and U2410 (N_2410,N_1802,N_1771);
and U2411 (N_2411,N_1657,N_1644);
xnor U2412 (N_2412,N_1727,N_1538);
nand U2413 (N_2413,N_1780,N_1818);
or U2414 (N_2414,N_1905,N_1503);
xnor U2415 (N_2415,N_1700,N_1874);
nand U2416 (N_2416,N_1548,N_1970);
nor U2417 (N_2417,N_1673,N_1856);
and U2418 (N_2418,N_1763,N_1711);
or U2419 (N_2419,N_1526,N_1994);
nor U2420 (N_2420,N_1505,N_1745);
nor U2421 (N_2421,N_1940,N_1963);
nor U2422 (N_2422,N_1771,N_1625);
and U2423 (N_2423,N_1928,N_1755);
or U2424 (N_2424,N_1935,N_1502);
nor U2425 (N_2425,N_1997,N_1528);
nor U2426 (N_2426,N_1767,N_1569);
nor U2427 (N_2427,N_1905,N_1805);
and U2428 (N_2428,N_1506,N_1822);
xnor U2429 (N_2429,N_1792,N_1706);
and U2430 (N_2430,N_1741,N_1981);
and U2431 (N_2431,N_1597,N_1559);
xnor U2432 (N_2432,N_1846,N_1565);
xor U2433 (N_2433,N_1986,N_1571);
nor U2434 (N_2434,N_1824,N_1572);
nor U2435 (N_2435,N_1950,N_1934);
and U2436 (N_2436,N_1530,N_1507);
nor U2437 (N_2437,N_1807,N_1705);
nand U2438 (N_2438,N_1503,N_1668);
xor U2439 (N_2439,N_1874,N_1595);
nand U2440 (N_2440,N_1851,N_1570);
nor U2441 (N_2441,N_1745,N_1860);
and U2442 (N_2442,N_1502,N_1869);
or U2443 (N_2443,N_1616,N_1973);
nand U2444 (N_2444,N_1848,N_1670);
nand U2445 (N_2445,N_1518,N_1769);
or U2446 (N_2446,N_1908,N_1657);
or U2447 (N_2447,N_1901,N_1755);
nand U2448 (N_2448,N_1777,N_1959);
nor U2449 (N_2449,N_1878,N_1591);
nand U2450 (N_2450,N_1749,N_1823);
nor U2451 (N_2451,N_1742,N_1520);
xnor U2452 (N_2452,N_1610,N_1946);
or U2453 (N_2453,N_1790,N_1829);
xor U2454 (N_2454,N_1863,N_1511);
or U2455 (N_2455,N_1702,N_1726);
and U2456 (N_2456,N_1527,N_1755);
nand U2457 (N_2457,N_1755,N_1764);
nand U2458 (N_2458,N_1818,N_1749);
xor U2459 (N_2459,N_1916,N_1965);
and U2460 (N_2460,N_1758,N_1595);
and U2461 (N_2461,N_1648,N_1661);
or U2462 (N_2462,N_1505,N_1928);
nand U2463 (N_2463,N_1945,N_1845);
or U2464 (N_2464,N_1967,N_1983);
xnor U2465 (N_2465,N_1895,N_1590);
nand U2466 (N_2466,N_1735,N_1679);
or U2467 (N_2467,N_1876,N_1536);
nor U2468 (N_2468,N_1960,N_1627);
nand U2469 (N_2469,N_1925,N_1554);
xor U2470 (N_2470,N_1637,N_1774);
or U2471 (N_2471,N_1657,N_1863);
xor U2472 (N_2472,N_1878,N_1999);
and U2473 (N_2473,N_1776,N_1888);
xor U2474 (N_2474,N_1754,N_1566);
and U2475 (N_2475,N_1960,N_1800);
xor U2476 (N_2476,N_1849,N_1646);
or U2477 (N_2477,N_1650,N_1737);
xnor U2478 (N_2478,N_1526,N_1690);
and U2479 (N_2479,N_1842,N_1575);
nor U2480 (N_2480,N_1713,N_1617);
or U2481 (N_2481,N_1841,N_1859);
nor U2482 (N_2482,N_1622,N_1867);
nand U2483 (N_2483,N_1650,N_1756);
nand U2484 (N_2484,N_1901,N_1571);
or U2485 (N_2485,N_1729,N_1630);
nand U2486 (N_2486,N_1917,N_1707);
nor U2487 (N_2487,N_1628,N_1798);
xor U2488 (N_2488,N_1730,N_1761);
xor U2489 (N_2489,N_1979,N_1865);
and U2490 (N_2490,N_1535,N_1762);
nor U2491 (N_2491,N_1992,N_1593);
or U2492 (N_2492,N_1980,N_1921);
nand U2493 (N_2493,N_1801,N_1947);
nor U2494 (N_2494,N_1617,N_1647);
and U2495 (N_2495,N_1814,N_1885);
nor U2496 (N_2496,N_1839,N_1561);
nor U2497 (N_2497,N_1510,N_1901);
xnor U2498 (N_2498,N_1549,N_1723);
xnor U2499 (N_2499,N_1935,N_1870);
and U2500 (N_2500,N_2189,N_2176);
and U2501 (N_2501,N_2033,N_2077);
nor U2502 (N_2502,N_2392,N_2095);
and U2503 (N_2503,N_2246,N_2313);
and U2504 (N_2504,N_2334,N_2405);
nand U2505 (N_2505,N_2396,N_2276);
nand U2506 (N_2506,N_2388,N_2387);
nor U2507 (N_2507,N_2252,N_2475);
and U2508 (N_2508,N_2328,N_2379);
and U2509 (N_2509,N_2274,N_2347);
xor U2510 (N_2510,N_2046,N_2195);
xnor U2511 (N_2511,N_2020,N_2182);
and U2512 (N_2512,N_2462,N_2266);
nor U2513 (N_2513,N_2237,N_2308);
or U2514 (N_2514,N_2065,N_2275);
nand U2515 (N_2515,N_2269,N_2148);
or U2516 (N_2516,N_2364,N_2226);
nor U2517 (N_2517,N_2497,N_2283);
and U2518 (N_2518,N_2419,N_2193);
or U2519 (N_2519,N_2224,N_2023);
nor U2520 (N_2520,N_2430,N_2265);
nor U2521 (N_2521,N_2410,N_2267);
nor U2522 (N_2522,N_2382,N_2102);
or U2523 (N_2523,N_2288,N_2422);
or U2524 (N_2524,N_2116,N_2407);
xor U2525 (N_2525,N_2397,N_2244);
and U2526 (N_2526,N_2446,N_2476);
nand U2527 (N_2527,N_2017,N_2317);
nor U2528 (N_2528,N_2425,N_2311);
nand U2529 (N_2529,N_2389,N_2473);
nor U2530 (N_2530,N_2232,N_2022);
and U2531 (N_2531,N_2486,N_2030);
nor U2532 (N_2532,N_2336,N_2432);
nand U2533 (N_2533,N_2147,N_2408);
xor U2534 (N_2534,N_2211,N_2270);
or U2535 (N_2535,N_2309,N_2412);
nor U2536 (N_2536,N_2135,N_2113);
and U2537 (N_2537,N_2036,N_2279);
xnor U2538 (N_2538,N_2361,N_2190);
and U2539 (N_2539,N_2345,N_2078);
or U2540 (N_2540,N_2039,N_2084);
nor U2541 (N_2541,N_2414,N_2088);
and U2542 (N_2542,N_2171,N_2447);
nor U2543 (N_2543,N_2292,N_2149);
xor U2544 (N_2544,N_2472,N_2185);
nand U2545 (N_2545,N_2324,N_2172);
xnor U2546 (N_2546,N_2398,N_2263);
or U2547 (N_2547,N_2483,N_2250);
or U2548 (N_2548,N_2289,N_2253);
nand U2549 (N_2549,N_2162,N_2247);
xor U2550 (N_2550,N_2134,N_2010);
or U2551 (N_2551,N_2071,N_2384);
nand U2552 (N_2552,N_2255,N_2471);
xnor U2553 (N_2553,N_2329,N_2212);
nor U2554 (N_2554,N_2107,N_2136);
nor U2555 (N_2555,N_2173,N_2346);
nand U2556 (N_2556,N_2340,N_2249);
nor U2557 (N_2557,N_2261,N_2111);
and U2558 (N_2558,N_2035,N_2458);
nor U2559 (N_2559,N_2062,N_2126);
or U2560 (N_2560,N_2366,N_2118);
nor U2561 (N_2561,N_2478,N_2394);
nor U2562 (N_2562,N_2153,N_2316);
nor U2563 (N_2563,N_2197,N_2395);
xor U2564 (N_2564,N_2174,N_2186);
and U2565 (N_2565,N_2068,N_2214);
nor U2566 (N_2566,N_2191,N_2012);
nor U2567 (N_2567,N_2409,N_2470);
and U2568 (N_2568,N_2386,N_2103);
nand U2569 (N_2569,N_2051,N_2303);
nand U2570 (N_2570,N_2202,N_2356);
xnor U2571 (N_2571,N_2128,N_2150);
or U2572 (N_2572,N_2312,N_2335);
or U2573 (N_2573,N_2056,N_2435);
xor U2574 (N_2574,N_2459,N_2119);
nand U2575 (N_2575,N_2307,N_2005);
nand U2576 (N_2576,N_2027,N_2445);
nor U2577 (N_2577,N_2254,N_2096);
or U2578 (N_2578,N_2058,N_2029);
xnor U2579 (N_2579,N_2165,N_2091);
or U2580 (N_2580,N_2122,N_2243);
nand U2581 (N_2581,N_2444,N_2025);
nand U2582 (N_2582,N_2110,N_2404);
xor U2583 (N_2583,N_2218,N_2198);
or U2584 (N_2584,N_2482,N_2293);
xor U2585 (N_2585,N_2146,N_2429);
nand U2586 (N_2586,N_2496,N_2424);
nand U2587 (N_2587,N_2448,N_2437);
nor U2588 (N_2588,N_2141,N_2373);
nand U2589 (N_2589,N_2491,N_2268);
and U2590 (N_2590,N_2325,N_2323);
or U2591 (N_2591,N_2367,N_2431);
nor U2592 (N_2592,N_2443,N_2248);
or U2593 (N_2593,N_2044,N_2264);
or U2594 (N_2594,N_2152,N_2402);
nor U2595 (N_2595,N_2348,N_2009);
nand U2596 (N_2596,N_2239,N_2390);
nor U2597 (N_2597,N_2105,N_2442);
xor U2598 (N_2598,N_2280,N_2489);
nand U2599 (N_2599,N_2210,N_2131);
nand U2600 (N_2600,N_2179,N_2238);
xor U2601 (N_2601,N_2042,N_2187);
xor U2602 (N_2602,N_2015,N_2217);
and U2603 (N_2603,N_2460,N_2495);
nand U2604 (N_2604,N_2188,N_2413);
nand U2605 (N_2605,N_2433,N_2351);
nand U2606 (N_2606,N_2260,N_2163);
and U2607 (N_2607,N_2003,N_2045);
nor U2608 (N_2608,N_2100,N_2485);
nor U2609 (N_2609,N_2206,N_2002);
nand U2610 (N_2610,N_2109,N_2256);
nor U2611 (N_2611,N_2011,N_2161);
or U2612 (N_2612,N_2441,N_2330);
xnor U2613 (N_2613,N_2204,N_2338);
and U2614 (N_2614,N_2021,N_2434);
or U2615 (N_2615,N_2142,N_2037);
nor U2616 (N_2616,N_2097,N_2298);
or U2617 (N_2617,N_2112,N_2220);
nor U2618 (N_2618,N_2456,N_2064);
and U2619 (N_2619,N_2257,N_2377);
nand U2620 (N_2620,N_2342,N_2498);
xnor U2621 (N_2621,N_2028,N_2259);
or U2622 (N_2622,N_2332,N_2032);
nand U2623 (N_2623,N_2201,N_2438);
and U2624 (N_2624,N_2199,N_2406);
xnor U2625 (N_2625,N_2296,N_2349);
nand U2626 (N_2626,N_2016,N_2468);
xor U2627 (N_2627,N_2284,N_2074);
and U2628 (N_2628,N_2183,N_2385);
nand U2629 (N_2629,N_2104,N_2125);
xor U2630 (N_2630,N_2075,N_2258);
xnor U2631 (N_2631,N_2216,N_2082);
and U2632 (N_2632,N_2467,N_2184);
xnor U2633 (N_2633,N_2219,N_2295);
nor U2634 (N_2634,N_2391,N_2155);
nor U2635 (N_2635,N_2207,N_2175);
or U2636 (N_2636,N_2166,N_2234);
or U2637 (N_2637,N_2227,N_2272);
xor U2638 (N_2638,N_2205,N_2494);
and U2639 (N_2639,N_2178,N_2233);
or U2640 (N_2640,N_2378,N_2203);
nand U2641 (N_2641,N_2297,N_2115);
xor U2642 (N_2642,N_2499,N_2094);
or U2643 (N_2643,N_2208,N_2121);
nand U2644 (N_2644,N_2123,N_2314);
xor U2645 (N_2645,N_2360,N_2354);
xor U2646 (N_2646,N_2477,N_2092);
or U2647 (N_2647,N_2060,N_2466);
and U2648 (N_2648,N_2426,N_2241);
or U2649 (N_2649,N_2215,N_2014);
or U2650 (N_2650,N_2371,N_2355);
nor U2651 (N_2651,N_2133,N_2120);
nand U2652 (N_2652,N_2353,N_2421);
or U2653 (N_2653,N_2273,N_2070);
nor U2654 (N_2654,N_2304,N_2352);
or U2655 (N_2655,N_2453,N_2140);
xnor U2656 (N_2656,N_2080,N_2240);
and U2657 (N_2657,N_2159,N_2306);
nand U2658 (N_2658,N_2436,N_2229);
xor U2659 (N_2659,N_2449,N_2180);
and U2660 (N_2660,N_2200,N_2461);
or U2661 (N_2661,N_2090,N_2374);
or U2662 (N_2662,N_2076,N_2117);
nand U2663 (N_2663,N_2222,N_2282);
nand U2664 (N_2664,N_2331,N_2411);
and U2665 (N_2665,N_2287,N_2363);
nor U2666 (N_2666,N_2209,N_2400);
or U2667 (N_2667,N_2291,N_2235);
xor U2668 (N_2668,N_2018,N_2488);
xor U2669 (N_2669,N_2106,N_2196);
nand U2670 (N_2670,N_2481,N_2061);
or U2671 (N_2671,N_2393,N_2008);
nor U2672 (N_2672,N_2359,N_2031);
and U2673 (N_2673,N_2127,N_2479);
or U2674 (N_2674,N_2415,N_2170);
xnor U2675 (N_2675,N_2108,N_2278);
nor U2676 (N_2676,N_2365,N_2139);
and U2677 (N_2677,N_2048,N_2164);
nand U2678 (N_2678,N_2177,N_2114);
and U2679 (N_2679,N_2333,N_2320);
xor U2680 (N_2680,N_2132,N_2375);
xnor U2681 (N_2681,N_2271,N_2228);
and U2682 (N_2682,N_2000,N_2192);
or U2683 (N_2683,N_2019,N_2047);
nor U2684 (N_2684,N_2428,N_2305);
nand U2685 (N_2685,N_2236,N_2053);
and U2686 (N_2686,N_2151,N_2381);
xor U2687 (N_2687,N_2055,N_2357);
nand U2688 (N_2688,N_2450,N_2144);
xnor U2689 (N_2689,N_2299,N_2006);
xor U2690 (N_2690,N_2083,N_2137);
nand U2691 (N_2691,N_2160,N_2423);
and U2692 (N_2692,N_2079,N_2368);
xor U2693 (N_2693,N_2073,N_2358);
and U2694 (N_2694,N_2063,N_2242);
nand U2695 (N_2695,N_2225,N_2052);
or U2696 (N_2696,N_2085,N_2337);
and U2697 (N_2697,N_2343,N_2167);
nand U2698 (N_2698,N_2315,N_2420);
or U2699 (N_2699,N_2465,N_2427);
xnor U2700 (N_2700,N_2154,N_2300);
nor U2701 (N_2701,N_2157,N_2451);
nand U2702 (N_2702,N_2286,N_2034);
nor U2703 (N_2703,N_2416,N_2493);
or U2704 (N_2704,N_2138,N_2327);
nor U2705 (N_2705,N_2004,N_2081);
nor U2706 (N_2706,N_2490,N_2454);
or U2707 (N_2707,N_2245,N_2455);
nor U2708 (N_2708,N_2087,N_2321);
nand U2709 (N_2709,N_2318,N_2362);
xnor U2710 (N_2710,N_2066,N_2440);
nand U2711 (N_2711,N_2294,N_2285);
nand U2712 (N_2712,N_2302,N_2370);
or U2713 (N_2713,N_2310,N_2043);
or U2714 (N_2714,N_2290,N_2399);
xnor U2715 (N_2715,N_2403,N_2376);
and U2716 (N_2716,N_2024,N_2181);
xnor U2717 (N_2717,N_2007,N_2072);
or U2718 (N_2718,N_2452,N_2099);
nand U2719 (N_2719,N_2372,N_2339);
and U2720 (N_2720,N_2383,N_2326);
and U2721 (N_2721,N_2143,N_2098);
or U2722 (N_2722,N_2487,N_2059);
and U2723 (N_2723,N_2168,N_2341);
and U2724 (N_2724,N_2380,N_2277);
or U2725 (N_2725,N_2484,N_2464);
and U2726 (N_2726,N_2457,N_2093);
nor U2727 (N_2727,N_2057,N_2319);
nand U2728 (N_2728,N_2350,N_2281);
xor U2729 (N_2729,N_2089,N_2145);
or U2730 (N_2730,N_2169,N_2469);
or U2731 (N_2731,N_2041,N_2417);
or U2732 (N_2732,N_2001,N_2344);
nand U2733 (N_2733,N_2401,N_2054);
and U2734 (N_2734,N_2069,N_2040);
xnor U2735 (N_2735,N_2086,N_2101);
or U2736 (N_2736,N_2230,N_2463);
nand U2737 (N_2737,N_2262,N_2480);
or U2738 (N_2738,N_2213,N_2050);
nand U2739 (N_2739,N_2221,N_2223);
and U2740 (N_2740,N_2251,N_2049);
or U2741 (N_2741,N_2418,N_2439);
nand U2742 (N_2742,N_2492,N_2129);
and U2743 (N_2743,N_2231,N_2038);
nand U2744 (N_2744,N_2322,N_2474);
and U2745 (N_2745,N_2013,N_2067);
or U2746 (N_2746,N_2124,N_2156);
nor U2747 (N_2747,N_2301,N_2130);
xnor U2748 (N_2748,N_2158,N_2194);
and U2749 (N_2749,N_2369,N_2026);
nand U2750 (N_2750,N_2414,N_2163);
or U2751 (N_2751,N_2397,N_2259);
xor U2752 (N_2752,N_2202,N_2187);
nor U2753 (N_2753,N_2149,N_2117);
xor U2754 (N_2754,N_2171,N_2358);
nor U2755 (N_2755,N_2211,N_2284);
or U2756 (N_2756,N_2310,N_2164);
nand U2757 (N_2757,N_2037,N_2309);
nand U2758 (N_2758,N_2318,N_2286);
xor U2759 (N_2759,N_2298,N_2360);
and U2760 (N_2760,N_2024,N_2201);
nor U2761 (N_2761,N_2301,N_2132);
nor U2762 (N_2762,N_2464,N_2431);
nor U2763 (N_2763,N_2296,N_2164);
nor U2764 (N_2764,N_2051,N_2156);
xor U2765 (N_2765,N_2280,N_2241);
nand U2766 (N_2766,N_2143,N_2246);
xor U2767 (N_2767,N_2356,N_2116);
xnor U2768 (N_2768,N_2052,N_2236);
nor U2769 (N_2769,N_2102,N_2030);
nor U2770 (N_2770,N_2122,N_2042);
or U2771 (N_2771,N_2355,N_2219);
nor U2772 (N_2772,N_2492,N_2458);
xnor U2773 (N_2773,N_2139,N_2354);
nor U2774 (N_2774,N_2151,N_2410);
nor U2775 (N_2775,N_2427,N_2030);
and U2776 (N_2776,N_2320,N_2270);
or U2777 (N_2777,N_2489,N_2296);
and U2778 (N_2778,N_2450,N_2222);
nor U2779 (N_2779,N_2436,N_2284);
xor U2780 (N_2780,N_2081,N_2043);
and U2781 (N_2781,N_2036,N_2208);
xnor U2782 (N_2782,N_2478,N_2437);
or U2783 (N_2783,N_2220,N_2001);
nor U2784 (N_2784,N_2481,N_2086);
nand U2785 (N_2785,N_2153,N_2369);
or U2786 (N_2786,N_2339,N_2122);
and U2787 (N_2787,N_2350,N_2062);
and U2788 (N_2788,N_2287,N_2219);
nand U2789 (N_2789,N_2236,N_2084);
nor U2790 (N_2790,N_2052,N_2263);
nand U2791 (N_2791,N_2212,N_2372);
and U2792 (N_2792,N_2284,N_2137);
and U2793 (N_2793,N_2002,N_2014);
nor U2794 (N_2794,N_2179,N_2389);
and U2795 (N_2795,N_2487,N_2190);
nand U2796 (N_2796,N_2150,N_2491);
nor U2797 (N_2797,N_2432,N_2040);
nand U2798 (N_2798,N_2057,N_2183);
and U2799 (N_2799,N_2132,N_2250);
nand U2800 (N_2800,N_2014,N_2416);
nor U2801 (N_2801,N_2289,N_2433);
or U2802 (N_2802,N_2206,N_2068);
nand U2803 (N_2803,N_2243,N_2489);
xor U2804 (N_2804,N_2253,N_2318);
and U2805 (N_2805,N_2328,N_2068);
xnor U2806 (N_2806,N_2014,N_2205);
nand U2807 (N_2807,N_2494,N_2001);
nor U2808 (N_2808,N_2012,N_2415);
nor U2809 (N_2809,N_2434,N_2152);
xor U2810 (N_2810,N_2102,N_2338);
nor U2811 (N_2811,N_2109,N_2487);
xnor U2812 (N_2812,N_2389,N_2400);
or U2813 (N_2813,N_2491,N_2450);
nor U2814 (N_2814,N_2060,N_2091);
nor U2815 (N_2815,N_2086,N_2424);
nand U2816 (N_2816,N_2316,N_2134);
nand U2817 (N_2817,N_2379,N_2101);
or U2818 (N_2818,N_2064,N_2421);
and U2819 (N_2819,N_2103,N_2450);
or U2820 (N_2820,N_2382,N_2052);
nand U2821 (N_2821,N_2027,N_2463);
nor U2822 (N_2822,N_2356,N_2255);
nor U2823 (N_2823,N_2448,N_2310);
or U2824 (N_2824,N_2304,N_2137);
and U2825 (N_2825,N_2213,N_2080);
or U2826 (N_2826,N_2446,N_2218);
or U2827 (N_2827,N_2359,N_2245);
nor U2828 (N_2828,N_2081,N_2179);
nor U2829 (N_2829,N_2203,N_2181);
nand U2830 (N_2830,N_2320,N_2454);
or U2831 (N_2831,N_2095,N_2045);
nor U2832 (N_2832,N_2017,N_2473);
xnor U2833 (N_2833,N_2129,N_2237);
nor U2834 (N_2834,N_2362,N_2240);
and U2835 (N_2835,N_2162,N_2259);
nor U2836 (N_2836,N_2094,N_2352);
nor U2837 (N_2837,N_2038,N_2077);
xnor U2838 (N_2838,N_2222,N_2241);
and U2839 (N_2839,N_2150,N_2088);
nand U2840 (N_2840,N_2259,N_2413);
and U2841 (N_2841,N_2113,N_2291);
and U2842 (N_2842,N_2147,N_2144);
or U2843 (N_2843,N_2438,N_2312);
and U2844 (N_2844,N_2460,N_2262);
or U2845 (N_2845,N_2019,N_2245);
or U2846 (N_2846,N_2078,N_2020);
or U2847 (N_2847,N_2390,N_2479);
nor U2848 (N_2848,N_2447,N_2301);
xnor U2849 (N_2849,N_2091,N_2451);
nand U2850 (N_2850,N_2144,N_2384);
and U2851 (N_2851,N_2164,N_2058);
and U2852 (N_2852,N_2194,N_2342);
nand U2853 (N_2853,N_2353,N_2275);
and U2854 (N_2854,N_2151,N_2277);
or U2855 (N_2855,N_2336,N_2204);
and U2856 (N_2856,N_2224,N_2439);
xor U2857 (N_2857,N_2338,N_2419);
or U2858 (N_2858,N_2399,N_2076);
nand U2859 (N_2859,N_2186,N_2379);
or U2860 (N_2860,N_2483,N_2268);
or U2861 (N_2861,N_2225,N_2425);
and U2862 (N_2862,N_2192,N_2086);
nand U2863 (N_2863,N_2042,N_2115);
nor U2864 (N_2864,N_2018,N_2072);
nand U2865 (N_2865,N_2263,N_2266);
nand U2866 (N_2866,N_2403,N_2174);
or U2867 (N_2867,N_2397,N_2061);
and U2868 (N_2868,N_2289,N_2209);
nor U2869 (N_2869,N_2203,N_2463);
or U2870 (N_2870,N_2390,N_2006);
xor U2871 (N_2871,N_2420,N_2346);
or U2872 (N_2872,N_2217,N_2436);
nor U2873 (N_2873,N_2144,N_2374);
xor U2874 (N_2874,N_2310,N_2414);
and U2875 (N_2875,N_2257,N_2361);
xor U2876 (N_2876,N_2422,N_2346);
and U2877 (N_2877,N_2005,N_2000);
nand U2878 (N_2878,N_2138,N_2074);
and U2879 (N_2879,N_2322,N_2356);
or U2880 (N_2880,N_2148,N_2278);
and U2881 (N_2881,N_2370,N_2017);
nand U2882 (N_2882,N_2437,N_2392);
or U2883 (N_2883,N_2432,N_2471);
and U2884 (N_2884,N_2010,N_2116);
nand U2885 (N_2885,N_2169,N_2111);
nor U2886 (N_2886,N_2253,N_2162);
xnor U2887 (N_2887,N_2238,N_2493);
and U2888 (N_2888,N_2246,N_2261);
and U2889 (N_2889,N_2039,N_2302);
and U2890 (N_2890,N_2486,N_2452);
xnor U2891 (N_2891,N_2474,N_2327);
nor U2892 (N_2892,N_2290,N_2270);
nor U2893 (N_2893,N_2317,N_2376);
nor U2894 (N_2894,N_2220,N_2191);
nor U2895 (N_2895,N_2070,N_2039);
or U2896 (N_2896,N_2322,N_2393);
xor U2897 (N_2897,N_2459,N_2310);
or U2898 (N_2898,N_2080,N_2215);
nand U2899 (N_2899,N_2490,N_2335);
xor U2900 (N_2900,N_2087,N_2142);
nor U2901 (N_2901,N_2495,N_2483);
or U2902 (N_2902,N_2405,N_2044);
nand U2903 (N_2903,N_2093,N_2228);
or U2904 (N_2904,N_2418,N_2123);
xnor U2905 (N_2905,N_2310,N_2224);
or U2906 (N_2906,N_2066,N_2051);
and U2907 (N_2907,N_2118,N_2163);
xor U2908 (N_2908,N_2181,N_2245);
xor U2909 (N_2909,N_2272,N_2090);
nand U2910 (N_2910,N_2164,N_2342);
or U2911 (N_2911,N_2320,N_2168);
nor U2912 (N_2912,N_2396,N_2045);
and U2913 (N_2913,N_2198,N_2099);
nand U2914 (N_2914,N_2145,N_2377);
nor U2915 (N_2915,N_2324,N_2193);
and U2916 (N_2916,N_2189,N_2499);
nor U2917 (N_2917,N_2410,N_2458);
xor U2918 (N_2918,N_2461,N_2492);
and U2919 (N_2919,N_2158,N_2046);
and U2920 (N_2920,N_2471,N_2253);
nor U2921 (N_2921,N_2035,N_2160);
and U2922 (N_2922,N_2491,N_2144);
or U2923 (N_2923,N_2438,N_2323);
and U2924 (N_2924,N_2315,N_2489);
nand U2925 (N_2925,N_2043,N_2420);
nand U2926 (N_2926,N_2326,N_2249);
xnor U2927 (N_2927,N_2339,N_2052);
xnor U2928 (N_2928,N_2377,N_2469);
and U2929 (N_2929,N_2305,N_2120);
and U2930 (N_2930,N_2242,N_2383);
or U2931 (N_2931,N_2232,N_2142);
xnor U2932 (N_2932,N_2321,N_2145);
nand U2933 (N_2933,N_2164,N_2233);
and U2934 (N_2934,N_2092,N_2390);
nand U2935 (N_2935,N_2223,N_2188);
xnor U2936 (N_2936,N_2122,N_2019);
nand U2937 (N_2937,N_2316,N_2358);
nand U2938 (N_2938,N_2478,N_2197);
xnor U2939 (N_2939,N_2357,N_2315);
nor U2940 (N_2940,N_2404,N_2364);
or U2941 (N_2941,N_2341,N_2091);
nand U2942 (N_2942,N_2357,N_2387);
nor U2943 (N_2943,N_2002,N_2258);
xor U2944 (N_2944,N_2203,N_2492);
and U2945 (N_2945,N_2204,N_2124);
and U2946 (N_2946,N_2486,N_2256);
nand U2947 (N_2947,N_2073,N_2479);
nor U2948 (N_2948,N_2155,N_2441);
or U2949 (N_2949,N_2116,N_2124);
xnor U2950 (N_2950,N_2333,N_2435);
or U2951 (N_2951,N_2272,N_2489);
or U2952 (N_2952,N_2309,N_2499);
nand U2953 (N_2953,N_2036,N_2093);
nand U2954 (N_2954,N_2219,N_2400);
nand U2955 (N_2955,N_2022,N_2252);
or U2956 (N_2956,N_2262,N_2361);
nand U2957 (N_2957,N_2206,N_2049);
nand U2958 (N_2958,N_2205,N_2115);
nor U2959 (N_2959,N_2413,N_2495);
nor U2960 (N_2960,N_2084,N_2495);
and U2961 (N_2961,N_2001,N_2457);
nor U2962 (N_2962,N_2222,N_2119);
or U2963 (N_2963,N_2104,N_2441);
nor U2964 (N_2964,N_2286,N_2272);
and U2965 (N_2965,N_2011,N_2363);
or U2966 (N_2966,N_2034,N_2014);
or U2967 (N_2967,N_2324,N_2291);
nor U2968 (N_2968,N_2474,N_2337);
xnor U2969 (N_2969,N_2142,N_2389);
or U2970 (N_2970,N_2142,N_2354);
or U2971 (N_2971,N_2159,N_2020);
xnor U2972 (N_2972,N_2300,N_2093);
nand U2973 (N_2973,N_2365,N_2284);
nor U2974 (N_2974,N_2088,N_2104);
nor U2975 (N_2975,N_2037,N_2026);
or U2976 (N_2976,N_2161,N_2433);
nor U2977 (N_2977,N_2128,N_2326);
xor U2978 (N_2978,N_2269,N_2003);
xnor U2979 (N_2979,N_2033,N_2107);
nand U2980 (N_2980,N_2103,N_2222);
nand U2981 (N_2981,N_2216,N_2013);
nor U2982 (N_2982,N_2297,N_2260);
and U2983 (N_2983,N_2110,N_2166);
xor U2984 (N_2984,N_2477,N_2085);
and U2985 (N_2985,N_2354,N_2106);
and U2986 (N_2986,N_2410,N_2144);
and U2987 (N_2987,N_2039,N_2102);
nand U2988 (N_2988,N_2158,N_2485);
xor U2989 (N_2989,N_2135,N_2452);
and U2990 (N_2990,N_2443,N_2470);
nand U2991 (N_2991,N_2257,N_2230);
nor U2992 (N_2992,N_2153,N_2198);
xor U2993 (N_2993,N_2429,N_2244);
and U2994 (N_2994,N_2331,N_2349);
nand U2995 (N_2995,N_2422,N_2231);
and U2996 (N_2996,N_2045,N_2382);
xnor U2997 (N_2997,N_2481,N_2059);
xor U2998 (N_2998,N_2033,N_2304);
or U2999 (N_2999,N_2197,N_2070);
and U3000 (N_3000,N_2658,N_2515);
xnor U3001 (N_3001,N_2587,N_2702);
xor U3002 (N_3002,N_2531,N_2568);
and U3003 (N_3003,N_2637,N_2780);
xor U3004 (N_3004,N_2633,N_2701);
or U3005 (N_3005,N_2916,N_2749);
nand U3006 (N_3006,N_2536,N_2902);
or U3007 (N_3007,N_2884,N_2646);
nor U3008 (N_3008,N_2887,N_2581);
xnor U3009 (N_3009,N_2662,N_2852);
nand U3010 (N_3010,N_2611,N_2886);
xnor U3011 (N_3011,N_2680,N_2904);
or U3012 (N_3012,N_2883,N_2817);
or U3013 (N_3013,N_2630,N_2871);
and U3014 (N_3014,N_2915,N_2641);
nor U3015 (N_3015,N_2688,N_2698);
xnor U3016 (N_3016,N_2726,N_2799);
or U3017 (N_3017,N_2789,N_2623);
or U3018 (N_3018,N_2982,N_2533);
nand U3019 (N_3019,N_2759,N_2717);
or U3020 (N_3020,N_2739,N_2559);
nor U3021 (N_3021,N_2931,N_2683);
nand U3022 (N_3022,N_2891,N_2919);
and U3023 (N_3023,N_2922,N_2737);
nor U3024 (N_3024,N_2728,N_2540);
nor U3025 (N_3025,N_2986,N_2797);
nand U3026 (N_3026,N_2996,N_2651);
and U3027 (N_3027,N_2750,N_2865);
xor U3028 (N_3028,N_2753,N_2825);
and U3029 (N_3029,N_2501,N_2649);
nand U3030 (N_3030,N_2804,N_2960);
nor U3031 (N_3031,N_2657,N_2732);
nor U3032 (N_3032,N_2861,N_2951);
and U3033 (N_3033,N_2744,N_2621);
or U3034 (N_3034,N_2577,N_2706);
or U3035 (N_3035,N_2517,N_2598);
xnor U3036 (N_3036,N_2670,N_2842);
or U3037 (N_3037,N_2578,N_2603);
nand U3038 (N_3038,N_2827,N_2970);
xor U3039 (N_3039,N_2714,N_2946);
and U3040 (N_3040,N_2859,N_2522);
nor U3041 (N_3041,N_2547,N_2542);
nand U3042 (N_3042,N_2729,N_2803);
or U3043 (N_3043,N_2513,N_2815);
nor U3044 (N_3044,N_2736,N_2609);
and U3045 (N_3045,N_2601,N_2634);
nand U3046 (N_3046,N_2932,N_2867);
nand U3047 (N_3047,N_2663,N_2597);
xor U3048 (N_3048,N_2795,N_2945);
and U3049 (N_3049,N_2622,N_2541);
or U3050 (N_3050,N_2711,N_2565);
and U3051 (N_3051,N_2537,N_2903);
xnor U3052 (N_3052,N_2573,N_2929);
or U3053 (N_3053,N_2880,N_2713);
xor U3054 (N_3054,N_2685,N_2920);
nand U3055 (N_3055,N_2735,N_2992);
and U3056 (N_3056,N_2776,N_2553);
xnor U3057 (N_3057,N_2707,N_2936);
or U3058 (N_3058,N_2505,N_2524);
nor U3059 (N_3059,N_2673,N_2740);
and U3060 (N_3060,N_2901,N_2695);
nand U3061 (N_3061,N_2636,N_2873);
or U3062 (N_3062,N_2864,N_2668);
and U3063 (N_3063,N_2585,N_2692);
and U3064 (N_3064,N_2907,N_2760);
nor U3065 (N_3065,N_2967,N_2521);
nor U3066 (N_3066,N_2660,N_2900);
xnor U3067 (N_3067,N_2975,N_2928);
xor U3068 (N_3068,N_2878,N_2872);
xor U3069 (N_3069,N_2669,N_2843);
or U3070 (N_3070,N_2790,N_2703);
nand U3071 (N_3071,N_2938,N_2857);
xnor U3072 (N_3072,N_2991,N_2994);
nand U3073 (N_3073,N_2972,N_2558);
or U3074 (N_3074,N_2767,N_2808);
or U3075 (N_3075,N_2911,N_2796);
and U3076 (N_3076,N_2869,N_2957);
xnor U3077 (N_3077,N_2503,N_2855);
nand U3078 (N_3078,N_2675,N_2882);
xor U3079 (N_3079,N_2560,N_2543);
and U3080 (N_3080,N_2627,N_2681);
and U3081 (N_3081,N_2580,N_2570);
nand U3082 (N_3082,N_2545,N_2950);
nor U3083 (N_3083,N_2774,N_2566);
xor U3084 (N_3084,N_2763,N_2879);
or U3085 (N_3085,N_2947,N_2672);
xor U3086 (N_3086,N_2571,N_2769);
nor U3087 (N_3087,N_2500,N_2518);
xor U3088 (N_3088,N_2617,N_2792);
or U3089 (N_3089,N_2514,N_2937);
nand U3090 (N_3090,N_2605,N_2958);
nor U3091 (N_3091,N_2550,N_2818);
xnor U3092 (N_3092,N_2574,N_2829);
nand U3093 (N_3093,N_2708,N_2775);
xor U3094 (N_3094,N_2602,N_2530);
nand U3095 (N_3095,N_2899,N_2794);
and U3096 (N_3096,N_2858,N_2716);
xnor U3097 (N_3097,N_2564,N_2665);
nor U3098 (N_3098,N_2511,N_2538);
xor U3099 (N_3099,N_2731,N_2823);
nor U3100 (N_3100,N_2826,N_2628);
nor U3101 (N_3101,N_2990,N_2892);
nor U3102 (N_3102,N_2752,N_2912);
nand U3103 (N_3103,N_2631,N_2983);
nand U3104 (N_3104,N_2913,N_2828);
or U3105 (N_3105,N_2582,N_2968);
xnor U3106 (N_3106,N_2730,N_2835);
and U3107 (N_3107,N_2906,N_2745);
or U3108 (N_3108,N_2589,N_2549);
and U3109 (N_3109,N_2607,N_2615);
xor U3110 (N_3110,N_2694,N_2898);
or U3111 (N_3111,N_2644,N_2691);
nand U3112 (N_3112,N_2625,N_2761);
or U3113 (N_3113,N_2682,N_2894);
nor U3114 (N_3114,N_2999,N_2594);
xor U3115 (N_3115,N_2684,N_2645);
or U3116 (N_3116,N_2526,N_2979);
xor U3117 (N_3117,N_2851,N_2697);
and U3118 (N_3118,N_2788,N_2838);
and U3119 (N_3119,N_2897,N_2941);
nor U3120 (N_3120,N_2596,N_2965);
nand U3121 (N_3121,N_2592,N_2870);
nor U3122 (N_3122,N_2525,N_2846);
or U3123 (N_3123,N_2943,N_2724);
or U3124 (N_3124,N_2926,N_2807);
xor U3125 (N_3125,N_2727,N_2757);
or U3126 (N_3126,N_2924,N_2743);
or U3127 (N_3127,N_2934,N_2802);
or U3128 (N_3128,N_2973,N_2954);
nor U3129 (N_3129,N_2600,N_2544);
xor U3130 (N_3130,N_2839,N_2719);
or U3131 (N_3131,N_2506,N_2569);
and U3132 (N_3132,N_2754,N_2532);
nand U3133 (N_3133,N_2656,N_2679);
nor U3134 (N_3134,N_2985,N_2908);
nor U3135 (N_3135,N_2624,N_2889);
or U3136 (N_3136,N_2678,N_2579);
xnor U3137 (N_3137,N_2770,N_2576);
nor U3138 (N_3138,N_2704,N_2654);
and U3139 (N_3139,N_2860,N_2626);
nand U3140 (N_3140,N_2925,N_2552);
nor U3141 (N_3141,N_2847,N_2667);
and U3142 (N_3142,N_2952,N_2755);
nor U3143 (N_3143,N_2746,N_2516);
nand U3144 (N_3144,N_2529,N_2953);
nand U3145 (N_3145,N_2554,N_2806);
or U3146 (N_3146,N_2987,N_2642);
and U3147 (N_3147,N_2567,N_2535);
or U3148 (N_3148,N_2664,N_2659);
nand U3149 (N_3149,N_2620,N_2791);
and U3150 (N_3150,N_2773,N_2647);
nor U3151 (N_3151,N_2853,N_2779);
and U3152 (N_3152,N_2787,N_2956);
nor U3153 (N_3153,N_2756,N_2885);
nor U3154 (N_3154,N_2995,N_2548);
nand U3155 (N_3155,N_2781,N_2961);
nor U3156 (N_3156,N_2921,N_2832);
or U3157 (N_3157,N_2700,N_2981);
and U3158 (N_3158,N_2896,N_2850);
and U3159 (N_3159,N_2862,N_2593);
nand U3160 (N_3160,N_2874,N_2639);
and U3161 (N_3161,N_2616,N_2762);
nor U3162 (N_3162,N_2635,N_2816);
nand U3163 (N_3163,N_2914,N_2748);
nand U3164 (N_3164,N_2557,N_2720);
and U3165 (N_3165,N_2980,N_2809);
or U3166 (N_3166,N_2689,N_2856);
nor U3167 (N_3167,N_2655,N_2638);
or U3168 (N_3168,N_2812,N_2722);
xnor U3169 (N_3169,N_2705,N_2822);
nand U3170 (N_3170,N_2877,N_2939);
or U3171 (N_3171,N_2562,N_2528);
nand U3172 (N_3172,N_2881,N_2507);
nand U3173 (N_3173,N_2805,N_2875);
or U3174 (N_3174,N_2629,N_2661);
nor U3175 (N_3175,N_2772,N_2813);
nand U3176 (N_3176,N_2677,N_2527);
or U3177 (N_3177,N_2844,N_2653);
and U3178 (N_3178,N_2801,N_2648);
xnor U3179 (N_3179,N_2786,N_2811);
or U3180 (N_3180,N_2502,N_2590);
and U3181 (N_3181,N_2863,N_2643);
and U3182 (N_3182,N_2833,N_2895);
xor U3183 (N_3183,N_2520,N_2930);
nor U3184 (N_3184,N_2509,N_2632);
and U3185 (N_3185,N_2854,N_2836);
xor U3186 (N_3186,N_2747,N_2519);
xor U3187 (N_3187,N_2523,N_2612);
and U3188 (N_3188,N_2741,N_2733);
or U3189 (N_3189,N_2588,N_2998);
xor U3190 (N_3190,N_2676,N_2510);
or U3191 (N_3191,N_2710,N_2765);
and U3192 (N_3192,N_2868,N_2821);
or U3193 (N_3193,N_2640,N_2652);
nor U3194 (N_3194,N_2686,N_2933);
nand U3195 (N_3195,N_2504,N_2546);
nand U3196 (N_3196,N_2604,N_2940);
nor U3197 (N_3197,N_2782,N_2534);
nand U3198 (N_3198,N_2935,N_2866);
xor U3199 (N_3199,N_2551,N_2778);
xor U3200 (N_3200,N_2610,N_2837);
xnor U3201 (N_3201,N_2959,N_2793);
nand U3202 (N_3202,N_2693,N_2712);
or U3203 (N_3203,N_2814,N_2595);
xor U3204 (N_3204,N_2845,N_2993);
or U3205 (N_3205,N_2619,N_2948);
and U3206 (N_3206,N_2674,N_2709);
nand U3207 (N_3207,N_2989,N_2783);
and U3208 (N_3208,N_2918,N_2555);
and U3209 (N_3209,N_2824,N_2966);
and U3210 (N_3210,N_2955,N_2810);
nand U3211 (N_3211,N_2909,N_2977);
xnor U3212 (N_3212,N_2650,N_2798);
nand U3213 (N_3213,N_2988,N_2890);
or U3214 (N_3214,N_2978,N_2888);
nand U3215 (N_3215,N_2841,N_2618);
xor U3216 (N_3216,N_2997,N_2949);
xor U3217 (N_3217,N_2819,N_2876);
and U3218 (N_3218,N_2751,N_2613);
and U3219 (N_3219,N_2599,N_2964);
or U3220 (N_3220,N_2563,N_2758);
or U3221 (N_3221,N_2738,N_2539);
or U3222 (N_3222,N_2784,N_2586);
nor U3223 (N_3223,N_2800,N_2893);
nor U3224 (N_3224,N_2831,N_2777);
or U3225 (N_3225,N_2984,N_2923);
and U3226 (N_3226,N_2764,N_2974);
nand U3227 (N_3227,N_2584,N_2976);
nand U3228 (N_3228,N_2768,N_2556);
xnor U3229 (N_3229,N_2671,N_2830);
nor U3230 (N_3230,N_2944,N_2606);
or U3231 (N_3231,N_2696,N_2848);
xor U3232 (N_3232,N_2512,N_2910);
xor U3233 (N_3233,N_2742,N_2771);
nand U3234 (N_3234,N_2840,N_2849);
and U3235 (N_3235,N_2561,N_2608);
and U3236 (N_3236,N_2969,N_2917);
nand U3237 (N_3237,N_2591,N_2725);
xnor U3238 (N_3238,N_2927,N_2905);
xor U3239 (N_3239,N_2666,N_2718);
nand U3240 (N_3240,N_2508,N_2687);
and U3241 (N_3241,N_2690,N_2962);
nor U3242 (N_3242,N_2699,N_2723);
xor U3243 (N_3243,N_2721,N_2766);
xor U3244 (N_3244,N_2614,N_2820);
nor U3245 (N_3245,N_2963,N_2834);
nor U3246 (N_3246,N_2971,N_2942);
and U3247 (N_3247,N_2734,N_2583);
nand U3248 (N_3248,N_2785,N_2715);
xor U3249 (N_3249,N_2572,N_2575);
nor U3250 (N_3250,N_2952,N_2830);
or U3251 (N_3251,N_2754,N_2563);
nor U3252 (N_3252,N_2597,N_2762);
xor U3253 (N_3253,N_2709,N_2551);
or U3254 (N_3254,N_2532,N_2737);
and U3255 (N_3255,N_2839,N_2916);
nand U3256 (N_3256,N_2879,N_2711);
xor U3257 (N_3257,N_2940,N_2612);
or U3258 (N_3258,N_2904,N_2799);
and U3259 (N_3259,N_2526,N_2574);
nand U3260 (N_3260,N_2892,N_2643);
nand U3261 (N_3261,N_2811,N_2793);
and U3262 (N_3262,N_2639,N_2753);
xor U3263 (N_3263,N_2688,N_2838);
xnor U3264 (N_3264,N_2612,N_2646);
nand U3265 (N_3265,N_2545,N_2782);
xor U3266 (N_3266,N_2983,N_2843);
or U3267 (N_3267,N_2723,N_2589);
xor U3268 (N_3268,N_2906,N_2945);
xor U3269 (N_3269,N_2505,N_2559);
and U3270 (N_3270,N_2781,N_2572);
nand U3271 (N_3271,N_2807,N_2860);
or U3272 (N_3272,N_2504,N_2838);
or U3273 (N_3273,N_2847,N_2805);
nor U3274 (N_3274,N_2832,N_2840);
nand U3275 (N_3275,N_2972,N_2876);
xor U3276 (N_3276,N_2553,N_2938);
and U3277 (N_3277,N_2953,N_2737);
or U3278 (N_3278,N_2947,N_2629);
nand U3279 (N_3279,N_2666,N_2576);
or U3280 (N_3280,N_2907,N_2608);
nand U3281 (N_3281,N_2885,N_2853);
nor U3282 (N_3282,N_2675,N_2966);
and U3283 (N_3283,N_2981,N_2684);
and U3284 (N_3284,N_2564,N_2759);
xnor U3285 (N_3285,N_2923,N_2595);
nor U3286 (N_3286,N_2738,N_2847);
xnor U3287 (N_3287,N_2905,N_2702);
nor U3288 (N_3288,N_2974,N_2860);
and U3289 (N_3289,N_2862,N_2741);
or U3290 (N_3290,N_2703,N_2658);
nand U3291 (N_3291,N_2678,N_2571);
nand U3292 (N_3292,N_2973,N_2623);
and U3293 (N_3293,N_2568,N_2726);
xor U3294 (N_3294,N_2947,N_2606);
or U3295 (N_3295,N_2601,N_2894);
and U3296 (N_3296,N_2591,N_2746);
and U3297 (N_3297,N_2887,N_2502);
and U3298 (N_3298,N_2514,N_2529);
nor U3299 (N_3299,N_2872,N_2740);
xor U3300 (N_3300,N_2524,N_2956);
xnor U3301 (N_3301,N_2594,N_2784);
or U3302 (N_3302,N_2959,N_2858);
or U3303 (N_3303,N_2817,N_2666);
nor U3304 (N_3304,N_2839,N_2589);
nor U3305 (N_3305,N_2978,N_2717);
xnor U3306 (N_3306,N_2672,N_2611);
or U3307 (N_3307,N_2611,N_2629);
and U3308 (N_3308,N_2897,N_2753);
or U3309 (N_3309,N_2675,N_2544);
xnor U3310 (N_3310,N_2794,N_2589);
and U3311 (N_3311,N_2886,N_2915);
or U3312 (N_3312,N_2749,N_2970);
and U3313 (N_3313,N_2850,N_2624);
nand U3314 (N_3314,N_2940,N_2510);
nand U3315 (N_3315,N_2780,N_2689);
or U3316 (N_3316,N_2523,N_2615);
or U3317 (N_3317,N_2500,N_2654);
nand U3318 (N_3318,N_2850,N_2564);
or U3319 (N_3319,N_2715,N_2555);
nor U3320 (N_3320,N_2758,N_2898);
nand U3321 (N_3321,N_2595,N_2695);
nand U3322 (N_3322,N_2905,N_2521);
and U3323 (N_3323,N_2839,N_2953);
nor U3324 (N_3324,N_2620,N_2872);
xnor U3325 (N_3325,N_2530,N_2794);
xnor U3326 (N_3326,N_2974,N_2752);
nor U3327 (N_3327,N_2717,N_2952);
or U3328 (N_3328,N_2706,N_2612);
or U3329 (N_3329,N_2797,N_2592);
xnor U3330 (N_3330,N_2586,N_2658);
and U3331 (N_3331,N_2846,N_2609);
nor U3332 (N_3332,N_2668,N_2897);
xnor U3333 (N_3333,N_2778,N_2621);
and U3334 (N_3334,N_2700,N_2580);
xnor U3335 (N_3335,N_2984,N_2706);
xor U3336 (N_3336,N_2958,N_2576);
or U3337 (N_3337,N_2881,N_2561);
xor U3338 (N_3338,N_2710,N_2670);
nor U3339 (N_3339,N_2743,N_2839);
xor U3340 (N_3340,N_2700,N_2898);
or U3341 (N_3341,N_2820,N_2507);
and U3342 (N_3342,N_2856,N_2670);
and U3343 (N_3343,N_2769,N_2674);
nor U3344 (N_3344,N_2911,N_2995);
nor U3345 (N_3345,N_2868,N_2567);
and U3346 (N_3346,N_2556,N_2693);
or U3347 (N_3347,N_2584,N_2992);
and U3348 (N_3348,N_2952,N_2923);
or U3349 (N_3349,N_2711,N_2833);
nor U3350 (N_3350,N_2937,N_2522);
nor U3351 (N_3351,N_2502,N_2638);
nand U3352 (N_3352,N_2663,N_2574);
xnor U3353 (N_3353,N_2994,N_2921);
nand U3354 (N_3354,N_2591,N_2900);
or U3355 (N_3355,N_2951,N_2972);
nor U3356 (N_3356,N_2863,N_2828);
nor U3357 (N_3357,N_2952,N_2630);
xnor U3358 (N_3358,N_2511,N_2677);
or U3359 (N_3359,N_2846,N_2631);
nand U3360 (N_3360,N_2967,N_2712);
and U3361 (N_3361,N_2838,N_2561);
xor U3362 (N_3362,N_2998,N_2709);
and U3363 (N_3363,N_2941,N_2621);
xnor U3364 (N_3364,N_2844,N_2615);
nand U3365 (N_3365,N_2990,N_2808);
or U3366 (N_3366,N_2681,N_2606);
nor U3367 (N_3367,N_2783,N_2860);
xnor U3368 (N_3368,N_2790,N_2972);
xnor U3369 (N_3369,N_2837,N_2557);
and U3370 (N_3370,N_2592,N_2684);
and U3371 (N_3371,N_2608,N_2984);
xnor U3372 (N_3372,N_2670,N_2646);
nand U3373 (N_3373,N_2767,N_2910);
nand U3374 (N_3374,N_2869,N_2669);
nand U3375 (N_3375,N_2501,N_2906);
nor U3376 (N_3376,N_2503,N_2841);
or U3377 (N_3377,N_2549,N_2968);
nor U3378 (N_3378,N_2542,N_2909);
and U3379 (N_3379,N_2642,N_2891);
xor U3380 (N_3380,N_2661,N_2845);
or U3381 (N_3381,N_2953,N_2889);
nand U3382 (N_3382,N_2988,N_2677);
nand U3383 (N_3383,N_2506,N_2568);
nor U3384 (N_3384,N_2720,N_2716);
nand U3385 (N_3385,N_2547,N_2564);
nand U3386 (N_3386,N_2761,N_2878);
xnor U3387 (N_3387,N_2875,N_2604);
nand U3388 (N_3388,N_2988,N_2754);
xnor U3389 (N_3389,N_2518,N_2630);
and U3390 (N_3390,N_2990,N_2744);
nand U3391 (N_3391,N_2670,N_2769);
nor U3392 (N_3392,N_2664,N_2515);
nand U3393 (N_3393,N_2859,N_2767);
nor U3394 (N_3394,N_2920,N_2584);
nor U3395 (N_3395,N_2654,N_2894);
xor U3396 (N_3396,N_2545,N_2744);
nand U3397 (N_3397,N_2557,N_2523);
nor U3398 (N_3398,N_2866,N_2791);
nor U3399 (N_3399,N_2975,N_2517);
nand U3400 (N_3400,N_2976,N_2599);
or U3401 (N_3401,N_2915,N_2818);
or U3402 (N_3402,N_2951,N_2532);
or U3403 (N_3403,N_2642,N_2679);
nand U3404 (N_3404,N_2688,N_2687);
xnor U3405 (N_3405,N_2583,N_2987);
nand U3406 (N_3406,N_2586,N_2703);
and U3407 (N_3407,N_2591,N_2748);
xor U3408 (N_3408,N_2816,N_2767);
nor U3409 (N_3409,N_2520,N_2543);
nand U3410 (N_3410,N_2577,N_2950);
nand U3411 (N_3411,N_2987,N_2758);
and U3412 (N_3412,N_2563,N_2669);
nor U3413 (N_3413,N_2691,N_2823);
or U3414 (N_3414,N_2997,N_2971);
or U3415 (N_3415,N_2999,N_2548);
xor U3416 (N_3416,N_2806,N_2564);
xor U3417 (N_3417,N_2640,N_2929);
or U3418 (N_3418,N_2867,N_2588);
or U3419 (N_3419,N_2986,N_2884);
xnor U3420 (N_3420,N_2691,N_2841);
xnor U3421 (N_3421,N_2787,N_2593);
nand U3422 (N_3422,N_2586,N_2746);
and U3423 (N_3423,N_2810,N_2674);
nor U3424 (N_3424,N_2626,N_2669);
nand U3425 (N_3425,N_2912,N_2614);
and U3426 (N_3426,N_2506,N_2525);
nand U3427 (N_3427,N_2501,N_2530);
or U3428 (N_3428,N_2885,N_2953);
nand U3429 (N_3429,N_2699,N_2820);
or U3430 (N_3430,N_2627,N_2871);
or U3431 (N_3431,N_2731,N_2873);
nand U3432 (N_3432,N_2743,N_2789);
nor U3433 (N_3433,N_2971,N_2881);
nand U3434 (N_3434,N_2650,N_2956);
nor U3435 (N_3435,N_2765,N_2697);
nor U3436 (N_3436,N_2673,N_2661);
nor U3437 (N_3437,N_2605,N_2785);
nor U3438 (N_3438,N_2697,N_2770);
nand U3439 (N_3439,N_2581,N_2551);
xor U3440 (N_3440,N_2694,N_2508);
xor U3441 (N_3441,N_2674,N_2682);
xnor U3442 (N_3442,N_2973,N_2501);
nor U3443 (N_3443,N_2909,N_2799);
nor U3444 (N_3444,N_2616,N_2665);
nor U3445 (N_3445,N_2730,N_2925);
nand U3446 (N_3446,N_2890,N_2756);
xor U3447 (N_3447,N_2807,N_2890);
nand U3448 (N_3448,N_2989,N_2952);
nand U3449 (N_3449,N_2724,N_2812);
nor U3450 (N_3450,N_2903,N_2723);
or U3451 (N_3451,N_2943,N_2770);
and U3452 (N_3452,N_2902,N_2747);
and U3453 (N_3453,N_2982,N_2526);
or U3454 (N_3454,N_2845,N_2651);
xnor U3455 (N_3455,N_2854,N_2754);
nand U3456 (N_3456,N_2904,N_2646);
nor U3457 (N_3457,N_2914,N_2981);
nand U3458 (N_3458,N_2868,N_2606);
or U3459 (N_3459,N_2865,N_2583);
nor U3460 (N_3460,N_2851,N_2661);
xor U3461 (N_3461,N_2673,N_2908);
xor U3462 (N_3462,N_2730,N_2676);
or U3463 (N_3463,N_2764,N_2783);
and U3464 (N_3464,N_2656,N_2743);
and U3465 (N_3465,N_2578,N_2557);
xor U3466 (N_3466,N_2717,N_2996);
nor U3467 (N_3467,N_2519,N_2762);
nand U3468 (N_3468,N_2960,N_2700);
or U3469 (N_3469,N_2829,N_2923);
and U3470 (N_3470,N_2887,N_2967);
and U3471 (N_3471,N_2669,N_2600);
or U3472 (N_3472,N_2753,N_2725);
and U3473 (N_3473,N_2642,N_2893);
and U3474 (N_3474,N_2897,N_2979);
nor U3475 (N_3475,N_2810,N_2864);
nand U3476 (N_3476,N_2688,N_2875);
or U3477 (N_3477,N_2795,N_2749);
xor U3478 (N_3478,N_2520,N_2560);
or U3479 (N_3479,N_2927,N_2536);
xnor U3480 (N_3480,N_2721,N_2725);
and U3481 (N_3481,N_2765,N_2790);
nor U3482 (N_3482,N_2902,N_2949);
and U3483 (N_3483,N_2818,N_2817);
nand U3484 (N_3484,N_2713,N_2942);
nor U3485 (N_3485,N_2856,N_2882);
or U3486 (N_3486,N_2522,N_2775);
xnor U3487 (N_3487,N_2923,N_2553);
nand U3488 (N_3488,N_2536,N_2510);
and U3489 (N_3489,N_2922,N_2989);
nor U3490 (N_3490,N_2727,N_2567);
or U3491 (N_3491,N_2694,N_2641);
or U3492 (N_3492,N_2914,N_2878);
nand U3493 (N_3493,N_2723,N_2952);
and U3494 (N_3494,N_2730,N_2642);
xnor U3495 (N_3495,N_2996,N_2935);
nor U3496 (N_3496,N_2841,N_2902);
xnor U3497 (N_3497,N_2914,N_2771);
nor U3498 (N_3498,N_2643,N_2880);
xor U3499 (N_3499,N_2598,N_2596);
nor U3500 (N_3500,N_3086,N_3420);
or U3501 (N_3501,N_3382,N_3324);
and U3502 (N_3502,N_3486,N_3255);
nor U3503 (N_3503,N_3146,N_3053);
or U3504 (N_3504,N_3311,N_3458);
nor U3505 (N_3505,N_3497,N_3263);
nor U3506 (N_3506,N_3366,N_3152);
nor U3507 (N_3507,N_3154,N_3401);
nor U3508 (N_3508,N_3171,N_3384);
nand U3509 (N_3509,N_3250,N_3249);
xor U3510 (N_3510,N_3134,N_3183);
or U3511 (N_3511,N_3432,N_3261);
or U3512 (N_3512,N_3169,N_3080);
nand U3513 (N_3513,N_3257,N_3399);
and U3514 (N_3514,N_3428,N_3270);
and U3515 (N_3515,N_3467,N_3403);
nor U3516 (N_3516,N_3296,N_3198);
or U3517 (N_3517,N_3179,N_3440);
nor U3518 (N_3518,N_3431,N_3021);
nor U3519 (N_3519,N_3306,N_3472);
and U3520 (N_3520,N_3278,N_3029);
nor U3521 (N_3521,N_3406,N_3030);
and U3522 (N_3522,N_3172,N_3065);
and U3523 (N_3523,N_3355,N_3484);
nor U3524 (N_3524,N_3004,N_3337);
nor U3525 (N_3525,N_3454,N_3387);
nand U3526 (N_3526,N_3412,N_3058);
nand U3527 (N_3527,N_3372,N_3248);
or U3528 (N_3528,N_3488,N_3364);
or U3529 (N_3529,N_3268,N_3000);
and U3530 (N_3530,N_3396,N_3465);
nor U3531 (N_3531,N_3457,N_3433);
nor U3532 (N_3532,N_3269,N_3499);
nor U3533 (N_3533,N_3425,N_3067);
nand U3534 (N_3534,N_3155,N_3208);
and U3535 (N_3535,N_3473,N_3277);
nand U3536 (N_3536,N_3418,N_3342);
nand U3537 (N_3537,N_3101,N_3343);
nor U3538 (N_3538,N_3104,N_3471);
nand U3539 (N_3539,N_3203,N_3416);
xor U3540 (N_3540,N_3056,N_3312);
xor U3541 (N_3541,N_3087,N_3247);
nand U3542 (N_3542,N_3421,N_3340);
nand U3543 (N_3543,N_3254,N_3411);
or U3544 (N_3544,N_3314,N_3037);
xor U3545 (N_3545,N_3327,N_3394);
nand U3546 (N_3546,N_3181,N_3307);
and U3547 (N_3547,N_3113,N_3218);
nand U3548 (N_3548,N_3444,N_3137);
nand U3549 (N_3549,N_3438,N_3336);
nand U3550 (N_3550,N_3066,N_3100);
nor U3551 (N_3551,N_3258,N_3455);
or U3552 (N_3552,N_3062,N_3196);
and U3553 (N_3553,N_3102,N_3069);
nand U3554 (N_3554,N_3129,N_3320);
nor U3555 (N_3555,N_3166,N_3359);
nor U3556 (N_3556,N_3015,N_3429);
nand U3557 (N_3557,N_3443,N_3220);
nand U3558 (N_3558,N_3132,N_3474);
nand U3559 (N_3559,N_3153,N_3392);
or U3560 (N_3560,N_3139,N_3106);
nand U3561 (N_3561,N_3151,N_3280);
or U3562 (N_3562,N_3447,N_3180);
xnor U3563 (N_3563,N_3121,N_3027);
or U3564 (N_3564,N_3093,N_3374);
xnor U3565 (N_3565,N_3301,N_3333);
nor U3566 (N_3566,N_3126,N_3468);
nand U3567 (N_3567,N_3223,N_3477);
nand U3568 (N_3568,N_3158,N_3334);
and U3569 (N_3569,N_3323,N_3259);
nand U3570 (N_3570,N_3291,N_3060);
xor U3571 (N_3571,N_3266,N_3008);
or U3572 (N_3572,N_3009,N_3271);
nor U3573 (N_3573,N_3043,N_3368);
or U3574 (N_3574,N_3156,N_3352);
xnor U3575 (N_3575,N_3245,N_3213);
and U3576 (N_3576,N_3483,N_3178);
nor U3577 (N_3577,N_3339,N_3222);
or U3578 (N_3578,N_3079,N_3174);
and U3579 (N_3579,N_3017,N_3480);
nand U3580 (N_3580,N_3300,N_3441);
xnor U3581 (N_3581,N_3304,N_3237);
nand U3582 (N_3582,N_3096,N_3138);
and U3583 (N_3583,N_3038,N_3191);
xor U3584 (N_3584,N_3319,N_3256);
xnor U3585 (N_3585,N_3348,N_3046);
nor U3586 (N_3586,N_3063,N_3185);
nand U3587 (N_3587,N_3439,N_3238);
and U3588 (N_3588,N_3493,N_3197);
or U3589 (N_3589,N_3175,N_3118);
nand U3590 (N_3590,N_3460,N_3184);
xnor U3591 (N_3591,N_3243,N_3089);
and U3592 (N_3592,N_3267,N_3083);
and U3593 (N_3593,N_3242,N_3281);
xnor U3594 (N_3594,N_3014,N_3305);
nor U3595 (N_3595,N_3285,N_3052);
xor U3596 (N_3596,N_3426,N_3091);
xor U3597 (N_3597,N_3230,N_3119);
xnor U3598 (N_3598,N_3316,N_3195);
or U3599 (N_3599,N_3075,N_3293);
xor U3600 (N_3600,N_3105,N_3451);
nor U3601 (N_3601,N_3356,N_3330);
or U3602 (N_3602,N_3313,N_3207);
and U3603 (N_3603,N_3456,N_3168);
nor U3604 (N_3604,N_3363,N_3033);
or U3605 (N_3605,N_3190,N_3288);
nand U3606 (N_3606,N_3408,N_3380);
xnor U3607 (N_3607,N_3244,N_3163);
nor U3608 (N_3608,N_3318,N_3369);
or U3609 (N_3609,N_3442,N_3262);
or U3610 (N_3610,N_3097,N_3236);
nand U3611 (N_3611,N_3260,N_3430);
and U3612 (N_3612,N_3001,N_3367);
nor U3613 (N_3613,N_3192,N_3354);
or U3614 (N_3614,N_3290,N_3231);
xnor U3615 (N_3615,N_3076,N_3272);
nand U3616 (N_3616,N_3322,N_3295);
nor U3617 (N_3617,N_3144,N_3020);
nand U3618 (N_3618,N_3461,N_3234);
nor U3619 (N_3619,N_3164,N_3481);
and U3620 (N_3620,N_3041,N_3498);
xor U3621 (N_3621,N_3048,N_3482);
or U3622 (N_3622,N_3331,N_3279);
or U3623 (N_3623,N_3404,N_3310);
nand U3624 (N_3624,N_3099,N_3379);
nor U3625 (N_3625,N_3240,N_3116);
or U3626 (N_3626,N_3286,N_3095);
and U3627 (N_3627,N_3026,N_3098);
xor U3628 (N_3628,N_3165,N_3189);
xnor U3629 (N_3629,N_3273,N_3315);
nand U3630 (N_3630,N_3298,N_3123);
nor U3631 (N_3631,N_3182,N_3159);
xnor U3632 (N_3632,N_3341,N_3167);
or U3633 (N_3633,N_3115,N_3003);
or U3634 (N_3634,N_3437,N_3393);
nand U3635 (N_3635,N_3452,N_3414);
and U3636 (N_3636,N_3206,N_3283);
and U3637 (N_3637,N_3410,N_3224);
nand U3638 (N_3638,N_3375,N_3358);
nor U3639 (N_3639,N_3317,N_3292);
and U3640 (N_3640,N_3332,N_3084);
or U3641 (N_3641,N_3040,N_3186);
and U3642 (N_3642,N_3459,N_3365);
nor U3643 (N_3643,N_3054,N_3199);
xnor U3644 (N_3644,N_3050,N_3219);
and U3645 (N_3645,N_3325,N_3391);
nand U3646 (N_3646,N_3162,N_3215);
nor U3647 (N_3647,N_3141,N_3055);
nor U3648 (N_3648,N_3214,N_3226);
or U3649 (N_3649,N_3494,N_3016);
xor U3650 (N_3650,N_3131,N_3326);
nor U3651 (N_3651,N_3209,N_3395);
nand U3652 (N_3652,N_3389,N_3059);
and U3653 (N_3653,N_3349,N_3350);
or U3654 (N_3654,N_3353,N_3338);
nor U3655 (N_3655,N_3303,N_3246);
xnor U3656 (N_3656,N_3487,N_3042);
and U3657 (N_3657,N_3485,N_3036);
or U3658 (N_3658,N_3034,N_3402);
and U3659 (N_3659,N_3361,N_3045);
and U3660 (N_3660,N_3405,N_3108);
nor U3661 (N_3661,N_3462,N_3227);
nand U3662 (N_3662,N_3204,N_3490);
nand U3663 (N_3663,N_3140,N_3413);
xnor U3664 (N_3664,N_3217,N_3085);
and U3665 (N_3665,N_3463,N_3229);
xnor U3666 (N_3666,N_3398,N_3212);
nand U3667 (N_3667,N_3148,N_3409);
xor U3668 (N_3668,N_3007,N_3188);
or U3669 (N_3669,N_3194,N_3479);
and U3670 (N_3670,N_3360,N_3039);
nand U3671 (N_3671,N_3423,N_3211);
or U3672 (N_3672,N_3176,N_3078);
nor U3673 (N_3673,N_3489,N_3068);
xor U3674 (N_3674,N_3057,N_3390);
or U3675 (N_3675,N_3415,N_3228);
or U3676 (N_3676,N_3233,N_3232);
and U3677 (N_3677,N_3371,N_3018);
nor U3678 (N_3678,N_3388,N_3193);
nor U3679 (N_3679,N_3170,N_3496);
nor U3680 (N_3680,N_3346,N_3107);
xnor U3681 (N_3681,N_3120,N_3299);
xnor U3682 (N_3682,N_3147,N_3135);
or U3683 (N_3683,N_3407,N_3061);
and U3684 (N_3684,N_3127,N_3377);
nor U3685 (N_3685,N_3435,N_3142);
xor U3686 (N_3686,N_3373,N_3210);
and U3687 (N_3687,N_3424,N_3145);
nor U3688 (N_3688,N_3202,N_3239);
nor U3689 (N_3689,N_3011,N_3276);
or U3690 (N_3690,N_3251,N_3157);
or U3691 (N_3691,N_3446,N_3434);
and U3692 (N_3692,N_3019,N_3449);
xnor U3693 (N_3693,N_3252,N_3397);
xor U3694 (N_3694,N_3370,N_3445);
nor U3695 (N_3695,N_3122,N_3200);
xnor U3696 (N_3696,N_3329,N_3072);
or U3697 (N_3697,N_3024,N_3351);
xor U3698 (N_3698,N_3235,N_3022);
nor U3699 (N_3699,N_3321,N_3453);
nor U3700 (N_3700,N_3112,N_3476);
nor U3701 (N_3701,N_3419,N_3284);
and U3702 (N_3702,N_3124,N_3309);
or U3703 (N_3703,N_3450,N_3297);
nand U3704 (N_3704,N_3225,N_3417);
nand U3705 (N_3705,N_3264,N_3469);
xor U3706 (N_3706,N_3287,N_3133);
nor U3707 (N_3707,N_3160,N_3241);
and U3708 (N_3708,N_3002,N_3077);
nor U3709 (N_3709,N_3010,N_3274);
xor U3710 (N_3710,N_3110,N_3023);
xnor U3711 (N_3711,N_3143,N_3308);
nor U3712 (N_3712,N_3221,N_3173);
nand U3713 (N_3713,N_3074,N_3470);
or U3714 (N_3714,N_3347,N_3094);
and U3715 (N_3715,N_3130,N_3117);
xor U3716 (N_3716,N_3109,N_3031);
or U3717 (N_3717,N_3073,N_3464);
or U3718 (N_3718,N_3025,N_3216);
or U3719 (N_3719,N_3253,N_3090);
xor U3720 (N_3720,N_3006,N_3161);
and U3721 (N_3721,N_3070,N_3344);
nor U3722 (N_3722,N_3044,N_3328);
or U3723 (N_3723,N_3128,N_3345);
nand U3724 (N_3724,N_3422,N_3381);
and U3725 (N_3725,N_3492,N_3071);
or U3726 (N_3726,N_3047,N_3362);
nor U3727 (N_3727,N_3378,N_3051);
and U3728 (N_3728,N_3205,N_3081);
or U3729 (N_3729,N_3376,N_3103);
nand U3730 (N_3730,N_3201,N_3032);
or U3731 (N_3731,N_3125,N_3427);
and U3732 (N_3732,N_3049,N_3335);
xor U3733 (N_3733,N_3064,N_3187);
and U3734 (N_3734,N_3092,N_3177);
and U3735 (N_3735,N_3012,N_3386);
nor U3736 (N_3736,N_3478,N_3136);
and U3737 (N_3737,N_3028,N_3357);
xor U3738 (N_3738,N_3150,N_3294);
and U3739 (N_3739,N_3491,N_3282);
or U3740 (N_3740,N_3114,N_3149);
or U3741 (N_3741,N_3111,N_3082);
nor U3742 (N_3742,N_3005,N_3436);
and U3743 (N_3743,N_3400,N_3495);
and U3744 (N_3744,N_3466,N_3035);
nand U3745 (N_3745,N_3302,N_3275);
nor U3746 (N_3746,N_3289,N_3265);
and U3747 (N_3747,N_3088,N_3448);
and U3748 (N_3748,N_3383,N_3475);
and U3749 (N_3749,N_3385,N_3013);
and U3750 (N_3750,N_3374,N_3129);
nand U3751 (N_3751,N_3119,N_3474);
nand U3752 (N_3752,N_3149,N_3078);
nand U3753 (N_3753,N_3292,N_3099);
or U3754 (N_3754,N_3079,N_3146);
or U3755 (N_3755,N_3372,N_3445);
and U3756 (N_3756,N_3064,N_3223);
and U3757 (N_3757,N_3357,N_3299);
or U3758 (N_3758,N_3367,N_3212);
nor U3759 (N_3759,N_3188,N_3250);
nand U3760 (N_3760,N_3047,N_3170);
xnor U3761 (N_3761,N_3256,N_3343);
and U3762 (N_3762,N_3227,N_3043);
and U3763 (N_3763,N_3247,N_3111);
and U3764 (N_3764,N_3221,N_3040);
nand U3765 (N_3765,N_3169,N_3121);
and U3766 (N_3766,N_3403,N_3087);
nand U3767 (N_3767,N_3382,N_3479);
nor U3768 (N_3768,N_3011,N_3399);
and U3769 (N_3769,N_3016,N_3131);
nand U3770 (N_3770,N_3402,N_3150);
nand U3771 (N_3771,N_3083,N_3461);
nand U3772 (N_3772,N_3221,N_3285);
nand U3773 (N_3773,N_3199,N_3011);
nor U3774 (N_3774,N_3018,N_3299);
and U3775 (N_3775,N_3183,N_3264);
or U3776 (N_3776,N_3048,N_3038);
and U3777 (N_3777,N_3486,N_3223);
or U3778 (N_3778,N_3027,N_3141);
xnor U3779 (N_3779,N_3327,N_3102);
xor U3780 (N_3780,N_3013,N_3077);
nand U3781 (N_3781,N_3424,N_3413);
xnor U3782 (N_3782,N_3361,N_3441);
xor U3783 (N_3783,N_3250,N_3423);
and U3784 (N_3784,N_3270,N_3341);
nand U3785 (N_3785,N_3386,N_3143);
or U3786 (N_3786,N_3142,N_3167);
nand U3787 (N_3787,N_3418,N_3125);
or U3788 (N_3788,N_3496,N_3293);
and U3789 (N_3789,N_3007,N_3340);
and U3790 (N_3790,N_3103,N_3444);
xnor U3791 (N_3791,N_3265,N_3067);
or U3792 (N_3792,N_3257,N_3467);
nand U3793 (N_3793,N_3475,N_3336);
nand U3794 (N_3794,N_3360,N_3204);
nand U3795 (N_3795,N_3383,N_3328);
nand U3796 (N_3796,N_3225,N_3263);
or U3797 (N_3797,N_3188,N_3322);
nand U3798 (N_3798,N_3153,N_3418);
nor U3799 (N_3799,N_3238,N_3354);
or U3800 (N_3800,N_3115,N_3151);
and U3801 (N_3801,N_3373,N_3461);
and U3802 (N_3802,N_3265,N_3019);
nor U3803 (N_3803,N_3221,N_3262);
nor U3804 (N_3804,N_3289,N_3356);
nor U3805 (N_3805,N_3103,N_3371);
nor U3806 (N_3806,N_3467,N_3202);
or U3807 (N_3807,N_3386,N_3342);
nor U3808 (N_3808,N_3106,N_3063);
nand U3809 (N_3809,N_3071,N_3024);
and U3810 (N_3810,N_3130,N_3022);
nor U3811 (N_3811,N_3245,N_3464);
nor U3812 (N_3812,N_3433,N_3180);
and U3813 (N_3813,N_3484,N_3205);
xnor U3814 (N_3814,N_3092,N_3202);
nand U3815 (N_3815,N_3286,N_3495);
xnor U3816 (N_3816,N_3230,N_3235);
nand U3817 (N_3817,N_3037,N_3262);
nand U3818 (N_3818,N_3064,N_3335);
nor U3819 (N_3819,N_3261,N_3439);
nand U3820 (N_3820,N_3499,N_3496);
nand U3821 (N_3821,N_3208,N_3479);
nand U3822 (N_3822,N_3032,N_3156);
nand U3823 (N_3823,N_3013,N_3483);
and U3824 (N_3824,N_3138,N_3270);
and U3825 (N_3825,N_3115,N_3060);
xnor U3826 (N_3826,N_3314,N_3099);
or U3827 (N_3827,N_3382,N_3325);
nand U3828 (N_3828,N_3267,N_3139);
and U3829 (N_3829,N_3317,N_3441);
nand U3830 (N_3830,N_3482,N_3270);
nand U3831 (N_3831,N_3229,N_3133);
nand U3832 (N_3832,N_3387,N_3040);
and U3833 (N_3833,N_3376,N_3451);
nor U3834 (N_3834,N_3150,N_3253);
or U3835 (N_3835,N_3176,N_3275);
or U3836 (N_3836,N_3494,N_3423);
xor U3837 (N_3837,N_3381,N_3255);
xor U3838 (N_3838,N_3000,N_3148);
and U3839 (N_3839,N_3292,N_3090);
xnor U3840 (N_3840,N_3221,N_3063);
or U3841 (N_3841,N_3105,N_3183);
or U3842 (N_3842,N_3455,N_3342);
xnor U3843 (N_3843,N_3227,N_3410);
nor U3844 (N_3844,N_3143,N_3306);
and U3845 (N_3845,N_3044,N_3307);
nand U3846 (N_3846,N_3083,N_3118);
xor U3847 (N_3847,N_3336,N_3160);
and U3848 (N_3848,N_3026,N_3376);
or U3849 (N_3849,N_3202,N_3149);
or U3850 (N_3850,N_3043,N_3232);
nor U3851 (N_3851,N_3045,N_3164);
xnor U3852 (N_3852,N_3273,N_3230);
and U3853 (N_3853,N_3463,N_3494);
nor U3854 (N_3854,N_3310,N_3033);
xnor U3855 (N_3855,N_3405,N_3400);
and U3856 (N_3856,N_3452,N_3287);
nand U3857 (N_3857,N_3146,N_3330);
nor U3858 (N_3858,N_3108,N_3303);
nand U3859 (N_3859,N_3081,N_3386);
nand U3860 (N_3860,N_3037,N_3150);
and U3861 (N_3861,N_3418,N_3447);
and U3862 (N_3862,N_3393,N_3340);
and U3863 (N_3863,N_3215,N_3029);
or U3864 (N_3864,N_3495,N_3391);
nor U3865 (N_3865,N_3470,N_3315);
nand U3866 (N_3866,N_3021,N_3268);
or U3867 (N_3867,N_3124,N_3383);
nand U3868 (N_3868,N_3463,N_3200);
xnor U3869 (N_3869,N_3261,N_3398);
nor U3870 (N_3870,N_3434,N_3176);
or U3871 (N_3871,N_3461,N_3430);
or U3872 (N_3872,N_3144,N_3031);
and U3873 (N_3873,N_3184,N_3334);
xnor U3874 (N_3874,N_3478,N_3033);
and U3875 (N_3875,N_3458,N_3091);
or U3876 (N_3876,N_3251,N_3435);
or U3877 (N_3877,N_3107,N_3278);
and U3878 (N_3878,N_3465,N_3248);
or U3879 (N_3879,N_3160,N_3174);
or U3880 (N_3880,N_3010,N_3279);
xnor U3881 (N_3881,N_3408,N_3118);
nand U3882 (N_3882,N_3098,N_3461);
or U3883 (N_3883,N_3320,N_3206);
nand U3884 (N_3884,N_3373,N_3069);
nor U3885 (N_3885,N_3191,N_3077);
or U3886 (N_3886,N_3318,N_3246);
and U3887 (N_3887,N_3103,N_3226);
or U3888 (N_3888,N_3119,N_3487);
nand U3889 (N_3889,N_3420,N_3337);
xor U3890 (N_3890,N_3175,N_3266);
or U3891 (N_3891,N_3197,N_3464);
xor U3892 (N_3892,N_3007,N_3216);
nor U3893 (N_3893,N_3400,N_3016);
nor U3894 (N_3894,N_3239,N_3297);
and U3895 (N_3895,N_3166,N_3204);
or U3896 (N_3896,N_3015,N_3276);
nor U3897 (N_3897,N_3116,N_3219);
or U3898 (N_3898,N_3282,N_3297);
nor U3899 (N_3899,N_3056,N_3456);
or U3900 (N_3900,N_3499,N_3096);
and U3901 (N_3901,N_3017,N_3470);
nand U3902 (N_3902,N_3361,N_3116);
nor U3903 (N_3903,N_3152,N_3163);
or U3904 (N_3904,N_3313,N_3422);
and U3905 (N_3905,N_3488,N_3424);
xor U3906 (N_3906,N_3102,N_3119);
nor U3907 (N_3907,N_3246,N_3208);
xor U3908 (N_3908,N_3150,N_3047);
and U3909 (N_3909,N_3030,N_3308);
nor U3910 (N_3910,N_3337,N_3027);
or U3911 (N_3911,N_3162,N_3436);
nand U3912 (N_3912,N_3483,N_3117);
nor U3913 (N_3913,N_3337,N_3240);
and U3914 (N_3914,N_3332,N_3018);
and U3915 (N_3915,N_3337,N_3339);
nor U3916 (N_3916,N_3358,N_3178);
or U3917 (N_3917,N_3382,N_3403);
nand U3918 (N_3918,N_3084,N_3118);
or U3919 (N_3919,N_3470,N_3381);
nand U3920 (N_3920,N_3025,N_3253);
and U3921 (N_3921,N_3410,N_3340);
nand U3922 (N_3922,N_3080,N_3351);
nor U3923 (N_3923,N_3383,N_3476);
nor U3924 (N_3924,N_3164,N_3028);
xor U3925 (N_3925,N_3157,N_3069);
and U3926 (N_3926,N_3438,N_3202);
xor U3927 (N_3927,N_3137,N_3160);
or U3928 (N_3928,N_3068,N_3229);
nand U3929 (N_3929,N_3451,N_3052);
and U3930 (N_3930,N_3180,N_3255);
xor U3931 (N_3931,N_3068,N_3402);
and U3932 (N_3932,N_3303,N_3296);
xor U3933 (N_3933,N_3241,N_3365);
and U3934 (N_3934,N_3472,N_3379);
nand U3935 (N_3935,N_3493,N_3133);
xnor U3936 (N_3936,N_3238,N_3357);
nand U3937 (N_3937,N_3276,N_3485);
nand U3938 (N_3938,N_3265,N_3364);
and U3939 (N_3939,N_3482,N_3078);
nor U3940 (N_3940,N_3049,N_3244);
nor U3941 (N_3941,N_3352,N_3402);
or U3942 (N_3942,N_3347,N_3318);
and U3943 (N_3943,N_3211,N_3174);
nand U3944 (N_3944,N_3234,N_3182);
nor U3945 (N_3945,N_3022,N_3115);
nor U3946 (N_3946,N_3015,N_3045);
nor U3947 (N_3947,N_3142,N_3447);
nor U3948 (N_3948,N_3451,N_3144);
nand U3949 (N_3949,N_3074,N_3256);
nor U3950 (N_3950,N_3436,N_3018);
and U3951 (N_3951,N_3232,N_3155);
nor U3952 (N_3952,N_3475,N_3248);
nand U3953 (N_3953,N_3117,N_3229);
nand U3954 (N_3954,N_3143,N_3122);
or U3955 (N_3955,N_3423,N_3159);
xor U3956 (N_3956,N_3223,N_3412);
and U3957 (N_3957,N_3208,N_3281);
nor U3958 (N_3958,N_3342,N_3308);
nand U3959 (N_3959,N_3081,N_3142);
or U3960 (N_3960,N_3355,N_3189);
nand U3961 (N_3961,N_3463,N_3302);
xnor U3962 (N_3962,N_3210,N_3241);
xnor U3963 (N_3963,N_3169,N_3145);
nand U3964 (N_3964,N_3309,N_3429);
or U3965 (N_3965,N_3299,N_3493);
nand U3966 (N_3966,N_3356,N_3396);
nor U3967 (N_3967,N_3048,N_3398);
nor U3968 (N_3968,N_3172,N_3349);
and U3969 (N_3969,N_3444,N_3490);
or U3970 (N_3970,N_3058,N_3302);
nand U3971 (N_3971,N_3145,N_3287);
or U3972 (N_3972,N_3381,N_3129);
xor U3973 (N_3973,N_3366,N_3215);
and U3974 (N_3974,N_3265,N_3112);
xor U3975 (N_3975,N_3069,N_3073);
nand U3976 (N_3976,N_3293,N_3182);
nor U3977 (N_3977,N_3258,N_3459);
nand U3978 (N_3978,N_3331,N_3288);
or U3979 (N_3979,N_3181,N_3496);
and U3980 (N_3980,N_3100,N_3174);
xnor U3981 (N_3981,N_3018,N_3314);
nand U3982 (N_3982,N_3390,N_3301);
nor U3983 (N_3983,N_3074,N_3475);
or U3984 (N_3984,N_3072,N_3179);
or U3985 (N_3985,N_3327,N_3426);
xnor U3986 (N_3986,N_3043,N_3163);
or U3987 (N_3987,N_3476,N_3473);
xor U3988 (N_3988,N_3470,N_3175);
or U3989 (N_3989,N_3243,N_3488);
and U3990 (N_3990,N_3336,N_3322);
nand U3991 (N_3991,N_3212,N_3297);
nor U3992 (N_3992,N_3157,N_3311);
nor U3993 (N_3993,N_3180,N_3036);
or U3994 (N_3994,N_3495,N_3265);
or U3995 (N_3995,N_3004,N_3189);
nor U3996 (N_3996,N_3099,N_3189);
nand U3997 (N_3997,N_3488,N_3154);
xor U3998 (N_3998,N_3164,N_3463);
xor U3999 (N_3999,N_3249,N_3447);
nor U4000 (N_4000,N_3521,N_3744);
and U4001 (N_4001,N_3801,N_3976);
nand U4002 (N_4002,N_3986,N_3648);
or U4003 (N_4003,N_3613,N_3653);
and U4004 (N_4004,N_3676,N_3852);
xnor U4005 (N_4005,N_3909,N_3752);
xor U4006 (N_4006,N_3687,N_3711);
nor U4007 (N_4007,N_3694,N_3951);
or U4008 (N_4008,N_3791,N_3634);
nand U4009 (N_4009,N_3566,N_3544);
nand U4010 (N_4010,N_3865,N_3778);
nand U4011 (N_4011,N_3656,N_3892);
nand U4012 (N_4012,N_3858,N_3912);
and U4013 (N_4013,N_3849,N_3954);
or U4014 (N_4014,N_3818,N_3925);
and U4015 (N_4015,N_3735,N_3949);
xnor U4016 (N_4016,N_3580,N_3828);
nand U4017 (N_4017,N_3884,N_3916);
or U4018 (N_4018,N_3804,N_3797);
and U4019 (N_4019,N_3957,N_3651);
and U4020 (N_4020,N_3635,N_3863);
xor U4021 (N_4021,N_3757,N_3528);
xor U4022 (N_4022,N_3713,N_3642);
nand U4023 (N_4023,N_3607,N_3817);
xnor U4024 (N_4024,N_3795,N_3866);
nor U4025 (N_4025,N_3641,N_3592);
or U4026 (N_4026,N_3888,N_3983);
xnor U4027 (N_4027,N_3738,N_3968);
xor U4028 (N_4028,N_3980,N_3591);
xnor U4029 (N_4029,N_3948,N_3990);
nor U4030 (N_4030,N_3924,N_3947);
xor U4031 (N_4031,N_3515,N_3511);
nor U4032 (N_4032,N_3869,N_3677);
or U4033 (N_4033,N_3771,N_3862);
and U4034 (N_4034,N_3729,N_3880);
nand U4035 (N_4035,N_3767,N_3549);
xor U4036 (N_4036,N_3820,N_3879);
or U4037 (N_4037,N_3628,N_3668);
nor U4038 (N_4038,N_3814,N_3576);
xnor U4039 (N_4039,N_3612,N_3736);
nor U4040 (N_4040,N_3906,N_3901);
nor U4041 (N_4041,N_3755,N_3546);
and U4042 (N_4042,N_3590,N_3898);
or U4043 (N_4043,N_3946,N_3522);
nor U4044 (N_4044,N_3977,N_3507);
nor U4045 (N_4045,N_3559,N_3971);
or U4046 (N_4046,N_3763,N_3710);
or U4047 (N_4047,N_3589,N_3835);
xor U4048 (N_4048,N_3688,N_3707);
or U4049 (N_4049,N_3984,N_3700);
or U4050 (N_4050,N_3856,N_3671);
nor U4051 (N_4051,N_3517,N_3706);
and U4052 (N_4052,N_3722,N_3867);
and U4053 (N_4053,N_3601,N_3913);
xor U4054 (N_4054,N_3701,N_3709);
nand U4055 (N_4055,N_3824,N_3626);
xor U4056 (N_4056,N_3810,N_3702);
and U4057 (N_4057,N_3734,N_3654);
and U4058 (N_4058,N_3508,N_3779);
and U4059 (N_4059,N_3667,N_3562);
and U4060 (N_4060,N_3800,N_3535);
and U4061 (N_4061,N_3605,N_3716);
or U4062 (N_4062,N_3991,N_3506);
nand U4063 (N_4063,N_3705,N_3583);
nor U4064 (N_4064,N_3708,N_3678);
nand U4065 (N_4065,N_3693,N_3882);
nor U4066 (N_4066,N_3561,N_3987);
nor U4067 (N_4067,N_3806,N_3611);
or U4068 (N_4068,N_3776,N_3629);
xor U4069 (N_4069,N_3900,N_3540);
nor U4070 (N_4070,N_3685,N_3740);
or U4071 (N_4071,N_3588,N_3930);
nand U4072 (N_4072,N_3550,N_3837);
nand U4073 (N_4073,N_3632,N_3855);
nor U4074 (N_4074,N_3899,N_3664);
nand U4075 (N_4075,N_3665,N_3772);
nand U4076 (N_4076,N_3773,N_3881);
and U4077 (N_4077,N_3682,N_3574);
and U4078 (N_4078,N_3696,N_3753);
xnor U4079 (N_4079,N_3934,N_3661);
nand U4080 (N_4080,N_3717,N_3860);
and U4081 (N_4081,N_3650,N_3802);
and U4082 (N_4082,N_3624,N_3789);
nand U4083 (N_4083,N_3578,N_3614);
nand U4084 (N_4084,N_3887,N_3695);
nand U4085 (N_4085,N_3812,N_3966);
or U4086 (N_4086,N_3754,N_3870);
nand U4087 (N_4087,N_3610,N_3878);
nand U4088 (N_4088,N_3907,N_3842);
and U4089 (N_4089,N_3638,N_3926);
or U4090 (N_4090,N_3952,N_3756);
and U4091 (N_4091,N_3942,N_3974);
xor U4092 (N_4092,N_3575,N_3564);
nor U4093 (N_4093,N_3644,N_3686);
nand U4094 (N_4094,N_3959,N_3568);
xnor U4095 (N_4095,N_3718,N_3785);
and U4096 (N_4096,N_3799,N_3973);
nor U4097 (N_4097,N_3875,N_3950);
or U4098 (N_4098,N_3895,N_3853);
nand U4099 (N_4099,N_3794,N_3847);
nor U4100 (N_4100,N_3584,N_3871);
and U4101 (N_4101,N_3739,N_3958);
nand U4102 (N_4102,N_3723,N_3816);
xor U4103 (N_4103,N_3874,N_3586);
and U4104 (N_4104,N_3827,N_3724);
nand U4105 (N_4105,N_3885,N_3750);
nor U4106 (N_4106,N_3598,N_3886);
and U4107 (N_4107,N_3620,N_3539);
and U4108 (N_4108,N_3793,N_3516);
xor U4109 (N_4109,N_3999,N_3536);
xnor U4110 (N_4110,N_3581,N_3903);
nor U4111 (N_4111,N_3808,N_3979);
xor U4112 (N_4112,N_3680,N_3981);
or U4113 (N_4113,N_3790,N_3531);
nor U4114 (N_4114,N_3989,N_3955);
and U4115 (N_4115,N_3727,N_3967);
nor U4116 (N_4116,N_3647,N_3525);
nand U4117 (N_4117,N_3622,N_3832);
nand U4118 (N_4118,N_3937,N_3572);
nor U4119 (N_4119,N_3645,N_3587);
nor U4120 (N_4120,N_3931,N_3652);
or U4121 (N_4121,N_3662,N_3555);
nor U4122 (N_4122,N_3965,N_3962);
xnor U4123 (N_4123,N_3944,N_3780);
nand U4124 (N_4124,N_3787,N_3530);
and U4125 (N_4125,N_3660,N_3501);
xnor U4126 (N_4126,N_3993,N_3692);
or U4127 (N_4127,N_3640,N_3631);
nor U4128 (N_4128,N_3670,N_3768);
nor U4129 (N_4129,N_3577,N_3963);
xor U4130 (N_4130,N_3741,N_3658);
or U4131 (N_4131,N_3932,N_3877);
nor U4132 (N_4132,N_3630,N_3594);
nand U4133 (N_4133,N_3714,N_3617);
nor U4134 (N_4134,N_3929,N_3836);
xor U4135 (N_4135,N_3585,N_3831);
nand U4136 (N_4136,N_3616,N_3503);
and U4137 (N_4137,N_3933,N_3745);
or U4138 (N_4138,N_3527,N_3659);
nand U4139 (N_4139,N_3910,N_3921);
and U4140 (N_4140,N_3915,N_3766);
nand U4141 (N_4141,N_3500,N_3759);
xor U4142 (N_4142,N_3758,N_3704);
xor U4143 (N_4143,N_3674,N_3784);
nand U4144 (N_4144,N_3938,N_3783);
xor U4145 (N_4145,N_3728,N_3819);
nand U4146 (N_4146,N_3883,N_3524);
or U4147 (N_4147,N_3571,N_3558);
or U4148 (N_4148,N_3529,N_3940);
and U4149 (N_4149,N_3737,N_3972);
nor U4150 (N_4150,N_3636,N_3803);
nand U4151 (N_4151,N_3551,N_3553);
and U4152 (N_4152,N_3994,N_3864);
or U4153 (N_4153,N_3838,N_3845);
or U4154 (N_4154,N_3821,N_3712);
nand U4155 (N_4155,N_3843,N_3719);
and U4156 (N_4156,N_3730,N_3597);
nand U4157 (N_4157,N_3859,N_3851);
nand U4158 (N_4158,N_3873,N_3945);
nor U4159 (N_4159,N_3770,N_3639);
or U4160 (N_4160,N_3788,N_3917);
xnor U4161 (N_4161,N_3606,N_3509);
or U4162 (N_4162,N_3563,N_3765);
or U4163 (N_4163,N_3512,N_3715);
and U4164 (N_4164,N_3978,N_3627);
or U4165 (N_4165,N_3593,N_3679);
and U4166 (N_4166,N_3775,N_3623);
and U4167 (N_4167,N_3518,N_3935);
or U4168 (N_4168,N_3997,N_3599);
and U4169 (N_4169,N_3513,N_3672);
or U4170 (N_4170,N_3643,N_3505);
xor U4171 (N_4171,N_3985,N_3996);
and U4172 (N_4172,N_3857,N_3618);
and U4173 (N_4173,N_3953,N_3699);
nor U4174 (N_4174,N_3602,N_3556);
nand U4175 (N_4175,N_3625,N_3896);
or U4176 (N_4176,N_3922,N_3840);
nand U4177 (N_4177,N_3582,N_3603);
nor U4178 (N_4178,N_3732,N_3600);
or U4179 (N_4179,N_3655,N_3960);
nand U4180 (N_4180,N_3782,N_3548);
nor U4181 (N_4181,N_3807,N_3547);
and U4182 (N_4182,N_3988,N_3746);
and U4183 (N_4183,N_3520,N_3519);
nand U4184 (N_4184,N_3846,N_3809);
and U4185 (N_4185,N_3684,N_3760);
and U4186 (N_4186,N_3908,N_3928);
nand U4187 (N_4187,N_3918,N_3905);
xor U4188 (N_4188,N_3904,N_3844);
nand U4189 (N_4189,N_3982,N_3764);
or U4190 (N_4190,N_3689,N_3646);
or U4191 (N_4191,N_3683,N_3811);
and U4192 (N_4192,N_3914,N_3839);
nor U4193 (N_4193,N_3927,N_3970);
and U4194 (N_4194,N_3663,N_3894);
nor U4195 (N_4195,N_3969,N_3786);
or U4196 (N_4196,N_3777,N_3579);
nor U4197 (N_4197,N_3830,N_3726);
nor U4198 (N_4198,N_3565,N_3554);
nand U4199 (N_4199,N_3537,N_3995);
or U4200 (N_4200,N_3541,N_3769);
nand U4201 (N_4201,N_3608,N_3825);
or U4202 (N_4202,N_3552,N_3813);
nor U4203 (N_4203,N_3649,N_3621);
and U4204 (N_4204,N_3720,N_3619);
nand U4205 (N_4205,N_3956,N_3889);
and U4206 (N_4206,N_3595,N_3911);
xnor U4207 (N_4207,N_3992,N_3543);
nor U4208 (N_4208,N_3854,N_3673);
and U4209 (N_4209,N_3538,N_3792);
nand U4210 (N_4210,N_3596,N_3573);
or U4211 (N_4211,N_3526,N_3703);
nand U4212 (N_4212,N_3633,N_3998);
nand U4213 (N_4213,N_3923,N_3781);
nor U4214 (N_4214,N_3961,N_3919);
or U4215 (N_4215,N_3534,N_3742);
or U4216 (N_4216,N_3681,N_3567);
xor U4217 (N_4217,N_3798,N_3848);
nand U4218 (N_4218,N_3569,N_3872);
or U4219 (N_4219,N_3691,N_3690);
nand U4220 (N_4220,N_3749,N_3721);
nand U4221 (N_4221,N_3666,N_3743);
and U4222 (N_4222,N_3975,N_3891);
nor U4223 (N_4223,N_3796,N_3523);
xor U4224 (N_4224,N_3560,N_3733);
nand U4225 (N_4225,N_3514,N_3897);
and U4226 (N_4226,N_3868,N_3941);
xnor U4227 (N_4227,N_3504,N_3604);
nor U4228 (N_4228,N_3805,N_3815);
or U4229 (N_4229,N_3747,N_3533);
and U4230 (N_4230,N_3964,N_3823);
nand U4231 (N_4231,N_3675,N_3669);
nor U4232 (N_4232,N_3890,N_3861);
or U4233 (N_4233,N_3725,N_3829);
and U4234 (N_4234,N_3850,N_3637);
or U4235 (N_4235,N_3902,N_3774);
nand U4236 (N_4236,N_3731,N_3609);
nor U4237 (N_4237,N_3920,N_3697);
nand U4238 (N_4238,N_3761,N_3657);
or U4239 (N_4239,N_3893,N_3542);
nand U4240 (N_4240,N_3826,N_3841);
xor U4241 (N_4241,N_3557,N_3833);
nand U4242 (N_4242,N_3532,N_3698);
and U4243 (N_4243,N_3943,N_3748);
and U4244 (N_4244,N_3615,N_3939);
or U4245 (N_4245,N_3510,N_3502);
nand U4246 (N_4246,N_3751,N_3876);
nor U4247 (N_4247,N_3822,N_3545);
or U4248 (N_4248,N_3762,N_3936);
and U4249 (N_4249,N_3570,N_3834);
nand U4250 (N_4250,N_3569,N_3684);
nand U4251 (N_4251,N_3834,N_3921);
nand U4252 (N_4252,N_3520,N_3743);
xor U4253 (N_4253,N_3969,N_3668);
xor U4254 (N_4254,N_3802,N_3963);
or U4255 (N_4255,N_3966,N_3904);
and U4256 (N_4256,N_3737,N_3509);
xnor U4257 (N_4257,N_3667,N_3693);
nor U4258 (N_4258,N_3780,N_3914);
or U4259 (N_4259,N_3705,N_3670);
and U4260 (N_4260,N_3547,N_3907);
xnor U4261 (N_4261,N_3512,N_3938);
and U4262 (N_4262,N_3643,N_3974);
xnor U4263 (N_4263,N_3997,N_3801);
and U4264 (N_4264,N_3708,N_3541);
and U4265 (N_4265,N_3672,N_3566);
nor U4266 (N_4266,N_3719,N_3805);
or U4267 (N_4267,N_3913,N_3800);
nor U4268 (N_4268,N_3520,N_3670);
and U4269 (N_4269,N_3745,N_3536);
nor U4270 (N_4270,N_3669,N_3836);
nor U4271 (N_4271,N_3892,N_3817);
and U4272 (N_4272,N_3769,N_3528);
nor U4273 (N_4273,N_3999,N_3880);
xnor U4274 (N_4274,N_3549,N_3975);
and U4275 (N_4275,N_3825,N_3749);
nand U4276 (N_4276,N_3898,N_3671);
and U4277 (N_4277,N_3918,N_3613);
or U4278 (N_4278,N_3730,N_3791);
nor U4279 (N_4279,N_3611,N_3994);
nand U4280 (N_4280,N_3512,N_3922);
xnor U4281 (N_4281,N_3636,N_3956);
or U4282 (N_4282,N_3989,N_3576);
xor U4283 (N_4283,N_3756,N_3961);
xor U4284 (N_4284,N_3575,N_3769);
and U4285 (N_4285,N_3819,N_3778);
or U4286 (N_4286,N_3590,N_3792);
nand U4287 (N_4287,N_3823,N_3805);
or U4288 (N_4288,N_3660,N_3645);
nor U4289 (N_4289,N_3639,N_3738);
or U4290 (N_4290,N_3785,N_3624);
xor U4291 (N_4291,N_3585,N_3994);
nand U4292 (N_4292,N_3695,N_3822);
or U4293 (N_4293,N_3820,N_3559);
and U4294 (N_4294,N_3675,N_3713);
and U4295 (N_4295,N_3520,N_3645);
and U4296 (N_4296,N_3938,N_3951);
nand U4297 (N_4297,N_3608,N_3875);
or U4298 (N_4298,N_3868,N_3776);
xnor U4299 (N_4299,N_3542,N_3829);
and U4300 (N_4300,N_3719,N_3521);
nand U4301 (N_4301,N_3935,N_3810);
xnor U4302 (N_4302,N_3898,N_3751);
or U4303 (N_4303,N_3577,N_3934);
xor U4304 (N_4304,N_3818,N_3639);
and U4305 (N_4305,N_3884,N_3516);
xnor U4306 (N_4306,N_3650,N_3675);
xnor U4307 (N_4307,N_3586,N_3916);
and U4308 (N_4308,N_3745,N_3541);
or U4309 (N_4309,N_3930,N_3608);
nor U4310 (N_4310,N_3696,N_3790);
xnor U4311 (N_4311,N_3803,N_3826);
nor U4312 (N_4312,N_3552,N_3827);
nor U4313 (N_4313,N_3565,N_3993);
or U4314 (N_4314,N_3738,N_3550);
xor U4315 (N_4315,N_3725,N_3992);
xor U4316 (N_4316,N_3535,N_3576);
xor U4317 (N_4317,N_3685,N_3604);
and U4318 (N_4318,N_3524,N_3636);
or U4319 (N_4319,N_3598,N_3558);
nand U4320 (N_4320,N_3806,N_3559);
and U4321 (N_4321,N_3556,N_3686);
and U4322 (N_4322,N_3542,N_3717);
and U4323 (N_4323,N_3598,N_3863);
and U4324 (N_4324,N_3627,N_3629);
and U4325 (N_4325,N_3902,N_3956);
nor U4326 (N_4326,N_3751,N_3605);
nand U4327 (N_4327,N_3985,N_3659);
nand U4328 (N_4328,N_3635,N_3929);
or U4329 (N_4329,N_3989,N_3818);
nand U4330 (N_4330,N_3677,N_3830);
or U4331 (N_4331,N_3573,N_3910);
nand U4332 (N_4332,N_3623,N_3642);
or U4333 (N_4333,N_3665,N_3982);
xor U4334 (N_4334,N_3756,N_3846);
nor U4335 (N_4335,N_3669,N_3982);
and U4336 (N_4336,N_3973,N_3564);
or U4337 (N_4337,N_3800,N_3936);
and U4338 (N_4338,N_3941,N_3807);
or U4339 (N_4339,N_3592,N_3848);
and U4340 (N_4340,N_3749,N_3914);
nor U4341 (N_4341,N_3534,N_3536);
or U4342 (N_4342,N_3820,N_3731);
xor U4343 (N_4343,N_3673,N_3963);
xnor U4344 (N_4344,N_3542,N_3880);
or U4345 (N_4345,N_3825,N_3606);
nand U4346 (N_4346,N_3873,N_3631);
and U4347 (N_4347,N_3695,N_3898);
xor U4348 (N_4348,N_3632,N_3870);
nand U4349 (N_4349,N_3674,N_3842);
nor U4350 (N_4350,N_3982,N_3535);
nor U4351 (N_4351,N_3542,N_3642);
nand U4352 (N_4352,N_3678,N_3667);
nor U4353 (N_4353,N_3893,N_3768);
or U4354 (N_4354,N_3615,N_3544);
nand U4355 (N_4355,N_3721,N_3940);
nor U4356 (N_4356,N_3826,N_3990);
nor U4357 (N_4357,N_3839,N_3519);
or U4358 (N_4358,N_3608,N_3657);
nor U4359 (N_4359,N_3583,N_3719);
xor U4360 (N_4360,N_3649,N_3596);
nand U4361 (N_4361,N_3868,N_3963);
nand U4362 (N_4362,N_3966,N_3737);
xnor U4363 (N_4363,N_3806,N_3643);
or U4364 (N_4364,N_3832,N_3594);
nand U4365 (N_4365,N_3669,N_3924);
nand U4366 (N_4366,N_3709,N_3922);
or U4367 (N_4367,N_3891,N_3881);
xnor U4368 (N_4368,N_3527,N_3567);
and U4369 (N_4369,N_3905,N_3528);
and U4370 (N_4370,N_3840,N_3509);
nor U4371 (N_4371,N_3984,N_3628);
or U4372 (N_4372,N_3554,N_3995);
nand U4373 (N_4373,N_3978,N_3516);
nand U4374 (N_4374,N_3666,N_3534);
and U4375 (N_4375,N_3727,N_3581);
or U4376 (N_4376,N_3679,N_3663);
or U4377 (N_4377,N_3626,N_3814);
nand U4378 (N_4378,N_3986,N_3565);
xnor U4379 (N_4379,N_3840,N_3554);
or U4380 (N_4380,N_3731,N_3997);
nand U4381 (N_4381,N_3672,N_3831);
nor U4382 (N_4382,N_3533,N_3966);
nand U4383 (N_4383,N_3895,N_3767);
nor U4384 (N_4384,N_3595,N_3898);
xor U4385 (N_4385,N_3514,N_3655);
or U4386 (N_4386,N_3766,N_3932);
or U4387 (N_4387,N_3604,N_3745);
nand U4388 (N_4388,N_3763,N_3972);
xnor U4389 (N_4389,N_3506,N_3684);
nor U4390 (N_4390,N_3852,N_3878);
or U4391 (N_4391,N_3931,N_3808);
or U4392 (N_4392,N_3890,N_3790);
nor U4393 (N_4393,N_3764,N_3625);
or U4394 (N_4394,N_3597,N_3713);
or U4395 (N_4395,N_3791,N_3971);
and U4396 (N_4396,N_3973,N_3937);
or U4397 (N_4397,N_3897,N_3775);
xor U4398 (N_4398,N_3598,N_3799);
nand U4399 (N_4399,N_3721,N_3547);
xor U4400 (N_4400,N_3537,N_3731);
and U4401 (N_4401,N_3592,N_3850);
nand U4402 (N_4402,N_3859,N_3768);
and U4403 (N_4403,N_3782,N_3522);
xnor U4404 (N_4404,N_3772,N_3736);
and U4405 (N_4405,N_3578,N_3527);
nor U4406 (N_4406,N_3889,N_3620);
and U4407 (N_4407,N_3859,N_3790);
xor U4408 (N_4408,N_3527,N_3504);
and U4409 (N_4409,N_3908,N_3528);
xnor U4410 (N_4410,N_3719,N_3540);
xor U4411 (N_4411,N_3685,N_3552);
or U4412 (N_4412,N_3686,N_3569);
and U4413 (N_4413,N_3808,N_3621);
and U4414 (N_4414,N_3904,N_3785);
nand U4415 (N_4415,N_3771,N_3519);
and U4416 (N_4416,N_3538,N_3624);
nor U4417 (N_4417,N_3790,N_3834);
xor U4418 (N_4418,N_3847,N_3821);
nor U4419 (N_4419,N_3824,N_3640);
xnor U4420 (N_4420,N_3998,N_3606);
nand U4421 (N_4421,N_3723,N_3745);
or U4422 (N_4422,N_3654,N_3787);
nor U4423 (N_4423,N_3593,N_3888);
and U4424 (N_4424,N_3871,N_3805);
and U4425 (N_4425,N_3771,N_3754);
nor U4426 (N_4426,N_3804,N_3636);
nand U4427 (N_4427,N_3935,N_3893);
nand U4428 (N_4428,N_3987,N_3655);
xnor U4429 (N_4429,N_3901,N_3776);
or U4430 (N_4430,N_3752,N_3742);
or U4431 (N_4431,N_3768,N_3764);
or U4432 (N_4432,N_3844,N_3639);
nor U4433 (N_4433,N_3971,N_3628);
and U4434 (N_4434,N_3546,N_3732);
nand U4435 (N_4435,N_3847,N_3787);
or U4436 (N_4436,N_3997,N_3878);
nand U4437 (N_4437,N_3950,N_3611);
or U4438 (N_4438,N_3917,N_3642);
nor U4439 (N_4439,N_3968,N_3574);
and U4440 (N_4440,N_3777,N_3580);
nand U4441 (N_4441,N_3683,N_3988);
nor U4442 (N_4442,N_3506,N_3937);
nor U4443 (N_4443,N_3596,N_3977);
nand U4444 (N_4444,N_3972,N_3603);
xor U4445 (N_4445,N_3558,N_3779);
or U4446 (N_4446,N_3754,N_3877);
xor U4447 (N_4447,N_3824,N_3541);
and U4448 (N_4448,N_3654,N_3778);
nand U4449 (N_4449,N_3509,N_3827);
and U4450 (N_4450,N_3968,N_3748);
nand U4451 (N_4451,N_3801,N_3533);
or U4452 (N_4452,N_3917,N_3502);
or U4453 (N_4453,N_3534,N_3589);
and U4454 (N_4454,N_3883,N_3661);
or U4455 (N_4455,N_3604,N_3874);
and U4456 (N_4456,N_3698,N_3768);
nand U4457 (N_4457,N_3924,N_3613);
nand U4458 (N_4458,N_3615,N_3585);
nor U4459 (N_4459,N_3898,N_3531);
nor U4460 (N_4460,N_3655,N_3762);
nand U4461 (N_4461,N_3794,N_3962);
and U4462 (N_4462,N_3781,N_3965);
or U4463 (N_4463,N_3715,N_3838);
nand U4464 (N_4464,N_3803,N_3629);
xor U4465 (N_4465,N_3592,N_3626);
xnor U4466 (N_4466,N_3786,N_3674);
xnor U4467 (N_4467,N_3893,N_3679);
or U4468 (N_4468,N_3744,N_3723);
or U4469 (N_4469,N_3565,N_3946);
and U4470 (N_4470,N_3685,N_3982);
or U4471 (N_4471,N_3708,N_3906);
nand U4472 (N_4472,N_3726,N_3505);
or U4473 (N_4473,N_3834,N_3805);
nor U4474 (N_4474,N_3607,N_3695);
or U4475 (N_4475,N_3538,N_3660);
and U4476 (N_4476,N_3748,N_3985);
or U4477 (N_4477,N_3565,N_3601);
and U4478 (N_4478,N_3627,N_3654);
and U4479 (N_4479,N_3840,N_3978);
or U4480 (N_4480,N_3999,N_3781);
or U4481 (N_4481,N_3516,N_3637);
nand U4482 (N_4482,N_3678,N_3608);
or U4483 (N_4483,N_3669,N_3840);
nor U4484 (N_4484,N_3648,N_3656);
nor U4485 (N_4485,N_3546,N_3905);
or U4486 (N_4486,N_3999,N_3502);
nor U4487 (N_4487,N_3772,N_3871);
nor U4488 (N_4488,N_3787,N_3842);
or U4489 (N_4489,N_3528,N_3569);
nor U4490 (N_4490,N_3665,N_3863);
nand U4491 (N_4491,N_3786,N_3645);
nor U4492 (N_4492,N_3851,N_3731);
and U4493 (N_4493,N_3676,N_3739);
or U4494 (N_4494,N_3611,N_3699);
nand U4495 (N_4495,N_3747,N_3687);
or U4496 (N_4496,N_3695,N_3998);
and U4497 (N_4497,N_3981,N_3579);
or U4498 (N_4498,N_3899,N_3559);
or U4499 (N_4499,N_3537,N_3911);
and U4500 (N_4500,N_4276,N_4372);
or U4501 (N_4501,N_4034,N_4026);
and U4502 (N_4502,N_4214,N_4209);
or U4503 (N_4503,N_4153,N_4006);
xnor U4504 (N_4504,N_4407,N_4130);
or U4505 (N_4505,N_4322,N_4236);
or U4506 (N_4506,N_4356,N_4043);
xor U4507 (N_4507,N_4001,N_4299);
xnor U4508 (N_4508,N_4012,N_4492);
xnor U4509 (N_4509,N_4449,N_4250);
or U4510 (N_4510,N_4191,N_4154);
or U4511 (N_4511,N_4383,N_4336);
xor U4512 (N_4512,N_4171,N_4499);
nor U4513 (N_4513,N_4457,N_4406);
xnor U4514 (N_4514,N_4025,N_4329);
nand U4515 (N_4515,N_4038,N_4082);
nand U4516 (N_4516,N_4291,N_4042);
xor U4517 (N_4517,N_4089,N_4371);
or U4518 (N_4518,N_4119,N_4247);
xor U4519 (N_4519,N_4105,N_4382);
and U4520 (N_4520,N_4249,N_4233);
nand U4521 (N_4521,N_4439,N_4289);
nor U4522 (N_4522,N_4108,N_4101);
nand U4523 (N_4523,N_4128,N_4441);
nand U4524 (N_4524,N_4041,N_4493);
xnor U4525 (N_4525,N_4053,N_4084);
and U4526 (N_4526,N_4496,N_4150);
nor U4527 (N_4527,N_4312,N_4033);
or U4528 (N_4528,N_4062,N_4109);
nor U4529 (N_4529,N_4264,N_4267);
and U4530 (N_4530,N_4181,N_4176);
nor U4531 (N_4531,N_4324,N_4189);
xnor U4532 (N_4532,N_4460,N_4092);
and U4533 (N_4533,N_4319,N_4418);
nor U4534 (N_4534,N_4323,N_4468);
nand U4535 (N_4535,N_4132,N_4451);
nand U4536 (N_4536,N_4081,N_4126);
or U4537 (N_4537,N_4431,N_4438);
nor U4538 (N_4538,N_4384,N_4167);
or U4539 (N_4539,N_4207,N_4203);
nand U4540 (N_4540,N_4278,N_4024);
nand U4541 (N_4541,N_4156,N_4088);
nand U4542 (N_4542,N_4437,N_4058);
and U4543 (N_4543,N_4087,N_4432);
xnor U4544 (N_4544,N_4458,N_4477);
and U4545 (N_4545,N_4466,N_4339);
nand U4546 (N_4546,N_4271,N_4448);
and U4547 (N_4547,N_4196,N_4444);
nor U4548 (N_4548,N_4143,N_4136);
and U4549 (N_4549,N_4164,N_4253);
xor U4550 (N_4550,N_4282,N_4193);
xnor U4551 (N_4551,N_4030,N_4399);
or U4552 (N_4552,N_4137,N_4442);
nand U4553 (N_4553,N_4227,N_4148);
or U4554 (N_4554,N_4144,N_4133);
or U4555 (N_4555,N_4295,N_4281);
nand U4556 (N_4556,N_4293,N_4314);
or U4557 (N_4557,N_4182,N_4317);
nor U4558 (N_4558,N_4335,N_4435);
and U4559 (N_4559,N_4232,N_4313);
nor U4560 (N_4560,N_4474,N_4443);
and U4561 (N_4561,N_4478,N_4211);
nand U4562 (N_4562,N_4301,N_4297);
and U4563 (N_4563,N_4219,N_4420);
nand U4564 (N_4564,N_4408,N_4085);
nand U4565 (N_4565,N_4117,N_4343);
nor U4566 (N_4566,N_4370,N_4131);
or U4567 (N_4567,N_4465,N_4255);
nor U4568 (N_4568,N_4402,N_4020);
xor U4569 (N_4569,N_4160,N_4455);
xor U4570 (N_4570,N_4254,N_4275);
or U4571 (N_4571,N_4142,N_4059);
or U4572 (N_4572,N_4036,N_4202);
and U4573 (N_4573,N_4204,N_4424);
or U4574 (N_4574,N_4332,N_4423);
nor U4575 (N_4575,N_4321,N_4390);
or U4576 (N_4576,N_4489,N_4450);
xor U4577 (N_4577,N_4306,N_4111);
xor U4578 (N_4578,N_4260,N_4225);
nand U4579 (N_4579,N_4309,N_4248);
nor U4580 (N_4580,N_4422,N_4378);
xor U4581 (N_4581,N_4057,N_4086);
and U4582 (N_4582,N_4228,N_4320);
xnor U4583 (N_4583,N_4326,N_4467);
nand U4584 (N_4584,N_4213,N_4364);
xor U4585 (N_4585,N_4123,N_4073);
xor U4586 (N_4586,N_4099,N_4484);
nand U4587 (N_4587,N_4486,N_4425);
nand U4588 (N_4588,N_4127,N_4051);
nand U4589 (N_4589,N_4464,N_4075);
or U4590 (N_4590,N_4284,N_4374);
and U4591 (N_4591,N_4031,N_4004);
nor U4592 (N_4592,N_4064,N_4269);
nor U4593 (N_4593,N_4338,N_4362);
nor U4594 (N_4594,N_4386,N_4172);
and U4595 (N_4595,N_4310,N_4060);
nor U4596 (N_4596,N_4273,N_4434);
or U4597 (N_4597,N_4162,N_4195);
or U4598 (N_4598,N_4433,N_4405);
nand U4599 (N_4599,N_4106,N_4185);
xor U4600 (N_4600,N_4107,N_4461);
nor U4601 (N_4601,N_4019,N_4256);
nand U4602 (N_4602,N_4151,N_4440);
nor U4603 (N_4603,N_4049,N_4165);
xor U4604 (N_4604,N_4363,N_4381);
or U4605 (N_4605,N_4394,N_4018);
nand U4606 (N_4606,N_4265,N_4471);
or U4607 (N_4607,N_4333,N_4459);
and U4608 (N_4608,N_4222,N_4104);
nand U4609 (N_4609,N_4199,N_4341);
or U4610 (N_4610,N_4452,N_4045);
or U4611 (N_4611,N_4277,N_4221);
nor U4612 (N_4612,N_4414,N_4140);
or U4613 (N_4613,N_4094,N_4472);
nand U4614 (N_4614,N_4490,N_4218);
nand U4615 (N_4615,N_4375,N_4129);
or U4616 (N_4616,N_4354,N_4103);
nand U4617 (N_4617,N_4463,N_4470);
or U4618 (N_4618,N_4047,N_4013);
nand U4619 (N_4619,N_4421,N_4102);
or U4620 (N_4620,N_4358,N_4266);
and U4621 (N_4621,N_4274,N_4331);
nand U4622 (N_4622,N_4398,N_4246);
and U4623 (N_4623,N_4392,N_4345);
nor U4624 (N_4624,N_4304,N_4428);
nand U4625 (N_4625,N_4240,N_4308);
and U4626 (N_4626,N_4122,N_4359);
and U4627 (N_4627,N_4046,N_4252);
xor U4628 (N_4628,N_4445,N_4328);
and U4629 (N_4629,N_4367,N_4070);
nor U4630 (N_4630,N_4279,N_4397);
nand U4631 (N_4631,N_4066,N_4347);
nand U4632 (N_4632,N_4003,N_4366);
xnor U4633 (N_4633,N_4145,N_4068);
and U4634 (N_4634,N_4487,N_4009);
nand U4635 (N_4635,N_4355,N_4453);
or U4636 (N_4636,N_4417,N_4174);
xor U4637 (N_4637,N_4226,N_4159);
nand U4638 (N_4638,N_4208,N_4014);
xnor U4639 (N_4639,N_4005,N_4237);
or U4640 (N_4640,N_4411,N_4169);
and U4641 (N_4641,N_4327,N_4404);
nor U4642 (N_4642,N_4395,N_4037);
xnor U4643 (N_4643,N_4098,N_4010);
and U4644 (N_4644,N_4179,N_4121);
and U4645 (N_4645,N_4180,N_4325);
and U4646 (N_4646,N_4419,N_4290);
or U4647 (N_4647,N_4100,N_4303);
nor U4648 (N_4648,N_4334,N_4488);
nor U4649 (N_4649,N_4285,N_4192);
nand U4650 (N_4650,N_4251,N_4065);
or U4651 (N_4651,N_4380,N_4044);
or U4652 (N_4652,N_4178,N_4096);
and U4653 (N_4653,N_4139,N_4436);
nor U4654 (N_4654,N_4258,N_4050);
or U4655 (N_4655,N_4166,N_4230);
or U4656 (N_4656,N_4239,N_4482);
and U4657 (N_4657,N_4002,N_4361);
and U4658 (N_4658,N_4353,N_4263);
xor U4659 (N_4659,N_4015,N_4346);
or U4660 (N_4660,N_4287,N_4124);
xor U4661 (N_4661,N_4023,N_4078);
nand U4662 (N_4662,N_4280,N_4305);
xnor U4663 (N_4663,N_4352,N_4022);
and U4664 (N_4664,N_4112,N_4152);
and U4665 (N_4665,N_4369,N_4307);
nand U4666 (N_4666,N_4495,N_4373);
or U4667 (N_4667,N_4120,N_4365);
nor U4668 (N_4668,N_4074,N_4091);
nand U4669 (N_4669,N_4157,N_4217);
and U4670 (N_4670,N_4077,N_4000);
and U4671 (N_4671,N_4447,N_4187);
nor U4672 (N_4672,N_4083,N_4008);
or U4673 (N_4673,N_4377,N_4200);
xnor U4674 (N_4674,N_4268,N_4235);
or U4675 (N_4675,N_4095,N_4243);
and U4676 (N_4676,N_4376,N_4387);
or U4677 (N_4677,N_4286,N_4224);
xor U4678 (N_4678,N_4048,N_4028);
xnor U4679 (N_4679,N_4300,N_4396);
and U4680 (N_4680,N_4011,N_4498);
nand U4681 (N_4681,N_4456,N_4186);
and U4682 (N_4682,N_4283,N_4462);
and U4683 (N_4683,N_4175,N_4400);
and U4684 (N_4684,N_4016,N_4294);
nand U4685 (N_4685,N_4097,N_4368);
nand U4686 (N_4686,N_4212,N_4412);
xor U4687 (N_4687,N_4481,N_4298);
nand U4688 (N_4688,N_4215,N_4446);
and U4689 (N_4689,N_4302,N_4110);
or U4690 (N_4690,N_4205,N_4125);
nand U4691 (N_4691,N_4072,N_4426);
nand U4692 (N_4692,N_4007,N_4344);
nor U4693 (N_4693,N_4076,N_4296);
and U4694 (N_4694,N_4403,N_4027);
nor U4695 (N_4695,N_4393,N_4491);
xor U4696 (N_4696,N_4223,N_4055);
xnor U4697 (N_4697,N_4259,N_4071);
and U4698 (N_4698,N_4454,N_4118);
or U4699 (N_4699,N_4430,N_4035);
xnor U4700 (N_4700,N_4311,N_4183);
or U4701 (N_4701,N_4184,N_4210);
and U4702 (N_4702,N_4155,N_4138);
nand U4703 (N_4703,N_4245,N_4229);
or U4704 (N_4704,N_4113,N_4272);
and U4705 (N_4705,N_4429,N_4134);
nor U4706 (N_4706,N_4340,N_4146);
nand U4707 (N_4707,N_4158,N_4234);
nand U4708 (N_4708,N_4473,N_4318);
nor U4709 (N_4709,N_4188,N_4220);
xor U4710 (N_4710,N_4337,N_4261);
and U4711 (N_4711,N_4017,N_4357);
nand U4712 (N_4712,N_4244,N_4497);
and U4713 (N_4713,N_4093,N_4168);
xor U4714 (N_4714,N_4040,N_4116);
nand U4715 (N_4715,N_4054,N_4315);
nor U4716 (N_4716,N_4316,N_4475);
nor U4717 (N_4717,N_4479,N_4348);
xnor U4718 (N_4718,N_4173,N_4231);
xor U4719 (N_4719,N_4201,N_4052);
nor U4720 (N_4720,N_4270,N_4135);
or U4721 (N_4721,N_4114,N_4494);
xor U4722 (N_4722,N_4389,N_4238);
xor U4723 (N_4723,N_4021,N_4351);
nand U4724 (N_4724,N_4039,N_4350);
nor U4725 (N_4725,N_4288,N_4469);
or U4726 (N_4726,N_4385,N_4360);
xnor U4727 (N_4727,N_4416,N_4480);
or U4728 (N_4728,N_4410,N_4067);
and U4729 (N_4729,N_4485,N_4197);
or U4730 (N_4730,N_4415,N_4198);
nand U4731 (N_4731,N_4483,N_4342);
and U4732 (N_4732,N_4194,N_4262);
nand U4733 (N_4733,N_4163,N_4061);
nor U4734 (N_4734,N_4149,N_4079);
xor U4735 (N_4735,N_4056,N_4069);
nand U4736 (N_4736,N_4391,N_4206);
nand U4737 (N_4737,N_4090,N_4257);
xnor U4738 (N_4738,N_4401,N_4063);
or U4739 (N_4739,N_4292,N_4177);
or U4740 (N_4740,N_4409,N_4029);
nor U4741 (N_4741,N_4427,N_4147);
xnor U4742 (N_4742,N_4115,N_4349);
nand U4743 (N_4743,N_4242,N_4388);
or U4744 (N_4744,N_4476,N_4141);
and U4745 (N_4745,N_4190,N_4080);
and U4746 (N_4746,N_4161,N_4413);
and U4747 (N_4747,N_4216,N_4241);
and U4748 (N_4748,N_4379,N_4170);
xnor U4749 (N_4749,N_4032,N_4330);
xor U4750 (N_4750,N_4308,N_4062);
and U4751 (N_4751,N_4419,N_4451);
and U4752 (N_4752,N_4127,N_4178);
or U4753 (N_4753,N_4209,N_4484);
or U4754 (N_4754,N_4305,N_4299);
nand U4755 (N_4755,N_4150,N_4057);
nand U4756 (N_4756,N_4131,N_4338);
xnor U4757 (N_4757,N_4412,N_4369);
and U4758 (N_4758,N_4261,N_4232);
and U4759 (N_4759,N_4226,N_4068);
nor U4760 (N_4760,N_4452,N_4446);
nor U4761 (N_4761,N_4147,N_4075);
nor U4762 (N_4762,N_4228,N_4353);
nor U4763 (N_4763,N_4264,N_4033);
and U4764 (N_4764,N_4295,N_4103);
or U4765 (N_4765,N_4171,N_4196);
or U4766 (N_4766,N_4498,N_4083);
nor U4767 (N_4767,N_4242,N_4466);
nand U4768 (N_4768,N_4232,N_4015);
or U4769 (N_4769,N_4044,N_4439);
xor U4770 (N_4770,N_4460,N_4242);
xor U4771 (N_4771,N_4103,N_4008);
or U4772 (N_4772,N_4443,N_4139);
nand U4773 (N_4773,N_4424,N_4056);
nor U4774 (N_4774,N_4423,N_4032);
xnor U4775 (N_4775,N_4285,N_4202);
nand U4776 (N_4776,N_4074,N_4077);
nand U4777 (N_4777,N_4325,N_4140);
and U4778 (N_4778,N_4141,N_4043);
xnor U4779 (N_4779,N_4364,N_4404);
xnor U4780 (N_4780,N_4222,N_4206);
or U4781 (N_4781,N_4404,N_4029);
xor U4782 (N_4782,N_4318,N_4447);
or U4783 (N_4783,N_4497,N_4456);
nor U4784 (N_4784,N_4046,N_4126);
xnor U4785 (N_4785,N_4177,N_4337);
nand U4786 (N_4786,N_4167,N_4059);
or U4787 (N_4787,N_4379,N_4446);
xnor U4788 (N_4788,N_4069,N_4291);
nor U4789 (N_4789,N_4454,N_4406);
xnor U4790 (N_4790,N_4314,N_4470);
nor U4791 (N_4791,N_4212,N_4005);
nor U4792 (N_4792,N_4404,N_4427);
nand U4793 (N_4793,N_4329,N_4161);
nor U4794 (N_4794,N_4019,N_4370);
nand U4795 (N_4795,N_4368,N_4149);
or U4796 (N_4796,N_4465,N_4263);
nor U4797 (N_4797,N_4062,N_4497);
xnor U4798 (N_4798,N_4471,N_4153);
nor U4799 (N_4799,N_4026,N_4110);
nand U4800 (N_4800,N_4102,N_4076);
xor U4801 (N_4801,N_4240,N_4325);
and U4802 (N_4802,N_4365,N_4211);
xor U4803 (N_4803,N_4398,N_4030);
and U4804 (N_4804,N_4191,N_4178);
or U4805 (N_4805,N_4225,N_4035);
xnor U4806 (N_4806,N_4150,N_4002);
or U4807 (N_4807,N_4124,N_4492);
nor U4808 (N_4808,N_4491,N_4287);
and U4809 (N_4809,N_4306,N_4206);
and U4810 (N_4810,N_4332,N_4066);
nor U4811 (N_4811,N_4167,N_4410);
nand U4812 (N_4812,N_4450,N_4371);
nand U4813 (N_4813,N_4339,N_4052);
nor U4814 (N_4814,N_4221,N_4231);
nor U4815 (N_4815,N_4380,N_4397);
nand U4816 (N_4816,N_4171,N_4140);
xnor U4817 (N_4817,N_4287,N_4263);
xor U4818 (N_4818,N_4143,N_4387);
or U4819 (N_4819,N_4154,N_4297);
nor U4820 (N_4820,N_4099,N_4234);
and U4821 (N_4821,N_4106,N_4225);
and U4822 (N_4822,N_4167,N_4312);
or U4823 (N_4823,N_4438,N_4016);
xor U4824 (N_4824,N_4253,N_4349);
and U4825 (N_4825,N_4325,N_4225);
and U4826 (N_4826,N_4496,N_4102);
xnor U4827 (N_4827,N_4358,N_4180);
nand U4828 (N_4828,N_4447,N_4026);
nor U4829 (N_4829,N_4497,N_4276);
xnor U4830 (N_4830,N_4111,N_4084);
nor U4831 (N_4831,N_4035,N_4392);
nand U4832 (N_4832,N_4373,N_4053);
nor U4833 (N_4833,N_4375,N_4494);
nor U4834 (N_4834,N_4251,N_4213);
and U4835 (N_4835,N_4160,N_4177);
nor U4836 (N_4836,N_4063,N_4339);
nor U4837 (N_4837,N_4239,N_4268);
xor U4838 (N_4838,N_4147,N_4215);
nand U4839 (N_4839,N_4444,N_4046);
nand U4840 (N_4840,N_4488,N_4395);
nor U4841 (N_4841,N_4057,N_4254);
nor U4842 (N_4842,N_4008,N_4427);
xnor U4843 (N_4843,N_4171,N_4247);
and U4844 (N_4844,N_4464,N_4170);
or U4845 (N_4845,N_4041,N_4117);
or U4846 (N_4846,N_4394,N_4412);
nor U4847 (N_4847,N_4258,N_4273);
nand U4848 (N_4848,N_4303,N_4402);
xor U4849 (N_4849,N_4483,N_4117);
xor U4850 (N_4850,N_4217,N_4495);
nor U4851 (N_4851,N_4397,N_4270);
xnor U4852 (N_4852,N_4345,N_4096);
and U4853 (N_4853,N_4323,N_4032);
nor U4854 (N_4854,N_4017,N_4363);
nor U4855 (N_4855,N_4037,N_4281);
xnor U4856 (N_4856,N_4417,N_4224);
nor U4857 (N_4857,N_4239,N_4058);
and U4858 (N_4858,N_4086,N_4024);
nand U4859 (N_4859,N_4305,N_4497);
nand U4860 (N_4860,N_4221,N_4160);
and U4861 (N_4861,N_4159,N_4198);
xor U4862 (N_4862,N_4072,N_4086);
and U4863 (N_4863,N_4246,N_4458);
xor U4864 (N_4864,N_4130,N_4037);
or U4865 (N_4865,N_4100,N_4278);
and U4866 (N_4866,N_4242,N_4172);
nand U4867 (N_4867,N_4095,N_4431);
nand U4868 (N_4868,N_4488,N_4356);
nand U4869 (N_4869,N_4222,N_4194);
xnor U4870 (N_4870,N_4031,N_4012);
and U4871 (N_4871,N_4208,N_4094);
and U4872 (N_4872,N_4272,N_4216);
nand U4873 (N_4873,N_4205,N_4346);
or U4874 (N_4874,N_4351,N_4428);
nand U4875 (N_4875,N_4064,N_4053);
and U4876 (N_4876,N_4431,N_4031);
nand U4877 (N_4877,N_4311,N_4356);
and U4878 (N_4878,N_4006,N_4160);
nand U4879 (N_4879,N_4076,N_4124);
or U4880 (N_4880,N_4070,N_4323);
nand U4881 (N_4881,N_4169,N_4230);
nor U4882 (N_4882,N_4325,N_4428);
or U4883 (N_4883,N_4041,N_4367);
and U4884 (N_4884,N_4253,N_4418);
xor U4885 (N_4885,N_4045,N_4342);
and U4886 (N_4886,N_4487,N_4395);
nand U4887 (N_4887,N_4050,N_4006);
nor U4888 (N_4888,N_4299,N_4371);
nand U4889 (N_4889,N_4258,N_4303);
nor U4890 (N_4890,N_4439,N_4485);
or U4891 (N_4891,N_4020,N_4288);
nand U4892 (N_4892,N_4104,N_4101);
xnor U4893 (N_4893,N_4328,N_4195);
and U4894 (N_4894,N_4285,N_4436);
xnor U4895 (N_4895,N_4354,N_4413);
nor U4896 (N_4896,N_4217,N_4427);
and U4897 (N_4897,N_4490,N_4458);
xnor U4898 (N_4898,N_4274,N_4288);
xor U4899 (N_4899,N_4252,N_4204);
or U4900 (N_4900,N_4010,N_4071);
nor U4901 (N_4901,N_4148,N_4478);
or U4902 (N_4902,N_4464,N_4496);
nor U4903 (N_4903,N_4227,N_4136);
nor U4904 (N_4904,N_4360,N_4139);
xnor U4905 (N_4905,N_4400,N_4264);
xor U4906 (N_4906,N_4160,N_4185);
and U4907 (N_4907,N_4433,N_4220);
and U4908 (N_4908,N_4000,N_4030);
or U4909 (N_4909,N_4343,N_4366);
nand U4910 (N_4910,N_4203,N_4470);
nor U4911 (N_4911,N_4074,N_4102);
or U4912 (N_4912,N_4440,N_4083);
xnor U4913 (N_4913,N_4155,N_4026);
and U4914 (N_4914,N_4266,N_4330);
and U4915 (N_4915,N_4443,N_4466);
or U4916 (N_4916,N_4115,N_4169);
and U4917 (N_4917,N_4217,N_4431);
or U4918 (N_4918,N_4201,N_4469);
nand U4919 (N_4919,N_4113,N_4069);
and U4920 (N_4920,N_4184,N_4408);
nand U4921 (N_4921,N_4187,N_4183);
xor U4922 (N_4922,N_4249,N_4217);
and U4923 (N_4923,N_4090,N_4041);
or U4924 (N_4924,N_4140,N_4202);
xor U4925 (N_4925,N_4346,N_4120);
or U4926 (N_4926,N_4371,N_4127);
or U4927 (N_4927,N_4338,N_4159);
nor U4928 (N_4928,N_4167,N_4381);
nand U4929 (N_4929,N_4010,N_4162);
nor U4930 (N_4930,N_4267,N_4433);
xnor U4931 (N_4931,N_4048,N_4290);
nor U4932 (N_4932,N_4264,N_4362);
nand U4933 (N_4933,N_4305,N_4005);
nand U4934 (N_4934,N_4339,N_4343);
nor U4935 (N_4935,N_4129,N_4328);
nor U4936 (N_4936,N_4057,N_4143);
or U4937 (N_4937,N_4149,N_4182);
and U4938 (N_4938,N_4321,N_4147);
nor U4939 (N_4939,N_4143,N_4157);
nand U4940 (N_4940,N_4338,N_4071);
nand U4941 (N_4941,N_4200,N_4323);
nand U4942 (N_4942,N_4353,N_4279);
or U4943 (N_4943,N_4198,N_4101);
nand U4944 (N_4944,N_4060,N_4026);
or U4945 (N_4945,N_4400,N_4367);
nand U4946 (N_4946,N_4134,N_4448);
nand U4947 (N_4947,N_4080,N_4059);
xnor U4948 (N_4948,N_4075,N_4259);
and U4949 (N_4949,N_4154,N_4204);
xnor U4950 (N_4950,N_4187,N_4321);
and U4951 (N_4951,N_4345,N_4123);
nand U4952 (N_4952,N_4065,N_4374);
nand U4953 (N_4953,N_4419,N_4194);
nor U4954 (N_4954,N_4022,N_4030);
or U4955 (N_4955,N_4397,N_4030);
and U4956 (N_4956,N_4040,N_4462);
nor U4957 (N_4957,N_4435,N_4142);
and U4958 (N_4958,N_4097,N_4290);
and U4959 (N_4959,N_4183,N_4091);
nor U4960 (N_4960,N_4352,N_4116);
or U4961 (N_4961,N_4251,N_4465);
xnor U4962 (N_4962,N_4312,N_4377);
nor U4963 (N_4963,N_4361,N_4444);
nand U4964 (N_4964,N_4055,N_4485);
nand U4965 (N_4965,N_4267,N_4139);
or U4966 (N_4966,N_4151,N_4451);
and U4967 (N_4967,N_4190,N_4341);
or U4968 (N_4968,N_4384,N_4135);
xnor U4969 (N_4969,N_4025,N_4482);
xnor U4970 (N_4970,N_4097,N_4231);
xor U4971 (N_4971,N_4036,N_4025);
and U4972 (N_4972,N_4200,N_4003);
nand U4973 (N_4973,N_4192,N_4489);
or U4974 (N_4974,N_4249,N_4486);
xor U4975 (N_4975,N_4438,N_4395);
or U4976 (N_4976,N_4156,N_4000);
xor U4977 (N_4977,N_4015,N_4080);
nor U4978 (N_4978,N_4265,N_4028);
and U4979 (N_4979,N_4481,N_4268);
and U4980 (N_4980,N_4248,N_4041);
or U4981 (N_4981,N_4431,N_4054);
nand U4982 (N_4982,N_4204,N_4244);
nor U4983 (N_4983,N_4221,N_4120);
xor U4984 (N_4984,N_4403,N_4209);
or U4985 (N_4985,N_4399,N_4184);
or U4986 (N_4986,N_4340,N_4039);
and U4987 (N_4987,N_4448,N_4431);
xnor U4988 (N_4988,N_4277,N_4326);
nand U4989 (N_4989,N_4350,N_4010);
xor U4990 (N_4990,N_4366,N_4026);
nor U4991 (N_4991,N_4394,N_4320);
xor U4992 (N_4992,N_4477,N_4137);
xor U4993 (N_4993,N_4037,N_4017);
xnor U4994 (N_4994,N_4102,N_4142);
nand U4995 (N_4995,N_4136,N_4062);
xor U4996 (N_4996,N_4421,N_4205);
or U4997 (N_4997,N_4116,N_4154);
and U4998 (N_4998,N_4130,N_4043);
nor U4999 (N_4999,N_4187,N_4034);
nand UO_0 (O_0,N_4552,N_4750);
nor UO_1 (O_1,N_4861,N_4948);
and UO_2 (O_2,N_4614,N_4915);
xor UO_3 (O_3,N_4865,N_4926);
xor UO_4 (O_4,N_4601,N_4687);
xnor UO_5 (O_5,N_4514,N_4918);
nand UO_6 (O_6,N_4658,N_4647);
and UO_7 (O_7,N_4795,N_4678);
nand UO_8 (O_8,N_4889,N_4866);
and UO_9 (O_9,N_4857,N_4877);
or UO_10 (O_10,N_4632,N_4810);
or UO_11 (O_11,N_4569,N_4923);
xor UO_12 (O_12,N_4711,N_4990);
nor UO_13 (O_13,N_4782,N_4738);
or UO_14 (O_14,N_4622,N_4972);
xor UO_15 (O_15,N_4920,N_4526);
nand UO_16 (O_16,N_4847,N_4586);
nor UO_17 (O_17,N_4595,N_4987);
xor UO_18 (O_18,N_4872,N_4502);
and UO_19 (O_19,N_4769,N_4742);
xor UO_20 (O_20,N_4648,N_4544);
or UO_21 (O_21,N_4639,N_4779);
or UO_22 (O_22,N_4954,N_4524);
xnor UO_23 (O_23,N_4612,N_4659);
xor UO_24 (O_24,N_4627,N_4628);
nand UO_25 (O_25,N_4697,N_4831);
xor UO_26 (O_26,N_4976,N_4559);
or UO_27 (O_27,N_4860,N_4778);
xnor UO_28 (O_28,N_4517,N_4969);
nor UO_29 (O_29,N_4820,N_4975);
nand UO_30 (O_30,N_4608,N_4638);
xor UO_31 (O_31,N_4564,N_4567);
nor UO_32 (O_32,N_4518,N_4940);
nand UO_33 (O_33,N_4930,N_4934);
nor UO_34 (O_34,N_4837,N_4688);
and UO_35 (O_35,N_4723,N_4533);
and UO_36 (O_36,N_4571,N_4618);
and UO_37 (O_37,N_4727,N_4830);
or UO_38 (O_38,N_4650,N_4551);
nor UO_39 (O_39,N_4853,N_4507);
nand UO_40 (O_40,N_4996,N_4561);
nor UO_41 (O_41,N_4719,N_4501);
and UO_42 (O_42,N_4675,N_4864);
nand UO_43 (O_43,N_4785,N_4797);
nor UO_44 (O_44,N_4731,N_4753);
xnor UO_45 (O_45,N_4717,N_4720);
or UO_46 (O_46,N_4671,N_4910);
nand UO_47 (O_47,N_4921,N_4806);
or UO_48 (O_48,N_4539,N_4899);
nor UO_49 (O_49,N_4781,N_4819);
and UO_50 (O_50,N_4832,N_4757);
xor UO_51 (O_51,N_4566,N_4884);
nand UO_52 (O_52,N_4540,N_4991);
xnor UO_53 (O_53,N_4621,N_4749);
nand UO_54 (O_54,N_4689,N_4662);
nand UO_55 (O_55,N_4525,N_4786);
nand UO_56 (O_56,N_4748,N_4611);
xnor UO_57 (O_57,N_4663,N_4791);
nand UO_58 (O_58,N_4962,N_4609);
and UO_59 (O_59,N_4883,N_4610);
nor UO_60 (O_60,N_4634,N_4796);
xnor UO_61 (O_61,N_4712,N_4503);
and UO_62 (O_62,N_4968,N_4955);
xnor UO_63 (O_63,N_4716,N_4957);
nor UO_64 (O_64,N_4766,N_4735);
or UO_65 (O_65,N_4936,N_4585);
nor UO_66 (O_66,N_4905,N_4841);
nor UO_67 (O_67,N_4932,N_4803);
nand UO_68 (O_68,N_4986,N_4509);
nand UO_69 (O_69,N_4730,N_4670);
nor UO_70 (O_70,N_4937,N_4762);
xnor UO_71 (O_71,N_4682,N_4994);
nand UO_72 (O_72,N_4535,N_4505);
and UO_73 (O_73,N_4553,N_4928);
nand UO_74 (O_74,N_4840,N_4655);
nand UO_75 (O_75,N_4563,N_4652);
or UO_76 (O_76,N_4939,N_4677);
nand UO_77 (O_77,N_4802,N_4759);
nor UO_78 (O_78,N_4617,N_4916);
or UO_79 (O_79,N_4699,N_4992);
nor UO_80 (O_80,N_4624,N_4587);
or UO_81 (O_81,N_4836,N_4822);
xor UO_82 (O_82,N_4772,N_4863);
and UO_83 (O_83,N_4683,N_4734);
or UO_84 (O_84,N_4900,N_4947);
nor UO_85 (O_85,N_4842,N_4744);
xor UO_86 (O_86,N_4834,N_4755);
nand UO_87 (O_87,N_4686,N_4593);
nor UO_88 (O_88,N_4620,N_4728);
nand UO_89 (O_89,N_4511,N_4747);
or UO_90 (O_90,N_4546,N_4823);
nor UO_91 (O_91,N_4589,N_4851);
nor UO_92 (O_92,N_4956,N_4927);
or UO_93 (O_93,N_4799,N_4530);
nor UO_94 (O_94,N_4824,N_4907);
and UO_95 (O_95,N_4952,N_4839);
nor UO_96 (O_96,N_4971,N_4945);
and UO_97 (O_97,N_4702,N_4560);
and UO_98 (O_98,N_4902,N_4718);
and UO_99 (O_99,N_4654,N_4911);
nand UO_100 (O_100,N_4653,N_4629);
nand UO_101 (O_101,N_4868,N_4771);
nand UO_102 (O_102,N_4674,N_4846);
nand UO_103 (O_103,N_4619,N_4873);
xor UO_104 (O_104,N_4685,N_4953);
and UO_105 (O_105,N_4856,N_4970);
nor UO_106 (O_106,N_4512,N_4967);
nand UO_107 (O_107,N_4713,N_4515);
and UO_108 (O_108,N_4903,N_4754);
nor UO_109 (O_109,N_4741,N_4579);
xnor UO_110 (O_110,N_4554,N_4510);
or UO_111 (O_111,N_4995,N_4989);
or UO_112 (O_112,N_4732,N_4974);
nand UO_113 (O_113,N_4850,N_4809);
and UO_114 (O_114,N_4878,N_4684);
nand UO_115 (O_115,N_4607,N_4740);
and UO_116 (O_116,N_4758,N_4642);
xnor UO_117 (O_117,N_4545,N_4881);
or UO_118 (O_118,N_4793,N_4931);
nor UO_119 (O_119,N_4774,N_4672);
nand UO_120 (O_120,N_4736,N_4644);
and UO_121 (O_121,N_4789,N_4690);
nor UO_122 (O_122,N_4603,N_4529);
xnor UO_123 (O_123,N_4984,N_4739);
and UO_124 (O_124,N_4929,N_4679);
and UO_125 (O_125,N_4555,N_4615);
nand UO_126 (O_126,N_4844,N_4998);
xor UO_127 (O_127,N_4891,N_4714);
or UO_128 (O_128,N_4890,N_4594);
nor UO_129 (O_129,N_4909,N_4722);
and UO_130 (O_130,N_4788,N_4604);
or UO_131 (O_131,N_4737,N_4807);
nor UO_132 (O_132,N_4917,N_4602);
xor UO_133 (O_133,N_4641,N_4549);
and UO_134 (O_134,N_4982,N_4775);
nand UO_135 (O_135,N_4800,N_4828);
xnor UO_136 (O_136,N_4838,N_4950);
and UO_137 (O_137,N_4924,N_4855);
or UO_138 (O_138,N_4783,N_4997);
nor UO_139 (O_139,N_4710,N_4827);
nand UO_140 (O_140,N_4849,N_4949);
nor UO_141 (O_141,N_4854,N_4763);
xor UO_142 (O_142,N_4888,N_4764);
xnor UO_143 (O_143,N_4547,N_4565);
xor UO_144 (O_144,N_4752,N_4983);
nand UO_145 (O_145,N_4943,N_4724);
nor UO_146 (O_146,N_4558,N_4574);
or UO_147 (O_147,N_4651,N_4625);
nor UO_148 (O_148,N_4506,N_4582);
and UO_149 (O_149,N_4787,N_4816);
xor UO_150 (O_150,N_4596,N_4695);
nor UO_151 (O_151,N_4798,N_4813);
nand UO_152 (O_152,N_4729,N_4904);
nand UO_153 (O_153,N_4829,N_4590);
or UO_154 (O_154,N_4532,N_4623);
or UO_155 (O_155,N_4528,N_4973);
nand UO_156 (O_156,N_4550,N_4726);
nor UO_157 (O_157,N_4696,N_4668);
and UO_158 (O_158,N_4906,N_4874);
or UO_159 (O_159,N_4692,N_4977);
nor UO_160 (O_160,N_4500,N_4848);
nor UO_161 (O_161,N_4698,N_4951);
and UO_162 (O_162,N_4591,N_4879);
or UO_163 (O_163,N_4541,N_4808);
or UO_164 (O_164,N_4805,N_4616);
xor UO_165 (O_165,N_4988,N_4573);
nand UO_166 (O_166,N_4568,N_4527);
and UO_167 (O_167,N_4667,N_4875);
or UO_168 (O_168,N_4600,N_4701);
and UO_169 (O_169,N_4656,N_4770);
or UO_170 (O_170,N_4703,N_4978);
or UO_171 (O_171,N_4531,N_4966);
and UO_172 (O_172,N_4913,N_4681);
nand UO_173 (O_173,N_4583,N_4876);
nor UO_174 (O_174,N_4598,N_4592);
xnor UO_175 (O_175,N_4942,N_4633);
xor UO_176 (O_176,N_4635,N_4880);
and UO_177 (O_177,N_4584,N_4818);
and UO_178 (O_178,N_4522,N_4745);
nand UO_179 (O_179,N_4790,N_4534);
and UO_180 (O_180,N_4985,N_4933);
or UO_181 (O_181,N_4768,N_4760);
xnor UO_182 (O_182,N_4925,N_4811);
xor UO_183 (O_183,N_4673,N_4508);
nand UO_184 (O_184,N_4756,N_4706);
and UO_185 (O_185,N_4557,N_4513);
or UO_186 (O_186,N_4751,N_4645);
nand UO_187 (O_187,N_4961,N_4665);
or UO_188 (O_188,N_4680,N_4938);
nand UO_189 (O_189,N_4538,N_4825);
nand UO_190 (O_190,N_4895,N_4519);
or UO_191 (O_191,N_4999,N_4700);
nor UO_192 (O_192,N_4892,N_4912);
and UO_193 (O_193,N_4817,N_4901);
xor UO_194 (O_194,N_4858,N_4649);
and UO_195 (O_195,N_4520,N_4777);
and UO_196 (O_196,N_4504,N_4814);
nand UO_197 (O_197,N_4708,N_4993);
nand UO_198 (O_198,N_4709,N_4542);
nand UO_199 (O_199,N_4852,N_4588);
and UO_200 (O_200,N_4661,N_4963);
xnor UO_201 (O_201,N_4669,N_4543);
nor UO_202 (O_202,N_4765,N_4867);
or UO_203 (O_203,N_4580,N_4761);
or UO_204 (O_204,N_4743,N_4922);
xnor UO_205 (O_205,N_4792,N_4964);
or UO_206 (O_206,N_4919,N_4715);
or UO_207 (O_207,N_4523,N_4887);
nand UO_208 (O_208,N_4958,N_4577);
nor UO_209 (O_209,N_4578,N_4606);
nand UO_210 (O_210,N_4637,N_4660);
or UO_211 (O_211,N_4897,N_4664);
or UO_212 (O_212,N_4960,N_4636);
nand UO_213 (O_213,N_4576,N_4871);
nand UO_214 (O_214,N_4640,N_4767);
nand UO_215 (O_215,N_4812,N_4893);
and UO_216 (O_216,N_4666,N_4801);
or UO_217 (O_217,N_4821,N_4885);
nand UO_218 (O_218,N_4980,N_4597);
and UO_219 (O_219,N_4894,N_4575);
or UO_220 (O_220,N_4944,N_4599);
or UO_221 (O_221,N_4914,N_4935);
and UO_222 (O_222,N_4862,N_4572);
and UO_223 (O_223,N_4843,N_4780);
xor UO_224 (O_224,N_4704,N_4613);
xnor UO_225 (O_225,N_4725,N_4859);
nand UO_226 (O_226,N_4721,N_4794);
and UO_227 (O_227,N_4815,N_4845);
or UO_228 (O_228,N_4657,N_4979);
or UO_229 (O_229,N_4981,N_4733);
or UO_230 (O_230,N_4896,N_4869);
nand UO_231 (O_231,N_4548,N_4946);
or UO_232 (O_232,N_4646,N_4908);
xor UO_233 (O_233,N_4691,N_4537);
and UO_234 (O_234,N_4882,N_4746);
or UO_235 (O_235,N_4826,N_4562);
or UO_236 (O_236,N_4631,N_4707);
xor UO_237 (O_237,N_4833,N_4516);
nand UO_238 (O_238,N_4605,N_4676);
nand UO_239 (O_239,N_4581,N_4521);
nor UO_240 (O_240,N_4626,N_4536);
nand UO_241 (O_241,N_4776,N_4835);
or UO_242 (O_242,N_4941,N_4643);
or UO_243 (O_243,N_4959,N_4694);
or UO_244 (O_244,N_4886,N_4693);
nor UO_245 (O_245,N_4705,N_4784);
nand UO_246 (O_246,N_4773,N_4556);
or UO_247 (O_247,N_4570,N_4965);
nor UO_248 (O_248,N_4870,N_4804);
and UO_249 (O_249,N_4630,N_4898);
nor UO_250 (O_250,N_4637,N_4641);
or UO_251 (O_251,N_4989,N_4734);
nor UO_252 (O_252,N_4715,N_4961);
or UO_253 (O_253,N_4614,N_4905);
nand UO_254 (O_254,N_4553,N_4837);
nor UO_255 (O_255,N_4953,N_4598);
or UO_256 (O_256,N_4671,N_4975);
xnor UO_257 (O_257,N_4560,N_4799);
nand UO_258 (O_258,N_4631,N_4647);
and UO_259 (O_259,N_4512,N_4645);
and UO_260 (O_260,N_4797,N_4970);
xor UO_261 (O_261,N_4574,N_4913);
nand UO_262 (O_262,N_4537,N_4673);
nor UO_263 (O_263,N_4753,N_4879);
and UO_264 (O_264,N_4588,N_4948);
xor UO_265 (O_265,N_4991,N_4690);
nand UO_266 (O_266,N_4730,N_4551);
xor UO_267 (O_267,N_4882,N_4562);
xnor UO_268 (O_268,N_4736,N_4560);
xor UO_269 (O_269,N_4741,N_4637);
nor UO_270 (O_270,N_4995,N_4659);
or UO_271 (O_271,N_4923,N_4961);
xnor UO_272 (O_272,N_4749,N_4886);
nand UO_273 (O_273,N_4746,N_4502);
nand UO_274 (O_274,N_4865,N_4721);
xor UO_275 (O_275,N_4783,N_4586);
and UO_276 (O_276,N_4603,N_4773);
xnor UO_277 (O_277,N_4611,N_4601);
or UO_278 (O_278,N_4659,N_4958);
or UO_279 (O_279,N_4565,N_4561);
nand UO_280 (O_280,N_4772,N_4815);
nand UO_281 (O_281,N_4986,N_4540);
nand UO_282 (O_282,N_4801,N_4849);
nand UO_283 (O_283,N_4867,N_4698);
xor UO_284 (O_284,N_4687,N_4817);
or UO_285 (O_285,N_4602,N_4784);
and UO_286 (O_286,N_4635,N_4839);
nor UO_287 (O_287,N_4790,N_4933);
xor UO_288 (O_288,N_4926,N_4724);
or UO_289 (O_289,N_4631,N_4884);
nor UO_290 (O_290,N_4971,N_4736);
and UO_291 (O_291,N_4917,N_4816);
nor UO_292 (O_292,N_4663,N_4512);
or UO_293 (O_293,N_4906,N_4644);
xor UO_294 (O_294,N_4934,N_4865);
and UO_295 (O_295,N_4558,N_4842);
xnor UO_296 (O_296,N_4989,N_4769);
nor UO_297 (O_297,N_4618,N_4501);
or UO_298 (O_298,N_4874,N_4607);
nor UO_299 (O_299,N_4949,N_4813);
nand UO_300 (O_300,N_4643,N_4617);
nand UO_301 (O_301,N_4992,N_4953);
xnor UO_302 (O_302,N_4785,N_4811);
nand UO_303 (O_303,N_4617,N_4657);
nor UO_304 (O_304,N_4845,N_4971);
or UO_305 (O_305,N_4943,N_4811);
nor UO_306 (O_306,N_4668,N_4815);
and UO_307 (O_307,N_4645,N_4920);
or UO_308 (O_308,N_4830,N_4880);
nand UO_309 (O_309,N_4715,N_4663);
nand UO_310 (O_310,N_4954,N_4820);
and UO_311 (O_311,N_4506,N_4572);
xor UO_312 (O_312,N_4664,N_4940);
and UO_313 (O_313,N_4929,N_4697);
xor UO_314 (O_314,N_4527,N_4839);
nor UO_315 (O_315,N_4785,N_4550);
and UO_316 (O_316,N_4529,N_4677);
and UO_317 (O_317,N_4876,N_4560);
nor UO_318 (O_318,N_4978,N_4828);
xnor UO_319 (O_319,N_4756,N_4987);
xnor UO_320 (O_320,N_4865,N_4891);
nand UO_321 (O_321,N_4807,N_4537);
or UO_322 (O_322,N_4637,N_4635);
nand UO_323 (O_323,N_4921,N_4914);
and UO_324 (O_324,N_4911,N_4889);
and UO_325 (O_325,N_4933,N_4721);
and UO_326 (O_326,N_4804,N_4934);
nor UO_327 (O_327,N_4510,N_4752);
nor UO_328 (O_328,N_4823,N_4965);
nand UO_329 (O_329,N_4915,N_4544);
xor UO_330 (O_330,N_4668,N_4537);
nor UO_331 (O_331,N_4554,N_4694);
nand UO_332 (O_332,N_4746,N_4641);
nand UO_333 (O_333,N_4936,N_4571);
nand UO_334 (O_334,N_4583,N_4617);
or UO_335 (O_335,N_4939,N_4679);
and UO_336 (O_336,N_4702,N_4622);
xor UO_337 (O_337,N_4737,N_4845);
and UO_338 (O_338,N_4549,N_4686);
nor UO_339 (O_339,N_4886,N_4523);
or UO_340 (O_340,N_4621,N_4970);
or UO_341 (O_341,N_4903,N_4911);
nand UO_342 (O_342,N_4664,N_4619);
or UO_343 (O_343,N_4856,N_4666);
nand UO_344 (O_344,N_4710,N_4601);
nand UO_345 (O_345,N_4676,N_4966);
and UO_346 (O_346,N_4771,N_4735);
or UO_347 (O_347,N_4907,N_4820);
and UO_348 (O_348,N_4753,N_4909);
xor UO_349 (O_349,N_4972,N_4944);
nor UO_350 (O_350,N_4854,N_4907);
and UO_351 (O_351,N_4673,N_4701);
nor UO_352 (O_352,N_4858,N_4938);
nand UO_353 (O_353,N_4727,N_4735);
and UO_354 (O_354,N_4526,N_4794);
nor UO_355 (O_355,N_4714,N_4705);
and UO_356 (O_356,N_4559,N_4702);
and UO_357 (O_357,N_4692,N_4530);
nand UO_358 (O_358,N_4836,N_4820);
or UO_359 (O_359,N_4866,N_4610);
nand UO_360 (O_360,N_4969,N_4520);
or UO_361 (O_361,N_4752,N_4931);
nand UO_362 (O_362,N_4779,N_4738);
or UO_363 (O_363,N_4969,N_4624);
xor UO_364 (O_364,N_4589,N_4655);
nor UO_365 (O_365,N_4616,N_4728);
and UO_366 (O_366,N_4953,N_4526);
or UO_367 (O_367,N_4997,N_4633);
and UO_368 (O_368,N_4558,N_4628);
nand UO_369 (O_369,N_4907,N_4845);
xnor UO_370 (O_370,N_4631,N_4518);
xnor UO_371 (O_371,N_4962,N_4564);
or UO_372 (O_372,N_4628,N_4527);
and UO_373 (O_373,N_4978,N_4881);
nor UO_374 (O_374,N_4620,N_4807);
and UO_375 (O_375,N_4832,N_4541);
nand UO_376 (O_376,N_4936,N_4668);
xor UO_377 (O_377,N_4598,N_4924);
or UO_378 (O_378,N_4760,N_4938);
and UO_379 (O_379,N_4921,N_4684);
nand UO_380 (O_380,N_4898,N_4587);
and UO_381 (O_381,N_4593,N_4741);
and UO_382 (O_382,N_4691,N_4614);
and UO_383 (O_383,N_4602,N_4795);
and UO_384 (O_384,N_4709,N_4620);
nor UO_385 (O_385,N_4597,N_4640);
xnor UO_386 (O_386,N_4748,N_4897);
and UO_387 (O_387,N_4887,N_4698);
nand UO_388 (O_388,N_4905,N_4909);
and UO_389 (O_389,N_4597,N_4516);
and UO_390 (O_390,N_4586,N_4527);
or UO_391 (O_391,N_4528,N_4634);
and UO_392 (O_392,N_4737,N_4932);
nand UO_393 (O_393,N_4572,N_4954);
nor UO_394 (O_394,N_4597,N_4878);
nand UO_395 (O_395,N_4790,N_4937);
xnor UO_396 (O_396,N_4695,N_4764);
nor UO_397 (O_397,N_4682,N_4874);
nand UO_398 (O_398,N_4801,N_4577);
nand UO_399 (O_399,N_4720,N_4774);
and UO_400 (O_400,N_4952,N_4873);
and UO_401 (O_401,N_4545,N_4633);
nor UO_402 (O_402,N_4779,N_4814);
nand UO_403 (O_403,N_4984,N_4892);
nand UO_404 (O_404,N_4973,N_4883);
xnor UO_405 (O_405,N_4939,N_4654);
nor UO_406 (O_406,N_4966,N_4827);
nand UO_407 (O_407,N_4662,N_4572);
nand UO_408 (O_408,N_4623,N_4772);
nand UO_409 (O_409,N_4727,N_4532);
nor UO_410 (O_410,N_4971,N_4699);
and UO_411 (O_411,N_4695,N_4570);
nand UO_412 (O_412,N_4751,N_4512);
xor UO_413 (O_413,N_4615,N_4935);
and UO_414 (O_414,N_4627,N_4501);
nand UO_415 (O_415,N_4717,N_4529);
and UO_416 (O_416,N_4915,N_4940);
xor UO_417 (O_417,N_4700,N_4909);
and UO_418 (O_418,N_4699,N_4524);
xnor UO_419 (O_419,N_4679,N_4819);
or UO_420 (O_420,N_4638,N_4563);
nor UO_421 (O_421,N_4656,N_4501);
nor UO_422 (O_422,N_4929,N_4778);
or UO_423 (O_423,N_4574,N_4898);
xor UO_424 (O_424,N_4617,N_4595);
nor UO_425 (O_425,N_4594,N_4742);
and UO_426 (O_426,N_4983,N_4508);
xnor UO_427 (O_427,N_4528,N_4970);
nand UO_428 (O_428,N_4588,N_4528);
nor UO_429 (O_429,N_4521,N_4559);
xnor UO_430 (O_430,N_4870,N_4779);
nand UO_431 (O_431,N_4738,N_4749);
nand UO_432 (O_432,N_4784,N_4854);
or UO_433 (O_433,N_4978,N_4877);
or UO_434 (O_434,N_4786,N_4636);
and UO_435 (O_435,N_4889,N_4686);
or UO_436 (O_436,N_4782,N_4893);
nand UO_437 (O_437,N_4933,N_4612);
and UO_438 (O_438,N_4817,N_4991);
and UO_439 (O_439,N_4791,N_4769);
and UO_440 (O_440,N_4800,N_4707);
nand UO_441 (O_441,N_4556,N_4849);
nand UO_442 (O_442,N_4984,N_4797);
xnor UO_443 (O_443,N_4731,N_4728);
nor UO_444 (O_444,N_4893,N_4814);
or UO_445 (O_445,N_4970,N_4836);
nand UO_446 (O_446,N_4816,N_4978);
and UO_447 (O_447,N_4596,N_4983);
or UO_448 (O_448,N_4996,N_4585);
or UO_449 (O_449,N_4530,N_4570);
or UO_450 (O_450,N_4627,N_4510);
or UO_451 (O_451,N_4599,N_4886);
nor UO_452 (O_452,N_4867,N_4572);
xor UO_453 (O_453,N_4921,N_4789);
and UO_454 (O_454,N_4612,N_4594);
nand UO_455 (O_455,N_4803,N_4726);
or UO_456 (O_456,N_4869,N_4595);
nand UO_457 (O_457,N_4969,N_4949);
and UO_458 (O_458,N_4965,N_4546);
nand UO_459 (O_459,N_4537,N_4734);
xnor UO_460 (O_460,N_4695,N_4981);
nor UO_461 (O_461,N_4835,N_4543);
xnor UO_462 (O_462,N_4907,N_4867);
nor UO_463 (O_463,N_4810,N_4512);
nor UO_464 (O_464,N_4761,N_4906);
xor UO_465 (O_465,N_4922,N_4662);
and UO_466 (O_466,N_4966,N_4880);
nor UO_467 (O_467,N_4695,N_4949);
nand UO_468 (O_468,N_4960,N_4562);
nand UO_469 (O_469,N_4609,N_4505);
or UO_470 (O_470,N_4728,N_4795);
nand UO_471 (O_471,N_4842,N_4636);
nor UO_472 (O_472,N_4574,N_4766);
or UO_473 (O_473,N_4987,N_4876);
nand UO_474 (O_474,N_4752,N_4660);
nor UO_475 (O_475,N_4917,N_4741);
xor UO_476 (O_476,N_4788,N_4786);
and UO_477 (O_477,N_4573,N_4583);
nor UO_478 (O_478,N_4928,N_4790);
and UO_479 (O_479,N_4965,N_4984);
nand UO_480 (O_480,N_4807,N_4741);
and UO_481 (O_481,N_4582,N_4552);
or UO_482 (O_482,N_4548,N_4642);
nand UO_483 (O_483,N_4517,N_4598);
nand UO_484 (O_484,N_4558,N_4617);
and UO_485 (O_485,N_4627,N_4955);
and UO_486 (O_486,N_4600,N_4687);
xor UO_487 (O_487,N_4792,N_4829);
nand UO_488 (O_488,N_4739,N_4502);
nand UO_489 (O_489,N_4862,N_4880);
or UO_490 (O_490,N_4957,N_4681);
and UO_491 (O_491,N_4590,N_4996);
and UO_492 (O_492,N_4513,N_4566);
xnor UO_493 (O_493,N_4927,N_4896);
and UO_494 (O_494,N_4981,N_4986);
and UO_495 (O_495,N_4690,N_4918);
or UO_496 (O_496,N_4732,N_4710);
xor UO_497 (O_497,N_4971,N_4988);
nand UO_498 (O_498,N_4912,N_4562);
xnor UO_499 (O_499,N_4553,N_4886);
or UO_500 (O_500,N_4638,N_4859);
nand UO_501 (O_501,N_4664,N_4827);
xnor UO_502 (O_502,N_4763,N_4652);
nand UO_503 (O_503,N_4864,N_4727);
nand UO_504 (O_504,N_4607,N_4917);
nand UO_505 (O_505,N_4963,N_4530);
and UO_506 (O_506,N_4611,N_4681);
or UO_507 (O_507,N_4824,N_4747);
and UO_508 (O_508,N_4950,N_4588);
nor UO_509 (O_509,N_4655,N_4947);
nor UO_510 (O_510,N_4721,N_4533);
xnor UO_511 (O_511,N_4821,N_4862);
nor UO_512 (O_512,N_4904,N_4556);
nand UO_513 (O_513,N_4785,N_4991);
xnor UO_514 (O_514,N_4974,N_4546);
nor UO_515 (O_515,N_4813,N_4529);
nand UO_516 (O_516,N_4753,N_4529);
and UO_517 (O_517,N_4934,N_4976);
or UO_518 (O_518,N_4511,N_4877);
or UO_519 (O_519,N_4826,N_4759);
and UO_520 (O_520,N_4801,N_4518);
or UO_521 (O_521,N_4896,N_4739);
nand UO_522 (O_522,N_4635,N_4677);
and UO_523 (O_523,N_4929,N_4819);
and UO_524 (O_524,N_4697,N_4568);
or UO_525 (O_525,N_4937,N_4585);
nand UO_526 (O_526,N_4945,N_4610);
nand UO_527 (O_527,N_4504,N_4723);
and UO_528 (O_528,N_4547,N_4632);
nand UO_529 (O_529,N_4540,N_4669);
and UO_530 (O_530,N_4705,N_4598);
and UO_531 (O_531,N_4503,N_4612);
xor UO_532 (O_532,N_4515,N_4870);
xnor UO_533 (O_533,N_4930,N_4524);
nor UO_534 (O_534,N_4747,N_4954);
xor UO_535 (O_535,N_4748,N_4556);
and UO_536 (O_536,N_4909,N_4600);
xnor UO_537 (O_537,N_4554,N_4953);
and UO_538 (O_538,N_4821,N_4590);
xor UO_539 (O_539,N_4728,N_4651);
xor UO_540 (O_540,N_4619,N_4947);
or UO_541 (O_541,N_4576,N_4957);
xor UO_542 (O_542,N_4602,N_4818);
xor UO_543 (O_543,N_4954,N_4860);
and UO_544 (O_544,N_4866,N_4586);
and UO_545 (O_545,N_4888,N_4840);
nand UO_546 (O_546,N_4839,N_4748);
nor UO_547 (O_547,N_4910,N_4615);
and UO_548 (O_548,N_4516,N_4781);
nor UO_549 (O_549,N_4705,N_4699);
or UO_550 (O_550,N_4818,N_4502);
or UO_551 (O_551,N_4745,N_4963);
nor UO_552 (O_552,N_4675,N_4770);
and UO_553 (O_553,N_4560,N_4987);
nor UO_554 (O_554,N_4934,N_4524);
nand UO_555 (O_555,N_4923,N_4845);
xor UO_556 (O_556,N_4747,N_4873);
xnor UO_557 (O_557,N_4726,N_4619);
or UO_558 (O_558,N_4720,N_4631);
or UO_559 (O_559,N_4546,N_4782);
nand UO_560 (O_560,N_4802,N_4868);
nor UO_561 (O_561,N_4678,N_4804);
and UO_562 (O_562,N_4559,N_4537);
or UO_563 (O_563,N_4883,N_4745);
and UO_564 (O_564,N_4655,N_4864);
xnor UO_565 (O_565,N_4545,N_4853);
or UO_566 (O_566,N_4690,N_4744);
or UO_567 (O_567,N_4754,N_4974);
nor UO_568 (O_568,N_4882,N_4575);
and UO_569 (O_569,N_4619,N_4743);
or UO_570 (O_570,N_4848,N_4578);
xnor UO_571 (O_571,N_4959,N_4787);
nor UO_572 (O_572,N_4864,N_4933);
and UO_573 (O_573,N_4705,N_4877);
nand UO_574 (O_574,N_4681,N_4901);
xnor UO_575 (O_575,N_4776,N_4819);
or UO_576 (O_576,N_4800,N_4769);
or UO_577 (O_577,N_4916,N_4771);
nand UO_578 (O_578,N_4504,N_4789);
or UO_579 (O_579,N_4810,N_4962);
nor UO_580 (O_580,N_4752,N_4607);
nand UO_581 (O_581,N_4686,N_4543);
nand UO_582 (O_582,N_4569,N_4986);
and UO_583 (O_583,N_4919,N_4544);
nor UO_584 (O_584,N_4580,N_4620);
nand UO_585 (O_585,N_4791,N_4803);
and UO_586 (O_586,N_4791,N_4774);
xor UO_587 (O_587,N_4685,N_4814);
or UO_588 (O_588,N_4760,N_4682);
xor UO_589 (O_589,N_4632,N_4902);
xnor UO_590 (O_590,N_4776,N_4890);
or UO_591 (O_591,N_4713,N_4930);
nor UO_592 (O_592,N_4873,N_4926);
xnor UO_593 (O_593,N_4742,N_4659);
nand UO_594 (O_594,N_4526,N_4892);
xnor UO_595 (O_595,N_4595,N_4622);
nand UO_596 (O_596,N_4816,N_4948);
nor UO_597 (O_597,N_4989,N_4848);
and UO_598 (O_598,N_4835,N_4947);
or UO_599 (O_599,N_4790,N_4995);
and UO_600 (O_600,N_4619,N_4571);
or UO_601 (O_601,N_4795,N_4623);
xor UO_602 (O_602,N_4933,N_4561);
nor UO_603 (O_603,N_4566,N_4831);
nand UO_604 (O_604,N_4707,N_4604);
xor UO_605 (O_605,N_4713,N_4984);
xor UO_606 (O_606,N_4992,N_4602);
and UO_607 (O_607,N_4828,N_4937);
nor UO_608 (O_608,N_4815,N_4779);
nand UO_609 (O_609,N_4652,N_4966);
nand UO_610 (O_610,N_4741,N_4930);
nand UO_611 (O_611,N_4893,N_4555);
xnor UO_612 (O_612,N_4577,N_4800);
and UO_613 (O_613,N_4667,N_4583);
nor UO_614 (O_614,N_4742,N_4909);
or UO_615 (O_615,N_4967,N_4537);
and UO_616 (O_616,N_4863,N_4710);
and UO_617 (O_617,N_4578,N_4562);
or UO_618 (O_618,N_4735,N_4717);
xnor UO_619 (O_619,N_4954,N_4556);
and UO_620 (O_620,N_4826,N_4671);
or UO_621 (O_621,N_4856,N_4857);
nand UO_622 (O_622,N_4624,N_4891);
or UO_623 (O_623,N_4814,N_4720);
and UO_624 (O_624,N_4937,N_4930);
and UO_625 (O_625,N_4504,N_4771);
xnor UO_626 (O_626,N_4885,N_4952);
xor UO_627 (O_627,N_4620,N_4893);
xor UO_628 (O_628,N_4637,N_4574);
nor UO_629 (O_629,N_4980,N_4646);
nor UO_630 (O_630,N_4801,N_4685);
xor UO_631 (O_631,N_4743,N_4827);
xnor UO_632 (O_632,N_4638,N_4992);
nand UO_633 (O_633,N_4821,N_4971);
xnor UO_634 (O_634,N_4855,N_4916);
and UO_635 (O_635,N_4792,N_4606);
nor UO_636 (O_636,N_4646,N_4693);
or UO_637 (O_637,N_4845,N_4717);
xor UO_638 (O_638,N_4941,N_4629);
nand UO_639 (O_639,N_4830,N_4545);
nand UO_640 (O_640,N_4894,N_4712);
or UO_641 (O_641,N_4560,N_4508);
and UO_642 (O_642,N_4653,N_4500);
or UO_643 (O_643,N_4590,N_4815);
xnor UO_644 (O_644,N_4930,N_4710);
and UO_645 (O_645,N_4606,N_4965);
nand UO_646 (O_646,N_4547,N_4594);
or UO_647 (O_647,N_4634,N_4895);
nand UO_648 (O_648,N_4778,N_4760);
nor UO_649 (O_649,N_4517,N_4516);
and UO_650 (O_650,N_4558,N_4662);
nor UO_651 (O_651,N_4506,N_4965);
nand UO_652 (O_652,N_4628,N_4503);
or UO_653 (O_653,N_4548,N_4964);
or UO_654 (O_654,N_4506,N_4759);
nand UO_655 (O_655,N_4785,N_4980);
nand UO_656 (O_656,N_4900,N_4860);
or UO_657 (O_657,N_4777,N_4841);
or UO_658 (O_658,N_4941,N_4663);
nor UO_659 (O_659,N_4524,N_4815);
nand UO_660 (O_660,N_4695,N_4858);
xor UO_661 (O_661,N_4874,N_4900);
and UO_662 (O_662,N_4666,N_4925);
xnor UO_663 (O_663,N_4561,N_4724);
nor UO_664 (O_664,N_4933,N_4700);
nor UO_665 (O_665,N_4917,N_4886);
nand UO_666 (O_666,N_4810,N_4598);
and UO_667 (O_667,N_4902,N_4510);
or UO_668 (O_668,N_4910,N_4516);
and UO_669 (O_669,N_4903,N_4820);
or UO_670 (O_670,N_4816,N_4869);
and UO_671 (O_671,N_4530,N_4603);
and UO_672 (O_672,N_4840,N_4824);
or UO_673 (O_673,N_4925,N_4635);
or UO_674 (O_674,N_4614,N_4653);
and UO_675 (O_675,N_4544,N_4808);
xor UO_676 (O_676,N_4647,N_4792);
nor UO_677 (O_677,N_4834,N_4905);
nor UO_678 (O_678,N_4863,N_4789);
or UO_679 (O_679,N_4572,N_4932);
nor UO_680 (O_680,N_4538,N_4762);
xnor UO_681 (O_681,N_4556,N_4984);
or UO_682 (O_682,N_4984,N_4599);
nor UO_683 (O_683,N_4785,N_4896);
xnor UO_684 (O_684,N_4564,N_4644);
and UO_685 (O_685,N_4672,N_4723);
nand UO_686 (O_686,N_4970,N_4578);
and UO_687 (O_687,N_4541,N_4702);
and UO_688 (O_688,N_4924,N_4594);
nand UO_689 (O_689,N_4942,N_4970);
or UO_690 (O_690,N_4747,N_4674);
nor UO_691 (O_691,N_4873,N_4687);
nand UO_692 (O_692,N_4801,N_4803);
and UO_693 (O_693,N_4674,N_4699);
nor UO_694 (O_694,N_4963,N_4666);
and UO_695 (O_695,N_4610,N_4561);
nand UO_696 (O_696,N_4763,N_4564);
and UO_697 (O_697,N_4623,N_4621);
or UO_698 (O_698,N_4674,N_4622);
and UO_699 (O_699,N_4994,N_4960);
and UO_700 (O_700,N_4515,N_4766);
nand UO_701 (O_701,N_4939,N_4632);
and UO_702 (O_702,N_4908,N_4670);
or UO_703 (O_703,N_4796,N_4757);
nor UO_704 (O_704,N_4594,N_4966);
and UO_705 (O_705,N_4976,N_4777);
nand UO_706 (O_706,N_4771,N_4639);
nand UO_707 (O_707,N_4579,N_4863);
nand UO_708 (O_708,N_4666,N_4875);
nand UO_709 (O_709,N_4978,N_4690);
and UO_710 (O_710,N_4929,N_4584);
or UO_711 (O_711,N_4952,N_4565);
xnor UO_712 (O_712,N_4633,N_4987);
and UO_713 (O_713,N_4912,N_4520);
xor UO_714 (O_714,N_4728,N_4580);
or UO_715 (O_715,N_4720,N_4794);
or UO_716 (O_716,N_4562,N_4968);
and UO_717 (O_717,N_4902,N_4727);
xnor UO_718 (O_718,N_4761,N_4655);
nor UO_719 (O_719,N_4911,N_4796);
and UO_720 (O_720,N_4657,N_4653);
and UO_721 (O_721,N_4762,N_4742);
or UO_722 (O_722,N_4500,N_4527);
and UO_723 (O_723,N_4593,N_4863);
and UO_724 (O_724,N_4635,N_4695);
nor UO_725 (O_725,N_4606,N_4660);
or UO_726 (O_726,N_4631,N_4956);
nor UO_727 (O_727,N_4772,N_4697);
nor UO_728 (O_728,N_4879,N_4640);
or UO_729 (O_729,N_4587,N_4635);
nor UO_730 (O_730,N_4699,N_4758);
xor UO_731 (O_731,N_4797,N_4733);
and UO_732 (O_732,N_4624,N_4878);
nand UO_733 (O_733,N_4824,N_4757);
xnor UO_734 (O_734,N_4976,N_4633);
xnor UO_735 (O_735,N_4941,N_4762);
or UO_736 (O_736,N_4719,N_4648);
or UO_737 (O_737,N_4570,N_4951);
nor UO_738 (O_738,N_4975,N_4986);
xnor UO_739 (O_739,N_4931,N_4943);
xnor UO_740 (O_740,N_4589,N_4748);
xor UO_741 (O_741,N_4731,N_4748);
or UO_742 (O_742,N_4590,N_4755);
xnor UO_743 (O_743,N_4852,N_4902);
or UO_744 (O_744,N_4804,N_4831);
or UO_745 (O_745,N_4815,N_4694);
nand UO_746 (O_746,N_4645,N_4821);
nand UO_747 (O_747,N_4614,N_4988);
nor UO_748 (O_748,N_4995,N_4556);
nand UO_749 (O_749,N_4709,N_4743);
and UO_750 (O_750,N_4855,N_4892);
or UO_751 (O_751,N_4727,N_4533);
and UO_752 (O_752,N_4743,N_4581);
nand UO_753 (O_753,N_4563,N_4703);
nor UO_754 (O_754,N_4633,N_4838);
and UO_755 (O_755,N_4984,N_4584);
xor UO_756 (O_756,N_4979,N_4711);
nand UO_757 (O_757,N_4518,N_4755);
nand UO_758 (O_758,N_4645,N_4649);
nand UO_759 (O_759,N_4841,N_4567);
nor UO_760 (O_760,N_4680,N_4586);
nand UO_761 (O_761,N_4936,N_4915);
xnor UO_762 (O_762,N_4600,N_4655);
xnor UO_763 (O_763,N_4681,N_4598);
nand UO_764 (O_764,N_4568,N_4836);
xor UO_765 (O_765,N_4840,N_4767);
and UO_766 (O_766,N_4925,N_4804);
or UO_767 (O_767,N_4955,N_4722);
nand UO_768 (O_768,N_4557,N_4567);
xnor UO_769 (O_769,N_4592,N_4924);
and UO_770 (O_770,N_4794,N_4986);
nor UO_771 (O_771,N_4801,N_4512);
nor UO_772 (O_772,N_4710,N_4806);
or UO_773 (O_773,N_4603,N_4564);
or UO_774 (O_774,N_4943,N_4571);
nand UO_775 (O_775,N_4754,N_4686);
nor UO_776 (O_776,N_4808,N_4810);
nand UO_777 (O_777,N_4646,N_4756);
and UO_778 (O_778,N_4620,N_4996);
and UO_779 (O_779,N_4926,N_4524);
and UO_780 (O_780,N_4683,N_4589);
or UO_781 (O_781,N_4577,N_4754);
nand UO_782 (O_782,N_4906,N_4636);
and UO_783 (O_783,N_4652,N_4504);
xor UO_784 (O_784,N_4965,N_4902);
nand UO_785 (O_785,N_4712,N_4996);
nand UO_786 (O_786,N_4709,N_4610);
nor UO_787 (O_787,N_4754,N_4596);
and UO_788 (O_788,N_4715,N_4894);
nor UO_789 (O_789,N_4581,N_4806);
nor UO_790 (O_790,N_4655,N_4682);
nand UO_791 (O_791,N_4794,N_4976);
nor UO_792 (O_792,N_4958,N_4591);
and UO_793 (O_793,N_4777,N_4908);
xnor UO_794 (O_794,N_4687,N_4694);
nand UO_795 (O_795,N_4598,N_4881);
nor UO_796 (O_796,N_4605,N_4750);
nor UO_797 (O_797,N_4776,N_4908);
nor UO_798 (O_798,N_4866,N_4994);
xnor UO_799 (O_799,N_4603,N_4636);
nor UO_800 (O_800,N_4553,N_4981);
xnor UO_801 (O_801,N_4823,N_4640);
nor UO_802 (O_802,N_4714,N_4837);
and UO_803 (O_803,N_4792,N_4818);
xor UO_804 (O_804,N_4923,N_4875);
xnor UO_805 (O_805,N_4617,N_4693);
nand UO_806 (O_806,N_4613,N_4658);
and UO_807 (O_807,N_4945,N_4893);
nor UO_808 (O_808,N_4736,N_4647);
nand UO_809 (O_809,N_4736,N_4789);
nand UO_810 (O_810,N_4860,N_4728);
nor UO_811 (O_811,N_4917,N_4755);
and UO_812 (O_812,N_4666,N_4626);
and UO_813 (O_813,N_4846,N_4928);
or UO_814 (O_814,N_4781,N_4613);
nand UO_815 (O_815,N_4564,N_4706);
nand UO_816 (O_816,N_4943,N_4916);
xor UO_817 (O_817,N_4864,N_4802);
xnor UO_818 (O_818,N_4932,N_4540);
or UO_819 (O_819,N_4572,N_4882);
nand UO_820 (O_820,N_4673,N_4618);
and UO_821 (O_821,N_4946,N_4714);
or UO_822 (O_822,N_4521,N_4625);
xor UO_823 (O_823,N_4863,N_4869);
nor UO_824 (O_824,N_4831,N_4765);
nor UO_825 (O_825,N_4699,N_4762);
nand UO_826 (O_826,N_4554,N_4672);
or UO_827 (O_827,N_4862,N_4684);
or UO_828 (O_828,N_4774,N_4895);
and UO_829 (O_829,N_4837,N_4952);
nor UO_830 (O_830,N_4616,N_4880);
xnor UO_831 (O_831,N_4557,N_4546);
nand UO_832 (O_832,N_4873,N_4786);
xor UO_833 (O_833,N_4500,N_4638);
nand UO_834 (O_834,N_4765,N_4943);
xnor UO_835 (O_835,N_4926,N_4568);
nand UO_836 (O_836,N_4738,N_4645);
or UO_837 (O_837,N_4624,N_4948);
or UO_838 (O_838,N_4840,N_4927);
and UO_839 (O_839,N_4680,N_4816);
or UO_840 (O_840,N_4685,N_4536);
and UO_841 (O_841,N_4990,N_4817);
or UO_842 (O_842,N_4880,N_4794);
xnor UO_843 (O_843,N_4769,N_4766);
or UO_844 (O_844,N_4772,N_4577);
nand UO_845 (O_845,N_4922,N_4742);
xor UO_846 (O_846,N_4727,N_4747);
nand UO_847 (O_847,N_4761,N_4799);
nor UO_848 (O_848,N_4608,N_4720);
nor UO_849 (O_849,N_4842,N_4756);
nand UO_850 (O_850,N_4694,N_4774);
nand UO_851 (O_851,N_4724,N_4529);
xnor UO_852 (O_852,N_4561,N_4568);
nor UO_853 (O_853,N_4789,N_4587);
and UO_854 (O_854,N_4723,N_4829);
or UO_855 (O_855,N_4730,N_4972);
xnor UO_856 (O_856,N_4898,N_4985);
xnor UO_857 (O_857,N_4743,N_4849);
or UO_858 (O_858,N_4763,N_4619);
nor UO_859 (O_859,N_4970,N_4568);
or UO_860 (O_860,N_4905,N_4927);
or UO_861 (O_861,N_4723,N_4505);
nor UO_862 (O_862,N_4716,N_4584);
nand UO_863 (O_863,N_4511,N_4927);
xnor UO_864 (O_864,N_4700,N_4782);
nand UO_865 (O_865,N_4686,N_4934);
or UO_866 (O_866,N_4696,N_4990);
nor UO_867 (O_867,N_4680,N_4512);
xor UO_868 (O_868,N_4716,N_4599);
or UO_869 (O_869,N_4645,N_4650);
or UO_870 (O_870,N_4727,N_4589);
and UO_871 (O_871,N_4788,N_4675);
or UO_872 (O_872,N_4599,N_4706);
and UO_873 (O_873,N_4762,N_4804);
nor UO_874 (O_874,N_4542,N_4947);
xnor UO_875 (O_875,N_4732,N_4546);
nand UO_876 (O_876,N_4858,N_4813);
or UO_877 (O_877,N_4576,N_4726);
nand UO_878 (O_878,N_4576,N_4611);
or UO_879 (O_879,N_4761,N_4502);
or UO_880 (O_880,N_4559,N_4531);
and UO_881 (O_881,N_4694,N_4616);
xor UO_882 (O_882,N_4745,N_4527);
nand UO_883 (O_883,N_4785,N_4879);
or UO_884 (O_884,N_4716,N_4981);
nor UO_885 (O_885,N_4510,N_4883);
xnor UO_886 (O_886,N_4859,N_4526);
xnor UO_887 (O_887,N_4602,N_4651);
nand UO_888 (O_888,N_4766,N_4619);
nand UO_889 (O_889,N_4712,N_4765);
xor UO_890 (O_890,N_4643,N_4733);
and UO_891 (O_891,N_4729,N_4664);
or UO_892 (O_892,N_4945,N_4736);
nor UO_893 (O_893,N_4892,N_4695);
and UO_894 (O_894,N_4677,N_4684);
xor UO_895 (O_895,N_4593,N_4601);
nand UO_896 (O_896,N_4539,N_4719);
or UO_897 (O_897,N_4738,N_4777);
nor UO_898 (O_898,N_4730,N_4614);
xnor UO_899 (O_899,N_4921,N_4802);
xor UO_900 (O_900,N_4606,N_4590);
nor UO_901 (O_901,N_4622,N_4885);
xnor UO_902 (O_902,N_4720,N_4634);
and UO_903 (O_903,N_4515,N_4659);
nor UO_904 (O_904,N_4778,N_4849);
xnor UO_905 (O_905,N_4728,N_4676);
xor UO_906 (O_906,N_4591,N_4757);
and UO_907 (O_907,N_4652,N_4971);
nor UO_908 (O_908,N_4733,N_4842);
nor UO_909 (O_909,N_4921,N_4865);
or UO_910 (O_910,N_4891,N_4955);
and UO_911 (O_911,N_4927,N_4573);
nor UO_912 (O_912,N_4799,N_4762);
xor UO_913 (O_913,N_4829,N_4593);
or UO_914 (O_914,N_4881,N_4854);
or UO_915 (O_915,N_4652,N_4783);
nor UO_916 (O_916,N_4750,N_4920);
nand UO_917 (O_917,N_4970,N_4566);
nand UO_918 (O_918,N_4780,N_4998);
nor UO_919 (O_919,N_4500,N_4745);
or UO_920 (O_920,N_4937,N_4738);
and UO_921 (O_921,N_4685,N_4638);
nor UO_922 (O_922,N_4914,N_4656);
xnor UO_923 (O_923,N_4698,N_4523);
xor UO_924 (O_924,N_4525,N_4566);
nor UO_925 (O_925,N_4517,N_4867);
nor UO_926 (O_926,N_4848,N_4903);
nand UO_927 (O_927,N_4804,N_4757);
or UO_928 (O_928,N_4560,N_4674);
or UO_929 (O_929,N_4900,N_4691);
or UO_930 (O_930,N_4739,N_4550);
nor UO_931 (O_931,N_4860,N_4894);
nand UO_932 (O_932,N_4793,N_4958);
nand UO_933 (O_933,N_4769,N_4816);
xnor UO_934 (O_934,N_4872,N_4677);
or UO_935 (O_935,N_4793,N_4848);
xor UO_936 (O_936,N_4968,N_4751);
nand UO_937 (O_937,N_4962,N_4575);
nand UO_938 (O_938,N_4664,N_4920);
xor UO_939 (O_939,N_4971,N_4910);
xor UO_940 (O_940,N_4544,N_4556);
and UO_941 (O_941,N_4851,N_4539);
and UO_942 (O_942,N_4974,N_4654);
nor UO_943 (O_943,N_4556,N_4846);
and UO_944 (O_944,N_4513,N_4766);
xnor UO_945 (O_945,N_4747,N_4887);
or UO_946 (O_946,N_4575,N_4584);
nand UO_947 (O_947,N_4632,N_4543);
xor UO_948 (O_948,N_4939,N_4785);
nand UO_949 (O_949,N_4575,N_4778);
and UO_950 (O_950,N_4658,N_4680);
nor UO_951 (O_951,N_4574,N_4686);
nand UO_952 (O_952,N_4682,N_4639);
nor UO_953 (O_953,N_4799,N_4748);
xor UO_954 (O_954,N_4780,N_4871);
nor UO_955 (O_955,N_4955,N_4736);
nand UO_956 (O_956,N_4759,N_4581);
nand UO_957 (O_957,N_4617,N_4654);
or UO_958 (O_958,N_4673,N_4602);
xor UO_959 (O_959,N_4914,N_4679);
nand UO_960 (O_960,N_4501,N_4922);
nand UO_961 (O_961,N_4691,N_4810);
or UO_962 (O_962,N_4564,N_4829);
or UO_963 (O_963,N_4884,N_4757);
or UO_964 (O_964,N_4521,N_4704);
nor UO_965 (O_965,N_4538,N_4500);
nand UO_966 (O_966,N_4805,N_4788);
or UO_967 (O_967,N_4767,N_4701);
nand UO_968 (O_968,N_4831,N_4879);
nor UO_969 (O_969,N_4667,N_4838);
xnor UO_970 (O_970,N_4877,N_4991);
nor UO_971 (O_971,N_4815,N_4686);
nand UO_972 (O_972,N_4754,N_4644);
and UO_973 (O_973,N_4644,N_4790);
and UO_974 (O_974,N_4548,N_4608);
nand UO_975 (O_975,N_4762,N_4831);
nand UO_976 (O_976,N_4985,N_4855);
or UO_977 (O_977,N_4777,N_4693);
nor UO_978 (O_978,N_4816,N_4559);
nor UO_979 (O_979,N_4823,N_4504);
and UO_980 (O_980,N_4512,N_4674);
nor UO_981 (O_981,N_4531,N_4798);
nand UO_982 (O_982,N_4839,N_4989);
and UO_983 (O_983,N_4631,N_4808);
nand UO_984 (O_984,N_4816,N_4619);
or UO_985 (O_985,N_4863,N_4795);
nor UO_986 (O_986,N_4687,N_4959);
and UO_987 (O_987,N_4730,N_4961);
and UO_988 (O_988,N_4600,N_4811);
xnor UO_989 (O_989,N_4556,N_4964);
and UO_990 (O_990,N_4659,N_4597);
nor UO_991 (O_991,N_4642,N_4570);
nand UO_992 (O_992,N_4916,N_4641);
and UO_993 (O_993,N_4691,N_4950);
or UO_994 (O_994,N_4715,N_4580);
or UO_995 (O_995,N_4704,N_4660);
or UO_996 (O_996,N_4944,N_4999);
nand UO_997 (O_997,N_4951,N_4962);
or UO_998 (O_998,N_4888,N_4801);
xor UO_999 (O_999,N_4689,N_4966);
endmodule