module basic_500_3000_500_50_levels_5xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nor U0 (N_0,In_331,In_232);
nor U1 (N_1,In_170,In_119);
or U2 (N_2,In_455,In_488);
nand U3 (N_3,In_79,In_147);
or U4 (N_4,In_402,In_54);
xor U5 (N_5,In_186,In_4);
and U6 (N_6,In_218,In_57);
nand U7 (N_7,In_83,In_230);
or U8 (N_8,In_258,In_233);
nand U9 (N_9,In_37,In_5);
or U10 (N_10,In_281,In_381);
and U11 (N_11,In_447,In_461);
and U12 (N_12,In_149,In_177);
nor U13 (N_13,In_131,In_209);
or U14 (N_14,In_460,In_264);
or U15 (N_15,In_397,In_457);
nand U16 (N_16,In_107,In_338);
nor U17 (N_17,In_221,In_354);
nand U18 (N_18,In_109,In_81);
and U19 (N_19,In_24,In_70);
nor U20 (N_20,In_395,In_432);
or U21 (N_21,In_55,In_326);
nand U22 (N_22,In_275,In_216);
nand U23 (N_23,In_392,In_439);
or U24 (N_24,In_296,In_433);
or U25 (N_25,In_316,In_219);
nand U26 (N_26,In_121,In_270);
nor U27 (N_27,In_476,In_104);
or U28 (N_28,In_239,In_375);
xor U29 (N_29,In_139,In_220);
or U30 (N_30,In_7,In_135);
or U31 (N_31,In_33,In_241);
nor U32 (N_32,In_98,In_47);
nor U33 (N_33,In_440,In_329);
or U34 (N_34,In_126,In_332);
and U35 (N_35,In_340,In_200);
nand U36 (N_36,In_134,In_297);
xor U37 (N_37,In_217,In_358);
and U38 (N_38,In_437,In_180);
xor U39 (N_39,In_388,In_94);
xor U40 (N_40,In_145,In_322);
and U41 (N_41,In_27,In_283);
or U42 (N_42,In_374,In_399);
nand U43 (N_43,In_11,In_409);
xor U44 (N_44,In_345,In_330);
nand U45 (N_45,In_84,In_159);
nand U46 (N_46,In_467,In_474);
and U47 (N_47,In_362,In_127);
and U48 (N_48,In_357,In_74);
and U49 (N_49,In_85,In_368);
nand U50 (N_50,In_334,In_295);
nand U51 (N_51,In_475,In_89);
nand U52 (N_52,In_192,In_44);
or U53 (N_53,In_367,In_304);
nor U54 (N_54,In_118,In_408);
or U55 (N_55,In_175,In_361);
nor U56 (N_56,In_15,In_208);
xor U57 (N_57,In_260,In_113);
and U58 (N_58,In_172,In_16);
or U59 (N_59,In_318,In_366);
nor U60 (N_60,In_224,In_41);
nor U61 (N_61,In_60,In_245);
and U62 (N_62,In_236,In_8);
nand U63 (N_63,In_133,In_88);
nand U64 (N_64,In_154,In_28);
xor U65 (N_65,In_396,In_491);
or U66 (N_66,In_273,In_34);
and U67 (N_67,In_306,In_10);
and U68 (N_68,In_337,In_76);
or U69 (N_69,In_77,In_243);
nor U70 (N_70,In_45,In_204);
xor U71 (N_71,In_314,N_45);
nand U72 (N_72,In_453,In_285);
nor U73 (N_73,In_406,In_495);
nand U74 (N_74,In_341,N_19);
xor U75 (N_75,In_259,In_184);
and U76 (N_76,In_417,In_385);
and U77 (N_77,In_282,In_312);
nand U78 (N_78,In_207,In_215);
and U79 (N_79,In_223,In_95);
nand U80 (N_80,In_487,In_317);
nand U81 (N_81,In_64,In_72);
or U82 (N_82,In_343,In_328);
nand U83 (N_83,In_101,In_496);
or U84 (N_84,In_468,In_155);
and U85 (N_85,In_268,In_80);
nor U86 (N_86,In_91,In_120);
nor U87 (N_87,In_364,In_344);
nand U88 (N_88,In_419,N_16);
nor U89 (N_89,In_48,In_480);
nor U90 (N_90,In_156,In_420);
or U91 (N_91,In_356,In_231);
nand U92 (N_92,N_6,In_188);
nand U93 (N_93,In_256,In_464);
xnor U94 (N_94,In_319,In_0);
nand U95 (N_95,In_189,In_249);
nand U96 (N_96,In_324,In_163);
and U97 (N_97,In_125,In_498);
and U98 (N_98,In_146,In_294);
nand U99 (N_99,N_47,In_214);
and U100 (N_100,In_53,In_247);
or U101 (N_101,In_376,In_50);
xor U102 (N_102,N_11,In_123);
nand U103 (N_103,In_255,In_31);
and U104 (N_104,In_383,In_242);
or U105 (N_105,In_181,In_140);
and U106 (N_106,In_234,In_473);
or U107 (N_107,In_213,In_211);
and U108 (N_108,N_14,N_21);
nor U109 (N_109,In_229,N_2);
nand U110 (N_110,N_29,In_350);
xor U111 (N_111,In_205,In_320);
nor U112 (N_112,In_179,N_7);
or U113 (N_113,In_286,In_450);
nand U114 (N_114,In_465,In_39);
and U115 (N_115,In_152,In_305);
nor U116 (N_116,In_478,In_132);
and U117 (N_117,In_19,N_33);
or U118 (N_118,In_416,In_142);
nand U119 (N_119,In_394,In_40);
nor U120 (N_120,In_427,In_150);
nand U121 (N_121,In_130,In_269);
nand U122 (N_122,In_17,N_86);
nand U123 (N_123,In_462,In_265);
and U124 (N_124,N_85,In_456);
nor U125 (N_125,N_30,N_0);
and U126 (N_126,N_63,N_73);
or U127 (N_127,In_448,In_3);
nand U128 (N_128,In_471,N_49);
nand U129 (N_129,N_62,N_94);
xnor U130 (N_130,In_244,In_203);
nand U131 (N_131,In_443,In_386);
or U132 (N_132,N_105,In_187);
or U133 (N_133,In_30,In_148);
or U134 (N_134,In_158,In_56);
nor U135 (N_135,In_171,In_261);
nor U136 (N_136,In_100,In_105);
nand U137 (N_137,In_373,N_81);
nand U138 (N_138,In_287,In_425);
nand U139 (N_139,N_44,In_289);
xor U140 (N_140,In_237,In_78);
or U141 (N_141,N_106,In_23);
nor U142 (N_142,In_407,In_38);
xor U143 (N_143,In_363,In_93);
nor U144 (N_144,In_35,N_57);
and U145 (N_145,N_65,In_62);
nor U146 (N_146,In_69,In_469);
or U147 (N_147,In_185,N_32);
or U148 (N_148,In_325,In_371);
nand U149 (N_149,N_84,In_235);
nand U150 (N_150,In_136,In_182);
xor U151 (N_151,In_400,N_88);
nand U152 (N_152,In_253,N_17);
nand U153 (N_153,N_116,In_372);
or U154 (N_154,In_360,In_404);
or U155 (N_155,N_31,N_9);
and U156 (N_156,In_497,In_138);
and U157 (N_157,In_102,In_199);
and U158 (N_158,N_113,N_12);
nand U159 (N_159,In_65,N_80);
nor U160 (N_160,In_477,In_90);
nor U161 (N_161,N_103,In_227);
nor U162 (N_162,In_277,In_52);
and U163 (N_163,In_106,N_110);
or U164 (N_164,In_418,In_302);
and U165 (N_165,In_403,In_202);
nor U166 (N_166,In_458,In_365);
nor U167 (N_167,In_251,In_293);
and U168 (N_168,In_14,In_25);
nor U169 (N_169,In_225,In_310);
xor U170 (N_170,N_10,In_387);
nor U171 (N_171,In_222,In_393);
xnor U172 (N_172,N_118,In_349);
nor U173 (N_173,N_53,In_82);
or U174 (N_174,In_196,In_68);
nor U175 (N_175,In_470,In_353);
and U176 (N_176,In_411,In_493);
nand U177 (N_177,In_494,In_129);
nor U178 (N_178,In_309,In_278);
and U179 (N_179,In_347,N_60);
xnor U180 (N_180,In_122,In_380);
and U181 (N_181,In_71,In_431);
nor U182 (N_182,In_114,N_117);
or U183 (N_183,In_342,N_38);
or U184 (N_184,In_482,In_162);
or U185 (N_185,In_32,In_311);
and U186 (N_186,N_74,In_414);
nand U187 (N_187,In_173,In_66);
and U188 (N_188,In_271,N_133);
nor U189 (N_189,In_246,In_201);
and U190 (N_190,In_301,N_69);
nor U191 (N_191,N_39,In_445);
or U192 (N_192,N_159,N_151);
nand U193 (N_193,N_3,N_166);
and U194 (N_194,In_288,N_79);
or U195 (N_195,In_111,In_191);
nand U196 (N_196,N_137,In_12);
or U197 (N_197,N_97,N_35);
nand U198 (N_198,N_141,N_158);
nand U199 (N_199,N_8,In_339);
or U200 (N_200,N_99,In_466);
and U201 (N_201,In_435,In_193);
or U202 (N_202,In_103,N_26);
nand U203 (N_203,In_436,In_124);
or U204 (N_204,In_59,N_121);
xnor U205 (N_205,In_303,In_198);
or U206 (N_206,N_104,N_170);
and U207 (N_207,In_99,In_161);
and U208 (N_208,N_132,In_292);
or U209 (N_209,N_75,In_290);
xnor U210 (N_210,N_15,N_129);
nor U211 (N_211,N_83,In_36);
xnor U212 (N_212,N_147,N_89);
nand U213 (N_213,In_108,In_280);
or U214 (N_214,In_454,N_161);
nor U215 (N_215,In_485,In_165);
xor U216 (N_216,In_26,N_98);
and U217 (N_217,N_101,In_20);
nor U218 (N_218,In_212,N_140);
nand U219 (N_219,N_59,In_438);
or U220 (N_220,N_66,In_206);
xor U221 (N_221,In_51,In_97);
nor U222 (N_222,N_90,In_2);
nand U223 (N_223,In_42,N_125);
nand U224 (N_224,N_77,N_145);
or U225 (N_225,In_307,In_43);
or U226 (N_226,In_391,N_111);
nand U227 (N_227,In_110,In_430);
nand U228 (N_228,N_144,In_335);
nor U229 (N_229,In_415,In_248);
nand U230 (N_230,In_238,In_263);
nor U231 (N_231,In_1,N_152);
nand U232 (N_232,N_1,N_164);
and U233 (N_233,In_377,N_22);
nand U234 (N_234,In_176,N_28);
nand U235 (N_235,In_421,In_226);
xnor U236 (N_236,N_138,In_298);
and U237 (N_237,N_23,In_21);
nor U238 (N_238,In_352,N_76);
or U239 (N_239,N_72,N_127);
and U240 (N_240,In_137,In_240);
nor U241 (N_241,In_446,In_313);
xnor U242 (N_242,In_490,In_267);
and U243 (N_243,N_174,N_207);
nor U244 (N_244,N_191,In_117);
or U245 (N_245,N_5,In_422);
and U246 (N_246,N_195,N_24);
or U247 (N_247,N_222,In_75);
or U248 (N_248,In_190,In_479);
and U249 (N_249,N_42,In_266);
nor U250 (N_250,In_429,In_315);
nor U251 (N_251,In_327,In_257);
nand U252 (N_252,In_276,N_169);
nand U253 (N_253,In_382,In_194);
nand U254 (N_254,N_206,N_100);
and U255 (N_255,In_167,N_136);
nand U256 (N_256,N_188,N_176);
and U257 (N_257,N_237,N_210);
nand U258 (N_258,N_115,N_229);
nand U259 (N_259,N_173,N_209);
xnor U260 (N_260,N_139,In_336);
nor U261 (N_261,N_18,N_192);
nand U262 (N_262,In_254,N_154);
nor U263 (N_263,In_96,In_413);
or U264 (N_264,N_148,In_169);
and U265 (N_265,N_185,N_155);
nand U266 (N_266,N_114,N_165);
and U267 (N_267,N_146,In_484);
nor U268 (N_268,In_128,In_166);
or U269 (N_269,N_67,In_410);
nand U270 (N_270,N_239,In_434);
or U271 (N_271,N_43,N_196);
and U272 (N_272,N_201,N_36);
nand U273 (N_273,N_202,In_369);
and U274 (N_274,N_13,In_197);
and U275 (N_275,N_216,N_96);
xnor U276 (N_276,In_274,N_234);
xnor U277 (N_277,N_219,N_182);
nor U278 (N_278,N_119,N_171);
nor U279 (N_279,In_144,N_56);
and U280 (N_280,In_183,N_197);
or U281 (N_281,In_489,In_442);
nand U282 (N_282,N_78,N_235);
or U283 (N_283,N_156,In_112);
and U284 (N_284,In_61,N_230);
xor U285 (N_285,N_93,In_73);
nor U286 (N_286,N_236,N_95);
nor U287 (N_287,N_51,N_70);
xor U288 (N_288,N_46,N_205);
xor U289 (N_289,In_299,N_168);
nor U290 (N_290,In_359,N_213);
or U291 (N_291,N_150,In_459);
or U292 (N_292,N_142,N_232);
and U293 (N_293,N_41,In_472);
or U294 (N_294,In_321,N_186);
or U295 (N_295,N_203,N_180);
nand U296 (N_296,In_164,In_424);
and U297 (N_297,N_225,In_463);
and U298 (N_298,N_40,In_13);
nand U299 (N_299,N_160,N_54);
and U300 (N_300,N_264,N_262);
nand U301 (N_301,N_178,In_49);
and U302 (N_302,In_262,In_210);
nand U303 (N_303,In_67,N_271);
nand U304 (N_304,N_143,N_265);
and U305 (N_305,In_153,N_130);
and U306 (N_306,In_323,N_228);
nor U307 (N_307,N_287,N_221);
or U308 (N_308,In_426,N_295);
or U309 (N_309,N_167,N_149);
xnor U310 (N_310,N_257,N_204);
or U311 (N_311,In_444,N_258);
or U312 (N_312,N_299,In_195);
nor U313 (N_313,In_157,N_184);
or U314 (N_314,N_263,N_120);
or U315 (N_315,N_153,In_481);
or U316 (N_316,N_208,N_162);
or U317 (N_317,N_134,In_300);
or U318 (N_318,N_102,N_172);
nor U319 (N_319,N_215,N_294);
and U320 (N_320,N_227,N_27);
xnor U321 (N_321,N_128,In_428);
nor U322 (N_322,N_157,N_268);
xnor U323 (N_323,In_252,N_286);
nor U324 (N_324,N_292,In_370);
and U325 (N_325,In_63,N_246);
and U326 (N_326,N_177,N_48);
and U327 (N_327,N_261,N_251);
or U328 (N_328,N_282,N_226);
and U329 (N_329,N_274,In_483);
nor U330 (N_330,N_279,In_449);
nor U331 (N_331,N_256,N_291);
and U332 (N_332,In_272,N_220);
and U333 (N_333,N_91,N_231);
and U334 (N_334,In_168,N_240);
nor U335 (N_335,N_58,N_20);
and U336 (N_336,N_289,N_183);
xor U337 (N_337,N_297,N_175);
and U338 (N_338,In_499,N_55);
nand U339 (N_339,N_126,In_441);
or U340 (N_340,N_298,In_87);
and U341 (N_341,In_92,N_248);
and U342 (N_342,N_87,In_384);
and U343 (N_343,N_123,N_267);
or U344 (N_344,N_243,In_116);
nand U345 (N_345,In_284,N_250);
and U346 (N_346,N_249,In_308);
and U347 (N_347,In_9,In_378);
nor U348 (N_348,N_124,N_92);
or U349 (N_349,N_193,N_181);
nor U350 (N_350,N_187,N_283);
nand U351 (N_351,In_178,N_163);
and U352 (N_352,N_272,N_290);
or U353 (N_353,In_355,N_25);
and U354 (N_354,N_212,N_223);
and U355 (N_355,N_244,In_398);
nand U356 (N_356,In_58,In_423);
nand U357 (N_357,N_200,N_135);
nor U358 (N_358,N_52,N_260);
nand U359 (N_359,In_379,N_198);
or U360 (N_360,N_259,N_314);
nor U361 (N_361,N_281,N_344);
and U362 (N_362,N_108,N_82);
or U363 (N_363,N_330,N_37);
and U364 (N_364,N_345,N_199);
nand U365 (N_365,In_351,In_486);
nor U366 (N_366,N_64,N_254);
nor U367 (N_367,In_151,N_301);
nor U368 (N_368,N_342,N_340);
nand U369 (N_369,N_332,N_321);
nor U370 (N_370,N_179,N_305);
nand U371 (N_371,N_359,N_309);
nor U372 (N_372,N_300,N_318);
or U373 (N_373,N_347,N_352);
or U374 (N_374,N_280,N_293);
and U375 (N_375,In_401,N_307);
or U376 (N_376,In_174,In_390);
nand U377 (N_377,N_61,In_228);
nor U378 (N_378,N_266,N_273);
or U379 (N_379,N_319,N_189);
nand U380 (N_380,In_492,N_4);
nand U381 (N_381,N_331,N_224);
nand U382 (N_382,N_317,N_335);
nand U383 (N_383,N_358,N_107);
nand U384 (N_384,N_326,N_308);
nor U385 (N_385,N_214,N_316);
nand U386 (N_386,N_310,N_313);
nor U387 (N_387,In_250,N_355);
nor U388 (N_388,N_349,N_306);
and U389 (N_389,N_320,N_71);
xor U390 (N_390,N_296,N_242);
xor U391 (N_391,In_160,In_143);
and U392 (N_392,N_50,N_336);
nor U393 (N_393,N_269,In_115);
nand U394 (N_394,N_339,N_312);
xor U395 (N_395,N_131,In_46);
and U396 (N_396,In_22,N_350);
nor U397 (N_397,N_194,N_245);
xor U398 (N_398,In_291,N_338);
nor U399 (N_399,N_253,N_34);
and U400 (N_400,N_238,In_346);
xnor U401 (N_401,In_451,N_343);
and U402 (N_402,In_452,N_302);
and U403 (N_403,N_278,N_354);
nor U404 (N_404,N_357,N_311);
nand U405 (N_405,N_276,In_18);
nor U406 (N_406,N_270,N_327);
or U407 (N_407,In_141,N_255);
xor U408 (N_408,N_303,N_315);
nand U409 (N_409,N_337,N_322);
nor U410 (N_410,N_190,N_275);
nand U411 (N_411,N_333,In_333);
or U412 (N_412,N_356,N_329);
nand U413 (N_413,N_247,N_241);
nor U414 (N_414,N_348,N_285);
or U415 (N_415,N_325,N_288);
and U416 (N_416,In_412,N_217);
or U417 (N_417,N_233,In_389);
or U418 (N_418,N_277,N_112);
nor U419 (N_419,In_279,N_252);
and U420 (N_420,N_122,In_29);
nand U421 (N_421,N_405,N_403);
or U422 (N_422,N_375,N_377);
and U423 (N_423,N_392,N_409);
or U424 (N_424,N_383,N_341);
nor U425 (N_425,N_397,N_390);
and U426 (N_426,N_382,N_410);
nand U427 (N_427,In_6,N_394);
xnor U428 (N_428,N_393,N_365);
nor U429 (N_429,N_398,N_401);
and U430 (N_430,N_109,N_389);
nand U431 (N_431,N_218,N_417);
nand U432 (N_432,N_391,N_395);
nand U433 (N_433,N_351,N_369);
nor U434 (N_434,N_396,N_304);
nand U435 (N_435,N_400,N_284);
xor U436 (N_436,N_371,N_361);
nor U437 (N_437,N_407,In_405);
or U438 (N_438,N_372,N_408);
or U439 (N_439,N_388,N_380);
or U440 (N_440,N_323,N_419);
nor U441 (N_441,N_411,N_402);
xnor U442 (N_442,N_211,N_363);
xnor U443 (N_443,N_399,N_386);
xnor U444 (N_444,N_360,N_416);
or U445 (N_445,N_404,N_414);
nand U446 (N_446,N_362,N_415);
nor U447 (N_447,N_376,N_324);
or U448 (N_448,N_406,N_346);
and U449 (N_449,N_412,N_418);
and U450 (N_450,In_348,N_367);
nor U451 (N_451,N_328,N_368);
or U452 (N_452,N_387,N_384);
or U453 (N_453,N_385,N_364);
nand U454 (N_454,N_374,N_334);
or U455 (N_455,In_86,N_370);
and U456 (N_456,N_353,N_366);
or U457 (N_457,N_413,N_373);
and U458 (N_458,N_378,N_381);
nor U459 (N_459,N_68,N_379);
nand U460 (N_460,N_382,N_377);
nand U461 (N_461,N_394,N_361);
or U462 (N_462,N_390,N_415);
nor U463 (N_463,N_381,N_391);
or U464 (N_464,N_404,N_409);
and U465 (N_465,N_351,N_334);
or U466 (N_466,N_416,N_328);
nor U467 (N_467,N_385,N_389);
and U468 (N_468,N_397,N_389);
nor U469 (N_469,N_364,N_386);
nor U470 (N_470,N_404,N_385);
nand U471 (N_471,N_378,N_369);
xor U472 (N_472,N_377,In_348);
and U473 (N_473,N_411,N_417);
and U474 (N_474,N_405,N_416);
xnor U475 (N_475,N_365,N_109);
nor U476 (N_476,N_413,N_386);
and U477 (N_477,N_409,N_365);
nand U478 (N_478,N_369,N_398);
nand U479 (N_479,N_411,N_412);
or U480 (N_480,N_467,N_462);
or U481 (N_481,N_439,N_465);
nand U482 (N_482,N_433,N_437);
nand U483 (N_483,N_473,N_479);
nand U484 (N_484,N_452,N_445);
nand U485 (N_485,N_444,N_453);
nor U486 (N_486,N_457,N_429);
and U487 (N_487,N_442,N_461);
xor U488 (N_488,N_460,N_470);
and U489 (N_489,N_449,N_441);
or U490 (N_490,N_458,N_464);
nand U491 (N_491,N_432,N_434);
nor U492 (N_492,N_438,N_466);
nor U493 (N_493,N_472,N_477);
nand U494 (N_494,N_450,N_456);
or U495 (N_495,N_446,N_469);
xor U496 (N_496,N_451,N_423);
and U497 (N_497,N_475,N_422);
and U498 (N_498,N_426,N_431);
xor U499 (N_499,N_448,N_430);
nor U500 (N_500,N_463,N_471);
nand U501 (N_501,N_428,N_454);
and U502 (N_502,N_468,N_440);
xor U503 (N_503,N_443,N_435);
and U504 (N_504,N_420,N_447);
nand U505 (N_505,N_424,N_455);
nand U506 (N_506,N_425,N_459);
and U507 (N_507,N_427,N_421);
and U508 (N_508,N_476,N_478);
nand U509 (N_509,N_474,N_436);
and U510 (N_510,N_469,N_479);
and U511 (N_511,N_469,N_450);
and U512 (N_512,N_465,N_445);
nand U513 (N_513,N_465,N_446);
and U514 (N_514,N_476,N_435);
nand U515 (N_515,N_430,N_424);
and U516 (N_516,N_440,N_459);
xnor U517 (N_517,N_436,N_425);
or U518 (N_518,N_456,N_468);
nand U519 (N_519,N_462,N_457);
or U520 (N_520,N_429,N_438);
and U521 (N_521,N_429,N_473);
or U522 (N_522,N_433,N_452);
xnor U523 (N_523,N_445,N_457);
nand U524 (N_524,N_443,N_440);
or U525 (N_525,N_479,N_470);
and U526 (N_526,N_464,N_472);
or U527 (N_527,N_473,N_444);
nor U528 (N_528,N_468,N_424);
nand U529 (N_529,N_465,N_455);
and U530 (N_530,N_420,N_469);
and U531 (N_531,N_448,N_438);
and U532 (N_532,N_447,N_460);
or U533 (N_533,N_427,N_462);
nand U534 (N_534,N_448,N_446);
nand U535 (N_535,N_421,N_464);
xnor U536 (N_536,N_435,N_459);
or U537 (N_537,N_479,N_436);
nand U538 (N_538,N_453,N_436);
and U539 (N_539,N_423,N_478);
nand U540 (N_540,N_536,N_506);
nor U541 (N_541,N_531,N_530);
nand U542 (N_542,N_539,N_484);
and U543 (N_543,N_511,N_491);
xor U544 (N_544,N_538,N_501);
and U545 (N_545,N_480,N_515);
and U546 (N_546,N_521,N_489);
or U547 (N_547,N_512,N_493);
nand U548 (N_548,N_482,N_492);
or U549 (N_549,N_487,N_534);
nor U550 (N_550,N_504,N_516);
nor U551 (N_551,N_537,N_522);
nor U552 (N_552,N_526,N_528);
and U553 (N_553,N_498,N_497);
nor U554 (N_554,N_486,N_525);
or U555 (N_555,N_535,N_509);
and U556 (N_556,N_481,N_510);
or U557 (N_557,N_499,N_494);
nor U558 (N_558,N_507,N_505);
and U559 (N_559,N_490,N_529);
nor U560 (N_560,N_508,N_503);
and U561 (N_561,N_519,N_483);
nand U562 (N_562,N_520,N_502);
nand U563 (N_563,N_513,N_514);
and U564 (N_564,N_523,N_485);
nand U565 (N_565,N_496,N_500);
nor U566 (N_566,N_517,N_524);
or U567 (N_567,N_488,N_518);
nand U568 (N_568,N_533,N_532);
or U569 (N_569,N_495,N_527);
xor U570 (N_570,N_514,N_539);
or U571 (N_571,N_534,N_523);
and U572 (N_572,N_518,N_524);
nor U573 (N_573,N_492,N_508);
or U574 (N_574,N_503,N_505);
and U575 (N_575,N_481,N_511);
or U576 (N_576,N_503,N_523);
nand U577 (N_577,N_537,N_528);
nand U578 (N_578,N_499,N_492);
nor U579 (N_579,N_490,N_518);
nand U580 (N_580,N_538,N_491);
nor U581 (N_581,N_515,N_535);
and U582 (N_582,N_537,N_531);
nand U583 (N_583,N_493,N_530);
nor U584 (N_584,N_515,N_527);
nor U585 (N_585,N_530,N_510);
xnor U586 (N_586,N_494,N_530);
and U587 (N_587,N_533,N_494);
nor U588 (N_588,N_524,N_490);
nor U589 (N_589,N_499,N_508);
and U590 (N_590,N_494,N_493);
or U591 (N_591,N_498,N_482);
nor U592 (N_592,N_527,N_503);
nor U593 (N_593,N_508,N_538);
nor U594 (N_594,N_525,N_504);
nor U595 (N_595,N_515,N_525);
and U596 (N_596,N_500,N_514);
nand U597 (N_597,N_530,N_514);
nand U598 (N_598,N_492,N_525);
nand U599 (N_599,N_529,N_523);
and U600 (N_600,N_554,N_596);
xor U601 (N_601,N_563,N_582);
nor U602 (N_602,N_584,N_572);
nand U603 (N_603,N_593,N_562);
xnor U604 (N_604,N_544,N_550);
nand U605 (N_605,N_595,N_568);
nand U606 (N_606,N_547,N_587);
xnor U607 (N_607,N_561,N_575);
and U608 (N_608,N_585,N_569);
or U609 (N_609,N_540,N_598);
and U610 (N_610,N_567,N_541);
nand U611 (N_611,N_565,N_591);
and U612 (N_612,N_557,N_586);
and U613 (N_613,N_588,N_576);
xnor U614 (N_614,N_597,N_549);
or U615 (N_615,N_564,N_560);
nand U616 (N_616,N_590,N_578);
and U617 (N_617,N_579,N_570);
or U618 (N_618,N_553,N_558);
xnor U619 (N_619,N_589,N_555);
or U620 (N_620,N_583,N_599);
nand U621 (N_621,N_545,N_592);
nor U622 (N_622,N_542,N_574);
nor U623 (N_623,N_543,N_594);
nand U624 (N_624,N_580,N_548);
or U625 (N_625,N_552,N_559);
or U626 (N_626,N_546,N_573);
or U627 (N_627,N_581,N_566);
or U628 (N_628,N_577,N_556);
or U629 (N_629,N_551,N_571);
and U630 (N_630,N_578,N_587);
and U631 (N_631,N_567,N_586);
nor U632 (N_632,N_552,N_598);
nor U633 (N_633,N_577,N_558);
nor U634 (N_634,N_567,N_540);
or U635 (N_635,N_573,N_590);
nand U636 (N_636,N_587,N_555);
xor U637 (N_637,N_581,N_594);
nand U638 (N_638,N_544,N_564);
and U639 (N_639,N_544,N_592);
nand U640 (N_640,N_596,N_587);
and U641 (N_641,N_550,N_574);
xnor U642 (N_642,N_542,N_571);
and U643 (N_643,N_592,N_562);
nand U644 (N_644,N_587,N_593);
nand U645 (N_645,N_564,N_547);
nor U646 (N_646,N_549,N_567);
nor U647 (N_647,N_564,N_561);
or U648 (N_648,N_589,N_541);
nand U649 (N_649,N_567,N_598);
nor U650 (N_650,N_586,N_589);
or U651 (N_651,N_548,N_561);
and U652 (N_652,N_589,N_593);
nand U653 (N_653,N_593,N_584);
and U654 (N_654,N_575,N_567);
nand U655 (N_655,N_554,N_571);
nor U656 (N_656,N_583,N_596);
nor U657 (N_657,N_541,N_578);
xor U658 (N_658,N_577,N_551);
nand U659 (N_659,N_560,N_589);
nand U660 (N_660,N_609,N_655);
and U661 (N_661,N_608,N_614);
nand U662 (N_662,N_643,N_616);
or U663 (N_663,N_640,N_623);
xor U664 (N_664,N_648,N_630);
and U665 (N_665,N_615,N_646);
and U666 (N_666,N_603,N_617);
nor U667 (N_667,N_629,N_627);
nor U668 (N_668,N_658,N_625);
nor U669 (N_669,N_620,N_631);
xor U670 (N_670,N_633,N_606);
nor U671 (N_671,N_645,N_635);
or U672 (N_672,N_602,N_610);
or U673 (N_673,N_618,N_644);
nor U674 (N_674,N_634,N_650);
or U675 (N_675,N_601,N_619);
or U676 (N_676,N_605,N_654);
nor U677 (N_677,N_612,N_628);
nor U678 (N_678,N_626,N_622);
or U679 (N_679,N_642,N_659);
nand U680 (N_680,N_649,N_613);
and U681 (N_681,N_647,N_652);
nand U682 (N_682,N_611,N_657);
nor U683 (N_683,N_653,N_636);
and U684 (N_684,N_637,N_656);
or U685 (N_685,N_638,N_604);
nand U686 (N_686,N_624,N_621);
or U687 (N_687,N_607,N_600);
and U688 (N_688,N_651,N_639);
nor U689 (N_689,N_641,N_632);
and U690 (N_690,N_657,N_608);
nand U691 (N_691,N_652,N_610);
xor U692 (N_692,N_620,N_624);
nand U693 (N_693,N_634,N_615);
and U694 (N_694,N_651,N_616);
nor U695 (N_695,N_630,N_606);
nand U696 (N_696,N_621,N_659);
nand U697 (N_697,N_605,N_633);
or U698 (N_698,N_605,N_600);
or U699 (N_699,N_623,N_637);
nand U700 (N_700,N_615,N_642);
nand U701 (N_701,N_643,N_622);
nand U702 (N_702,N_649,N_652);
xnor U703 (N_703,N_600,N_609);
or U704 (N_704,N_649,N_648);
nand U705 (N_705,N_637,N_625);
or U706 (N_706,N_600,N_637);
and U707 (N_707,N_612,N_655);
nor U708 (N_708,N_613,N_617);
and U709 (N_709,N_602,N_626);
and U710 (N_710,N_604,N_621);
or U711 (N_711,N_659,N_641);
and U712 (N_712,N_608,N_647);
and U713 (N_713,N_622,N_645);
and U714 (N_714,N_639,N_608);
and U715 (N_715,N_624,N_642);
and U716 (N_716,N_609,N_645);
nor U717 (N_717,N_613,N_614);
nor U718 (N_718,N_600,N_652);
xor U719 (N_719,N_626,N_629);
and U720 (N_720,N_708,N_668);
or U721 (N_721,N_682,N_711);
nor U722 (N_722,N_675,N_719);
nand U723 (N_723,N_667,N_685);
or U724 (N_724,N_690,N_704);
or U725 (N_725,N_705,N_709);
or U726 (N_726,N_706,N_679);
nor U727 (N_727,N_702,N_665);
nor U728 (N_728,N_686,N_714);
xnor U729 (N_729,N_663,N_662);
xnor U730 (N_730,N_694,N_681);
or U731 (N_731,N_698,N_674);
and U732 (N_732,N_717,N_707);
and U733 (N_733,N_673,N_669);
or U734 (N_734,N_677,N_660);
nor U735 (N_735,N_683,N_689);
or U736 (N_736,N_688,N_691);
or U737 (N_737,N_692,N_676);
xor U738 (N_738,N_666,N_700);
nor U739 (N_739,N_710,N_672);
or U740 (N_740,N_684,N_678);
and U741 (N_741,N_696,N_664);
and U742 (N_742,N_703,N_661);
nor U743 (N_743,N_718,N_697);
xor U744 (N_744,N_712,N_701);
or U745 (N_745,N_680,N_687);
nor U746 (N_746,N_699,N_713);
and U747 (N_747,N_670,N_695);
and U748 (N_748,N_715,N_671);
or U749 (N_749,N_693,N_716);
and U750 (N_750,N_673,N_708);
nor U751 (N_751,N_707,N_713);
or U752 (N_752,N_668,N_686);
nor U753 (N_753,N_691,N_716);
nor U754 (N_754,N_714,N_671);
nand U755 (N_755,N_707,N_660);
or U756 (N_756,N_671,N_666);
nor U757 (N_757,N_699,N_702);
xor U758 (N_758,N_710,N_661);
nand U759 (N_759,N_681,N_716);
and U760 (N_760,N_680,N_691);
and U761 (N_761,N_703,N_702);
nand U762 (N_762,N_670,N_717);
nand U763 (N_763,N_671,N_668);
or U764 (N_764,N_687,N_697);
and U765 (N_765,N_714,N_669);
nor U766 (N_766,N_661,N_673);
and U767 (N_767,N_691,N_718);
nand U768 (N_768,N_681,N_715);
nand U769 (N_769,N_680,N_688);
or U770 (N_770,N_688,N_696);
nand U771 (N_771,N_664,N_677);
nand U772 (N_772,N_671,N_673);
or U773 (N_773,N_688,N_670);
xor U774 (N_774,N_718,N_660);
nand U775 (N_775,N_716,N_692);
xor U776 (N_776,N_711,N_692);
nand U777 (N_777,N_695,N_686);
and U778 (N_778,N_698,N_679);
nor U779 (N_779,N_675,N_685);
nand U780 (N_780,N_754,N_724);
nand U781 (N_781,N_721,N_727);
or U782 (N_782,N_766,N_760);
and U783 (N_783,N_745,N_767);
nor U784 (N_784,N_776,N_758);
or U785 (N_785,N_750,N_774);
and U786 (N_786,N_746,N_756);
xor U787 (N_787,N_743,N_771);
xor U788 (N_788,N_733,N_734);
and U789 (N_789,N_777,N_757);
and U790 (N_790,N_740,N_731);
nand U791 (N_791,N_751,N_775);
xnor U792 (N_792,N_741,N_749);
and U793 (N_793,N_759,N_744);
and U794 (N_794,N_723,N_720);
and U795 (N_795,N_742,N_752);
nand U796 (N_796,N_735,N_778);
and U797 (N_797,N_769,N_728);
and U798 (N_798,N_729,N_748);
nor U799 (N_799,N_730,N_779);
nand U800 (N_800,N_722,N_773);
xor U801 (N_801,N_725,N_737);
nor U802 (N_802,N_761,N_753);
nand U803 (N_803,N_755,N_768);
or U804 (N_804,N_770,N_726);
or U805 (N_805,N_732,N_739);
and U806 (N_806,N_747,N_772);
or U807 (N_807,N_762,N_764);
nor U808 (N_808,N_765,N_763);
or U809 (N_809,N_738,N_736);
or U810 (N_810,N_741,N_731);
or U811 (N_811,N_759,N_724);
and U812 (N_812,N_753,N_768);
and U813 (N_813,N_723,N_728);
and U814 (N_814,N_772,N_746);
and U815 (N_815,N_744,N_747);
nand U816 (N_816,N_765,N_773);
and U817 (N_817,N_743,N_720);
nor U818 (N_818,N_737,N_734);
nand U819 (N_819,N_721,N_777);
and U820 (N_820,N_725,N_723);
or U821 (N_821,N_731,N_752);
or U822 (N_822,N_739,N_745);
nand U823 (N_823,N_746,N_769);
or U824 (N_824,N_733,N_725);
nor U825 (N_825,N_773,N_730);
nor U826 (N_826,N_742,N_779);
and U827 (N_827,N_721,N_765);
nor U828 (N_828,N_771,N_745);
nand U829 (N_829,N_722,N_723);
or U830 (N_830,N_750,N_779);
xnor U831 (N_831,N_737,N_771);
nor U832 (N_832,N_721,N_756);
and U833 (N_833,N_770,N_769);
and U834 (N_834,N_722,N_753);
and U835 (N_835,N_723,N_753);
xor U836 (N_836,N_755,N_758);
nand U837 (N_837,N_745,N_742);
xnor U838 (N_838,N_769,N_730);
nand U839 (N_839,N_764,N_752);
nor U840 (N_840,N_780,N_792);
or U841 (N_841,N_810,N_794);
nor U842 (N_842,N_813,N_837);
or U843 (N_843,N_799,N_805);
nand U844 (N_844,N_800,N_819);
nor U845 (N_845,N_797,N_798);
and U846 (N_846,N_826,N_785);
or U847 (N_847,N_788,N_835);
nand U848 (N_848,N_806,N_809);
nand U849 (N_849,N_823,N_828);
and U850 (N_850,N_814,N_802);
nor U851 (N_851,N_833,N_815);
or U852 (N_852,N_796,N_812);
and U853 (N_853,N_831,N_816);
nand U854 (N_854,N_827,N_808);
or U855 (N_855,N_784,N_832);
nor U856 (N_856,N_824,N_817);
nand U857 (N_857,N_793,N_821);
nor U858 (N_858,N_783,N_786);
or U859 (N_859,N_818,N_834);
xor U860 (N_860,N_790,N_804);
or U861 (N_861,N_782,N_789);
nor U862 (N_862,N_825,N_829);
xnor U863 (N_863,N_787,N_807);
and U864 (N_864,N_811,N_791);
nand U865 (N_865,N_822,N_801);
or U866 (N_866,N_820,N_838);
nand U867 (N_867,N_781,N_839);
nor U868 (N_868,N_795,N_830);
nor U869 (N_869,N_803,N_836);
and U870 (N_870,N_829,N_801);
nand U871 (N_871,N_783,N_823);
nor U872 (N_872,N_799,N_828);
nand U873 (N_873,N_811,N_801);
or U874 (N_874,N_823,N_812);
nand U875 (N_875,N_781,N_831);
xor U876 (N_876,N_792,N_819);
and U877 (N_877,N_787,N_813);
nor U878 (N_878,N_798,N_812);
nand U879 (N_879,N_829,N_822);
or U880 (N_880,N_829,N_823);
or U881 (N_881,N_831,N_792);
and U882 (N_882,N_821,N_796);
nor U883 (N_883,N_837,N_798);
nor U884 (N_884,N_782,N_797);
nor U885 (N_885,N_798,N_789);
nor U886 (N_886,N_811,N_792);
and U887 (N_887,N_829,N_833);
and U888 (N_888,N_811,N_794);
nor U889 (N_889,N_796,N_787);
xor U890 (N_890,N_801,N_817);
nor U891 (N_891,N_791,N_828);
nand U892 (N_892,N_809,N_832);
or U893 (N_893,N_792,N_816);
xor U894 (N_894,N_789,N_794);
nor U895 (N_895,N_829,N_805);
or U896 (N_896,N_833,N_822);
nor U897 (N_897,N_806,N_838);
or U898 (N_898,N_786,N_821);
or U899 (N_899,N_797,N_794);
xor U900 (N_900,N_866,N_851);
nor U901 (N_901,N_885,N_850);
nand U902 (N_902,N_845,N_858);
or U903 (N_903,N_864,N_887);
nor U904 (N_904,N_862,N_863);
and U905 (N_905,N_844,N_874);
xor U906 (N_906,N_849,N_883);
or U907 (N_907,N_893,N_856);
nor U908 (N_908,N_843,N_853);
xor U909 (N_909,N_868,N_877);
nand U910 (N_910,N_891,N_899);
and U911 (N_911,N_872,N_869);
nand U912 (N_912,N_881,N_855);
nand U913 (N_913,N_896,N_879);
nor U914 (N_914,N_870,N_890);
nand U915 (N_915,N_882,N_842);
nor U916 (N_916,N_880,N_871);
nor U917 (N_917,N_892,N_875);
or U918 (N_918,N_847,N_857);
nand U919 (N_919,N_840,N_861);
nand U920 (N_920,N_859,N_846);
or U921 (N_921,N_854,N_888);
or U922 (N_922,N_889,N_884);
and U923 (N_923,N_867,N_898);
nor U924 (N_924,N_848,N_878);
xor U925 (N_925,N_841,N_860);
nand U926 (N_926,N_895,N_865);
nand U927 (N_927,N_876,N_886);
nand U928 (N_928,N_894,N_873);
nor U929 (N_929,N_852,N_897);
nand U930 (N_930,N_850,N_894);
and U931 (N_931,N_888,N_853);
or U932 (N_932,N_843,N_899);
nand U933 (N_933,N_882,N_885);
and U934 (N_934,N_880,N_896);
nor U935 (N_935,N_843,N_858);
nor U936 (N_936,N_863,N_866);
and U937 (N_937,N_868,N_889);
nor U938 (N_938,N_842,N_856);
nor U939 (N_939,N_880,N_874);
nand U940 (N_940,N_863,N_868);
and U941 (N_941,N_884,N_859);
or U942 (N_942,N_847,N_865);
nand U943 (N_943,N_859,N_868);
or U944 (N_944,N_877,N_857);
nand U945 (N_945,N_865,N_881);
xnor U946 (N_946,N_853,N_878);
nor U947 (N_947,N_869,N_852);
xor U948 (N_948,N_889,N_857);
nor U949 (N_949,N_872,N_850);
and U950 (N_950,N_877,N_840);
nand U951 (N_951,N_852,N_864);
nand U952 (N_952,N_890,N_865);
and U953 (N_953,N_841,N_842);
and U954 (N_954,N_854,N_897);
or U955 (N_955,N_864,N_849);
nor U956 (N_956,N_895,N_859);
nor U957 (N_957,N_880,N_844);
xor U958 (N_958,N_854,N_872);
or U959 (N_959,N_884,N_863);
and U960 (N_960,N_937,N_958);
nand U961 (N_961,N_930,N_945);
or U962 (N_962,N_907,N_926);
nor U963 (N_963,N_909,N_935);
nand U964 (N_964,N_957,N_908);
or U965 (N_965,N_938,N_951);
or U966 (N_966,N_950,N_940);
and U967 (N_967,N_949,N_925);
or U968 (N_968,N_906,N_918);
nor U969 (N_969,N_944,N_956);
nand U970 (N_970,N_932,N_919);
nand U971 (N_971,N_952,N_911);
xnor U972 (N_972,N_917,N_959);
nand U973 (N_973,N_928,N_914);
or U974 (N_974,N_900,N_933);
and U975 (N_975,N_927,N_943);
nor U976 (N_976,N_934,N_905);
nand U977 (N_977,N_913,N_936);
and U978 (N_978,N_904,N_924);
nor U979 (N_979,N_903,N_912);
nor U980 (N_980,N_954,N_931);
nor U981 (N_981,N_901,N_955);
or U982 (N_982,N_902,N_948);
nor U983 (N_983,N_921,N_915);
nand U984 (N_984,N_922,N_941);
or U985 (N_985,N_910,N_946);
nor U986 (N_986,N_916,N_947);
nand U987 (N_987,N_942,N_920);
nor U988 (N_988,N_939,N_923);
nand U989 (N_989,N_929,N_953);
xor U990 (N_990,N_906,N_914);
or U991 (N_991,N_950,N_904);
and U992 (N_992,N_901,N_923);
or U993 (N_993,N_912,N_948);
nor U994 (N_994,N_934,N_909);
and U995 (N_995,N_914,N_901);
nand U996 (N_996,N_902,N_908);
nand U997 (N_997,N_954,N_959);
or U998 (N_998,N_940,N_917);
nor U999 (N_999,N_918,N_946);
and U1000 (N_1000,N_926,N_904);
nand U1001 (N_1001,N_908,N_955);
and U1002 (N_1002,N_922,N_943);
or U1003 (N_1003,N_936,N_956);
and U1004 (N_1004,N_909,N_933);
nor U1005 (N_1005,N_916,N_935);
nor U1006 (N_1006,N_938,N_949);
xnor U1007 (N_1007,N_930,N_919);
or U1008 (N_1008,N_905,N_906);
or U1009 (N_1009,N_956,N_943);
nor U1010 (N_1010,N_910,N_925);
xnor U1011 (N_1011,N_932,N_916);
nand U1012 (N_1012,N_904,N_948);
nand U1013 (N_1013,N_908,N_959);
nor U1014 (N_1014,N_919,N_908);
nor U1015 (N_1015,N_914,N_938);
and U1016 (N_1016,N_906,N_923);
nand U1017 (N_1017,N_949,N_954);
or U1018 (N_1018,N_927,N_905);
or U1019 (N_1019,N_957,N_956);
or U1020 (N_1020,N_1000,N_980);
or U1021 (N_1021,N_967,N_1001);
or U1022 (N_1022,N_986,N_977);
or U1023 (N_1023,N_962,N_963);
nor U1024 (N_1024,N_1011,N_999);
nand U1025 (N_1025,N_1012,N_966);
or U1026 (N_1026,N_1015,N_1019);
nand U1027 (N_1027,N_1007,N_975);
xnor U1028 (N_1028,N_997,N_983);
xor U1029 (N_1029,N_985,N_969);
xnor U1030 (N_1030,N_976,N_1006);
xor U1031 (N_1031,N_1009,N_972);
or U1032 (N_1032,N_1005,N_973);
or U1033 (N_1033,N_1002,N_1017);
or U1034 (N_1034,N_965,N_1010);
nor U1035 (N_1035,N_990,N_991);
and U1036 (N_1036,N_993,N_995);
and U1037 (N_1037,N_968,N_978);
and U1038 (N_1038,N_1013,N_1014);
or U1039 (N_1039,N_1008,N_971);
nor U1040 (N_1040,N_1003,N_992);
nor U1041 (N_1041,N_1004,N_961);
and U1042 (N_1042,N_994,N_964);
xnor U1043 (N_1043,N_1016,N_987);
nor U1044 (N_1044,N_970,N_974);
nand U1045 (N_1045,N_989,N_982);
or U1046 (N_1046,N_988,N_979);
nand U1047 (N_1047,N_998,N_996);
nand U1048 (N_1048,N_960,N_1018);
and U1049 (N_1049,N_984,N_981);
nor U1050 (N_1050,N_984,N_1014);
or U1051 (N_1051,N_1001,N_1009);
nand U1052 (N_1052,N_1002,N_973);
or U1053 (N_1053,N_978,N_1017);
or U1054 (N_1054,N_994,N_1017);
nor U1055 (N_1055,N_1011,N_979);
or U1056 (N_1056,N_969,N_995);
or U1057 (N_1057,N_977,N_990);
nand U1058 (N_1058,N_981,N_977);
and U1059 (N_1059,N_976,N_1017);
and U1060 (N_1060,N_996,N_960);
nand U1061 (N_1061,N_987,N_984);
and U1062 (N_1062,N_963,N_989);
nand U1063 (N_1063,N_1010,N_987);
nor U1064 (N_1064,N_966,N_1010);
or U1065 (N_1065,N_963,N_969);
nor U1066 (N_1066,N_965,N_993);
nand U1067 (N_1067,N_982,N_992);
and U1068 (N_1068,N_1019,N_1000);
and U1069 (N_1069,N_985,N_986);
nor U1070 (N_1070,N_1009,N_1013);
or U1071 (N_1071,N_978,N_985);
nor U1072 (N_1072,N_1005,N_965);
nor U1073 (N_1073,N_1004,N_975);
nor U1074 (N_1074,N_988,N_962);
or U1075 (N_1075,N_983,N_988);
xnor U1076 (N_1076,N_1011,N_1018);
and U1077 (N_1077,N_972,N_973);
nor U1078 (N_1078,N_966,N_1016);
nor U1079 (N_1079,N_960,N_991);
xnor U1080 (N_1080,N_1063,N_1040);
nand U1081 (N_1081,N_1025,N_1071);
nand U1082 (N_1082,N_1038,N_1059);
nand U1083 (N_1083,N_1026,N_1045);
or U1084 (N_1084,N_1069,N_1041);
and U1085 (N_1085,N_1078,N_1053);
or U1086 (N_1086,N_1022,N_1079);
or U1087 (N_1087,N_1034,N_1021);
and U1088 (N_1088,N_1029,N_1070);
nor U1089 (N_1089,N_1051,N_1030);
nor U1090 (N_1090,N_1048,N_1077);
nor U1091 (N_1091,N_1046,N_1060);
or U1092 (N_1092,N_1031,N_1054);
nand U1093 (N_1093,N_1074,N_1028);
nor U1094 (N_1094,N_1047,N_1036);
nor U1095 (N_1095,N_1064,N_1073);
nand U1096 (N_1096,N_1044,N_1032);
and U1097 (N_1097,N_1052,N_1076);
nor U1098 (N_1098,N_1075,N_1068);
nand U1099 (N_1099,N_1027,N_1049);
nor U1100 (N_1100,N_1056,N_1023);
and U1101 (N_1101,N_1043,N_1042);
or U1102 (N_1102,N_1065,N_1039);
nor U1103 (N_1103,N_1062,N_1020);
nor U1104 (N_1104,N_1061,N_1058);
and U1105 (N_1105,N_1066,N_1055);
nor U1106 (N_1106,N_1057,N_1037);
nor U1107 (N_1107,N_1035,N_1067);
or U1108 (N_1108,N_1024,N_1033);
nor U1109 (N_1109,N_1072,N_1050);
nor U1110 (N_1110,N_1073,N_1041);
nor U1111 (N_1111,N_1050,N_1056);
or U1112 (N_1112,N_1040,N_1035);
and U1113 (N_1113,N_1030,N_1057);
nor U1114 (N_1114,N_1067,N_1061);
nor U1115 (N_1115,N_1063,N_1020);
nor U1116 (N_1116,N_1041,N_1051);
or U1117 (N_1117,N_1046,N_1041);
and U1118 (N_1118,N_1032,N_1028);
or U1119 (N_1119,N_1072,N_1023);
or U1120 (N_1120,N_1046,N_1067);
nand U1121 (N_1121,N_1021,N_1048);
and U1122 (N_1122,N_1038,N_1079);
nand U1123 (N_1123,N_1049,N_1048);
nand U1124 (N_1124,N_1065,N_1023);
nor U1125 (N_1125,N_1049,N_1054);
or U1126 (N_1126,N_1020,N_1022);
and U1127 (N_1127,N_1052,N_1079);
nor U1128 (N_1128,N_1078,N_1027);
and U1129 (N_1129,N_1056,N_1026);
nor U1130 (N_1130,N_1032,N_1072);
or U1131 (N_1131,N_1069,N_1062);
or U1132 (N_1132,N_1066,N_1051);
nor U1133 (N_1133,N_1070,N_1047);
and U1134 (N_1134,N_1055,N_1073);
or U1135 (N_1135,N_1021,N_1046);
nand U1136 (N_1136,N_1025,N_1052);
and U1137 (N_1137,N_1044,N_1026);
or U1138 (N_1138,N_1067,N_1040);
nor U1139 (N_1139,N_1053,N_1030);
nor U1140 (N_1140,N_1113,N_1106);
nand U1141 (N_1141,N_1128,N_1133);
and U1142 (N_1142,N_1111,N_1096);
nand U1143 (N_1143,N_1130,N_1132);
nor U1144 (N_1144,N_1087,N_1129);
or U1145 (N_1145,N_1104,N_1083);
and U1146 (N_1146,N_1095,N_1136);
nor U1147 (N_1147,N_1135,N_1108);
or U1148 (N_1148,N_1137,N_1086);
or U1149 (N_1149,N_1120,N_1085);
nand U1150 (N_1150,N_1126,N_1121);
nor U1151 (N_1151,N_1114,N_1105);
xnor U1152 (N_1152,N_1088,N_1102);
nand U1153 (N_1153,N_1082,N_1080);
xor U1154 (N_1154,N_1101,N_1123);
nor U1155 (N_1155,N_1100,N_1138);
xor U1156 (N_1156,N_1116,N_1122);
xor U1157 (N_1157,N_1112,N_1091);
nand U1158 (N_1158,N_1117,N_1115);
or U1159 (N_1159,N_1127,N_1118);
or U1160 (N_1160,N_1099,N_1092);
or U1161 (N_1161,N_1107,N_1093);
nand U1162 (N_1162,N_1131,N_1098);
and U1163 (N_1163,N_1109,N_1097);
nor U1164 (N_1164,N_1124,N_1094);
xor U1165 (N_1165,N_1139,N_1119);
and U1166 (N_1166,N_1081,N_1134);
or U1167 (N_1167,N_1110,N_1089);
or U1168 (N_1168,N_1103,N_1090);
nor U1169 (N_1169,N_1125,N_1084);
and U1170 (N_1170,N_1083,N_1123);
or U1171 (N_1171,N_1138,N_1139);
nand U1172 (N_1172,N_1115,N_1099);
or U1173 (N_1173,N_1135,N_1118);
xor U1174 (N_1174,N_1101,N_1080);
nand U1175 (N_1175,N_1100,N_1129);
and U1176 (N_1176,N_1087,N_1120);
nand U1177 (N_1177,N_1088,N_1134);
nor U1178 (N_1178,N_1083,N_1137);
nand U1179 (N_1179,N_1130,N_1115);
and U1180 (N_1180,N_1105,N_1095);
nor U1181 (N_1181,N_1112,N_1127);
or U1182 (N_1182,N_1094,N_1126);
nand U1183 (N_1183,N_1102,N_1108);
xnor U1184 (N_1184,N_1102,N_1124);
and U1185 (N_1185,N_1084,N_1131);
and U1186 (N_1186,N_1115,N_1134);
nand U1187 (N_1187,N_1089,N_1138);
nand U1188 (N_1188,N_1101,N_1112);
or U1189 (N_1189,N_1104,N_1088);
and U1190 (N_1190,N_1097,N_1135);
xnor U1191 (N_1191,N_1117,N_1108);
and U1192 (N_1192,N_1100,N_1110);
and U1193 (N_1193,N_1084,N_1117);
nand U1194 (N_1194,N_1100,N_1093);
and U1195 (N_1195,N_1112,N_1106);
and U1196 (N_1196,N_1133,N_1086);
xor U1197 (N_1197,N_1131,N_1132);
nand U1198 (N_1198,N_1089,N_1130);
xnor U1199 (N_1199,N_1099,N_1131);
and U1200 (N_1200,N_1156,N_1181);
and U1201 (N_1201,N_1168,N_1154);
nand U1202 (N_1202,N_1191,N_1147);
nand U1203 (N_1203,N_1159,N_1193);
or U1204 (N_1204,N_1174,N_1183);
xnor U1205 (N_1205,N_1184,N_1176);
nand U1206 (N_1206,N_1195,N_1175);
and U1207 (N_1207,N_1149,N_1165);
or U1208 (N_1208,N_1150,N_1167);
nand U1209 (N_1209,N_1171,N_1164);
and U1210 (N_1210,N_1148,N_1197);
nand U1211 (N_1211,N_1199,N_1186);
xor U1212 (N_1212,N_1151,N_1163);
nor U1213 (N_1213,N_1194,N_1141);
nor U1214 (N_1214,N_1157,N_1153);
nand U1215 (N_1215,N_1196,N_1145);
nor U1216 (N_1216,N_1169,N_1192);
xor U1217 (N_1217,N_1161,N_1162);
and U1218 (N_1218,N_1189,N_1143);
and U1219 (N_1219,N_1198,N_1178);
nand U1220 (N_1220,N_1188,N_1144);
and U1221 (N_1221,N_1160,N_1177);
or U1222 (N_1222,N_1182,N_1172);
nand U1223 (N_1223,N_1152,N_1179);
nor U1224 (N_1224,N_1190,N_1155);
nand U1225 (N_1225,N_1170,N_1142);
and U1226 (N_1226,N_1173,N_1187);
nand U1227 (N_1227,N_1166,N_1180);
nand U1228 (N_1228,N_1146,N_1158);
nor U1229 (N_1229,N_1185,N_1140);
nand U1230 (N_1230,N_1145,N_1160);
nor U1231 (N_1231,N_1148,N_1150);
and U1232 (N_1232,N_1155,N_1148);
nor U1233 (N_1233,N_1146,N_1195);
nor U1234 (N_1234,N_1147,N_1145);
or U1235 (N_1235,N_1199,N_1193);
or U1236 (N_1236,N_1172,N_1190);
and U1237 (N_1237,N_1192,N_1159);
and U1238 (N_1238,N_1168,N_1153);
nor U1239 (N_1239,N_1149,N_1151);
or U1240 (N_1240,N_1170,N_1145);
nand U1241 (N_1241,N_1158,N_1170);
xnor U1242 (N_1242,N_1145,N_1154);
and U1243 (N_1243,N_1187,N_1174);
and U1244 (N_1244,N_1179,N_1180);
nor U1245 (N_1245,N_1192,N_1195);
nor U1246 (N_1246,N_1142,N_1174);
xor U1247 (N_1247,N_1179,N_1188);
nand U1248 (N_1248,N_1179,N_1197);
nor U1249 (N_1249,N_1182,N_1143);
and U1250 (N_1250,N_1146,N_1190);
nor U1251 (N_1251,N_1192,N_1170);
nor U1252 (N_1252,N_1165,N_1144);
and U1253 (N_1253,N_1189,N_1173);
nor U1254 (N_1254,N_1143,N_1150);
nor U1255 (N_1255,N_1183,N_1156);
nand U1256 (N_1256,N_1156,N_1145);
and U1257 (N_1257,N_1188,N_1160);
xnor U1258 (N_1258,N_1160,N_1174);
nor U1259 (N_1259,N_1161,N_1146);
and U1260 (N_1260,N_1202,N_1236);
or U1261 (N_1261,N_1247,N_1256);
nand U1262 (N_1262,N_1203,N_1206);
or U1263 (N_1263,N_1238,N_1220);
nor U1264 (N_1264,N_1234,N_1241);
nor U1265 (N_1265,N_1246,N_1233);
nand U1266 (N_1266,N_1222,N_1215);
and U1267 (N_1267,N_1210,N_1227);
and U1268 (N_1268,N_1218,N_1212);
nand U1269 (N_1269,N_1253,N_1205);
and U1270 (N_1270,N_1243,N_1245);
and U1271 (N_1271,N_1255,N_1211);
nand U1272 (N_1272,N_1250,N_1225);
or U1273 (N_1273,N_1221,N_1209);
and U1274 (N_1274,N_1240,N_1231);
and U1275 (N_1275,N_1200,N_1214);
xor U1276 (N_1276,N_1248,N_1251);
xnor U1277 (N_1277,N_1242,N_1239);
nand U1278 (N_1278,N_1223,N_1213);
and U1279 (N_1279,N_1219,N_1244);
and U1280 (N_1280,N_1259,N_1232);
nor U1281 (N_1281,N_1229,N_1252);
nand U1282 (N_1282,N_1207,N_1228);
and U1283 (N_1283,N_1249,N_1230);
nand U1284 (N_1284,N_1208,N_1201);
and U1285 (N_1285,N_1216,N_1237);
and U1286 (N_1286,N_1235,N_1254);
nor U1287 (N_1287,N_1204,N_1217);
and U1288 (N_1288,N_1257,N_1224);
and U1289 (N_1289,N_1258,N_1226);
nor U1290 (N_1290,N_1215,N_1250);
nor U1291 (N_1291,N_1219,N_1216);
nor U1292 (N_1292,N_1216,N_1207);
xor U1293 (N_1293,N_1234,N_1233);
or U1294 (N_1294,N_1246,N_1206);
xnor U1295 (N_1295,N_1222,N_1216);
or U1296 (N_1296,N_1200,N_1238);
nor U1297 (N_1297,N_1252,N_1212);
nor U1298 (N_1298,N_1232,N_1219);
nor U1299 (N_1299,N_1230,N_1240);
and U1300 (N_1300,N_1241,N_1223);
xnor U1301 (N_1301,N_1234,N_1210);
or U1302 (N_1302,N_1213,N_1210);
nor U1303 (N_1303,N_1217,N_1256);
and U1304 (N_1304,N_1228,N_1232);
nor U1305 (N_1305,N_1220,N_1250);
or U1306 (N_1306,N_1235,N_1249);
and U1307 (N_1307,N_1211,N_1231);
and U1308 (N_1308,N_1236,N_1254);
or U1309 (N_1309,N_1214,N_1239);
nand U1310 (N_1310,N_1214,N_1233);
or U1311 (N_1311,N_1235,N_1200);
nand U1312 (N_1312,N_1200,N_1227);
nor U1313 (N_1313,N_1202,N_1228);
nor U1314 (N_1314,N_1214,N_1250);
or U1315 (N_1315,N_1211,N_1247);
nand U1316 (N_1316,N_1211,N_1213);
nor U1317 (N_1317,N_1245,N_1217);
and U1318 (N_1318,N_1219,N_1237);
nor U1319 (N_1319,N_1220,N_1232);
and U1320 (N_1320,N_1317,N_1300);
nor U1321 (N_1321,N_1301,N_1277);
nor U1322 (N_1322,N_1308,N_1261);
nor U1323 (N_1323,N_1311,N_1278);
nand U1324 (N_1324,N_1292,N_1318);
and U1325 (N_1325,N_1295,N_1279);
and U1326 (N_1326,N_1265,N_1298);
and U1327 (N_1327,N_1306,N_1299);
nand U1328 (N_1328,N_1316,N_1313);
and U1329 (N_1329,N_1266,N_1309);
or U1330 (N_1330,N_1304,N_1283);
nand U1331 (N_1331,N_1273,N_1269);
nor U1332 (N_1332,N_1267,N_1281);
nand U1333 (N_1333,N_1268,N_1275);
nand U1334 (N_1334,N_1312,N_1280);
or U1335 (N_1335,N_1260,N_1284);
nand U1336 (N_1336,N_1307,N_1286);
and U1337 (N_1337,N_1288,N_1263);
nor U1338 (N_1338,N_1282,N_1287);
nand U1339 (N_1339,N_1271,N_1315);
nor U1340 (N_1340,N_1302,N_1303);
and U1341 (N_1341,N_1314,N_1293);
and U1342 (N_1342,N_1264,N_1270);
or U1343 (N_1343,N_1291,N_1276);
and U1344 (N_1344,N_1272,N_1305);
xor U1345 (N_1345,N_1262,N_1290);
xor U1346 (N_1346,N_1296,N_1289);
nor U1347 (N_1347,N_1319,N_1285);
nor U1348 (N_1348,N_1294,N_1310);
or U1349 (N_1349,N_1274,N_1297);
xnor U1350 (N_1350,N_1289,N_1317);
nand U1351 (N_1351,N_1263,N_1260);
or U1352 (N_1352,N_1300,N_1262);
or U1353 (N_1353,N_1289,N_1287);
nor U1354 (N_1354,N_1295,N_1316);
nor U1355 (N_1355,N_1303,N_1273);
and U1356 (N_1356,N_1261,N_1310);
or U1357 (N_1357,N_1293,N_1263);
or U1358 (N_1358,N_1296,N_1278);
and U1359 (N_1359,N_1287,N_1283);
nand U1360 (N_1360,N_1296,N_1275);
nor U1361 (N_1361,N_1280,N_1272);
or U1362 (N_1362,N_1270,N_1287);
nand U1363 (N_1363,N_1298,N_1273);
nand U1364 (N_1364,N_1262,N_1315);
or U1365 (N_1365,N_1277,N_1267);
nor U1366 (N_1366,N_1265,N_1301);
nand U1367 (N_1367,N_1296,N_1271);
nand U1368 (N_1368,N_1266,N_1298);
or U1369 (N_1369,N_1263,N_1277);
nor U1370 (N_1370,N_1285,N_1296);
nor U1371 (N_1371,N_1275,N_1287);
and U1372 (N_1372,N_1318,N_1260);
xor U1373 (N_1373,N_1317,N_1301);
or U1374 (N_1374,N_1284,N_1283);
nor U1375 (N_1375,N_1272,N_1269);
or U1376 (N_1376,N_1288,N_1299);
xnor U1377 (N_1377,N_1260,N_1309);
nor U1378 (N_1378,N_1303,N_1271);
or U1379 (N_1379,N_1301,N_1267);
or U1380 (N_1380,N_1377,N_1364);
nand U1381 (N_1381,N_1323,N_1351);
or U1382 (N_1382,N_1369,N_1354);
nand U1383 (N_1383,N_1334,N_1336);
nand U1384 (N_1384,N_1376,N_1347);
nor U1385 (N_1385,N_1345,N_1322);
nand U1386 (N_1386,N_1325,N_1329);
and U1387 (N_1387,N_1324,N_1365);
nor U1388 (N_1388,N_1338,N_1367);
xnor U1389 (N_1389,N_1356,N_1320);
or U1390 (N_1390,N_1344,N_1363);
or U1391 (N_1391,N_1371,N_1366);
and U1392 (N_1392,N_1339,N_1346);
xnor U1393 (N_1393,N_1360,N_1352);
nor U1394 (N_1394,N_1330,N_1337);
or U1395 (N_1395,N_1321,N_1373);
xor U1396 (N_1396,N_1357,N_1362);
nand U1397 (N_1397,N_1350,N_1368);
nand U1398 (N_1398,N_1359,N_1331);
or U1399 (N_1399,N_1361,N_1327);
and U1400 (N_1400,N_1326,N_1374);
or U1401 (N_1401,N_1379,N_1335);
and U1402 (N_1402,N_1372,N_1343);
nand U1403 (N_1403,N_1340,N_1348);
and U1404 (N_1404,N_1332,N_1370);
nand U1405 (N_1405,N_1328,N_1378);
or U1406 (N_1406,N_1341,N_1333);
and U1407 (N_1407,N_1355,N_1358);
nand U1408 (N_1408,N_1375,N_1353);
xnor U1409 (N_1409,N_1342,N_1349);
nand U1410 (N_1410,N_1353,N_1359);
nor U1411 (N_1411,N_1334,N_1376);
nand U1412 (N_1412,N_1337,N_1367);
nand U1413 (N_1413,N_1366,N_1360);
or U1414 (N_1414,N_1332,N_1362);
nand U1415 (N_1415,N_1346,N_1320);
xnor U1416 (N_1416,N_1375,N_1344);
and U1417 (N_1417,N_1342,N_1336);
and U1418 (N_1418,N_1331,N_1353);
xor U1419 (N_1419,N_1348,N_1352);
nor U1420 (N_1420,N_1341,N_1345);
or U1421 (N_1421,N_1369,N_1367);
or U1422 (N_1422,N_1337,N_1328);
xnor U1423 (N_1423,N_1350,N_1348);
or U1424 (N_1424,N_1370,N_1342);
or U1425 (N_1425,N_1378,N_1340);
nor U1426 (N_1426,N_1352,N_1347);
xnor U1427 (N_1427,N_1369,N_1331);
or U1428 (N_1428,N_1342,N_1367);
or U1429 (N_1429,N_1334,N_1378);
nor U1430 (N_1430,N_1354,N_1344);
nand U1431 (N_1431,N_1341,N_1340);
xor U1432 (N_1432,N_1350,N_1331);
nand U1433 (N_1433,N_1376,N_1353);
nand U1434 (N_1434,N_1352,N_1331);
nand U1435 (N_1435,N_1351,N_1341);
or U1436 (N_1436,N_1369,N_1368);
or U1437 (N_1437,N_1322,N_1321);
and U1438 (N_1438,N_1346,N_1372);
nor U1439 (N_1439,N_1364,N_1351);
xnor U1440 (N_1440,N_1389,N_1417);
nand U1441 (N_1441,N_1407,N_1388);
nor U1442 (N_1442,N_1434,N_1435);
or U1443 (N_1443,N_1381,N_1432);
and U1444 (N_1444,N_1409,N_1396);
nand U1445 (N_1445,N_1433,N_1419);
or U1446 (N_1446,N_1382,N_1393);
xnor U1447 (N_1447,N_1415,N_1424);
or U1448 (N_1448,N_1383,N_1384);
and U1449 (N_1449,N_1427,N_1431);
nand U1450 (N_1450,N_1385,N_1413);
nand U1451 (N_1451,N_1399,N_1423);
and U1452 (N_1452,N_1400,N_1436);
and U1453 (N_1453,N_1416,N_1408);
and U1454 (N_1454,N_1426,N_1410);
nor U1455 (N_1455,N_1397,N_1404);
or U1456 (N_1456,N_1390,N_1395);
nor U1457 (N_1457,N_1414,N_1402);
or U1458 (N_1458,N_1391,N_1422);
or U1459 (N_1459,N_1401,N_1428);
nor U1460 (N_1460,N_1420,N_1429);
xnor U1461 (N_1461,N_1406,N_1418);
and U1462 (N_1462,N_1387,N_1425);
and U1463 (N_1463,N_1439,N_1412);
nand U1464 (N_1464,N_1392,N_1394);
nand U1465 (N_1465,N_1405,N_1398);
nand U1466 (N_1466,N_1386,N_1437);
or U1467 (N_1467,N_1403,N_1380);
or U1468 (N_1468,N_1411,N_1438);
and U1469 (N_1469,N_1430,N_1421);
nand U1470 (N_1470,N_1429,N_1434);
nor U1471 (N_1471,N_1396,N_1406);
nor U1472 (N_1472,N_1407,N_1416);
nor U1473 (N_1473,N_1420,N_1387);
nor U1474 (N_1474,N_1396,N_1398);
and U1475 (N_1475,N_1423,N_1403);
and U1476 (N_1476,N_1395,N_1392);
nor U1477 (N_1477,N_1427,N_1411);
and U1478 (N_1478,N_1423,N_1404);
xnor U1479 (N_1479,N_1404,N_1389);
and U1480 (N_1480,N_1439,N_1405);
nor U1481 (N_1481,N_1399,N_1411);
nor U1482 (N_1482,N_1394,N_1400);
nor U1483 (N_1483,N_1390,N_1427);
and U1484 (N_1484,N_1421,N_1412);
nand U1485 (N_1485,N_1431,N_1422);
nor U1486 (N_1486,N_1424,N_1380);
nor U1487 (N_1487,N_1408,N_1422);
nand U1488 (N_1488,N_1429,N_1386);
or U1489 (N_1489,N_1432,N_1438);
nand U1490 (N_1490,N_1385,N_1397);
nand U1491 (N_1491,N_1394,N_1387);
nand U1492 (N_1492,N_1403,N_1412);
nor U1493 (N_1493,N_1425,N_1422);
nor U1494 (N_1494,N_1439,N_1430);
nand U1495 (N_1495,N_1421,N_1385);
nand U1496 (N_1496,N_1397,N_1438);
and U1497 (N_1497,N_1432,N_1398);
and U1498 (N_1498,N_1422,N_1388);
and U1499 (N_1499,N_1393,N_1436);
or U1500 (N_1500,N_1498,N_1492);
or U1501 (N_1501,N_1493,N_1468);
nor U1502 (N_1502,N_1450,N_1477);
and U1503 (N_1503,N_1496,N_1489);
nor U1504 (N_1504,N_1453,N_1469);
nand U1505 (N_1505,N_1466,N_1451);
or U1506 (N_1506,N_1480,N_1471);
or U1507 (N_1507,N_1476,N_1486);
nand U1508 (N_1508,N_1481,N_1454);
and U1509 (N_1509,N_1457,N_1452);
xnor U1510 (N_1510,N_1499,N_1485);
nor U1511 (N_1511,N_1473,N_1487);
and U1512 (N_1512,N_1483,N_1478);
or U1513 (N_1513,N_1475,N_1467);
and U1514 (N_1514,N_1488,N_1440);
xor U1515 (N_1515,N_1456,N_1444);
and U1516 (N_1516,N_1455,N_1462);
nor U1517 (N_1517,N_1446,N_1445);
nor U1518 (N_1518,N_1494,N_1463);
and U1519 (N_1519,N_1490,N_1447);
nor U1520 (N_1520,N_1474,N_1442);
or U1521 (N_1521,N_1448,N_1495);
nand U1522 (N_1522,N_1443,N_1461);
nor U1523 (N_1523,N_1460,N_1491);
nand U1524 (N_1524,N_1470,N_1472);
and U1525 (N_1525,N_1465,N_1464);
and U1526 (N_1526,N_1458,N_1449);
or U1527 (N_1527,N_1482,N_1459);
xor U1528 (N_1528,N_1441,N_1479);
nand U1529 (N_1529,N_1484,N_1497);
nand U1530 (N_1530,N_1483,N_1466);
xor U1531 (N_1531,N_1478,N_1445);
nand U1532 (N_1532,N_1440,N_1467);
nor U1533 (N_1533,N_1466,N_1473);
and U1534 (N_1534,N_1447,N_1465);
or U1535 (N_1535,N_1475,N_1480);
xnor U1536 (N_1536,N_1449,N_1473);
nor U1537 (N_1537,N_1486,N_1453);
nor U1538 (N_1538,N_1499,N_1470);
nand U1539 (N_1539,N_1451,N_1491);
nor U1540 (N_1540,N_1466,N_1457);
or U1541 (N_1541,N_1481,N_1496);
or U1542 (N_1542,N_1462,N_1488);
nor U1543 (N_1543,N_1482,N_1481);
nor U1544 (N_1544,N_1441,N_1486);
nand U1545 (N_1545,N_1451,N_1485);
nand U1546 (N_1546,N_1451,N_1462);
or U1547 (N_1547,N_1463,N_1493);
and U1548 (N_1548,N_1499,N_1480);
xor U1549 (N_1549,N_1480,N_1450);
or U1550 (N_1550,N_1464,N_1480);
nor U1551 (N_1551,N_1456,N_1446);
xnor U1552 (N_1552,N_1465,N_1493);
nor U1553 (N_1553,N_1448,N_1476);
or U1554 (N_1554,N_1460,N_1465);
nand U1555 (N_1555,N_1493,N_1443);
nor U1556 (N_1556,N_1458,N_1476);
nor U1557 (N_1557,N_1486,N_1495);
xnor U1558 (N_1558,N_1492,N_1483);
nand U1559 (N_1559,N_1450,N_1481);
nand U1560 (N_1560,N_1516,N_1517);
and U1561 (N_1561,N_1506,N_1514);
nand U1562 (N_1562,N_1528,N_1515);
nor U1563 (N_1563,N_1541,N_1518);
xor U1564 (N_1564,N_1508,N_1525);
nand U1565 (N_1565,N_1556,N_1533);
and U1566 (N_1566,N_1552,N_1546);
nand U1567 (N_1567,N_1548,N_1531);
and U1568 (N_1568,N_1536,N_1526);
nor U1569 (N_1569,N_1554,N_1523);
xor U1570 (N_1570,N_1555,N_1527);
and U1571 (N_1571,N_1524,N_1513);
or U1572 (N_1572,N_1509,N_1503);
and U1573 (N_1573,N_1539,N_1540);
nor U1574 (N_1574,N_1545,N_1547);
nand U1575 (N_1575,N_1504,N_1542);
or U1576 (N_1576,N_1519,N_1532);
and U1577 (N_1577,N_1511,N_1501);
and U1578 (N_1578,N_1558,N_1507);
and U1579 (N_1579,N_1535,N_1549);
and U1580 (N_1580,N_1550,N_1521);
or U1581 (N_1581,N_1544,N_1529);
nand U1582 (N_1582,N_1538,N_1534);
nand U1583 (N_1583,N_1512,N_1505);
nand U1584 (N_1584,N_1510,N_1543);
nand U1585 (N_1585,N_1553,N_1520);
nor U1586 (N_1586,N_1522,N_1537);
and U1587 (N_1587,N_1551,N_1500);
xor U1588 (N_1588,N_1502,N_1559);
xor U1589 (N_1589,N_1530,N_1557);
xor U1590 (N_1590,N_1523,N_1537);
or U1591 (N_1591,N_1501,N_1510);
or U1592 (N_1592,N_1549,N_1508);
and U1593 (N_1593,N_1526,N_1538);
and U1594 (N_1594,N_1551,N_1512);
xor U1595 (N_1595,N_1529,N_1535);
xor U1596 (N_1596,N_1537,N_1546);
nor U1597 (N_1597,N_1528,N_1555);
xor U1598 (N_1598,N_1517,N_1509);
or U1599 (N_1599,N_1512,N_1534);
nor U1600 (N_1600,N_1530,N_1552);
xnor U1601 (N_1601,N_1554,N_1526);
and U1602 (N_1602,N_1508,N_1559);
nand U1603 (N_1603,N_1511,N_1547);
and U1604 (N_1604,N_1539,N_1538);
nand U1605 (N_1605,N_1523,N_1544);
nor U1606 (N_1606,N_1516,N_1538);
nand U1607 (N_1607,N_1533,N_1501);
or U1608 (N_1608,N_1550,N_1507);
or U1609 (N_1609,N_1537,N_1513);
nand U1610 (N_1610,N_1507,N_1515);
xnor U1611 (N_1611,N_1508,N_1521);
xnor U1612 (N_1612,N_1507,N_1541);
nor U1613 (N_1613,N_1525,N_1548);
or U1614 (N_1614,N_1534,N_1539);
nand U1615 (N_1615,N_1548,N_1521);
xnor U1616 (N_1616,N_1527,N_1549);
and U1617 (N_1617,N_1518,N_1532);
nand U1618 (N_1618,N_1513,N_1526);
or U1619 (N_1619,N_1551,N_1531);
or U1620 (N_1620,N_1587,N_1568);
nand U1621 (N_1621,N_1605,N_1564);
or U1622 (N_1622,N_1574,N_1601);
or U1623 (N_1623,N_1610,N_1583);
and U1624 (N_1624,N_1565,N_1592);
xor U1625 (N_1625,N_1613,N_1595);
or U1626 (N_1626,N_1575,N_1563);
or U1627 (N_1627,N_1617,N_1566);
and U1628 (N_1628,N_1593,N_1599);
and U1629 (N_1629,N_1591,N_1609);
nor U1630 (N_1630,N_1604,N_1608);
xnor U1631 (N_1631,N_1615,N_1612);
and U1632 (N_1632,N_1619,N_1561);
nand U1633 (N_1633,N_1584,N_1562);
and U1634 (N_1634,N_1569,N_1600);
nand U1635 (N_1635,N_1576,N_1606);
and U1636 (N_1636,N_1572,N_1567);
or U1637 (N_1637,N_1607,N_1586);
xor U1638 (N_1638,N_1580,N_1594);
or U1639 (N_1639,N_1614,N_1618);
and U1640 (N_1640,N_1588,N_1579);
xnor U1641 (N_1641,N_1602,N_1571);
nor U1642 (N_1642,N_1598,N_1560);
nor U1643 (N_1643,N_1611,N_1597);
nor U1644 (N_1644,N_1603,N_1590);
xor U1645 (N_1645,N_1585,N_1581);
and U1646 (N_1646,N_1577,N_1573);
nor U1647 (N_1647,N_1578,N_1570);
nand U1648 (N_1648,N_1596,N_1582);
or U1649 (N_1649,N_1589,N_1616);
nand U1650 (N_1650,N_1583,N_1586);
nand U1651 (N_1651,N_1617,N_1590);
nor U1652 (N_1652,N_1580,N_1561);
xnor U1653 (N_1653,N_1564,N_1582);
xor U1654 (N_1654,N_1604,N_1616);
nor U1655 (N_1655,N_1615,N_1594);
or U1656 (N_1656,N_1577,N_1599);
or U1657 (N_1657,N_1598,N_1602);
or U1658 (N_1658,N_1575,N_1592);
nand U1659 (N_1659,N_1597,N_1582);
nor U1660 (N_1660,N_1614,N_1580);
and U1661 (N_1661,N_1619,N_1609);
or U1662 (N_1662,N_1581,N_1608);
or U1663 (N_1663,N_1588,N_1616);
and U1664 (N_1664,N_1609,N_1602);
nand U1665 (N_1665,N_1572,N_1609);
or U1666 (N_1666,N_1575,N_1576);
xor U1667 (N_1667,N_1599,N_1605);
nor U1668 (N_1668,N_1602,N_1582);
nand U1669 (N_1669,N_1619,N_1578);
and U1670 (N_1670,N_1599,N_1616);
nor U1671 (N_1671,N_1568,N_1591);
nand U1672 (N_1672,N_1594,N_1608);
nor U1673 (N_1673,N_1590,N_1598);
nor U1674 (N_1674,N_1583,N_1564);
nor U1675 (N_1675,N_1563,N_1617);
nand U1676 (N_1676,N_1613,N_1561);
and U1677 (N_1677,N_1574,N_1596);
xor U1678 (N_1678,N_1605,N_1596);
xor U1679 (N_1679,N_1571,N_1616);
nand U1680 (N_1680,N_1659,N_1653);
and U1681 (N_1681,N_1644,N_1679);
nand U1682 (N_1682,N_1669,N_1677);
xor U1683 (N_1683,N_1662,N_1664);
or U1684 (N_1684,N_1646,N_1672);
or U1685 (N_1685,N_1642,N_1636);
nand U1686 (N_1686,N_1660,N_1633);
and U1687 (N_1687,N_1622,N_1621);
nand U1688 (N_1688,N_1638,N_1626);
and U1689 (N_1689,N_1651,N_1668);
nor U1690 (N_1690,N_1674,N_1661);
and U1691 (N_1691,N_1673,N_1649);
or U1692 (N_1692,N_1654,N_1657);
nand U1693 (N_1693,N_1665,N_1620);
nor U1694 (N_1694,N_1648,N_1627);
or U1695 (N_1695,N_1666,N_1634);
and U1696 (N_1696,N_1624,N_1623);
nor U1697 (N_1697,N_1631,N_1645);
nor U1698 (N_1698,N_1641,N_1663);
nand U1699 (N_1699,N_1656,N_1652);
xnor U1700 (N_1700,N_1635,N_1639);
nor U1701 (N_1701,N_1676,N_1667);
and U1702 (N_1702,N_1628,N_1650);
nor U1703 (N_1703,N_1670,N_1640);
nor U1704 (N_1704,N_1630,N_1629);
nor U1705 (N_1705,N_1675,N_1655);
or U1706 (N_1706,N_1671,N_1678);
or U1707 (N_1707,N_1637,N_1632);
and U1708 (N_1708,N_1647,N_1625);
nand U1709 (N_1709,N_1643,N_1658);
nand U1710 (N_1710,N_1635,N_1641);
or U1711 (N_1711,N_1655,N_1648);
and U1712 (N_1712,N_1628,N_1660);
or U1713 (N_1713,N_1637,N_1661);
nor U1714 (N_1714,N_1622,N_1679);
nand U1715 (N_1715,N_1645,N_1629);
or U1716 (N_1716,N_1624,N_1626);
nor U1717 (N_1717,N_1671,N_1631);
and U1718 (N_1718,N_1626,N_1675);
nand U1719 (N_1719,N_1657,N_1674);
and U1720 (N_1720,N_1675,N_1646);
nand U1721 (N_1721,N_1625,N_1621);
and U1722 (N_1722,N_1660,N_1632);
and U1723 (N_1723,N_1671,N_1662);
or U1724 (N_1724,N_1665,N_1631);
nor U1725 (N_1725,N_1636,N_1645);
nand U1726 (N_1726,N_1640,N_1655);
nor U1727 (N_1727,N_1642,N_1668);
nand U1728 (N_1728,N_1666,N_1672);
and U1729 (N_1729,N_1636,N_1671);
nor U1730 (N_1730,N_1652,N_1621);
nand U1731 (N_1731,N_1637,N_1662);
nand U1732 (N_1732,N_1632,N_1663);
or U1733 (N_1733,N_1621,N_1675);
nand U1734 (N_1734,N_1664,N_1624);
and U1735 (N_1735,N_1668,N_1627);
and U1736 (N_1736,N_1644,N_1638);
nor U1737 (N_1737,N_1665,N_1650);
and U1738 (N_1738,N_1677,N_1629);
nor U1739 (N_1739,N_1645,N_1651);
nand U1740 (N_1740,N_1694,N_1693);
or U1741 (N_1741,N_1720,N_1703);
nand U1742 (N_1742,N_1715,N_1736);
nand U1743 (N_1743,N_1725,N_1733);
nand U1744 (N_1744,N_1681,N_1716);
or U1745 (N_1745,N_1726,N_1739);
nand U1746 (N_1746,N_1713,N_1712);
or U1747 (N_1747,N_1737,N_1682);
or U1748 (N_1748,N_1688,N_1696);
nand U1749 (N_1749,N_1707,N_1731);
nor U1750 (N_1750,N_1689,N_1687);
or U1751 (N_1751,N_1710,N_1708);
xnor U1752 (N_1752,N_1721,N_1711);
nand U1753 (N_1753,N_1686,N_1718);
nor U1754 (N_1754,N_1729,N_1705);
or U1755 (N_1755,N_1697,N_1704);
nand U1756 (N_1756,N_1724,N_1700);
nor U1757 (N_1757,N_1719,N_1727);
and U1758 (N_1758,N_1717,N_1691);
xor U1759 (N_1759,N_1701,N_1702);
nor U1760 (N_1760,N_1730,N_1734);
nor U1761 (N_1761,N_1732,N_1722);
nand U1762 (N_1762,N_1709,N_1680);
or U1763 (N_1763,N_1690,N_1738);
nor U1764 (N_1764,N_1684,N_1685);
or U1765 (N_1765,N_1735,N_1728);
and U1766 (N_1766,N_1698,N_1699);
and U1767 (N_1767,N_1695,N_1714);
nor U1768 (N_1768,N_1692,N_1723);
and U1769 (N_1769,N_1683,N_1706);
xnor U1770 (N_1770,N_1729,N_1715);
nand U1771 (N_1771,N_1699,N_1680);
or U1772 (N_1772,N_1710,N_1735);
or U1773 (N_1773,N_1693,N_1718);
nand U1774 (N_1774,N_1708,N_1689);
nor U1775 (N_1775,N_1738,N_1722);
nor U1776 (N_1776,N_1715,N_1734);
or U1777 (N_1777,N_1717,N_1728);
or U1778 (N_1778,N_1680,N_1691);
or U1779 (N_1779,N_1732,N_1689);
and U1780 (N_1780,N_1683,N_1726);
or U1781 (N_1781,N_1725,N_1704);
and U1782 (N_1782,N_1710,N_1682);
nand U1783 (N_1783,N_1687,N_1680);
xor U1784 (N_1784,N_1702,N_1700);
xnor U1785 (N_1785,N_1680,N_1731);
or U1786 (N_1786,N_1730,N_1701);
and U1787 (N_1787,N_1692,N_1701);
xnor U1788 (N_1788,N_1705,N_1715);
nand U1789 (N_1789,N_1703,N_1716);
nand U1790 (N_1790,N_1720,N_1714);
nor U1791 (N_1791,N_1738,N_1708);
and U1792 (N_1792,N_1723,N_1680);
and U1793 (N_1793,N_1689,N_1717);
and U1794 (N_1794,N_1689,N_1690);
or U1795 (N_1795,N_1720,N_1693);
nor U1796 (N_1796,N_1707,N_1718);
and U1797 (N_1797,N_1693,N_1735);
nor U1798 (N_1798,N_1691,N_1725);
nand U1799 (N_1799,N_1733,N_1704);
nand U1800 (N_1800,N_1790,N_1758);
nor U1801 (N_1801,N_1787,N_1746);
nor U1802 (N_1802,N_1764,N_1777);
and U1803 (N_1803,N_1761,N_1770);
and U1804 (N_1804,N_1765,N_1771);
and U1805 (N_1805,N_1745,N_1748);
nor U1806 (N_1806,N_1742,N_1754);
nand U1807 (N_1807,N_1798,N_1749);
or U1808 (N_1808,N_1795,N_1782);
nor U1809 (N_1809,N_1776,N_1769);
nand U1810 (N_1810,N_1778,N_1775);
and U1811 (N_1811,N_1760,N_1780);
xnor U1812 (N_1812,N_1779,N_1772);
and U1813 (N_1813,N_1763,N_1741);
or U1814 (N_1814,N_1793,N_1796);
nor U1815 (N_1815,N_1768,N_1752);
nand U1816 (N_1816,N_1784,N_1757);
and U1817 (N_1817,N_1786,N_1789);
and U1818 (N_1818,N_1792,N_1744);
or U1819 (N_1819,N_1774,N_1785);
xor U1820 (N_1820,N_1750,N_1781);
nor U1821 (N_1821,N_1767,N_1740);
xor U1822 (N_1822,N_1756,N_1799);
or U1823 (N_1823,N_1783,N_1753);
and U1824 (N_1824,N_1788,N_1773);
xor U1825 (N_1825,N_1755,N_1797);
nor U1826 (N_1826,N_1759,N_1751);
nand U1827 (N_1827,N_1747,N_1762);
and U1828 (N_1828,N_1766,N_1794);
and U1829 (N_1829,N_1743,N_1791);
nand U1830 (N_1830,N_1742,N_1744);
nor U1831 (N_1831,N_1787,N_1789);
xor U1832 (N_1832,N_1792,N_1756);
nor U1833 (N_1833,N_1790,N_1741);
nor U1834 (N_1834,N_1771,N_1748);
xor U1835 (N_1835,N_1778,N_1744);
nor U1836 (N_1836,N_1769,N_1766);
and U1837 (N_1837,N_1795,N_1754);
nand U1838 (N_1838,N_1797,N_1751);
or U1839 (N_1839,N_1766,N_1784);
or U1840 (N_1840,N_1796,N_1773);
nor U1841 (N_1841,N_1762,N_1743);
nand U1842 (N_1842,N_1749,N_1757);
or U1843 (N_1843,N_1740,N_1750);
nor U1844 (N_1844,N_1762,N_1790);
or U1845 (N_1845,N_1754,N_1776);
and U1846 (N_1846,N_1775,N_1797);
nor U1847 (N_1847,N_1767,N_1777);
nor U1848 (N_1848,N_1789,N_1770);
nor U1849 (N_1849,N_1781,N_1798);
nand U1850 (N_1850,N_1755,N_1776);
and U1851 (N_1851,N_1746,N_1791);
nand U1852 (N_1852,N_1789,N_1748);
nand U1853 (N_1853,N_1755,N_1768);
nor U1854 (N_1854,N_1760,N_1755);
or U1855 (N_1855,N_1765,N_1749);
xor U1856 (N_1856,N_1748,N_1786);
nor U1857 (N_1857,N_1749,N_1796);
and U1858 (N_1858,N_1748,N_1755);
nand U1859 (N_1859,N_1742,N_1770);
nand U1860 (N_1860,N_1837,N_1800);
nor U1861 (N_1861,N_1827,N_1836);
or U1862 (N_1862,N_1814,N_1846);
xnor U1863 (N_1863,N_1803,N_1849);
or U1864 (N_1864,N_1824,N_1847);
nand U1865 (N_1865,N_1808,N_1828);
nor U1866 (N_1866,N_1804,N_1819);
nand U1867 (N_1867,N_1810,N_1829);
nand U1868 (N_1868,N_1816,N_1833);
or U1869 (N_1869,N_1859,N_1813);
or U1870 (N_1870,N_1839,N_1806);
xnor U1871 (N_1871,N_1821,N_1805);
nand U1872 (N_1872,N_1854,N_1855);
xor U1873 (N_1873,N_1838,N_1843);
nand U1874 (N_1874,N_1851,N_1802);
nand U1875 (N_1875,N_1809,N_1823);
nand U1876 (N_1876,N_1835,N_1820);
nand U1877 (N_1877,N_1811,N_1801);
and U1878 (N_1878,N_1812,N_1848);
and U1879 (N_1879,N_1844,N_1834);
and U1880 (N_1880,N_1826,N_1807);
xnor U1881 (N_1881,N_1853,N_1818);
or U1882 (N_1882,N_1857,N_1831);
or U1883 (N_1883,N_1817,N_1841);
nor U1884 (N_1884,N_1815,N_1852);
nor U1885 (N_1885,N_1856,N_1842);
nor U1886 (N_1886,N_1822,N_1825);
and U1887 (N_1887,N_1858,N_1840);
or U1888 (N_1888,N_1832,N_1850);
nand U1889 (N_1889,N_1830,N_1845);
xor U1890 (N_1890,N_1800,N_1804);
nand U1891 (N_1891,N_1815,N_1849);
and U1892 (N_1892,N_1811,N_1854);
nand U1893 (N_1893,N_1855,N_1817);
nor U1894 (N_1894,N_1855,N_1816);
and U1895 (N_1895,N_1856,N_1813);
or U1896 (N_1896,N_1825,N_1817);
nor U1897 (N_1897,N_1823,N_1845);
xor U1898 (N_1898,N_1839,N_1858);
or U1899 (N_1899,N_1817,N_1837);
or U1900 (N_1900,N_1830,N_1807);
xor U1901 (N_1901,N_1857,N_1829);
nor U1902 (N_1902,N_1837,N_1816);
and U1903 (N_1903,N_1852,N_1845);
nand U1904 (N_1904,N_1835,N_1828);
xnor U1905 (N_1905,N_1807,N_1818);
and U1906 (N_1906,N_1845,N_1810);
nand U1907 (N_1907,N_1821,N_1825);
nor U1908 (N_1908,N_1817,N_1851);
or U1909 (N_1909,N_1811,N_1802);
and U1910 (N_1910,N_1819,N_1849);
or U1911 (N_1911,N_1823,N_1838);
nand U1912 (N_1912,N_1827,N_1859);
nand U1913 (N_1913,N_1846,N_1847);
nor U1914 (N_1914,N_1821,N_1844);
and U1915 (N_1915,N_1819,N_1857);
nand U1916 (N_1916,N_1839,N_1851);
nand U1917 (N_1917,N_1848,N_1850);
or U1918 (N_1918,N_1839,N_1833);
nor U1919 (N_1919,N_1829,N_1807);
nand U1920 (N_1920,N_1890,N_1887);
or U1921 (N_1921,N_1905,N_1892);
xnor U1922 (N_1922,N_1878,N_1912);
and U1923 (N_1923,N_1863,N_1910);
and U1924 (N_1924,N_1862,N_1893);
nand U1925 (N_1925,N_1885,N_1867);
nand U1926 (N_1926,N_1876,N_1868);
or U1927 (N_1927,N_1874,N_1879);
nor U1928 (N_1928,N_1914,N_1888);
nor U1929 (N_1929,N_1903,N_1891);
nand U1930 (N_1930,N_1907,N_1869);
or U1931 (N_1931,N_1864,N_1906);
and U1932 (N_1932,N_1880,N_1909);
nand U1933 (N_1933,N_1919,N_1889);
or U1934 (N_1934,N_1896,N_1902);
and U1935 (N_1935,N_1908,N_1882);
nand U1936 (N_1936,N_1877,N_1861);
or U1937 (N_1937,N_1870,N_1898);
and U1938 (N_1938,N_1897,N_1884);
nand U1939 (N_1939,N_1916,N_1895);
xor U1940 (N_1940,N_1865,N_1901);
and U1941 (N_1941,N_1873,N_1883);
nand U1942 (N_1942,N_1866,N_1904);
nand U1943 (N_1943,N_1899,N_1915);
xor U1944 (N_1944,N_1894,N_1871);
nand U1945 (N_1945,N_1872,N_1900);
nand U1946 (N_1946,N_1860,N_1886);
xnor U1947 (N_1947,N_1911,N_1875);
nand U1948 (N_1948,N_1918,N_1917);
and U1949 (N_1949,N_1913,N_1881);
nand U1950 (N_1950,N_1906,N_1905);
or U1951 (N_1951,N_1904,N_1896);
nor U1952 (N_1952,N_1887,N_1903);
xor U1953 (N_1953,N_1883,N_1894);
or U1954 (N_1954,N_1918,N_1899);
nor U1955 (N_1955,N_1884,N_1909);
nor U1956 (N_1956,N_1878,N_1862);
or U1957 (N_1957,N_1900,N_1918);
or U1958 (N_1958,N_1919,N_1891);
or U1959 (N_1959,N_1882,N_1869);
and U1960 (N_1960,N_1917,N_1892);
nor U1961 (N_1961,N_1892,N_1873);
nor U1962 (N_1962,N_1866,N_1891);
nand U1963 (N_1963,N_1879,N_1863);
or U1964 (N_1964,N_1897,N_1860);
nor U1965 (N_1965,N_1883,N_1876);
and U1966 (N_1966,N_1879,N_1916);
nand U1967 (N_1967,N_1887,N_1893);
xor U1968 (N_1968,N_1883,N_1871);
nand U1969 (N_1969,N_1878,N_1917);
and U1970 (N_1970,N_1862,N_1918);
nand U1971 (N_1971,N_1915,N_1901);
and U1972 (N_1972,N_1902,N_1863);
nor U1973 (N_1973,N_1885,N_1908);
or U1974 (N_1974,N_1907,N_1894);
nor U1975 (N_1975,N_1918,N_1913);
nor U1976 (N_1976,N_1884,N_1916);
nor U1977 (N_1977,N_1861,N_1874);
nand U1978 (N_1978,N_1895,N_1881);
xnor U1979 (N_1979,N_1908,N_1862);
nor U1980 (N_1980,N_1930,N_1956);
and U1981 (N_1981,N_1939,N_1937);
xor U1982 (N_1982,N_1969,N_1973);
or U1983 (N_1983,N_1946,N_1943);
nand U1984 (N_1984,N_1931,N_1934);
and U1985 (N_1985,N_1944,N_1971);
nor U1986 (N_1986,N_1923,N_1965);
nor U1987 (N_1987,N_1932,N_1960);
nand U1988 (N_1988,N_1955,N_1967);
xor U1989 (N_1989,N_1940,N_1975);
xor U1990 (N_1990,N_1963,N_1959);
or U1991 (N_1991,N_1929,N_1972);
or U1992 (N_1992,N_1962,N_1950);
nand U1993 (N_1993,N_1925,N_1938);
nor U1994 (N_1994,N_1948,N_1979);
xor U1995 (N_1995,N_1966,N_1926);
xnor U1996 (N_1996,N_1953,N_1954);
and U1997 (N_1997,N_1957,N_1964);
and U1998 (N_1998,N_1935,N_1968);
or U1999 (N_1999,N_1945,N_1928);
nand U2000 (N_2000,N_1936,N_1922);
nor U2001 (N_2001,N_1924,N_1977);
nand U2002 (N_2002,N_1941,N_1927);
xnor U2003 (N_2003,N_1921,N_1920);
nor U2004 (N_2004,N_1942,N_1951);
xor U2005 (N_2005,N_1952,N_1933);
or U2006 (N_2006,N_1974,N_1958);
or U2007 (N_2007,N_1978,N_1970);
or U2008 (N_2008,N_1976,N_1947);
or U2009 (N_2009,N_1961,N_1949);
xor U2010 (N_2010,N_1935,N_1962);
nand U2011 (N_2011,N_1959,N_1973);
xnor U2012 (N_2012,N_1963,N_1977);
xnor U2013 (N_2013,N_1952,N_1922);
xnor U2014 (N_2014,N_1937,N_1958);
xnor U2015 (N_2015,N_1969,N_1929);
nor U2016 (N_2016,N_1962,N_1976);
nand U2017 (N_2017,N_1947,N_1937);
nand U2018 (N_2018,N_1957,N_1969);
nand U2019 (N_2019,N_1953,N_1932);
and U2020 (N_2020,N_1951,N_1963);
and U2021 (N_2021,N_1966,N_1945);
and U2022 (N_2022,N_1979,N_1960);
nand U2023 (N_2023,N_1933,N_1963);
or U2024 (N_2024,N_1938,N_1921);
or U2025 (N_2025,N_1965,N_1962);
xnor U2026 (N_2026,N_1978,N_1940);
and U2027 (N_2027,N_1957,N_1947);
or U2028 (N_2028,N_1940,N_1970);
xor U2029 (N_2029,N_1938,N_1932);
nor U2030 (N_2030,N_1950,N_1939);
nand U2031 (N_2031,N_1951,N_1949);
nor U2032 (N_2032,N_1955,N_1941);
and U2033 (N_2033,N_1948,N_1958);
nor U2034 (N_2034,N_1933,N_1961);
or U2035 (N_2035,N_1961,N_1930);
nor U2036 (N_2036,N_1920,N_1949);
or U2037 (N_2037,N_1932,N_1930);
or U2038 (N_2038,N_1958,N_1922);
and U2039 (N_2039,N_1963,N_1936);
nand U2040 (N_2040,N_2003,N_2026);
xnor U2041 (N_2041,N_1990,N_2016);
and U2042 (N_2042,N_2032,N_1987);
and U2043 (N_2043,N_1997,N_1994);
and U2044 (N_2044,N_2018,N_1984);
and U2045 (N_2045,N_2021,N_2025);
nand U2046 (N_2046,N_2015,N_2035);
nand U2047 (N_2047,N_1980,N_2033);
nor U2048 (N_2048,N_2004,N_2039);
and U2049 (N_2049,N_1983,N_2000);
and U2050 (N_2050,N_1991,N_1989);
xnor U2051 (N_2051,N_2014,N_2031);
or U2052 (N_2052,N_1992,N_2023);
nand U2053 (N_2053,N_2006,N_2027);
or U2054 (N_2054,N_2037,N_2024);
or U2055 (N_2055,N_1985,N_1996);
and U2056 (N_2056,N_2002,N_2022);
or U2057 (N_2057,N_2011,N_1993);
and U2058 (N_2058,N_1982,N_2012);
nor U2059 (N_2059,N_2019,N_1981);
and U2060 (N_2060,N_1998,N_1995);
nor U2061 (N_2061,N_2036,N_2020);
and U2062 (N_2062,N_2030,N_2001);
nand U2063 (N_2063,N_2038,N_1986);
nand U2064 (N_2064,N_2009,N_2034);
or U2065 (N_2065,N_2017,N_1999);
nor U2066 (N_2066,N_1988,N_2010);
and U2067 (N_2067,N_2028,N_2007);
nor U2068 (N_2068,N_2029,N_2008);
or U2069 (N_2069,N_2013,N_2005);
nand U2070 (N_2070,N_1987,N_2035);
nand U2071 (N_2071,N_1990,N_1995);
nand U2072 (N_2072,N_2014,N_2020);
and U2073 (N_2073,N_2025,N_2020);
nand U2074 (N_2074,N_1990,N_2026);
nand U2075 (N_2075,N_2000,N_1998);
nand U2076 (N_2076,N_2024,N_1997);
xor U2077 (N_2077,N_1981,N_2039);
nor U2078 (N_2078,N_2001,N_2033);
xor U2079 (N_2079,N_2015,N_2030);
nor U2080 (N_2080,N_1994,N_1980);
and U2081 (N_2081,N_2023,N_2006);
nand U2082 (N_2082,N_2000,N_2008);
nand U2083 (N_2083,N_1985,N_2005);
xor U2084 (N_2084,N_2006,N_1995);
xnor U2085 (N_2085,N_2034,N_2012);
and U2086 (N_2086,N_2006,N_2009);
nor U2087 (N_2087,N_2023,N_2010);
nand U2088 (N_2088,N_2031,N_1984);
nand U2089 (N_2089,N_1990,N_2036);
and U2090 (N_2090,N_2004,N_2036);
nand U2091 (N_2091,N_2000,N_2033);
nand U2092 (N_2092,N_1983,N_2022);
and U2093 (N_2093,N_2031,N_2038);
nand U2094 (N_2094,N_2022,N_2020);
nor U2095 (N_2095,N_2000,N_2005);
nor U2096 (N_2096,N_2027,N_2039);
and U2097 (N_2097,N_1999,N_2037);
nand U2098 (N_2098,N_1995,N_2005);
nor U2099 (N_2099,N_2028,N_2013);
xnor U2100 (N_2100,N_2071,N_2088);
or U2101 (N_2101,N_2048,N_2051);
or U2102 (N_2102,N_2064,N_2077);
and U2103 (N_2103,N_2043,N_2082);
and U2104 (N_2104,N_2044,N_2079);
and U2105 (N_2105,N_2075,N_2089);
and U2106 (N_2106,N_2068,N_2084);
xor U2107 (N_2107,N_2041,N_2085);
and U2108 (N_2108,N_2078,N_2093);
and U2109 (N_2109,N_2097,N_2061);
nand U2110 (N_2110,N_2049,N_2076);
or U2111 (N_2111,N_2094,N_2060);
or U2112 (N_2112,N_2056,N_2091);
nor U2113 (N_2113,N_2081,N_2086);
nand U2114 (N_2114,N_2059,N_2058);
xnor U2115 (N_2115,N_2057,N_2072);
or U2116 (N_2116,N_2090,N_2047);
and U2117 (N_2117,N_2080,N_2070);
or U2118 (N_2118,N_2065,N_2096);
or U2119 (N_2119,N_2050,N_2095);
nand U2120 (N_2120,N_2099,N_2054);
and U2121 (N_2121,N_2067,N_2046);
nor U2122 (N_2122,N_2052,N_2074);
nand U2123 (N_2123,N_2053,N_2062);
and U2124 (N_2124,N_2040,N_2098);
or U2125 (N_2125,N_2092,N_2087);
or U2126 (N_2126,N_2073,N_2042);
or U2127 (N_2127,N_2066,N_2083);
xor U2128 (N_2128,N_2055,N_2069);
nand U2129 (N_2129,N_2045,N_2063);
nor U2130 (N_2130,N_2076,N_2075);
and U2131 (N_2131,N_2043,N_2058);
nand U2132 (N_2132,N_2084,N_2059);
nand U2133 (N_2133,N_2081,N_2042);
nand U2134 (N_2134,N_2090,N_2071);
xnor U2135 (N_2135,N_2045,N_2071);
and U2136 (N_2136,N_2079,N_2062);
and U2137 (N_2137,N_2045,N_2091);
or U2138 (N_2138,N_2072,N_2086);
nand U2139 (N_2139,N_2055,N_2091);
nand U2140 (N_2140,N_2091,N_2064);
or U2141 (N_2141,N_2060,N_2093);
nand U2142 (N_2142,N_2096,N_2055);
nor U2143 (N_2143,N_2086,N_2056);
nand U2144 (N_2144,N_2066,N_2094);
or U2145 (N_2145,N_2041,N_2099);
xor U2146 (N_2146,N_2061,N_2068);
and U2147 (N_2147,N_2040,N_2085);
and U2148 (N_2148,N_2058,N_2099);
or U2149 (N_2149,N_2063,N_2087);
and U2150 (N_2150,N_2042,N_2090);
and U2151 (N_2151,N_2064,N_2072);
or U2152 (N_2152,N_2077,N_2095);
or U2153 (N_2153,N_2086,N_2068);
or U2154 (N_2154,N_2077,N_2056);
and U2155 (N_2155,N_2076,N_2059);
nand U2156 (N_2156,N_2069,N_2053);
and U2157 (N_2157,N_2063,N_2054);
nor U2158 (N_2158,N_2077,N_2076);
nor U2159 (N_2159,N_2048,N_2081);
or U2160 (N_2160,N_2123,N_2138);
nor U2161 (N_2161,N_2151,N_2132);
nor U2162 (N_2162,N_2150,N_2122);
or U2163 (N_2163,N_2120,N_2107);
and U2164 (N_2164,N_2140,N_2121);
or U2165 (N_2165,N_2152,N_2125);
nand U2166 (N_2166,N_2112,N_2144);
nand U2167 (N_2167,N_2127,N_2139);
xor U2168 (N_2168,N_2100,N_2117);
nand U2169 (N_2169,N_2126,N_2156);
nand U2170 (N_2170,N_2124,N_2111);
and U2171 (N_2171,N_2119,N_2159);
nand U2172 (N_2172,N_2135,N_2110);
and U2173 (N_2173,N_2157,N_2115);
nor U2174 (N_2174,N_2103,N_2149);
nor U2175 (N_2175,N_2116,N_2104);
nand U2176 (N_2176,N_2114,N_2146);
nor U2177 (N_2177,N_2109,N_2113);
and U2178 (N_2178,N_2108,N_2137);
or U2179 (N_2179,N_2147,N_2106);
nor U2180 (N_2180,N_2105,N_2142);
or U2181 (N_2181,N_2118,N_2148);
nor U2182 (N_2182,N_2155,N_2128);
and U2183 (N_2183,N_2136,N_2145);
or U2184 (N_2184,N_2143,N_2141);
nor U2185 (N_2185,N_2129,N_2154);
and U2186 (N_2186,N_2133,N_2131);
nand U2187 (N_2187,N_2101,N_2130);
nand U2188 (N_2188,N_2153,N_2102);
and U2189 (N_2189,N_2158,N_2134);
and U2190 (N_2190,N_2138,N_2111);
or U2191 (N_2191,N_2155,N_2135);
xnor U2192 (N_2192,N_2131,N_2144);
or U2193 (N_2193,N_2129,N_2119);
nor U2194 (N_2194,N_2127,N_2136);
nor U2195 (N_2195,N_2154,N_2150);
or U2196 (N_2196,N_2105,N_2132);
and U2197 (N_2197,N_2108,N_2106);
nor U2198 (N_2198,N_2149,N_2152);
nand U2199 (N_2199,N_2130,N_2149);
nand U2200 (N_2200,N_2152,N_2137);
and U2201 (N_2201,N_2158,N_2103);
and U2202 (N_2202,N_2125,N_2133);
nor U2203 (N_2203,N_2159,N_2133);
nor U2204 (N_2204,N_2122,N_2132);
and U2205 (N_2205,N_2145,N_2124);
nand U2206 (N_2206,N_2136,N_2157);
xnor U2207 (N_2207,N_2109,N_2121);
nor U2208 (N_2208,N_2142,N_2138);
nand U2209 (N_2209,N_2105,N_2146);
or U2210 (N_2210,N_2134,N_2157);
and U2211 (N_2211,N_2158,N_2121);
and U2212 (N_2212,N_2114,N_2148);
and U2213 (N_2213,N_2147,N_2155);
nor U2214 (N_2214,N_2109,N_2115);
xor U2215 (N_2215,N_2114,N_2106);
and U2216 (N_2216,N_2105,N_2125);
or U2217 (N_2217,N_2146,N_2139);
and U2218 (N_2218,N_2148,N_2126);
nand U2219 (N_2219,N_2155,N_2150);
and U2220 (N_2220,N_2170,N_2163);
and U2221 (N_2221,N_2165,N_2161);
xnor U2222 (N_2222,N_2187,N_2166);
or U2223 (N_2223,N_2198,N_2202);
or U2224 (N_2224,N_2218,N_2191);
and U2225 (N_2225,N_2211,N_2196);
nand U2226 (N_2226,N_2197,N_2216);
or U2227 (N_2227,N_2164,N_2175);
or U2228 (N_2228,N_2212,N_2190);
and U2229 (N_2229,N_2219,N_2173);
nand U2230 (N_2230,N_2199,N_2179);
or U2231 (N_2231,N_2180,N_2186);
and U2232 (N_2232,N_2169,N_2160);
or U2233 (N_2233,N_2185,N_2205);
or U2234 (N_2234,N_2181,N_2207);
and U2235 (N_2235,N_2168,N_2209);
nand U2236 (N_2236,N_2178,N_2189);
nor U2237 (N_2237,N_2208,N_2217);
or U2238 (N_2238,N_2184,N_2200);
nand U2239 (N_2239,N_2177,N_2188);
nand U2240 (N_2240,N_2214,N_2176);
and U2241 (N_2241,N_2210,N_2171);
and U2242 (N_2242,N_2195,N_2162);
and U2243 (N_2243,N_2183,N_2203);
nand U2244 (N_2244,N_2194,N_2193);
or U2245 (N_2245,N_2182,N_2213);
nand U2246 (N_2246,N_2167,N_2172);
and U2247 (N_2247,N_2204,N_2206);
nand U2248 (N_2248,N_2174,N_2201);
nand U2249 (N_2249,N_2215,N_2192);
or U2250 (N_2250,N_2210,N_2164);
nor U2251 (N_2251,N_2173,N_2164);
nor U2252 (N_2252,N_2205,N_2190);
nand U2253 (N_2253,N_2205,N_2198);
or U2254 (N_2254,N_2218,N_2195);
nand U2255 (N_2255,N_2189,N_2191);
and U2256 (N_2256,N_2197,N_2180);
nor U2257 (N_2257,N_2209,N_2164);
xnor U2258 (N_2258,N_2187,N_2203);
nand U2259 (N_2259,N_2177,N_2219);
nor U2260 (N_2260,N_2164,N_2185);
or U2261 (N_2261,N_2185,N_2214);
or U2262 (N_2262,N_2205,N_2202);
nor U2263 (N_2263,N_2180,N_2177);
nand U2264 (N_2264,N_2184,N_2217);
nand U2265 (N_2265,N_2193,N_2208);
nand U2266 (N_2266,N_2205,N_2171);
and U2267 (N_2267,N_2165,N_2164);
nor U2268 (N_2268,N_2200,N_2177);
xor U2269 (N_2269,N_2177,N_2216);
nor U2270 (N_2270,N_2211,N_2182);
nor U2271 (N_2271,N_2161,N_2188);
nand U2272 (N_2272,N_2208,N_2173);
or U2273 (N_2273,N_2180,N_2187);
or U2274 (N_2274,N_2191,N_2186);
and U2275 (N_2275,N_2171,N_2162);
and U2276 (N_2276,N_2160,N_2207);
nand U2277 (N_2277,N_2202,N_2165);
nand U2278 (N_2278,N_2187,N_2168);
nand U2279 (N_2279,N_2173,N_2205);
and U2280 (N_2280,N_2232,N_2260);
and U2281 (N_2281,N_2235,N_2241);
nand U2282 (N_2282,N_2258,N_2261);
and U2283 (N_2283,N_2275,N_2267);
nor U2284 (N_2284,N_2254,N_2247);
or U2285 (N_2285,N_2262,N_2251);
xnor U2286 (N_2286,N_2278,N_2277);
nor U2287 (N_2287,N_2243,N_2255);
nor U2288 (N_2288,N_2242,N_2264);
and U2289 (N_2289,N_2245,N_2225);
or U2290 (N_2290,N_2220,N_2253);
and U2291 (N_2291,N_2263,N_2231);
nor U2292 (N_2292,N_2250,N_2273);
nor U2293 (N_2293,N_2265,N_2256);
and U2294 (N_2294,N_2276,N_2223);
and U2295 (N_2295,N_2272,N_2268);
and U2296 (N_2296,N_2246,N_2271);
nor U2297 (N_2297,N_2240,N_2238);
or U2298 (N_2298,N_2269,N_2233);
and U2299 (N_2299,N_2226,N_2229);
xor U2300 (N_2300,N_2221,N_2252);
xnor U2301 (N_2301,N_2237,N_2274);
xor U2302 (N_2302,N_2228,N_2236);
nand U2303 (N_2303,N_2222,N_2230);
and U2304 (N_2304,N_2266,N_2244);
xor U2305 (N_2305,N_2249,N_2234);
nor U2306 (N_2306,N_2259,N_2279);
nor U2307 (N_2307,N_2270,N_2248);
or U2308 (N_2308,N_2257,N_2224);
nor U2309 (N_2309,N_2239,N_2227);
and U2310 (N_2310,N_2257,N_2228);
or U2311 (N_2311,N_2259,N_2264);
nand U2312 (N_2312,N_2223,N_2222);
nor U2313 (N_2313,N_2241,N_2224);
nand U2314 (N_2314,N_2258,N_2222);
nand U2315 (N_2315,N_2235,N_2262);
and U2316 (N_2316,N_2271,N_2241);
nor U2317 (N_2317,N_2261,N_2241);
or U2318 (N_2318,N_2239,N_2271);
xnor U2319 (N_2319,N_2226,N_2266);
and U2320 (N_2320,N_2227,N_2231);
or U2321 (N_2321,N_2278,N_2262);
and U2322 (N_2322,N_2259,N_2273);
nand U2323 (N_2323,N_2259,N_2246);
nand U2324 (N_2324,N_2243,N_2228);
and U2325 (N_2325,N_2255,N_2256);
or U2326 (N_2326,N_2267,N_2259);
nand U2327 (N_2327,N_2248,N_2227);
nand U2328 (N_2328,N_2255,N_2223);
nand U2329 (N_2329,N_2232,N_2239);
nand U2330 (N_2330,N_2241,N_2240);
nand U2331 (N_2331,N_2267,N_2269);
or U2332 (N_2332,N_2260,N_2222);
or U2333 (N_2333,N_2270,N_2228);
nand U2334 (N_2334,N_2237,N_2270);
nor U2335 (N_2335,N_2254,N_2274);
nor U2336 (N_2336,N_2225,N_2229);
nand U2337 (N_2337,N_2237,N_2255);
and U2338 (N_2338,N_2261,N_2263);
or U2339 (N_2339,N_2254,N_2245);
nand U2340 (N_2340,N_2291,N_2290);
nor U2341 (N_2341,N_2330,N_2310);
nor U2342 (N_2342,N_2309,N_2337);
nand U2343 (N_2343,N_2298,N_2320);
nor U2344 (N_2344,N_2305,N_2302);
nand U2345 (N_2345,N_2293,N_2303);
nand U2346 (N_2346,N_2294,N_2283);
or U2347 (N_2347,N_2327,N_2334);
or U2348 (N_2348,N_2286,N_2331);
and U2349 (N_2349,N_2299,N_2329);
and U2350 (N_2350,N_2335,N_2317);
and U2351 (N_2351,N_2297,N_2314);
nor U2352 (N_2352,N_2339,N_2326);
xnor U2353 (N_2353,N_2312,N_2292);
or U2354 (N_2354,N_2336,N_2281);
xnor U2355 (N_2355,N_2322,N_2319);
or U2356 (N_2356,N_2301,N_2285);
and U2357 (N_2357,N_2289,N_2311);
xnor U2358 (N_2358,N_2333,N_2313);
nor U2359 (N_2359,N_2295,N_2332);
xnor U2360 (N_2360,N_2284,N_2296);
and U2361 (N_2361,N_2282,N_2338);
nor U2362 (N_2362,N_2280,N_2315);
nor U2363 (N_2363,N_2307,N_2300);
and U2364 (N_2364,N_2321,N_2318);
or U2365 (N_2365,N_2308,N_2328);
nand U2366 (N_2366,N_2316,N_2324);
nand U2367 (N_2367,N_2288,N_2304);
nor U2368 (N_2368,N_2287,N_2306);
or U2369 (N_2369,N_2325,N_2323);
xnor U2370 (N_2370,N_2313,N_2332);
nand U2371 (N_2371,N_2324,N_2320);
or U2372 (N_2372,N_2319,N_2330);
nor U2373 (N_2373,N_2281,N_2299);
and U2374 (N_2374,N_2297,N_2333);
nor U2375 (N_2375,N_2323,N_2328);
and U2376 (N_2376,N_2331,N_2318);
nor U2377 (N_2377,N_2319,N_2312);
nand U2378 (N_2378,N_2317,N_2303);
and U2379 (N_2379,N_2288,N_2311);
nand U2380 (N_2380,N_2300,N_2289);
nor U2381 (N_2381,N_2296,N_2316);
and U2382 (N_2382,N_2286,N_2334);
and U2383 (N_2383,N_2334,N_2317);
nand U2384 (N_2384,N_2306,N_2326);
and U2385 (N_2385,N_2334,N_2280);
nor U2386 (N_2386,N_2313,N_2325);
nand U2387 (N_2387,N_2334,N_2318);
and U2388 (N_2388,N_2334,N_2311);
nand U2389 (N_2389,N_2314,N_2308);
and U2390 (N_2390,N_2290,N_2296);
nor U2391 (N_2391,N_2328,N_2332);
or U2392 (N_2392,N_2331,N_2313);
or U2393 (N_2393,N_2290,N_2324);
and U2394 (N_2394,N_2334,N_2332);
nor U2395 (N_2395,N_2326,N_2296);
nand U2396 (N_2396,N_2327,N_2300);
or U2397 (N_2397,N_2306,N_2286);
nand U2398 (N_2398,N_2338,N_2323);
and U2399 (N_2399,N_2304,N_2305);
nand U2400 (N_2400,N_2393,N_2342);
nor U2401 (N_2401,N_2367,N_2354);
nand U2402 (N_2402,N_2340,N_2384);
nand U2403 (N_2403,N_2345,N_2379);
nand U2404 (N_2404,N_2351,N_2383);
and U2405 (N_2405,N_2362,N_2378);
nand U2406 (N_2406,N_2364,N_2398);
or U2407 (N_2407,N_2370,N_2353);
or U2408 (N_2408,N_2391,N_2394);
or U2409 (N_2409,N_2352,N_2372);
and U2410 (N_2410,N_2366,N_2390);
and U2411 (N_2411,N_2344,N_2361);
and U2412 (N_2412,N_2382,N_2399);
nor U2413 (N_2413,N_2358,N_2395);
nor U2414 (N_2414,N_2348,N_2392);
nand U2415 (N_2415,N_2369,N_2377);
and U2416 (N_2416,N_2375,N_2371);
nor U2417 (N_2417,N_2381,N_2386);
or U2418 (N_2418,N_2368,N_2385);
or U2419 (N_2419,N_2396,N_2397);
or U2420 (N_2420,N_2376,N_2356);
or U2421 (N_2421,N_2359,N_2341);
and U2422 (N_2422,N_2373,N_2355);
nand U2423 (N_2423,N_2346,N_2389);
and U2424 (N_2424,N_2387,N_2380);
or U2425 (N_2425,N_2349,N_2374);
xor U2426 (N_2426,N_2347,N_2365);
nand U2427 (N_2427,N_2350,N_2388);
nand U2428 (N_2428,N_2363,N_2360);
and U2429 (N_2429,N_2357,N_2343);
or U2430 (N_2430,N_2368,N_2361);
or U2431 (N_2431,N_2348,N_2342);
nor U2432 (N_2432,N_2393,N_2367);
or U2433 (N_2433,N_2379,N_2390);
and U2434 (N_2434,N_2356,N_2367);
nor U2435 (N_2435,N_2353,N_2391);
or U2436 (N_2436,N_2399,N_2367);
xnor U2437 (N_2437,N_2398,N_2341);
nand U2438 (N_2438,N_2392,N_2341);
nand U2439 (N_2439,N_2384,N_2342);
nor U2440 (N_2440,N_2363,N_2366);
and U2441 (N_2441,N_2355,N_2347);
and U2442 (N_2442,N_2399,N_2351);
and U2443 (N_2443,N_2376,N_2385);
nor U2444 (N_2444,N_2362,N_2341);
or U2445 (N_2445,N_2343,N_2350);
and U2446 (N_2446,N_2361,N_2370);
nand U2447 (N_2447,N_2361,N_2391);
nor U2448 (N_2448,N_2388,N_2395);
nor U2449 (N_2449,N_2367,N_2359);
and U2450 (N_2450,N_2376,N_2366);
and U2451 (N_2451,N_2386,N_2354);
or U2452 (N_2452,N_2366,N_2383);
or U2453 (N_2453,N_2379,N_2395);
nor U2454 (N_2454,N_2349,N_2375);
and U2455 (N_2455,N_2349,N_2358);
nor U2456 (N_2456,N_2341,N_2378);
or U2457 (N_2457,N_2379,N_2393);
nor U2458 (N_2458,N_2383,N_2347);
nor U2459 (N_2459,N_2380,N_2368);
and U2460 (N_2460,N_2445,N_2446);
nand U2461 (N_2461,N_2404,N_2405);
xor U2462 (N_2462,N_2436,N_2418);
nand U2463 (N_2463,N_2434,N_2428);
and U2464 (N_2464,N_2424,N_2437);
nand U2465 (N_2465,N_2401,N_2421);
xnor U2466 (N_2466,N_2451,N_2453);
xor U2467 (N_2467,N_2407,N_2430);
nor U2468 (N_2468,N_2416,N_2402);
and U2469 (N_2469,N_2456,N_2406);
xor U2470 (N_2470,N_2400,N_2454);
and U2471 (N_2471,N_2414,N_2423);
and U2472 (N_2472,N_2420,N_2408);
and U2473 (N_2473,N_2455,N_2452);
or U2474 (N_2474,N_2425,N_2459);
nand U2475 (N_2475,N_2440,N_2449);
and U2476 (N_2476,N_2411,N_2429);
and U2477 (N_2477,N_2403,N_2442);
xnor U2478 (N_2478,N_2447,N_2410);
nand U2479 (N_2479,N_2412,N_2415);
and U2480 (N_2480,N_2431,N_2439);
and U2481 (N_2481,N_2432,N_2444);
nand U2482 (N_2482,N_2450,N_2457);
nor U2483 (N_2483,N_2422,N_2433);
nand U2484 (N_2484,N_2426,N_2419);
xor U2485 (N_2485,N_2438,N_2435);
and U2486 (N_2486,N_2417,N_2441);
and U2487 (N_2487,N_2427,N_2409);
or U2488 (N_2488,N_2413,N_2458);
nor U2489 (N_2489,N_2443,N_2448);
xor U2490 (N_2490,N_2437,N_2421);
nor U2491 (N_2491,N_2424,N_2451);
nand U2492 (N_2492,N_2447,N_2427);
and U2493 (N_2493,N_2401,N_2416);
xnor U2494 (N_2494,N_2414,N_2443);
nor U2495 (N_2495,N_2438,N_2422);
or U2496 (N_2496,N_2442,N_2448);
and U2497 (N_2497,N_2401,N_2403);
and U2498 (N_2498,N_2422,N_2435);
xnor U2499 (N_2499,N_2452,N_2447);
or U2500 (N_2500,N_2442,N_2438);
or U2501 (N_2501,N_2413,N_2451);
nand U2502 (N_2502,N_2445,N_2428);
nand U2503 (N_2503,N_2440,N_2410);
nor U2504 (N_2504,N_2441,N_2452);
or U2505 (N_2505,N_2436,N_2443);
nand U2506 (N_2506,N_2439,N_2412);
or U2507 (N_2507,N_2430,N_2403);
or U2508 (N_2508,N_2441,N_2437);
nor U2509 (N_2509,N_2414,N_2429);
and U2510 (N_2510,N_2429,N_2406);
nand U2511 (N_2511,N_2436,N_2400);
nor U2512 (N_2512,N_2424,N_2445);
or U2513 (N_2513,N_2408,N_2404);
nor U2514 (N_2514,N_2404,N_2406);
and U2515 (N_2515,N_2456,N_2432);
and U2516 (N_2516,N_2447,N_2411);
nand U2517 (N_2517,N_2435,N_2425);
nand U2518 (N_2518,N_2449,N_2448);
nor U2519 (N_2519,N_2439,N_2401);
nor U2520 (N_2520,N_2481,N_2480);
or U2521 (N_2521,N_2517,N_2485);
nand U2522 (N_2522,N_2515,N_2497);
nor U2523 (N_2523,N_2474,N_2500);
nor U2524 (N_2524,N_2513,N_2504);
xor U2525 (N_2525,N_2508,N_2503);
or U2526 (N_2526,N_2471,N_2483);
or U2527 (N_2527,N_2490,N_2494);
and U2528 (N_2528,N_2478,N_2479);
and U2529 (N_2529,N_2491,N_2477);
nand U2530 (N_2530,N_2467,N_2470);
or U2531 (N_2531,N_2489,N_2492);
or U2532 (N_2532,N_2502,N_2518);
nor U2533 (N_2533,N_2505,N_2506);
or U2534 (N_2534,N_2493,N_2501);
nand U2535 (N_2535,N_2499,N_2496);
nand U2536 (N_2536,N_2488,N_2509);
or U2537 (N_2537,N_2462,N_2487);
nor U2538 (N_2538,N_2461,N_2468);
and U2539 (N_2539,N_2473,N_2463);
and U2540 (N_2540,N_2511,N_2514);
nand U2541 (N_2541,N_2486,N_2460);
xnor U2542 (N_2542,N_2472,N_2495);
and U2543 (N_2543,N_2484,N_2519);
and U2544 (N_2544,N_2516,N_2498);
nand U2545 (N_2545,N_2469,N_2476);
and U2546 (N_2546,N_2475,N_2466);
nor U2547 (N_2547,N_2512,N_2507);
or U2548 (N_2548,N_2465,N_2510);
nand U2549 (N_2549,N_2482,N_2464);
nand U2550 (N_2550,N_2512,N_2468);
nand U2551 (N_2551,N_2472,N_2468);
xor U2552 (N_2552,N_2491,N_2474);
nor U2553 (N_2553,N_2467,N_2482);
or U2554 (N_2554,N_2509,N_2507);
xnor U2555 (N_2555,N_2482,N_2466);
and U2556 (N_2556,N_2469,N_2511);
or U2557 (N_2557,N_2481,N_2500);
nand U2558 (N_2558,N_2480,N_2515);
or U2559 (N_2559,N_2498,N_2481);
and U2560 (N_2560,N_2512,N_2493);
and U2561 (N_2561,N_2460,N_2495);
xor U2562 (N_2562,N_2495,N_2475);
nor U2563 (N_2563,N_2500,N_2479);
and U2564 (N_2564,N_2464,N_2513);
or U2565 (N_2565,N_2515,N_2478);
or U2566 (N_2566,N_2483,N_2496);
nor U2567 (N_2567,N_2485,N_2460);
nor U2568 (N_2568,N_2518,N_2473);
nand U2569 (N_2569,N_2518,N_2485);
nand U2570 (N_2570,N_2518,N_2470);
xnor U2571 (N_2571,N_2481,N_2482);
and U2572 (N_2572,N_2484,N_2474);
or U2573 (N_2573,N_2516,N_2506);
nor U2574 (N_2574,N_2478,N_2486);
xnor U2575 (N_2575,N_2486,N_2505);
nor U2576 (N_2576,N_2467,N_2492);
or U2577 (N_2577,N_2486,N_2482);
and U2578 (N_2578,N_2476,N_2490);
xnor U2579 (N_2579,N_2514,N_2461);
nand U2580 (N_2580,N_2564,N_2556);
and U2581 (N_2581,N_2546,N_2537);
and U2582 (N_2582,N_2545,N_2538);
nor U2583 (N_2583,N_2548,N_2573);
nor U2584 (N_2584,N_2572,N_2523);
nand U2585 (N_2585,N_2560,N_2547);
xnor U2586 (N_2586,N_2525,N_2531);
or U2587 (N_2587,N_2575,N_2561);
nor U2588 (N_2588,N_2577,N_2578);
nor U2589 (N_2589,N_2535,N_2549);
nor U2590 (N_2590,N_2576,N_2521);
xor U2591 (N_2591,N_2567,N_2532);
xnor U2592 (N_2592,N_2524,N_2554);
and U2593 (N_2593,N_2536,N_2555);
nor U2594 (N_2594,N_2544,N_2522);
or U2595 (N_2595,N_2541,N_2569);
nand U2596 (N_2596,N_2566,N_2533);
or U2597 (N_2597,N_2570,N_2565);
or U2598 (N_2598,N_2558,N_2529);
nor U2599 (N_2599,N_2540,N_2571);
nand U2600 (N_2600,N_2527,N_2568);
xnor U2601 (N_2601,N_2552,N_2550);
and U2602 (N_2602,N_2562,N_2520);
nor U2603 (N_2603,N_2579,N_2551);
nand U2604 (N_2604,N_2542,N_2534);
and U2605 (N_2605,N_2530,N_2574);
nand U2606 (N_2606,N_2563,N_2543);
nor U2607 (N_2607,N_2539,N_2557);
nor U2608 (N_2608,N_2553,N_2528);
or U2609 (N_2609,N_2526,N_2559);
and U2610 (N_2610,N_2570,N_2573);
or U2611 (N_2611,N_2536,N_2542);
or U2612 (N_2612,N_2544,N_2566);
or U2613 (N_2613,N_2531,N_2565);
or U2614 (N_2614,N_2530,N_2533);
nor U2615 (N_2615,N_2569,N_2520);
or U2616 (N_2616,N_2579,N_2556);
nand U2617 (N_2617,N_2524,N_2573);
nor U2618 (N_2618,N_2535,N_2523);
or U2619 (N_2619,N_2523,N_2564);
and U2620 (N_2620,N_2570,N_2554);
nand U2621 (N_2621,N_2558,N_2577);
and U2622 (N_2622,N_2538,N_2540);
and U2623 (N_2623,N_2564,N_2566);
and U2624 (N_2624,N_2566,N_2560);
nand U2625 (N_2625,N_2534,N_2556);
and U2626 (N_2626,N_2523,N_2576);
nand U2627 (N_2627,N_2566,N_2557);
or U2628 (N_2628,N_2534,N_2525);
xnor U2629 (N_2629,N_2547,N_2538);
nand U2630 (N_2630,N_2527,N_2549);
or U2631 (N_2631,N_2526,N_2552);
nand U2632 (N_2632,N_2578,N_2573);
or U2633 (N_2633,N_2575,N_2568);
nor U2634 (N_2634,N_2547,N_2554);
or U2635 (N_2635,N_2542,N_2530);
nor U2636 (N_2636,N_2579,N_2557);
and U2637 (N_2637,N_2526,N_2577);
or U2638 (N_2638,N_2558,N_2562);
nor U2639 (N_2639,N_2521,N_2569);
nand U2640 (N_2640,N_2630,N_2607);
nor U2641 (N_2641,N_2584,N_2612);
nor U2642 (N_2642,N_2606,N_2627);
nor U2643 (N_2643,N_2621,N_2611);
or U2644 (N_2644,N_2596,N_2599);
or U2645 (N_2645,N_2631,N_2602);
nand U2646 (N_2646,N_2598,N_2605);
nor U2647 (N_2647,N_2600,N_2585);
or U2648 (N_2648,N_2615,N_2583);
nand U2649 (N_2649,N_2619,N_2592);
xnor U2650 (N_2650,N_2586,N_2609);
nor U2651 (N_2651,N_2625,N_2601);
or U2652 (N_2652,N_2622,N_2614);
xor U2653 (N_2653,N_2632,N_2595);
xor U2654 (N_2654,N_2639,N_2624);
xnor U2655 (N_2655,N_2638,N_2637);
nor U2656 (N_2656,N_2580,N_2618);
xnor U2657 (N_2657,N_2597,N_2589);
xor U2658 (N_2658,N_2613,N_2590);
and U2659 (N_2659,N_2591,N_2633);
and U2660 (N_2660,N_2636,N_2629);
nor U2661 (N_2661,N_2604,N_2620);
or U2662 (N_2662,N_2581,N_2608);
xor U2663 (N_2663,N_2634,N_2603);
nor U2664 (N_2664,N_2623,N_2616);
nor U2665 (N_2665,N_2617,N_2594);
nor U2666 (N_2666,N_2635,N_2587);
or U2667 (N_2667,N_2593,N_2626);
xor U2668 (N_2668,N_2582,N_2628);
nand U2669 (N_2669,N_2588,N_2610);
or U2670 (N_2670,N_2607,N_2619);
nand U2671 (N_2671,N_2603,N_2589);
and U2672 (N_2672,N_2637,N_2619);
or U2673 (N_2673,N_2622,N_2602);
nand U2674 (N_2674,N_2599,N_2607);
nor U2675 (N_2675,N_2628,N_2612);
and U2676 (N_2676,N_2629,N_2626);
or U2677 (N_2677,N_2584,N_2628);
or U2678 (N_2678,N_2636,N_2622);
nor U2679 (N_2679,N_2633,N_2599);
nand U2680 (N_2680,N_2591,N_2603);
nand U2681 (N_2681,N_2614,N_2609);
or U2682 (N_2682,N_2611,N_2593);
nor U2683 (N_2683,N_2582,N_2634);
nand U2684 (N_2684,N_2580,N_2611);
nand U2685 (N_2685,N_2581,N_2634);
and U2686 (N_2686,N_2585,N_2582);
or U2687 (N_2687,N_2621,N_2639);
nor U2688 (N_2688,N_2582,N_2586);
nand U2689 (N_2689,N_2599,N_2586);
nor U2690 (N_2690,N_2607,N_2603);
nand U2691 (N_2691,N_2630,N_2636);
nor U2692 (N_2692,N_2605,N_2603);
and U2693 (N_2693,N_2597,N_2582);
xnor U2694 (N_2694,N_2617,N_2588);
nand U2695 (N_2695,N_2605,N_2580);
xor U2696 (N_2696,N_2607,N_2617);
nor U2697 (N_2697,N_2611,N_2606);
nand U2698 (N_2698,N_2602,N_2593);
nor U2699 (N_2699,N_2599,N_2634);
and U2700 (N_2700,N_2693,N_2647);
and U2701 (N_2701,N_2688,N_2694);
nand U2702 (N_2702,N_2654,N_2643);
and U2703 (N_2703,N_2670,N_2689);
and U2704 (N_2704,N_2671,N_2696);
or U2705 (N_2705,N_2660,N_2642);
and U2706 (N_2706,N_2691,N_2658);
and U2707 (N_2707,N_2675,N_2697);
nor U2708 (N_2708,N_2672,N_2653);
or U2709 (N_2709,N_2668,N_2687);
nand U2710 (N_2710,N_2699,N_2678);
and U2711 (N_2711,N_2679,N_2649);
nor U2712 (N_2712,N_2666,N_2656);
and U2713 (N_2713,N_2695,N_2661);
and U2714 (N_2714,N_2677,N_2648);
nand U2715 (N_2715,N_2684,N_2673);
nor U2716 (N_2716,N_2674,N_2690);
xor U2717 (N_2717,N_2644,N_2657);
or U2718 (N_2718,N_2640,N_2682);
and U2719 (N_2719,N_2652,N_2667);
and U2720 (N_2720,N_2683,N_2664);
and U2721 (N_2721,N_2698,N_2665);
nand U2722 (N_2722,N_2686,N_2676);
and U2723 (N_2723,N_2650,N_2645);
or U2724 (N_2724,N_2680,N_2659);
nand U2725 (N_2725,N_2651,N_2669);
nor U2726 (N_2726,N_2641,N_2663);
nand U2727 (N_2727,N_2685,N_2655);
nand U2728 (N_2728,N_2662,N_2646);
or U2729 (N_2729,N_2692,N_2681);
nand U2730 (N_2730,N_2673,N_2689);
and U2731 (N_2731,N_2659,N_2665);
nand U2732 (N_2732,N_2644,N_2653);
and U2733 (N_2733,N_2640,N_2686);
and U2734 (N_2734,N_2663,N_2675);
xnor U2735 (N_2735,N_2697,N_2694);
or U2736 (N_2736,N_2686,N_2679);
nor U2737 (N_2737,N_2650,N_2659);
or U2738 (N_2738,N_2672,N_2695);
nand U2739 (N_2739,N_2668,N_2692);
or U2740 (N_2740,N_2655,N_2684);
nand U2741 (N_2741,N_2685,N_2660);
or U2742 (N_2742,N_2654,N_2697);
nor U2743 (N_2743,N_2678,N_2656);
nand U2744 (N_2744,N_2655,N_2686);
and U2745 (N_2745,N_2664,N_2680);
and U2746 (N_2746,N_2695,N_2670);
or U2747 (N_2747,N_2651,N_2696);
nand U2748 (N_2748,N_2647,N_2645);
nand U2749 (N_2749,N_2687,N_2666);
xor U2750 (N_2750,N_2651,N_2693);
or U2751 (N_2751,N_2671,N_2658);
nand U2752 (N_2752,N_2647,N_2656);
nor U2753 (N_2753,N_2661,N_2696);
and U2754 (N_2754,N_2664,N_2671);
or U2755 (N_2755,N_2641,N_2640);
and U2756 (N_2756,N_2681,N_2697);
nor U2757 (N_2757,N_2662,N_2645);
and U2758 (N_2758,N_2663,N_2689);
and U2759 (N_2759,N_2652,N_2697);
nand U2760 (N_2760,N_2717,N_2728);
nor U2761 (N_2761,N_2734,N_2753);
nor U2762 (N_2762,N_2716,N_2703);
or U2763 (N_2763,N_2743,N_2732);
nor U2764 (N_2764,N_2713,N_2710);
or U2765 (N_2765,N_2715,N_2720);
or U2766 (N_2766,N_2714,N_2744);
nand U2767 (N_2767,N_2757,N_2724);
nand U2768 (N_2768,N_2736,N_2739);
nand U2769 (N_2769,N_2731,N_2701);
nor U2770 (N_2770,N_2705,N_2706);
xnor U2771 (N_2771,N_2725,N_2750);
nand U2772 (N_2772,N_2704,N_2723);
and U2773 (N_2773,N_2748,N_2747);
and U2774 (N_2774,N_2737,N_2730);
nor U2775 (N_2775,N_2708,N_2756);
nand U2776 (N_2776,N_2742,N_2722);
and U2777 (N_2777,N_2727,N_2745);
nand U2778 (N_2778,N_2759,N_2735);
and U2779 (N_2779,N_2709,N_2733);
nor U2780 (N_2780,N_2712,N_2721);
or U2781 (N_2781,N_2740,N_2749);
nor U2782 (N_2782,N_2738,N_2758);
or U2783 (N_2783,N_2741,N_2711);
and U2784 (N_2784,N_2719,N_2752);
and U2785 (N_2785,N_2746,N_2718);
nand U2786 (N_2786,N_2754,N_2707);
or U2787 (N_2787,N_2700,N_2726);
nand U2788 (N_2788,N_2729,N_2755);
or U2789 (N_2789,N_2751,N_2702);
nor U2790 (N_2790,N_2710,N_2742);
or U2791 (N_2791,N_2720,N_2705);
xnor U2792 (N_2792,N_2700,N_2718);
nand U2793 (N_2793,N_2707,N_2742);
and U2794 (N_2794,N_2723,N_2736);
and U2795 (N_2795,N_2736,N_2722);
or U2796 (N_2796,N_2729,N_2758);
xnor U2797 (N_2797,N_2728,N_2750);
xor U2798 (N_2798,N_2707,N_2724);
nor U2799 (N_2799,N_2753,N_2751);
nand U2800 (N_2800,N_2747,N_2740);
nor U2801 (N_2801,N_2702,N_2708);
nand U2802 (N_2802,N_2701,N_2717);
nand U2803 (N_2803,N_2745,N_2705);
xnor U2804 (N_2804,N_2725,N_2758);
and U2805 (N_2805,N_2756,N_2723);
nor U2806 (N_2806,N_2711,N_2731);
or U2807 (N_2807,N_2720,N_2732);
nand U2808 (N_2808,N_2743,N_2717);
nor U2809 (N_2809,N_2730,N_2750);
nand U2810 (N_2810,N_2704,N_2707);
or U2811 (N_2811,N_2741,N_2742);
or U2812 (N_2812,N_2732,N_2737);
xnor U2813 (N_2813,N_2752,N_2712);
and U2814 (N_2814,N_2753,N_2737);
and U2815 (N_2815,N_2735,N_2728);
or U2816 (N_2816,N_2726,N_2702);
and U2817 (N_2817,N_2705,N_2737);
and U2818 (N_2818,N_2714,N_2741);
xnor U2819 (N_2819,N_2709,N_2741);
nand U2820 (N_2820,N_2819,N_2762);
nor U2821 (N_2821,N_2784,N_2805);
nand U2822 (N_2822,N_2812,N_2763);
or U2823 (N_2823,N_2800,N_2801);
nand U2824 (N_2824,N_2792,N_2780);
and U2825 (N_2825,N_2798,N_2782);
or U2826 (N_2826,N_2767,N_2799);
and U2827 (N_2827,N_2776,N_2808);
nor U2828 (N_2828,N_2771,N_2788);
nand U2829 (N_2829,N_2768,N_2765);
or U2830 (N_2830,N_2789,N_2806);
or U2831 (N_2831,N_2809,N_2794);
nor U2832 (N_2832,N_2786,N_2764);
nor U2833 (N_2833,N_2773,N_2760);
nor U2834 (N_2834,N_2811,N_2775);
nor U2835 (N_2835,N_2791,N_2796);
nor U2836 (N_2836,N_2797,N_2787);
and U2837 (N_2837,N_2774,N_2779);
and U2838 (N_2838,N_2810,N_2790);
nand U2839 (N_2839,N_2814,N_2766);
or U2840 (N_2840,N_2815,N_2802);
nor U2841 (N_2841,N_2803,N_2785);
nand U2842 (N_2842,N_2816,N_2761);
nor U2843 (N_2843,N_2793,N_2813);
or U2844 (N_2844,N_2804,N_2777);
nor U2845 (N_2845,N_2772,N_2769);
or U2846 (N_2846,N_2818,N_2778);
or U2847 (N_2847,N_2781,N_2795);
or U2848 (N_2848,N_2783,N_2770);
and U2849 (N_2849,N_2817,N_2807);
and U2850 (N_2850,N_2777,N_2784);
nor U2851 (N_2851,N_2811,N_2774);
or U2852 (N_2852,N_2780,N_2788);
nor U2853 (N_2853,N_2770,N_2790);
and U2854 (N_2854,N_2770,N_2784);
nand U2855 (N_2855,N_2795,N_2780);
nand U2856 (N_2856,N_2797,N_2786);
xnor U2857 (N_2857,N_2767,N_2813);
nand U2858 (N_2858,N_2792,N_2760);
xor U2859 (N_2859,N_2764,N_2807);
xnor U2860 (N_2860,N_2763,N_2767);
xnor U2861 (N_2861,N_2811,N_2766);
and U2862 (N_2862,N_2811,N_2802);
nor U2863 (N_2863,N_2794,N_2790);
nor U2864 (N_2864,N_2800,N_2799);
nor U2865 (N_2865,N_2819,N_2778);
or U2866 (N_2866,N_2784,N_2819);
or U2867 (N_2867,N_2814,N_2804);
and U2868 (N_2868,N_2763,N_2811);
xor U2869 (N_2869,N_2816,N_2800);
or U2870 (N_2870,N_2818,N_2776);
nor U2871 (N_2871,N_2770,N_2762);
or U2872 (N_2872,N_2809,N_2795);
nor U2873 (N_2873,N_2804,N_2762);
and U2874 (N_2874,N_2781,N_2806);
nand U2875 (N_2875,N_2781,N_2811);
nand U2876 (N_2876,N_2773,N_2809);
xnor U2877 (N_2877,N_2806,N_2809);
nand U2878 (N_2878,N_2781,N_2810);
nor U2879 (N_2879,N_2794,N_2800);
or U2880 (N_2880,N_2842,N_2872);
and U2881 (N_2881,N_2844,N_2853);
nor U2882 (N_2882,N_2865,N_2825);
nor U2883 (N_2883,N_2849,N_2831);
nor U2884 (N_2884,N_2834,N_2877);
nor U2885 (N_2885,N_2862,N_2871);
nand U2886 (N_2886,N_2873,N_2870);
nor U2887 (N_2887,N_2829,N_2852);
nor U2888 (N_2888,N_2826,N_2838);
and U2889 (N_2889,N_2824,N_2843);
nor U2890 (N_2890,N_2866,N_2821);
or U2891 (N_2891,N_2860,N_2837);
or U2892 (N_2892,N_2878,N_2869);
and U2893 (N_2893,N_2845,N_2840);
xor U2894 (N_2894,N_2836,N_2830);
or U2895 (N_2895,N_2854,N_2876);
and U2896 (N_2896,N_2848,N_2851);
or U2897 (N_2897,N_2863,N_2879);
and U2898 (N_2898,N_2833,N_2850);
nor U2899 (N_2899,N_2827,N_2864);
or U2900 (N_2900,N_2846,N_2839);
or U2901 (N_2901,N_2868,N_2822);
xnor U2902 (N_2902,N_2859,N_2856);
xnor U2903 (N_2903,N_2832,N_2874);
nand U2904 (N_2904,N_2847,N_2858);
nor U2905 (N_2905,N_2823,N_2857);
or U2906 (N_2906,N_2835,N_2875);
xnor U2907 (N_2907,N_2828,N_2820);
and U2908 (N_2908,N_2867,N_2861);
nand U2909 (N_2909,N_2855,N_2841);
xnor U2910 (N_2910,N_2825,N_2856);
xnor U2911 (N_2911,N_2849,N_2832);
or U2912 (N_2912,N_2839,N_2844);
or U2913 (N_2913,N_2826,N_2820);
or U2914 (N_2914,N_2879,N_2843);
xnor U2915 (N_2915,N_2873,N_2826);
nor U2916 (N_2916,N_2831,N_2848);
nor U2917 (N_2917,N_2825,N_2826);
nor U2918 (N_2918,N_2868,N_2854);
and U2919 (N_2919,N_2829,N_2878);
nand U2920 (N_2920,N_2834,N_2825);
nand U2921 (N_2921,N_2834,N_2822);
or U2922 (N_2922,N_2823,N_2855);
xor U2923 (N_2923,N_2838,N_2833);
or U2924 (N_2924,N_2864,N_2853);
or U2925 (N_2925,N_2843,N_2839);
and U2926 (N_2926,N_2875,N_2822);
nor U2927 (N_2927,N_2876,N_2873);
or U2928 (N_2928,N_2854,N_2840);
xor U2929 (N_2929,N_2832,N_2838);
xor U2930 (N_2930,N_2853,N_2850);
nor U2931 (N_2931,N_2871,N_2857);
nor U2932 (N_2932,N_2830,N_2842);
nor U2933 (N_2933,N_2840,N_2841);
nand U2934 (N_2934,N_2850,N_2855);
xor U2935 (N_2935,N_2849,N_2824);
and U2936 (N_2936,N_2834,N_2867);
nand U2937 (N_2937,N_2866,N_2860);
nand U2938 (N_2938,N_2866,N_2861);
and U2939 (N_2939,N_2820,N_2846);
nand U2940 (N_2940,N_2929,N_2903);
nor U2941 (N_2941,N_2939,N_2881);
xnor U2942 (N_2942,N_2924,N_2913);
nor U2943 (N_2943,N_2914,N_2917);
xor U2944 (N_2944,N_2911,N_2933);
or U2945 (N_2945,N_2899,N_2921);
nor U2946 (N_2946,N_2885,N_2928);
or U2947 (N_2947,N_2935,N_2906);
and U2948 (N_2948,N_2915,N_2931);
nand U2949 (N_2949,N_2888,N_2904);
and U2950 (N_2950,N_2920,N_2891);
or U2951 (N_2951,N_2934,N_2884);
and U2952 (N_2952,N_2883,N_2907);
or U2953 (N_2953,N_2901,N_2930);
nor U2954 (N_2954,N_2896,N_2938);
xor U2955 (N_2955,N_2910,N_2894);
or U2956 (N_2956,N_2926,N_2909);
nand U2957 (N_2957,N_2889,N_2895);
nor U2958 (N_2958,N_2922,N_2900);
xor U2959 (N_2959,N_2925,N_2927);
nand U2960 (N_2960,N_2905,N_2897);
and U2961 (N_2961,N_2937,N_2892);
nor U2962 (N_2962,N_2918,N_2893);
nand U2963 (N_2963,N_2898,N_2919);
nand U2964 (N_2964,N_2887,N_2908);
nor U2965 (N_2965,N_2932,N_2882);
and U2966 (N_2966,N_2880,N_2902);
nor U2967 (N_2967,N_2912,N_2916);
xnor U2968 (N_2968,N_2890,N_2936);
nor U2969 (N_2969,N_2923,N_2886);
or U2970 (N_2970,N_2901,N_2922);
and U2971 (N_2971,N_2913,N_2889);
or U2972 (N_2972,N_2896,N_2927);
nand U2973 (N_2973,N_2934,N_2922);
or U2974 (N_2974,N_2926,N_2923);
or U2975 (N_2975,N_2931,N_2939);
nand U2976 (N_2976,N_2934,N_2917);
and U2977 (N_2977,N_2937,N_2888);
nor U2978 (N_2978,N_2930,N_2893);
nor U2979 (N_2979,N_2922,N_2906);
or U2980 (N_2980,N_2922,N_2910);
nor U2981 (N_2981,N_2885,N_2933);
or U2982 (N_2982,N_2913,N_2887);
nand U2983 (N_2983,N_2885,N_2935);
nand U2984 (N_2984,N_2927,N_2917);
nand U2985 (N_2985,N_2885,N_2900);
or U2986 (N_2986,N_2920,N_2909);
nor U2987 (N_2987,N_2937,N_2903);
and U2988 (N_2988,N_2902,N_2916);
or U2989 (N_2989,N_2886,N_2936);
nor U2990 (N_2990,N_2900,N_2907);
or U2991 (N_2991,N_2907,N_2885);
and U2992 (N_2992,N_2917,N_2919);
nor U2993 (N_2993,N_2905,N_2888);
and U2994 (N_2994,N_2937,N_2897);
xnor U2995 (N_2995,N_2936,N_2928);
nand U2996 (N_2996,N_2895,N_2904);
nor U2997 (N_2997,N_2914,N_2920);
nor U2998 (N_2998,N_2920,N_2921);
nor U2999 (N_2999,N_2919,N_2899);
or UO_0 (O_0,N_2999,N_2983);
and UO_1 (O_1,N_2945,N_2963);
and UO_2 (O_2,N_2940,N_2993);
nand UO_3 (O_3,N_2946,N_2949);
nor UO_4 (O_4,N_2997,N_2978);
nor UO_5 (O_5,N_2960,N_2972);
and UO_6 (O_6,N_2962,N_2968);
xor UO_7 (O_7,N_2959,N_2988);
and UO_8 (O_8,N_2954,N_2966);
or UO_9 (O_9,N_2984,N_2969);
nor UO_10 (O_10,N_2977,N_2958);
nor UO_11 (O_11,N_2951,N_2957);
nor UO_12 (O_12,N_2961,N_2989);
and UO_13 (O_13,N_2976,N_2944);
xor UO_14 (O_14,N_2992,N_2975);
or UO_15 (O_15,N_2985,N_2967);
xnor UO_16 (O_16,N_2979,N_2995);
nand UO_17 (O_17,N_2964,N_2998);
nor UO_18 (O_18,N_2994,N_2956);
nor UO_19 (O_19,N_2986,N_2970);
nand UO_20 (O_20,N_2953,N_2981);
or UO_21 (O_21,N_2941,N_2942);
or UO_22 (O_22,N_2974,N_2943);
nand UO_23 (O_23,N_2965,N_2990);
and UO_24 (O_24,N_2948,N_2996);
xnor UO_25 (O_25,N_2955,N_2947);
nand UO_26 (O_26,N_2973,N_2982);
nand UO_27 (O_27,N_2987,N_2952);
nand UO_28 (O_28,N_2971,N_2991);
and UO_29 (O_29,N_2980,N_2950);
and UO_30 (O_30,N_2947,N_2992);
xor UO_31 (O_31,N_2992,N_2945);
nor UO_32 (O_32,N_2974,N_2961);
and UO_33 (O_33,N_2967,N_2964);
nand UO_34 (O_34,N_2963,N_2997);
nor UO_35 (O_35,N_2961,N_2979);
nor UO_36 (O_36,N_2940,N_2969);
or UO_37 (O_37,N_2964,N_2953);
and UO_38 (O_38,N_2987,N_2961);
nand UO_39 (O_39,N_2958,N_2968);
and UO_40 (O_40,N_2948,N_2940);
and UO_41 (O_41,N_2951,N_2968);
nand UO_42 (O_42,N_2970,N_2995);
and UO_43 (O_43,N_2992,N_2967);
and UO_44 (O_44,N_2970,N_2999);
nand UO_45 (O_45,N_2954,N_2985);
and UO_46 (O_46,N_2997,N_2979);
and UO_47 (O_47,N_2961,N_2973);
or UO_48 (O_48,N_2947,N_2984);
nor UO_49 (O_49,N_2980,N_2994);
and UO_50 (O_50,N_2978,N_2941);
nand UO_51 (O_51,N_2981,N_2987);
nand UO_52 (O_52,N_2943,N_2971);
nand UO_53 (O_53,N_2952,N_2947);
and UO_54 (O_54,N_2986,N_2951);
and UO_55 (O_55,N_2947,N_2990);
nor UO_56 (O_56,N_2956,N_2995);
and UO_57 (O_57,N_2993,N_2996);
or UO_58 (O_58,N_2968,N_2960);
nor UO_59 (O_59,N_2964,N_2965);
and UO_60 (O_60,N_2951,N_2979);
nor UO_61 (O_61,N_2998,N_2940);
or UO_62 (O_62,N_2966,N_2994);
nand UO_63 (O_63,N_2971,N_2968);
nand UO_64 (O_64,N_2980,N_2963);
or UO_65 (O_65,N_2961,N_2941);
and UO_66 (O_66,N_2971,N_2956);
nand UO_67 (O_67,N_2972,N_2995);
nor UO_68 (O_68,N_2943,N_2969);
xor UO_69 (O_69,N_2948,N_2977);
xnor UO_70 (O_70,N_2955,N_2970);
or UO_71 (O_71,N_2949,N_2974);
nor UO_72 (O_72,N_2990,N_2951);
or UO_73 (O_73,N_2966,N_2944);
nor UO_74 (O_74,N_2963,N_2966);
nand UO_75 (O_75,N_2979,N_2949);
nand UO_76 (O_76,N_2993,N_2966);
or UO_77 (O_77,N_2975,N_2959);
and UO_78 (O_78,N_2979,N_2993);
nand UO_79 (O_79,N_2940,N_2999);
nand UO_80 (O_80,N_2944,N_2946);
nand UO_81 (O_81,N_2983,N_2971);
nand UO_82 (O_82,N_2962,N_2959);
and UO_83 (O_83,N_2978,N_2952);
and UO_84 (O_84,N_2963,N_2975);
or UO_85 (O_85,N_2955,N_2998);
nor UO_86 (O_86,N_2975,N_2999);
nand UO_87 (O_87,N_2953,N_2957);
nand UO_88 (O_88,N_2976,N_2947);
or UO_89 (O_89,N_2947,N_2973);
nor UO_90 (O_90,N_2950,N_2978);
or UO_91 (O_91,N_2976,N_2972);
or UO_92 (O_92,N_2955,N_2985);
xor UO_93 (O_93,N_2951,N_2988);
and UO_94 (O_94,N_2958,N_2944);
or UO_95 (O_95,N_2949,N_2970);
or UO_96 (O_96,N_2964,N_2988);
and UO_97 (O_97,N_2957,N_2954);
nor UO_98 (O_98,N_2982,N_2993);
and UO_99 (O_99,N_2998,N_2970);
nor UO_100 (O_100,N_2961,N_2968);
nand UO_101 (O_101,N_2996,N_2997);
nand UO_102 (O_102,N_2980,N_2962);
xnor UO_103 (O_103,N_2972,N_2977);
or UO_104 (O_104,N_2949,N_2948);
nor UO_105 (O_105,N_2990,N_2950);
or UO_106 (O_106,N_2954,N_2992);
or UO_107 (O_107,N_2987,N_2971);
nor UO_108 (O_108,N_2991,N_2949);
or UO_109 (O_109,N_2954,N_2956);
or UO_110 (O_110,N_2975,N_2997);
nor UO_111 (O_111,N_2981,N_2988);
nor UO_112 (O_112,N_2942,N_2964);
and UO_113 (O_113,N_2978,N_2957);
nand UO_114 (O_114,N_2994,N_2957);
and UO_115 (O_115,N_2961,N_2970);
and UO_116 (O_116,N_2952,N_2982);
nor UO_117 (O_117,N_2985,N_2943);
xnor UO_118 (O_118,N_2962,N_2946);
or UO_119 (O_119,N_2943,N_2978);
xnor UO_120 (O_120,N_2953,N_2954);
and UO_121 (O_121,N_2998,N_2946);
nand UO_122 (O_122,N_2952,N_2968);
nand UO_123 (O_123,N_2970,N_2980);
xnor UO_124 (O_124,N_2972,N_2957);
xor UO_125 (O_125,N_2960,N_2981);
nor UO_126 (O_126,N_2994,N_2960);
nand UO_127 (O_127,N_2958,N_2986);
or UO_128 (O_128,N_2945,N_2974);
xnor UO_129 (O_129,N_2985,N_2960);
nor UO_130 (O_130,N_2972,N_2987);
xnor UO_131 (O_131,N_2997,N_2941);
or UO_132 (O_132,N_2970,N_2987);
nand UO_133 (O_133,N_2955,N_2956);
nand UO_134 (O_134,N_2969,N_2944);
or UO_135 (O_135,N_2973,N_2976);
and UO_136 (O_136,N_2944,N_2964);
nand UO_137 (O_137,N_2982,N_2994);
nor UO_138 (O_138,N_2988,N_2945);
nand UO_139 (O_139,N_2955,N_2944);
and UO_140 (O_140,N_2971,N_2965);
nand UO_141 (O_141,N_2989,N_2950);
or UO_142 (O_142,N_2954,N_2969);
or UO_143 (O_143,N_2986,N_2954);
nor UO_144 (O_144,N_2957,N_2968);
and UO_145 (O_145,N_2944,N_2947);
xor UO_146 (O_146,N_2964,N_2961);
and UO_147 (O_147,N_2955,N_2980);
nand UO_148 (O_148,N_2962,N_2960);
and UO_149 (O_149,N_2944,N_2975);
nor UO_150 (O_150,N_2966,N_2952);
nor UO_151 (O_151,N_2956,N_2952);
and UO_152 (O_152,N_2947,N_2968);
or UO_153 (O_153,N_2999,N_2947);
or UO_154 (O_154,N_2952,N_2985);
nand UO_155 (O_155,N_2981,N_2951);
xnor UO_156 (O_156,N_2992,N_2963);
or UO_157 (O_157,N_2985,N_2941);
or UO_158 (O_158,N_2959,N_2992);
nor UO_159 (O_159,N_2956,N_2997);
or UO_160 (O_160,N_2977,N_2990);
nor UO_161 (O_161,N_2983,N_2987);
or UO_162 (O_162,N_2955,N_2984);
nor UO_163 (O_163,N_2992,N_2942);
nor UO_164 (O_164,N_2950,N_2968);
nor UO_165 (O_165,N_2972,N_2965);
or UO_166 (O_166,N_2968,N_2949);
or UO_167 (O_167,N_2962,N_2986);
and UO_168 (O_168,N_2949,N_2955);
or UO_169 (O_169,N_2953,N_2998);
nor UO_170 (O_170,N_2986,N_2974);
and UO_171 (O_171,N_2948,N_2946);
nor UO_172 (O_172,N_2982,N_2972);
nor UO_173 (O_173,N_2954,N_2979);
or UO_174 (O_174,N_2975,N_2960);
nand UO_175 (O_175,N_2944,N_2942);
xor UO_176 (O_176,N_2964,N_2983);
and UO_177 (O_177,N_2940,N_2996);
and UO_178 (O_178,N_2965,N_2947);
nand UO_179 (O_179,N_2945,N_2972);
nor UO_180 (O_180,N_2958,N_2963);
nor UO_181 (O_181,N_2983,N_2998);
or UO_182 (O_182,N_2972,N_2978);
nor UO_183 (O_183,N_2999,N_2964);
nand UO_184 (O_184,N_2975,N_2988);
nor UO_185 (O_185,N_2974,N_2983);
xnor UO_186 (O_186,N_2968,N_2975);
or UO_187 (O_187,N_2987,N_2956);
or UO_188 (O_188,N_2991,N_2966);
xnor UO_189 (O_189,N_2956,N_2981);
nand UO_190 (O_190,N_2941,N_2967);
or UO_191 (O_191,N_2983,N_2991);
or UO_192 (O_192,N_2962,N_2947);
nor UO_193 (O_193,N_2948,N_2981);
nand UO_194 (O_194,N_2941,N_2944);
nand UO_195 (O_195,N_2949,N_2992);
nor UO_196 (O_196,N_2963,N_2978);
and UO_197 (O_197,N_2986,N_2961);
nand UO_198 (O_198,N_2986,N_2978);
or UO_199 (O_199,N_2991,N_2998);
or UO_200 (O_200,N_2969,N_2994);
and UO_201 (O_201,N_2956,N_2943);
nor UO_202 (O_202,N_2981,N_2970);
nand UO_203 (O_203,N_2968,N_2948);
or UO_204 (O_204,N_2979,N_2965);
and UO_205 (O_205,N_2941,N_2994);
nand UO_206 (O_206,N_2942,N_2959);
and UO_207 (O_207,N_2981,N_2991);
and UO_208 (O_208,N_2964,N_2962);
xnor UO_209 (O_209,N_2945,N_2977);
nand UO_210 (O_210,N_2993,N_2949);
nor UO_211 (O_211,N_2970,N_2959);
and UO_212 (O_212,N_2974,N_2979);
and UO_213 (O_213,N_2986,N_2989);
or UO_214 (O_214,N_2965,N_2945);
nand UO_215 (O_215,N_2999,N_2984);
xor UO_216 (O_216,N_2986,N_2988);
nor UO_217 (O_217,N_2995,N_2971);
and UO_218 (O_218,N_2951,N_2989);
or UO_219 (O_219,N_2995,N_2989);
and UO_220 (O_220,N_2988,N_2952);
or UO_221 (O_221,N_2998,N_2952);
and UO_222 (O_222,N_2947,N_2988);
nand UO_223 (O_223,N_2982,N_2988);
or UO_224 (O_224,N_2973,N_2959);
nor UO_225 (O_225,N_2984,N_2974);
or UO_226 (O_226,N_2988,N_2962);
or UO_227 (O_227,N_2969,N_2997);
xnor UO_228 (O_228,N_2963,N_2954);
nand UO_229 (O_229,N_2968,N_2959);
or UO_230 (O_230,N_2994,N_2947);
nand UO_231 (O_231,N_2963,N_2994);
and UO_232 (O_232,N_2964,N_2952);
nor UO_233 (O_233,N_2990,N_2998);
or UO_234 (O_234,N_2977,N_2980);
and UO_235 (O_235,N_2961,N_2955);
nand UO_236 (O_236,N_2981,N_2998);
nand UO_237 (O_237,N_2966,N_2980);
nand UO_238 (O_238,N_2996,N_2961);
nand UO_239 (O_239,N_2995,N_2994);
and UO_240 (O_240,N_2967,N_2960);
nor UO_241 (O_241,N_2995,N_2990);
and UO_242 (O_242,N_2992,N_2971);
or UO_243 (O_243,N_2977,N_2964);
and UO_244 (O_244,N_2978,N_2968);
nand UO_245 (O_245,N_2997,N_2955);
nor UO_246 (O_246,N_2944,N_2984);
nor UO_247 (O_247,N_2946,N_2977);
and UO_248 (O_248,N_2961,N_2959);
xnor UO_249 (O_249,N_2999,N_2954);
or UO_250 (O_250,N_2985,N_2946);
and UO_251 (O_251,N_2972,N_2956);
nand UO_252 (O_252,N_2958,N_2940);
nor UO_253 (O_253,N_2944,N_2963);
nand UO_254 (O_254,N_2967,N_2949);
and UO_255 (O_255,N_2997,N_2972);
nor UO_256 (O_256,N_2959,N_2998);
or UO_257 (O_257,N_2995,N_2959);
or UO_258 (O_258,N_2995,N_2986);
xnor UO_259 (O_259,N_2997,N_2940);
or UO_260 (O_260,N_2973,N_2979);
or UO_261 (O_261,N_2998,N_2996);
nor UO_262 (O_262,N_2991,N_2996);
or UO_263 (O_263,N_2943,N_2960);
or UO_264 (O_264,N_2986,N_2976);
nor UO_265 (O_265,N_2972,N_2942);
nor UO_266 (O_266,N_2999,N_2950);
nor UO_267 (O_267,N_2992,N_2972);
nand UO_268 (O_268,N_2970,N_2957);
nand UO_269 (O_269,N_2953,N_2989);
or UO_270 (O_270,N_2985,N_2963);
nand UO_271 (O_271,N_2949,N_2997);
nand UO_272 (O_272,N_2981,N_2952);
and UO_273 (O_273,N_2954,N_2962);
or UO_274 (O_274,N_2987,N_2963);
nand UO_275 (O_275,N_2953,N_2946);
or UO_276 (O_276,N_2942,N_2997);
and UO_277 (O_277,N_2968,N_2967);
nand UO_278 (O_278,N_2977,N_2965);
or UO_279 (O_279,N_2994,N_2946);
xor UO_280 (O_280,N_2984,N_2981);
and UO_281 (O_281,N_2945,N_2949);
nor UO_282 (O_282,N_2958,N_2997);
nor UO_283 (O_283,N_2951,N_2971);
nand UO_284 (O_284,N_2941,N_2964);
nand UO_285 (O_285,N_2956,N_2977);
nand UO_286 (O_286,N_2954,N_2945);
or UO_287 (O_287,N_2966,N_2964);
and UO_288 (O_288,N_2985,N_2957);
and UO_289 (O_289,N_2974,N_2995);
or UO_290 (O_290,N_2975,N_2957);
xor UO_291 (O_291,N_2948,N_2986);
and UO_292 (O_292,N_2948,N_2972);
or UO_293 (O_293,N_2957,N_2991);
nor UO_294 (O_294,N_2955,N_2946);
nand UO_295 (O_295,N_2991,N_2999);
nand UO_296 (O_296,N_2953,N_2977);
or UO_297 (O_297,N_2983,N_2954);
nor UO_298 (O_298,N_2982,N_2940);
or UO_299 (O_299,N_2970,N_2992);
xnor UO_300 (O_300,N_2958,N_2948);
or UO_301 (O_301,N_2992,N_2998);
or UO_302 (O_302,N_2975,N_2954);
and UO_303 (O_303,N_2946,N_2999);
nand UO_304 (O_304,N_2982,N_2986);
nand UO_305 (O_305,N_2952,N_2967);
nor UO_306 (O_306,N_2983,N_2941);
and UO_307 (O_307,N_2959,N_2967);
or UO_308 (O_308,N_2998,N_2945);
or UO_309 (O_309,N_2994,N_2958);
nand UO_310 (O_310,N_2978,N_2947);
or UO_311 (O_311,N_2977,N_2984);
nor UO_312 (O_312,N_2949,N_2990);
nor UO_313 (O_313,N_2971,N_2999);
xnor UO_314 (O_314,N_2990,N_2961);
and UO_315 (O_315,N_2964,N_2960);
nor UO_316 (O_316,N_2957,N_2948);
nor UO_317 (O_317,N_2971,N_2996);
nand UO_318 (O_318,N_2960,N_2956);
and UO_319 (O_319,N_2987,N_2982);
nor UO_320 (O_320,N_2978,N_2969);
and UO_321 (O_321,N_2973,N_2989);
or UO_322 (O_322,N_2977,N_2969);
or UO_323 (O_323,N_2987,N_2993);
or UO_324 (O_324,N_2974,N_2994);
or UO_325 (O_325,N_2990,N_2992);
xor UO_326 (O_326,N_2949,N_2956);
xor UO_327 (O_327,N_2961,N_2997);
and UO_328 (O_328,N_2974,N_2989);
and UO_329 (O_329,N_2964,N_2958);
or UO_330 (O_330,N_2956,N_2941);
or UO_331 (O_331,N_2941,N_2958);
xnor UO_332 (O_332,N_2958,N_2983);
nor UO_333 (O_333,N_2974,N_2952);
xor UO_334 (O_334,N_2997,N_2993);
and UO_335 (O_335,N_2960,N_2989);
nand UO_336 (O_336,N_2945,N_2950);
nand UO_337 (O_337,N_2954,N_2998);
nand UO_338 (O_338,N_2982,N_2958);
and UO_339 (O_339,N_2964,N_2978);
and UO_340 (O_340,N_2966,N_2953);
and UO_341 (O_341,N_2978,N_2960);
and UO_342 (O_342,N_2997,N_2986);
and UO_343 (O_343,N_2980,N_2952);
or UO_344 (O_344,N_2944,N_2979);
xor UO_345 (O_345,N_2978,N_2953);
nor UO_346 (O_346,N_2965,N_2946);
nor UO_347 (O_347,N_2971,N_2955);
nand UO_348 (O_348,N_2949,N_2986);
nor UO_349 (O_349,N_2976,N_2971);
and UO_350 (O_350,N_2965,N_2957);
or UO_351 (O_351,N_2956,N_2942);
nand UO_352 (O_352,N_2940,N_2992);
nor UO_353 (O_353,N_2966,N_2987);
or UO_354 (O_354,N_2951,N_2950);
nand UO_355 (O_355,N_2984,N_2997);
nand UO_356 (O_356,N_2961,N_2992);
nor UO_357 (O_357,N_2991,N_2987);
nor UO_358 (O_358,N_2996,N_2949);
nor UO_359 (O_359,N_2989,N_2978);
or UO_360 (O_360,N_2953,N_2979);
nor UO_361 (O_361,N_2967,N_2978);
or UO_362 (O_362,N_2991,N_2997);
or UO_363 (O_363,N_2972,N_2944);
and UO_364 (O_364,N_2971,N_2974);
or UO_365 (O_365,N_2986,N_2944);
or UO_366 (O_366,N_2940,N_2976);
or UO_367 (O_367,N_2990,N_2973);
xor UO_368 (O_368,N_2943,N_2970);
and UO_369 (O_369,N_2990,N_2981);
and UO_370 (O_370,N_2959,N_2994);
nor UO_371 (O_371,N_2985,N_2951);
and UO_372 (O_372,N_2992,N_2964);
or UO_373 (O_373,N_2993,N_2981);
or UO_374 (O_374,N_2946,N_2943);
and UO_375 (O_375,N_2951,N_2999);
or UO_376 (O_376,N_2954,N_2978);
xor UO_377 (O_377,N_2985,N_2995);
nor UO_378 (O_378,N_2945,N_2964);
nor UO_379 (O_379,N_2968,N_2986);
and UO_380 (O_380,N_2947,N_2980);
and UO_381 (O_381,N_2998,N_2961);
nand UO_382 (O_382,N_2995,N_2998);
xnor UO_383 (O_383,N_2956,N_2984);
nor UO_384 (O_384,N_2962,N_2989);
and UO_385 (O_385,N_2987,N_2959);
and UO_386 (O_386,N_2970,N_2985);
or UO_387 (O_387,N_2994,N_2984);
nand UO_388 (O_388,N_2945,N_2980);
nor UO_389 (O_389,N_2983,N_2966);
or UO_390 (O_390,N_2967,N_2980);
nor UO_391 (O_391,N_2993,N_2973);
and UO_392 (O_392,N_2977,N_2973);
and UO_393 (O_393,N_2954,N_2989);
nand UO_394 (O_394,N_2954,N_2991);
and UO_395 (O_395,N_2987,N_2968);
nor UO_396 (O_396,N_2991,N_2964);
or UO_397 (O_397,N_2981,N_2964);
or UO_398 (O_398,N_2990,N_2959);
nand UO_399 (O_399,N_2947,N_2979);
and UO_400 (O_400,N_2947,N_2986);
nand UO_401 (O_401,N_2995,N_2987);
or UO_402 (O_402,N_2949,N_2947);
xnor UO_403 (O_403,N_2943,N_2979);
or UO_404 (O_404,N_2999,N_2997);
nor UO_405 (O_405,N_2972,N_2973);
nor UO_406 (O_406,N_2977,N_2940);
nor UO_407 (O_407,N_2953,N_2996);
nand UO_408 (O_408,N_2973,N_2997);
xnor UO_409 (O_409,N_2954,N_2984);
nor UO_410 (O_410,N_2940,N_2984);
nand UO_411 (O_411,N_2990,N_2968);
and UO_412 (O_412,N_2992,N_2958);
nor UO_413 (O_413,N_2943,N_2998);
or UO_414 (O_414,N_2946,N_2958);
or UO_415 (O_415,N_2944,N_2983);
nor UO_416 (O_416,N_2961,N_2958);
or UO_417 (O_417,N_2944,N_2998);
nand UO_418 (O_418,N_2973,N_2954);
or UO_419 (O_419,N_2952,N_2999);
xnor UO_420 (O_420,N_2970,N_2967);
and UO_421 (O_421,N_2950,N_2948);
or UO_422 (O_422,N_2955,N_2979);
xnor UO_423 (O_423,N_2977,N_2941);
nand UO_424 (O_424,N_2958,N_2945);
and UO_425 (O_425,N_2980,N_2984);
nand UO_426 (O_426,N_2979,N_2999);
and UO_427 (O_427,N_2950,N_2944);
nand UO_428 (O_428,N_2962,N_2953);
and UO_429 (O_429,N_2949,N_2950);
or UO_430 (O_430,N_2976,N_2996);
nor UO_431 (O_431,N_2995,N_2960);
nor UO_432 (O_432,N_2988,N_2943);
xnor UO_433 (O_433,N_2997,N_2950);
and UO_434 (O_434,N_2977,N_2995);
nand UO_435 (O_435,N_2943,N_2955);
nand UO_436 (O_436,N_2963,N_2943);
nor UO_437 (O_437,N_2943,N_2984);
nor UO_438 (O_438,N_2963,N_2947);
nor UO_439 (O_439,N_2970,N_2964);
nor UO_440 (O_440,N_2952,N_2953);
or UO_441 (O_441,N_2987,N_2998);
or UO_442 (O_442,N_2947,N_2966);
or UO_443 (O_443,N_2976,N_2969);
nor UO_444 (O_444,N_2970,N_2975);
nand UO_445 (O_445,N_2996,N_2985);
and UO_446 (O_446,N_2948,N_2982);
nand UO_447 (O_447,N_2948,N_2945);
nor UO_448 (O_448,N_2966,N_2977);
xnor UO_449 (O_449,N_2962,N_2975);
or UO_450 (O_450,N_2988,N_2944);
and UO_451 (O_451,N_2959,N_2965);
and UO_452 (O_452,N_2948,N_2942);
and UO_453 (O_453,N_2985,N_2976);
nor UO_454 (O_454,N_2950,N_2970);
or UO_455 (O_455,N_2999,N_2985);
nor UO_456 (O_456,N_2999,N_2981);
nor UO_457 (O_457,N_2966,N_2960);
nor UO_458 (O_458,N_2991,N_2992);
nand UO_459 (O_459,N_2954,N_2987);
and UO_460 (O_460,N_2981,N_2977);
and UO_461 (O_461,N_2999,N_2960);
nor UO_462 (O_462,N_2941,N_2974);
nand UO_463 (O_463,N_2983,N_2981);
nor UO_464 (O_464,N_2978,N_2961);
nand UO_465 (O_465,N_2984,N_2963);
nand UO_466 (O_466,N_2969,N_2991);
xnor UO_467 (O_467,N_2966,N_2969);
or UO_468 (O_468,N_2972,N_2954);
nor UO_469 (O_469,N_2995,N_2948);
and UO_470 (O_470,N_2950,N_2987);
nor UO_471 (O_471,N_2998,N_2982);
nor UO_472 (O_472,N_2989,N_2990);
nor UO_473 (O_473,N_2961,N_2949);
nand UO_474 (O_474,N_2942,N_2999);
or UO_475 (O_475,N_2956,N_2962);
or UO_476 (O_476,N_2968,N_2955);
or UO_477 (O_477,N_2965,N_2948);
xor UO_478 (O_478,N_2961,N_2962);
xnor UO_479 (O_479,N_2969,N_2945);
nor UO_480 (O_480,N_2985,N_2978);
or UO_481 (O_481,N_2965,N_2974);
or UO_482 (O_482,N_2951,N_2965);
nand UO_483 (O_483,N_2982,N_2977);
nor UO_484 (O_484,N_2983,N_2943);
or UO_485 (O_485,N_2940,N_2983);
nand UO_486 (O_486,N_2981,N_2954);
xor UO_487 (O_487,N_2956,N_2944);
or UO_488 (O_488,N_2996,N_2959);
nor UO_489 (O_489,N_2966,N_2972);
or UO_490 (O_490,N_2980,N_2965);
or UO_491 (O_491,N_2947,N_2971);
nand UO_492 (O_492,N_2989,N_2998);
nand UO_493 (O_493,N_2947,N_2961);
or UO_494 (O_494,N_2974,N_2958);
or UO_495 (O_495,N_2966,N_2946);
xnor UO_496 (O_496,N_2976,N_2984);
nand UO_497 (O_497,N_2992,N_2983);
or UO_498 (O_498,N_2988,N_2940);
or UO_499 (O_499,N_2950,N_2964);
endmodule