module basic_1000_10000_1500_4_levels_10xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
xor U0 (N_0,In_690,In_162);
xor U1 (N_1,In_369,In_395);
or U2 (N_2,In_186,In_916);
xnor U3 (N_3,In_294,In_919);
xnor U4 (N_4,In_967,In_798);
or U5 (N_5,In_229,In_138);
nand U6 (N_6,In_361,In_340);
and U7 (N_7,In_167,In_911);
xnor U8 (N_8,In_292,In_713);
xnor U9 (N_9,In_654,In_929);
and U10 (N_10,In_195,In_758);
nor U11 (N_11,In_693,In_691);
and U12 (N_12,In_778,In_549);
and U13 (N_13,In_100,In_663);
nand U14 (N_14,In_692,In_764);
nand U15 (N_15,In_850,In_187);
nand U16 (N_16,In_446,In_683);
nor U17 (N_17,In_439,In_180);
nand U18 (N_18,In_134,In_62);
nand U19 (N_19,In_587,In_259);
nor U20 (N_20,In_770,In_814);
xor U21 (N_21,In_788,In_556);
xor U22 (N_22,In_91,In_989);
and U23 (N_23,In_241,In_791);
and U24 (N_24,In_226,In_102);
xor U25 (N_25,In_511,In_615);
nand U26 (N_26,In_506,In_812);
and U27 (N_27,In_321,In_430);
nor U28 (N_28,In_390,In_284);
and U29 (N_29,In_961,In_22);
nand U30 (N_30,In_290,In_279);
xor U31 (N_31,In_924,In_86);
nand U32 (N_32,In_732,In_478);
nand U33 (N_33,In_101,In_740);
nor U34 (N_34,In_533,In_816);
nand U35 (N_35,In_640,In_135);
nand U36 (N_36,In_328,In_928);
xor U37 (N_37,In_391,In_348);
nand U38 (N_38,In_76,In_116);
and U39 (N_39,In_394,In_819);
or U40 (N_40,In_917,In_69);
and U41 (N_41,In_337,In_273);
nand U42 (N_42,In_119,In_277);
and U43 (N_43,In_23,In_425);
xnor U44 (N_44,In_884,In_742);
xor U45 (N_45,In_635,In_811);
and U46 (N_46,In_753,In_338);
nor U47 (N_47,In_293,In_659);
xor U48 (N_48,In_623,In_28);
nor U49 (N_49,In_146,In_652);
or U50 (N_50,In_926,In_530);
or U51 (N_51,In_107,In_60);
nand U52 (N_52,In_589,In_233);
or U53 (N_53,In_963,In_952);
nor U54 (N_54,In_477,In_730);
xor U55 (N_55,In_359,In_260);
nand U56 (N_56,In_156,In_970);
nor U57 (N_57,In_888,In_795);
nor U58 (N_58,In_974,In_143);
or U59 (N_59,In_876,In_120);
nor U60 (N_60,In_262,In_643);
xnor U61 (N_61,In_196,In_968);
xor U62 (N_62,In_527,In_131);
and U63 (N_63,In_422,In_224);
nand U64 (N_64,In_96,In_631);
nor U65 (N_65,In_859,In_936);
nand U66 (N_66,In_949,In_65);
and U67 (N_67,In_784,In_649);
xor U68 (N_68,In_786,In_345);
xor U69 (N_69,In_848,In_665);
nand U70 (N_70,In_809,In_699);
xor U71 (N_71,In_695,In_87);
and U72 (N_72,In_492,In_948);
xor U73 (N_73,In_160,In_433);
and U74 (N_74,In_800,In_801);
or U75 (N_75,In_611,In_452);
and U76 (N_76,In_53,In_144);
or U77 (N_77,In_985,In_573);
or U78 (N_78,In_435,In_902);
nor U79 (N_79,In_577,In_36);
and U80 (N_80,In_222,In_515);
nor U81 (N_81,In_310,In_320);
or U82 (N_82,In_839,In_669);
or U83 (N_83,In_227,In_341);
nand U84 (N_84,In_548,In_558);
nand U85 (N_85,In_810,In_593);
nor U86 (N_86,In_317,In_873);
xor U87 (N_87,In_373,In_955);
or U88 (N_88,In_567,In_600);
xnor U89 (N_89,In_921,In_214);
nand U90 (N_90,In_104,In_736);
xor U91 (N_91,In_90,In_257);
nor U92 (N_92,In_271,In_482);
or U93 (N_93,In_35,In_426);
and U94 (N_94,In_891,In_918);
xnor U95 (N_95,In_37,In_441);
nand U96 (N_96,In_325,In_163);
and U97 (N_97,In_804,In_721);
xnor U98 (N_98,In_516,In_201);
and U99 (N_99,In_415,In_639);
xnor U100 (N_100,In_507,In_137);
nand U101 (N_101,In_582,In_268);
nor U102 (N_102,In_109,In_75);
and U103 (N_103,In_825,In_49);
nor U104 (N_104,In_706,In_702);
nand U105 (N_105,In_776,In_152);
or U106 (N_106,In_124,In_51);
and U107 (N_107,In_269,In_574);
nor U108 (N_108,In_553,In_579);
nand U109 (N_109,In_202,In_913);
nand U110 (N_110,In_738,In_563);
nand U111 (N_111,In_746,In_755);
xnor U112 (N_112,In_841,In_89);
or U113 (N_113,In_40,In_765);
xnor U114 (N_114,In_779,In_541);
and U115 (N_115,In_38,In_844);
or U116 (N_116,In_523,In_774);
nand U117 (N_117,In_991,In_469);
nor U118 (N_118,In_200,In_980);
nor U119 (N_119,In_302,In_8);
or U120 (N_120,In_676,In_629);
nand U121 (N_121,In_0,In_757);
xor U122 (N_122,In_169,In_912);
xor U123 (N_123,In_191,In_367);
xor U124 (N_124,In_904,In_682);
and U125 (N_125,In_455,In_34);
nor U126 (N_126,In_684,In_552);
or U127 (N_127,In_19,In_243);
nor U128 (N_128,In_418,In_951);
and U129 (N_129,In_865,In_495);
and U130 (N_130,In_215,In_80);
nand U131 (N_131,In_771,In_655);
nand U132 (N_132,In_164,In_990);
nand U133 (N_133,In_249,In_493);
xor U134 (N_134,In_539,In_641);
or U135 (N_135,In_524,In_638);
and U136 (N_136,In_922,In_324);
xor U137 (N_137,In_940,In_650);
nand U138 (N_138,In_608,In_339);
nor U139 (N_139,In_939,In_453);
or U140 (N_140,In_451,In_205);
and U141 (N_141,In_898,In_383);
nand U142 (N_142,In_569,In_729);
and U143 (N_143,In_303,In_956);
nand U144 (N_144,In_977,In_725);
xnor U145 (N_145,In_591,In_762);
nor U146 (N_146,In_806,In_993);
and U147 (N_147,In_688,In_835);
or U148 (N_148,In_709,In_518);
nor U149 (N_149,In_845,In_385);
or U150 (N_150,In_463,In_905);
nand U151 (N_151,In_712,In_342);
and U152 (N_152,In_934,In_356);
and U153 (N_153,In_68,In_7);
xnor U154 (N_154,In_467,In_903);
nor U155 (N_155,In_796,In_698);
xnor U156 (N_156,In_807,In_25);
or U157 (N_157,In_946,In_246);
nand U158 (N_158,In_216,In_722);
nor U159 (N_159,In_618,In_603);
nor U160 (N_160,In_283,In_71);
nand U161 (N_161,In_554,In_16);
xnor U162 (N_162,In_645,In_999);
nor U163 (N_163,In_672,In_941);
xor U164 (N_164,In_781,In_166);
nand U165 (N_165,In_609,In_741);
nor U166 (N_166,In_14,In_363);
or U167 (N_167,In_975,In_769);
and U168 (N_168,In_247,In_937);
nor U169 (N_169,In_947,In_127);
nand U170 (N_170,In_250,In_847);
or U171 (N_171,In_123,In_910);
and U172 (N_172,In_923,In_59);
and U173 (N_173,In_174,In_330);
nand U174 (N_174,In_994,In_756);
and U175 (N_175,In_909,In_719);
or U176 (N_176,In_128,In_856);
nor U177 (N_177,In_365,In_677);
nor U178 (N_178,In_67,In_57);
nor U179 (N_179,In_536,In_766);
and U180 (N_180,In_381,In_235);
xnor U181 (N_181,In_817,In_846);
or U182 (N_182,In_431,In_126);
nor U183 (N_183,In_759,In_983);
nor U184 (N_184,In_625,In_595);
nor U185 (N_185,In_48,In_175);
nor U186 (N_186,In_851,In_136);
and U187 (N_187,In_319,In_84);
and U188 (N_188,In_462,In_565);
and U189 (N_189,In_354,In_972);
or U190 (N_190,In_318,In_583);
nor U191 (N_191,In_855,In_378);
nand U192 (N_192,In_838,In_397);
or U193 (N_193,In_417,In_94);
and U194 (N_194,In_464,In_761);
nand U195 (N_195,In_636,In_969);
nand U196 (N_196,In_519,In_237);
nand U197 (N_197,In_456,In_885);
or U198 (N_198,In_334,In_327);
nor U199 (N_199,In_475,In_529);
or U200 (N_200,In_785,In_935);
nor U201 (N_201,In_389,In_125);
nor U202 (N_202,In_520,In_476);
or U203 (N_203,In_863,In_590);
or U204 (N_204,In_960,In_624);
or U205 (N_205,In_617,In_945);
or U206 (N_206,In_468,In_177);
nand U207 (N_207,In_872,In_188);
nor U208 (N_208,In_943,In_184);
and U209 (N_209,In_564,In_305);
xnor U210 (N_210,In_353,In_117);
nand U211 (N_211,In_570,In_255);
and U212 (N_212,In_165,In_656);
or U213 (N_213,In_933,In_559);
and U214 (N_214,In_2,In_323);
and U215 (N_215,In_723,In_352);
and U216 (N_216,In_890,In_209);
xor U217 (N_217,In_998,In_280);
xnor U218 (N_218,In_108,In_388);
or U219 (N_219,In_958,In_878);
nor U220 (N_220,In_39,In_364);
xnor U221 (N_221,In_379,In_82);
nand U222 (N_222,In_472,In_555);
or U223 (N_223,In_634,In_295);
xor U224 (N_224,In_883,In_997);
or U225 (N_225,In_981,In_500);
nand U226 (N_226,In_460,In_704);
nor U227 (N_227,In_687,In_892);
nand U228 (N_228,In_276,In_501);
and U229 (N_229,In_21,In_139);
and U230 (N_230,In_103,In_517);
or U231 (N_231,In_289,In_427);
or U232 (N_232,In_63,In_802);
xor U233 (N_233,In_147,In_987);
nor U234 (N_234,In_489,In_457);
and U235 (N_235,In_833,In_777);
xor U236 (N_236,In_199,In_572);
nor U237 (N_237,In_627,In_782);
nand U238 (N_238,In_930,In_11);
nand U239 (N_239,In_560,In_278);
xnor U240 (N_240,In_964,In_313);
or U241 (N_241,In_794,In_874);
and U242 (N_242,In_444,In_258);
nand U243 (N_243,In_207,In_375);
nor U244 (N_244,In_6,In_576);
or U245 (N_245,In_894,In_537);
or U246 (N_246,In_331,In_680);
xor U247 (N_247,In_543,In_773);
nand U248 (N_248,In_132,In_424);
nor U249 (N_249,In_410,In_965);
and U250 (N_250,In_689,In_944);
xor U251 (N_251,In_97,In_20);
and U252 (N_252,In_263,In_950);
nor U253 (N_253,In_105,In_648);
and U254 (N_254,In_308,In_868);
and U255 (N_255,In_896,In_72);
nand U256 (N_256,In_604,In_13);
xor U257 (N_257,In_402,In_172);
or U258 (N_258,In_953,In_571);
or U259 (N_259,In_971,In_920);
and U260 (N_260,In_984,In_74);
nor U261 (N_261,In_895,In_301);
nand U262 (N_262,In_875,In_106);
and U263 (N_263,In_628,In_822);
xor U264 (N_264,In_178,In_612);
nor U265 (N_265,In_133,In_538);
nand U266 (N_266,In_646,In_190);
or U267 (N_267,In_197,In_957);
and U268 (N_268,In_889,In_403);
and U269 (N_269,In_907,In_27);
nand U270 (N_270,In_157,In_244);
xor U271 (N_271,In_607,In_661);
xor U272 (N_272,In_803,In_154);
nor U273 (N_273,In_853,In_580);
nand U274 (N_274,In_220,In_252);
xor U275 (N_275,In_219,In_182);
xor U276 (N_276,In_854,In_508);
and U277 (N_277,In_33,In_843);
or U278 (N_278,In_540,In_978);
nand U279 (N_279,In_392,In_708);
and U280 (N_280,In_414,In_743);
nand U281 (N_281,In_266,In_221);
nand U282 (N_282,In_85,In_597);
xnor U283 (N_283,In_931,In_5);
xnor U284 (N_284,In_73,In_445);
nor U285 (N_285,In_396,In_992);
nand U286 (N_286,In_996,In_438);
nand U287 (N_287,In_808,In_360);
or U288 (N_288,In_61,In_897);
or U289 (N_289,In_31,In_528);
xnor U290 (N_290,In_401,In_473);
xnor U291 (N_291,In_670,In_561);
xnor U292 (N_292,In_52,In_783);
or U293 (N_293,In_288,In_265);
and U294 (N_294,In_578,In_599);
and U295 (N_295,In_179,In_357);
xnor U296 (N_296,In_588,In_299);
nor U297 (N_297,In_432,In_459);
and U298 (N_298,In_717,In_314);
xor U299 (N_299,In_678,In_881);
nand U300 (N_300,In_551,In_17);
nor U301 (N_301,In_88,In_275);
xnor U302 (N_302,In_306,In_867);
and U303 (N_303,In_54,In_355);
nand U304 (N_304,In_830,In_217);
nand U305 (N_305,In_542,In_685);
and U306 (N_306,In_606,In_58);
nand U307 (N_307,In_242,In_510);
or U308 (N_308,In_1,In_793);
xnor U309 (N_309,In_824,In_316);
nor U310 (N_310,In_236,In_218);
nor U311 (N_311,In_701,In_925);
xnor U312 (N_312,In_821,In_416);
xor U313 (N_313,In_50,In_512);
nor U314 (N_314,In_326,In_601);
nand U315 (N_315,In_142,In_705);
xor U316 (N_316,In_679,In_248);
and U317 (N_317,In_448,In_716);
nand U318 (N_318,In_210,In_155);
and U319 (N_319,In_387,In_836);
or U320 (N_320,In_181,In_532);
nand U321 (N_321,In_789,In_747);
nand U322 (N_322,In_272,In_366);
xor U323 (N_323,In_647,In_291);
or U324 (N_324,In_203,In_79);
nand U325 (N_325,In_681,In_882);
nand U326 (N_326,In_380,In_4);
and U327 (N_327,In_828,In_77);
or U328 (N_328,In_813,In_942);
nor U329 (N_329,In_792,In_421);
and U330 (N_330,In_976,In_899);
or U331 (N_331,In_474,In_129);
or U332 (N_332,In_485,In_377);
and U333 (N_333,In_727,In_95);
nand U334 (N_334,In_228,In_660);
or U335 (N_335,In_498,In_461);
and U336 (N_336,In_534,In_98);
nor U337 (N_337,In_823,In_232);
and U338 (N_338,In_915,In_644);
nand U339 (N_339,In_393,In_158);
and U340 (N_340,In_906,In_121);
nor U341 (N_341,In_592,In_491);
and U342 (N_342,In_488,In_546);
nand U343 (N_343,In_711,In_99);
nand U344 (N_344,In_633,In_862);
xor U345 (N_345,In_440,In_333);
nor U346 (N_346,In_988,In_55);
nand U347 (N_347,In_406,In_70);
xor U348 (N_348,In_322,In_151);
xnor U349 (N_349,In_986,In_831);
or U350 (N_350,In_503,In_442);
or U351 (N_351,In_304,In_637);
and U352 (N_352,In_42,In_535);
nand U353 (N_353,In_479,In_173);
nor U354 (N_354,In_145,In_256);
or U355 (N_355,In_733,In_531);
nor U356 (N_356,In_651,In_505);
or U357 (N_357,In_307,In_797);
and U358 (N_358,In_760,In_194);
nand U359 (N_359,In_312,In_487);
and U360 (N_360,In_398,In_412);
and U361 (N_361,In_858,In_621);
and U362 (N_362,In_657,In_871);
or U363 (N_363,In_545,In_526);
or U364 (N_364,In_471,In_9);
nor U365 (N_365,In_349,In_399);
nand U366 (N_366,In_213,In_668);
and U367 (N_367,In_168,In_893);
or U368 (N_368,In_544,In_336);
and U369 (N_369,In_632,In_423);
xnor U370 (N_370,In_286,In_613);
or U371 (N_371,In_726,In_602);
xnor U372 (N_372,In_724,In_92);
xnor U373 (N_373,In_409,In_66);
nor U374 (N_374,In_18,In_739);
nand U375 (N_375,In_400,In_877);
nor U376 (N_376,In_405,In_522);
or U377 (N_377,In_973,In_763);
or U378 (N_378,In_658,In_490);
or U379 (N_379,In_300,In_297);
or U380 (N_380,In_240,In_829);
nor U381 (N_381,In_56,In_112);
or U382 (N_382,In_370,In_662);
nand U383 (N_383,In_745,In_212);
or U384 (N_384,In_696,In_620);
nand U385 (N_385,In_787,In_118);
or U386 (N_386,In_26,In_447);
xnor U387 (N_387,In_581,In_768);
and U388 (N_388,In_914,In_234);
and U389 (N_389,In_857,In_486);
nand U390 (N_390,In_799,In_64);
and U391 (N_391,In_332,In_481);
nand U392 (N_392,In_864,In_496);
xnor U393 (N_393,In_351,In_932);
xor U394 (N_394,In_413,In_206);
nand U395 (N_395,In_767,In_170);
nor U396 (N_396,In_982,In_251);
nand U397 (N_397,In_115,In_282);
nor U398 (N_398,In_211,In_509);
nand U399 (N_399,In_616,In_605);
xnor U400 (N_400,In_586,In_750);
nand U401 (N_401,In_153,In_285);
or U402 (N_402,In_962,In_230);
xnor U403 (N_403,In_870,In_887);
nor U404 (N_404,In_737,In_880);
nand U405 (N_405,In_466,In_826);
nor U406 (N_406,In_513,In_562);
xnor U407 (N_407,In_264,In_208);
nor U408 (N_408,In_497,In_827);
nand U409 (N_409,In_347,In_450);
or U410 (N_410,In_484,In_130);
xor U411 (N_411,In_630,In_869);
nor U412 (N_412,In_386,In_666);
or U413 (N_413,In_12,In_309);
and U414 (N_414,In_24,In_959);
nand U415 (N_415,In_81,In_350);
nor U416 (N_416,In_780,In_614);
or U417 (N_417,In_966,In_298);
nor U418 (N_418,In_734,In_483);
xnor U419 (N_419,In_346,In_596);
or U420 (N_420,In_458,In_674);
and U421 (N_421,In_584,In_449);
nor U422 (N_422,In_594,In_411);
or U423 (N_423,In_335,In_470);
or U424 (N_424,In_311,In_428);
nor U425 (N_425,In_110,In_749);
or U426 (N_426,In_382,In_502);
or U427 (N_427,In_225,In_30);
nor U428 (N_428,In_707,In_642);
and U429 (N_429,In_566,In_610);
and U430 (N_430,In_671,In_720);
and U431 (N_431,In_267,In_113);
and U432 (N_432,In_374,In_710);
nor U433 (N_433,In_254,In_407);
nand U434 (N_434,In_368,In_238);
nand U435 (N_435,In_815,In_751);
or U436 (N_436,In_694,In_46);
or U437 (N_437,In_748,In_420);
nor U438 (N_438,In_122,In_183);
xnor U439 (N_439,In_189,In_287);
and U440 (N_440,In_901,In_735);
or U441 (N_441,In_731,In_465);
and U442 (N_442,In_192,In_329);
or U443 (N_443,In_419,In_198);
and U444 (N_444,In_772,In_840);
and U445 (N_445,In_842,In_626);
nor U446 (N_446,In_32,In_111);
or U447 (N_447,In_775,In_820);
or U448 (N_448,In_886,In_852);
nor U449 (N_449,In_45,In_622);
or U450 (N_450,In_41,In_667);
nand U451 (N_451,In_480,In_752);
and U452 (N_452,In_141,In_499);
xor U453 (N_453,In_979,In_140);
and U454 (N_454,In_550,In_525);
and U455 (N_455,In_404,In_832);
nor U456 (N_456,In_47,In_714);
nand U457 (N_457,In_700,In_673);
and U458 (N_458,In_575,In_239);
or U459 (N_459,In_185,In_245);
or U460 (N_460,In_664,In_204);
nor U461 (N_461,In_270,In_900);
xnor U462 (N_462,In_860,In_557);
xnor U463 (N_463,In_274,In_149);
or U464 (N_464,In_866,In_231);
nand U465 (N_465,In_568,In_429);
xnor U466 (N_466,In_261,In_78);
nand U467 (N_467,In_454,In_150);
and U468 (N_468,In_83,In_44);
and U469 (N_469,In_315,In_927);
nor U470 (N_470,In_954,In_43);
xnor U471 (N_471,In_514,In_358);
and U472 (N_472,In_504,In_3);
and U473 (N_473,In_818,In_223);
nor U474 (N_474,In_371,In_908);
nor U475 (N_475,In_408,In_10);
xor U476 (N_476,In_653,In_703);
or U477 (N_477,In_861,In_15);
nand U478 (N_478,In_343,In_879);
or U479 (N_479,In_494,In_376);
or U480 (N_480,In_114,In_718);
and U481 (N_481,In_344,In_754);
xnor U482 (N_482,In_715,In_790);
xor U483 (N_483,In_437,In_686);
nand U484 (N_484,In_521,In_362);
nor U485 (N_485,In_938,In_598);
and U486 (N_486,In_436,In_744);
nand U487 (N_487,In_161,In_434);
nand U488 (N_488,In_171,In_296);
and U489 (N_489,In_805,In_193);
nor U490 (N_490,In_29,In_585);
and U491 (N_491,In_253,In_148);
nand U492 (N_492,In_176,In_728);
or U493 (N_493,In_372,In_159);
and U494 (N_494,In_547,In_697);
nand U495 (N_495,In_849,In_93);
or U496 (N_496,In_619,In_281);
or U497 (N_497,In_837,In_443);
or U498 (N_498,In_384,In_834);
nand U499 (N_499,In_995,In_675);
and U500 (N_500,In_913,In_517);
nand U501 (N_501,In_698,In_443);
nor U502 (N_502,In_836,In_634);
xor U503 (N_503,In_459,In_682);
nor U504 (N_504,In_969,In_517);
or U505 (N_505,In_194,In_728);
or U506 (N_506,In_49,In_805);
nor U507 (N_507,In_355,In_551);
xnor U508 (N_508,In_721,In_538);
or U509 (N_509,In_155,In_778);
or U510 (N_510,In_109,In_669);
nor U511 (N_511,In_707,In_797);
and U512 (N_512,In_121,In_341);
and U513 (N_513,In_182,In_260);
nor U514 (N_514,In_908,In_287);
xor U515 (N_515,In_637,In_711);
xnor U516 (N_516,In_391,In_320);
or U517 (N_517,In_989,In_42);
and U518 (N_518,In_321,In_343);
or U519 (N_519,In_367,In_530);
nor U520 (N_520,In_535,In_751);
nand U521 (N_521,In_596,In_40);
nand U522 (N_522,In_265,In_980);
and U523 (N_523,In_183,In_753);
nor U524 (N_524,In_579,In_915);
or U525 (N_525,In_764,In_704);
xnor U526 (N_526,In_696,In_416);
xor U527 (N_527,In_833,In_824);
and U528 (N_528,In_878,In_471);
and U529 (N_529,In_381,In_4);
nor U530 (N_530,In_543,In_53);
or U531 (N_531,In_553,In_250);
nand U532 (N_532,In_322,In_853);
xnor U533 (N_533,In_15,In_340);
xor U534 (N_534,In_986,In_538);
nor U535 (N_535,In_286,In_827);
xor U536 (N_536,In_598,In_610);
nand U537 (N_537,In_458,In_810);
xnor U538 (N_538,In_23,In_9);
xor U539 (N_539,In_593,In_659);
nand U540 (N_540,In_400,In_195);
and U541 (N_541,In_959,In_91);
nand U542 (N_542,In_879,In_314);
nor U543 (N_543,In_315,In_286);
xnor U544 (N_544,In_849,In_971);
xnor U545 (N_545,In_925,In_801);
and U546 (N_546,In_906,In_823);
nand U547 (N_547,In_479,In_106);
and U548 (N_548,In_825,In_942);
or U549 (N_549,In_32,In_593);
or U550 (N_550,In_740,In_310);
and U551 (N_551,In_634,In_77);
and U552 (N_552,In_247,In_942);
and U553 (N_553,In_195,In_454);
nor U554 (N_554,In_811,In_117);
nand U555 (N_555,In_172,In_65);
xor U556 (N_556,In_700,In_417);
and U557 (N_557,In_855,In_141);
xor U558 (N_558,In_67,In_96);
or U559 (N_559,In_518,In_794);
xor U560 (N_560,In_936,In_764);
or U561 (N_561,In_103,In_361);
xnor U562 (N_562,In_109,In_470);
or U563 (N_563,In_260,In_570);
nor U564 (N_564,In_14,In_359);
and U565 (N_565,In_179,In_899);
nor U566 (N_566,In_181,In_255);
or U567 (N_567,In_587,In_498);
and U568 (N_568,In_850,In_252);
nor U569 (N_569,In_969,In_340);
xnor U570 (N_570,In_21,In_102);
nand U571 (N_571,In_785,In_267);
or U572 (N_572,In_426,In_706);
nor U573 (N_573,In_955,In_308);
nor U574 (N_574,In_446,In_356);
xnor U575 (N_575,In_671,In_46);
and U576 (N_576,In_462,In_19);
nor U577 (N_577,In_9,In_145);
or U578 (N_578,In_437,In_661);
or U579 (N_579,In_667,In_401);
nor U580 (N_580,In_202,In_363);
or U581 (N_581,In_19,In_201);
and U582 (N_582,In_264,In_868);
and U583 (N_583,In_214,In_349);
nand U584 (N_584,In_974,In_278);
nor U585 (N_585,In_411,In_912);
nor U586 (N_586,In_668,In_960);
and U587 (N_587,In_477,In_868);
or U588 (N_588,In_252,In_95);
and U589 (N_589,In_402,In_595);
nand U590 (N_590,In_785,In_683);
or U591 (N_591,In_576,In_500);
nor U592 (N_592,In_834,In_461);
nand U593 (N_593,In_621,In_709);
or U594 (N_594,In_550,In_641);
nand U595 (N_595,In_928,In_615);
or U596 (N_596,In_498,In_895);
or U597 (N_597,In_74,In_878);
nor U598 (N_598,In_665,In_316);
nor U599 (N_599,In_878,In_880);
nand U600 (N_600,In_803,In_783);
nand U601 (N_601,In_312,In_13);
and U602 (N_602,In_550,In_769);
nand U603 (N_603,In_371,In_107);
nand U604 (N_604,In_284,In_95);
nor U605 (N_605,In_10,In_212);
nand U606 (N_606,In_972,In_15);
or U607 (N_607,In_11,In_394);
and U608 (N_608,In_215,In_286);
nor U609 (N_609,In_739,In_377);
or U610 (N_610,In_418,In_929);
and U611 (N_611,In_900,In_603);
nor U612 (N_612,In_773,In_304);
xor U613 (N_613,In_454,In_172);
nand U614 (N_614,In_902,In_626);
xnor U615 (N_615,In_626,In_931);
nand U616 (N_616,In_572,In_708);
or U617 (N_617,In_955,In_918);
xnor U618 (N_618,In_34,In_82);
xnor U619 (N_619,In_463,In_654);
xor U620 (N_620,In_227,In_137);
nor U621 (N_621,In_900,In_806);
xor U622 (N_622,In_203,In_211);
nor U623 (N_623,In_608,In_705);
nand U624 (N_624,In_391,In_706);
and U625 (N_625,In_76,In_379);
nor U626 (N_626,In_926,In_510);
nor U627 (N_627,In_991,In_503);
xnor U628 (N_628,In_327,In_430);
nor U629 (N_629,In_152,In_765);
xor U630 (N_630,In_726,In_905);
xor U631 (N_631,In_900,In_980);
nor U632 (N_632,In_412,In_667);
nor U633 (N_633,In_372,In_150);
and U634 (N_634,In_731,In_78);
nand U635 (N_635,In_649,In_740);
xor U636 (N_636,In_73,In_508);
nand U637 (N_637,In_322,In_947);
xor U638 (N_638,In_195,In_457);
nand U639 (N_639,In_154,In_281);
nor U640 (N_640,In_843,In_611);
nor U641 (N_641,In_924,In_138);
nor U642 (N_642,In_168,In_518);
and U643 (N_643,In_119,In_453);
nor U644 (N_644,In_284,In_401);
nand U645 (N_645,In_777,In_338);
nand U646 (N_646,In_907,In_867);
and U647 (N_647,In_747,In_543);
or U648 (N_648,In_427,In_39);
nor U649 (N_649,In_690,In_225);
and U650 (N_650,In_970,In_977);
nor U651 (N_651,In_950,In_962);
nor U652 (N_652,In_490,In_876);
xnor U653 (N_653,In_944,In_883);
and U654 (N_654,In_721,In_510);
and U655 (N_655,In_240,In_192);
or U656 (N_656,In_581,In_532);
or U657 (N_657,In_332,In_570);
nand U658 (N_658,In_219,In_649);
or U659 (N_659,In_704,In_302);
and U660 (N_660,In_904,In_391);
or U661 (N_661,In_73,In_836);
nor U662 (N_662,In_411,In_787);
xor U663 (N_663,In_811,In_472);
xor U664 (N_664,In_866,In_327);
nor U665 (N_665,In_724,In_930);
xor U666 (N_666,In_70,In_939);
or U667 (N_667,In_833,In_637);
nor U668 (N_668,In_777,In_464);
or U669 (N_669,In_628,In_87);
nor U670 (N_670,In_166,In_61);
or U671 (N_671,In_889,In_557);
xor U672 (N_672,In_265,In_282);
or U673 (N_673,In_118,In_69);
nor U674 (N_674,In_959,In_639);
and U675 (N_675,In_623,In_908);
and U676 (N_676,In_272,In_277);
or U677 (N_677,In_0,In_141);
and U678 (N_678,In_343,In_519);
and U679 (N_679,In_982,In_168);
or U680 (N_680,In_29,In_239);
xnor U681 (N_681,In_451,In_994);
or U682 (N_682,In_699,In_26);
xor U683 (N_683,In_326,In_463);
nand U684 (N_684,In_353,In_507);
and U685 (N_685,In_190,In_609);
nor U686 (N_686,In_665,In_500);
xor U687 (N_687,In_977,In_277);
nand U688 (N_688,In_617,In_94);
nor U689 (N_689,In_311,In_415);
xnor U690 (N_690,In_981,In_20);
or U691 (N_691,In_988,In_936);
and U692 (N_692,In_360,In_950);
nor U693 (N_693,In_693,In_549);
and U694 (N_694,In_183,In_441);
or U695 (N_695,In_83,In_458);
and U696 (N_696,In_83,In_982);
nor U697 (N_697,In_156,In_633);
or U698 (N_698,In_595,In_409);
and U699 (N_699,In_197,In_296);
nor U700 (N_700,In_107,In_684);
or U701 (N_701,In_2,In_5);
and U702 (N_702,In_461,In_985);
nand U703 (N_703,In_446,In_543);
or U704 (N_704,In_689,In_153);
and U705 (N_705,In_978,In_591);
nor U706 (N_706,In_814,In_553);
and U707 (N_707,In_575,In_815);
nor U708 (N_708,In_747,In_859);
or U709 (N_709,In_716,In_39);
and U710 (N_710,In_101,In_133);
or U711 (N_711,In_920,In_962);
or U712 (N_712,In_201,In_664);
and U713 (N_713,In_447,In_706);
xor U714 (N_714,In_34,In_589);
xor U715 (N_715,In_795,In_313);
nand U716 (N_716,In_878,In_279);
and U717 (N_717,In_752,In_679);
and U718 (N_718,In_443,In_5);
nor U719 (N_719,In_966,In_192);
and U720 (N_720,In_853,In_613);
nand U721 (N_721,In_162,In_933);
or U722 (N_722,In_112,In_870);
xor U723 (N_723,In_775,In_17);
nor U724 (N_724,In_373,In_191);
nand U725 (N_725,In_630,In_938);
nand U726 (N_726,In_685,In_539);
nand U727 (N_727,In_15,In_226);
nor U728 (N_728,In_915,In_530);
nor U729 (N_729,In_856,In_506);
and U730 (N_730,In_80,In_480);
and U731 (N_731,In_614,In_588);
nand U732 (N_732,In_475,In_660);
or U733 (N_733,In_783,In_453);
or U734 (N_734,In_119,In_589);
or U735 (N_735,In_621,In_815);
nor U736 (N_736,In_947,In_191);
and U737 (N_737,In_952,In_106);
nand U738 (N_738,In_252,In_674);
xnor U739 (N_739,In_133,In_405);
nor U740 (N_740,In_597,In_154);
or U741 (N_741,In_695,In_33);
and U742 (N_742,In_65,In_518);
xnor U743 (N_743,In_677,In_595);
xor U744 (N_744,In_793,In_391);
and U745 (N_745,In_353,In_914);
or U746 (N_746,In_195,In_227);
or U747 (N_747,In_799,In_804);
nor U748 (N_748,In_348,In_396);
and U749 (N_749,In_211,In_681);
or U750 (N_750,In_215,In_5);
xnor U751 (N_751,In_347,In_61);
nor U752 (N_752,In_742,In_24);
nor U753 (N_753,In_387,In_304);
or U754 (N_754,In_343,In_643);
nand U755 (N_755,In_599,In_846);
xor U756 (N_756,In_62,In_810);
xnor U757 (N_757,In_448,In_296);
and U758 (N_758,In_580,In_982);
nand U759 (N_759,In_145,In_760);
or U760 (N_760,In_655,In_565);
and U761 (N_761,In_734,In_101);
nand U762 (N_762,In_613,In_39);
and U763 (N_763,In_319,In_865);
or U764 (N_764,In_404,In_584);
and U765 (N_765,In_662,In_757);
and U766 (N_766,In_118,In_115);
or U767 (N_767,In_940,In_328);
xnor U768 (N_768,In_247,In_804);
xor U769 (N_769,In_144,In_15);
xor U770 (N_770,In_659,In_978);
nand U771 (N_771,In_678,In_560);
nor U772 (N_772,In_166,In_734);
or U773 (N_773,In_448,In_372);
nand U774 (N_774,In_860,In_102);
and U775 (N_775,In_872,In_346);
nor U776 (N_776,In_874,In_531);
nor U777 (N_777,In_261,In_327);
nor U778 (N_778,In_76,In_454);
nand U779 (N_779,In_408,In_905);
xnor U780 (N_780,In_255,In_377);
nor U781 (N_781,In_738,In_699);
xor U782 (N_782,In_89,In_840);
nor U783 (N_783,In_239,In_255);
nand U784 (N_784,In_120,In_547);
and U785 (N_785,In_793,In_223);
and U786 (N_786,In_180,In_752);
nor U787 (N_787,In_963,In_695);
xnor U788 (N_788,In_324,In_567);
nor U789 (N_789,In_73,In_37);
and U790 (N_790,In_686,In_826);
nand U791 (N_791,In_749,In_514);
and U792 (N_792,In_308,In_36);
nor U793 (N_793,In_871,In_543);
and U794 (N_794,In_494,In_831);
or U795 (N_795,In_226,In_13);
nor U796 (N_796,In_296,In_607);
and U797 (N_797,In_301,In_149);
or U798 (N_798,In_192,In_838);
and U799 (N_799,In_711,In_101);
nor U800 (N_800,In_747,In_194);
or U801 (N_801,In_281,In_673);
or U802 (N_802,In_92,In_817);
or U803 (N_803,In_816,In_679);
nand U804 (N_804,In_204,In_771);
and U805 (N_805,In_630,In_151);
nor U806 (N_806,In_383,In_449);
nor U807 (N_807,In_440,In_809);
and U808 (N_808,In_886,In_490);
nand U809 (N_809,In_296,In_587);
or U810 (N_810,In_191,In_926);
or U811 (N_811,In_149,In_263);
and U812 (N_812,In_639,In_373);
nor U813 (N_813,In_260,In_698);
nand U814 (N_814,In_532,In_324);
or U815 (N_815,In_101,In_679);
or U816 (N_816,In_445,In_122);
and U817 (N_817,In_272,In_869);
xnor U818 (N_818,In_633,In_253);
nand U819 (N_819,In_189,In_250);
nand U820 (N_820,In_927,In_665);
xnor U821 (N_821,In_501,In_545);
nand U822 (N_822,In_627,In_469);
xor U823 (N_823,In_872,In_350);
or U824 (N_824,In_20,In_644);
xor U825 (N_825,In_251,In_438);
nor U826 (N_826,In_628,In_263);
nand U827 (N_827,In_352,In_415);
and U828 (N_828,In_389,In_128);
and U829 (N_829,In_114,In_522);
nor U830 (N_830,In_597,In_684);
xnor U831 (N_831,In_643,In_964);
nand U832 (N_832,In_784,In_822);
or U833 (N_833,In_309,In_135);
or U834 (N_834,In_653,In_556);
or U835 (N_835,In_792,In_94);
nand U836 (N_836,In_416,In_118);
nor U837 (N_837,In_211,In_290);
xnor U838 (N_838,In_329,In_959);
and U839 (N_839,In_645,In_871);
nand U840 (N_840,In_8,In_991);
or U841 (N_841,In_641,In_123);
nor U842 (N_842,In_507,In_0);
or U843 (N_843,In_16,In_381);
nand U844 (N_844,In_733,In_190);
nor U845 (N_845,In_55,In_471);
and U846 (N_846,In_42,In_943);
or U847 (N_847,In_538,In_368);
xnor U848 (N_848,In_253,In_400);
xnor U849 (N_849,In_519,In_861);
nand U850 (N_850,In_605,In_33);
and U851 (N_851,In_703,In_179);
and U852 (N_852,In_343,In_168);
and U853 (N_853,In_135,In_606);
or U854 (N_854,In_979,In_610);
and U855 (N_855,In_196,In_988);
nand U856 (N_856,In_760,In_468);
xnor U857 (N_857,In_625,In_692);
nand U858 (N_858,In_394,In_170);
xor U859 (N_859,In_435,In_171);
nand U860 (N_860,In_198,In_499);
xnor U861 (N_861,In_897,In_63);
nand U862 (N_862,In_944,In_80);
and U863 (N_863,In_489,In_971);
nand U864 (N_864,In_955,In_395);
nor U865 (N_865,In_839,In_224);
or U866 (N_866,In_255,In_435);
nand U867 (N_867,In_486,In_833);
xor U868 (N_868,In_472,In_349);
nor U869 (N_869,In_6,In_471);
nand U870 (N_870,In_386,In_130);
nor U871 (N_871,In_298,In_258);
and U872 (N_872,In_689,In_141);
or U873 (N_873,In_337,In_743);
nor U874 (N_874,In_547,In_706);
nand U875 (N_875,In_175,In_456);
or U876 (N_876,In_498,In_677);
and U877 (N_877,In_197,In_930);
or U878 (N_878,In_689,In_285);
and U879 (N_879,In_255,In_294);
xor U880 (N_880,In_572,In_40);
nand U881 (N_881,In_516,In_740);
nand U882 (N_882,In_765,In_919);
nand U883 (N_883,In_469,In_551);
nand U884 (N_884,In_925,In_582);
and U885 (N_885,In_891,In_591);
or U886 (N_886,In_394,In_281);
nor U887 (N_887,In_751,In_729);
nor U888 (N_888,In_424,In_887);
nor U889 (N_889,In_242,In_177);
nand U890 (N_890,In_562,In_821);
xnor U891 (N_891,In_115,In_257);
nor U892 (N_892,In_308,In_142);
nand U893 (N_893,In_912,In_592);
or U894 (N_894,In_396,In_118);
and U895 (N_895,In_180,In_243);
nand U896 (N_896,In_28,In_549);
nand U897 (N_897,In_127,In_791);
nand U898 (N_898,In_216,In_542);
xor U899 (N_899,In_593,In_338);
or U900 (N_900,In_563,In_543);
or U901 (N_901,In_516,In_312);
xnor U902 (N_902,In_329,In_358);
and U903 (N_903,In_636,In_607);
and U904 (N_904,In_721,In_281);
or U905 (N_905,In_137,In_487);
and U906 (N_906,In_854,In_269);
or U907 (N_907,In_879,In_283);
xnor U908 (N_908,In_445,In_367);
xnor U909 (N_909,In_590,In_310);
xnor U910 (N_910,In_584,In_20);
or U911 (N_911,In_79,In_941);
nor U912 (N_912,In_206,In_456);
and U913 (N_913,In_463,In_871);
and U914 (N_914,In_483,In_501);
or U915 (N_915,In_243,In_257);
or U916 (N_916,In_552,In_395);
nor U917 (N_917,In_495,In_447);
nand U918 (N_918,In_575,In_600);
and U919 (N_919,In_425,In_698);
nand U920 (N_920,In_677,In_828);
and U921 (N_921,In_351,In_613);
nor U922 (N_922,In_703,In_570);
and U923 (N_923,In_957,In_388);
nand U924 (N_924,In_80,In_892);
nand U925 (N_925,In_46,In_446);
and U926 (N_926,In_796,In_133);
or U927 (N_927,In_425,In_842);
nand U928 (N_928,In_650,In_926);
or U929 (N_929,In_558,In_601);
nor U930 (N_930,In_43,In_285);
nor U931 (N_931,In_348,In_158);
and U932 (N_932,In_213,In_648);
and U933 (N_933,In_647,In_567);
and U934 (N_934,In_534,In_399);
and U935 (N_935,In_339,In_917);
and U936 (N_936,In_343,In_567);
nand U937 (N_937,In_978,In_55);
or U938 (N_938,In_757,In_456);
xnor U939 (N_939,In_149,In_64);
or U940 (N_940,In_194,In_400);
nor U941 (N_941,In_446,In_621);
nor U942 (N_942,In_784,In_715);
nand U943 (N_943,In_900,In_822);
and U944 (N_944,In_116,In_675);
xor U945 (N_945,In_111,In_658);
or U946 (N_946,In_255,In_188);
nand U947 (N_947,In_858,In_347);
and U948 (N_948,In_770,In_310);
or U949 (N_949,In_280,In_89);
nor U950 (N_950,In_6,In_831);
xnor U951 (N_951,In_122,In_287);
or U952 (N_952,In_200,In_343);
and U953 (N_953,In_256,In_314);
xnor U954 (N_954,In_925,In_359);
xnor U955 (N_955,In_642,In_459);
or U956 (N_956,In_58,In_292);
and U957 (N_957,In_517,In_663);
nand U958 (N_958,In_892,In_732);
nand U959 (N_959,In_927,In_173);
nand U960 (N_960,In_646,In_743);
or U961 (N_961,In_634,In_676);
xnor U962 (N_962,In_426,In_793);
xnor U963 (N_963,In_971,In_435);
xor U964 (N_964,In_908,In_526);
and U965 (N_965,In_783,In_923);
nand U966 (N_966,In_471,In_304);
nand U967 (N_967,In_613,In_547);
or U968 (N_968,In_116,In_752);
and U969 (N_969,In_87,In_311);
nand U970 (N_970,In_570,In_200);
xnor U971 (N_971,In_431,In_898);
or U972 (N_972,In_171,In_299);
and U973 (N_973,In_547,In_700);
and U974 (N_974,In_786,In_360);
or U975 (N_975,In_729,In_585);
or U976 (N_976,In_2,In_659);
or U977 (N_977,In_643,In_358);
nand U978 (N_978,In_692,In_830);
xnor U979 (N_979,In_670,In_788);
or U980 (N_980,In_764,In_458);
nor U981 (N_981,In_763,In_250);
or U982 (N_982,In_237,In_94);
nor U983 (N_983,In_161,In_281);
or U984 (N_984,In_672,In_984);
or U985 (N_985,In_874,In_112);
or U986 (N_986,In_486,In_75);
xnor U987 (N_987,In_936,In_835);
or U988 (N_988,In_340,In_295);
nand U989 (N_989,In_440,In_369);
nand U990 (N_990,In_169,In_746);
nand U991 (N_991,In_832,In_411);
nor U992 (N_992,In_16,In_872);
or U993 (N_993,In_93,In_621);
nor U994 (N_994,In_474,In_281);
or U995 (N_995,In_63,In_156);
nand U996 (N_996,In_239,In_267);
and U997 (N_997,In_621,In_735);
nand U998 (N_998,In_152,In_957);
xor U999 (N_999,In_593,In_358);
xor U1000 (N_1000,In_926,In_255);
or U1001 (N_1001,In_310,In_913);
nor U1002 (N_1002,In_618,In_909);
xor U1003 (N_1003,In_863,In_73);
or U1004 (N_1004,In_737,In_412);
xor U1005 (N_1005,In_632,In_189);
or U1006 (N_1006,In_381,In_245);
or U1007 (N_1007,In_481,In_424);
nand U1008 (N_1008,In_233,In_600);
xor U1009 (N_1009,In_599,In_225);
nand U1010 (N_1010,In_279,In_716);
and U1011 (N_1011,In_734,In_345);
nor U1012 (N_1012,In_922,In_673);
nor U1013 (N_1013,In_434,In_863);
xor U1014 (N_1014,In_521,In_886);
nand U1015 (N_1015,In_582,In_311);
and U1016 (N_1016,In_773,In_393);
nand U1017 (N_1017,In_924,In_326);
or U1018 (N_1018,In_362,In_617);
and U1019 (N_1019,In_225,In_416);
nand U1020 (N_1020,In_1,In_43);
or U1021 (N_1021,In_529,In_389);
or U1022 (N_1022,In_386,In_387);
xor U1023 (N_1023,In_541,In_333);
and U1024 (N_1024,In_964,In_167);
nor U1025 (N_1025,In_362,In_698);
or U1026 (N_1026,In_814,In_595);
nor U1027 (N_1027,In_156,In_501);
xor U1028 (N_1028,In_316,In_951);
nor U1029 (N_1029,In_185,In_907);
or U1030 (N_1030,In_90,In_887);
or U1031 (N_1031,In_448,In_263);
and U1032 (N_1032,In_378,In_108);
or U1033 (N_1033,In_329,In_914);
xor U1034 (N_1034,In_122,In_411);
nand U1035 (N_1035,In_628,In_227);
and U1036 (N_1036,In_440,In_971);
nor U1037 (N_1037,In_620,In_909);
nand U1038 (N_1038,In_621,In_813);
xnor U1039 (N_1039,In_850,In_291);
xor U1040 (N_1040,In_263,In_52);
or U1041 (N_1041,In_324,In_718);
or U1042 (N_1042,In_41,In_457);
or U1043 (N_1043,In_637,In_187);
and U1044 (N_1044,In_604,In_246);
xnor U1045 (N_1045,In_570,In_295);
and U1046 (N_1046,In_511,In_811);
nor U1047 (N_1047,In_662,In_246);
nand U1048 (N_1048,In_44,In_861);
nor U1049 (N_1049,In_705,In_445);
nand U1050 (N_1050,In_708,In_971);
nand U1051 (N_1051,In_503,In_382);
and U1052 (N_1052,In_555,In_301);
xor U1053 (N_1053,In_814,In_69);
or U1054 (N_1054,In_518,In_375);
nand U1055 (N_1055,In_49,In_251);
or U1056 (N_1056,In_258,In_880);
and U1057 (N_1057,In_384,In_279);
and U1058 (N_1058,In_601,In_479);
and U1059 (N_1059,In_48,In_441);
or U1060 (N_1060,In_400,In_282);
nand U1061 (N_1061,In_316,In_771);
or U1062 (N_1062,In_685,In_234);
and U1063 (N_1063,In_221,In_613);
or U1064 (N_1064,In_17,In_179);
or U1065 (N_1065,In_840,In_888);
or U1066 (N_1066,In_406,In_533);
and U1067 (N_1067,In_109,In_634);
nor U1068 (N_1068,In_498,In_986);
nand U1069 (N_1069,In_896,In_5);
and U1070 (N_1070,In_664,In_914);
xor U1071 (N_1071,In_742,In_118);
nor U1072 (N_1072,In_502,In_223);
nor U1073 (N_1073,In_490,In_176);
nand U1074 (N_1074,In_319,In_243);
nor U1075 (N_1075,In_23,In_135);
nor U1076 (N_1076,In_535,In_941);
nand U1077 (N_1077,In_368,In_903);
or U1078 (N_1078,In_546,In_854);
and U1079 (N_1079,In_816,In_365);
nand U1080 (N_1080,In_957,In_452);
xor U1081 (N_1081,In_939,In_148);
xnor U1082 (N_1082,In_221,In_511);
nor U1083 (N_1083,In_5,In_222);
nand U1084 (N_1084,In_166,In_811);
nor U1085 (N_1085,In_436,In_879);
or U1086 (N_1086,In_324,In_66);
nor U1087 (N_1087,In_833,In_123);
xor U1088 (N_1088,In_799,In_121);
and U1089 (N_1089,In_339,In_275);
nor U1090 (N_1090,In_692,In_383);
or U1091 (N_1091,In_418,In_659);
nor U1092 (N_1092,In_294,In_197);
xor U1093 (N_1093,In_676,In_235);
nor U1094 (N_1094,In_275,In_260);
or U1095 (N_1095,In_371,In_499);
nor U1096 (N_1096,In_287,In_403);
or U1097 (N_1097,In_4,In_122);
or U1098 (N_1098,In_700,In_729);
nand U1099 (N_1099,In_829,In_24);
nand U1100 (N_1100,In_334,In_7);
and U1101 (N_1101,In_391,In_764);
xor U1102 (N_1102,In_352,In_559);
and U1103 (N_1103,In_522,In_88);
xnor U1104 (N_1104,In_689,In_161);
nand U1105 (N_1105,In_234,In_466);
or U1106 (N_1106,In_223,In_838);
nand U1107 (N_1107,In_825,In_351);
xnor U1108 (N_1108,In_227,In_226);
xnor U1109 (N_1109,In_832,In_781);
or U1110 (N_1110,In_521,In_753);
nand U1111 (N_1111,In_877,In_339);
or U1112 (N_1112,In_822,In_979);
nor U1113 (N_1113,In_781,In_352);
nand U1114 (N_1114,In_13,In_457);
and U1115 (N_1115,In_506,In_59);
nor U1116 (N_1116,In_19,In_127);
nand U1117 (N_1117,In_220,In_153);
nand U1118 (N_1118,In_169,In_938);
or U1119 (N_1119,In_585,In_393);
nor U1120 (N_1120,In_470,In_785);
nand U1121 (N_1121,In_413,In_544);
nor U1122 (N_1122,In_392,In_48);
nor U1123 (N_1123,In_571,In_864);
or U1124 (N_1124,In_330,In_862);
xnor U1125 (N_1125,In_191,In_208);
and U1126 (N_1126,In_800,In_370);
xnor U1127 (N_1127,In_7,In_709);
nand U1128 (N_1128,In_973,In_211);
nor U1129 (N_1129,In_19,In_878);
nor U1130 (N_1130,In_671,In_775);
and U1131 (N_1131,In_983,In_772);
nand U1132 (N_1132,In_229,In_581);
and U1133 (N_1133,In_330,In_522);
and U1134 (N_1134,In_865,In_197);
or U1135 (N_1135,In_91,In_92);
xor U1136 (N_1136,In_522,In_555);
nand U1137 (N_1137,In_711,In_58);
or U1138 (N_1138,In_592,In_443);
nand U1139 (N_1139,In_131,In_395);
or U1140 (N_1140,In_240,In_310);
or U1141 (N_1141,In_675,In_498);
nand U1142 (N_1142,In_860,In_95);
nor U1143 (N_1143,In_975,In_619);
nor U1144 (N_1144,In_170,In_932);
nand U1145 (N_1145,In_70,In_639);
nor U1146 (N_1146,In_679,In_305);
nor U1147 (N_1147,In_293,In_110);
and U1148 (N_1148,In_386,In_725);
nor U1149 (N_1149,In_667,In_503);
nand U1150 (N_1150,In_354,In_146);
or U1151 (N_1151,In_644,In_702);
nor U1152 (N_1152,In_905,In_599);
xnor U1153 (N_1153,In_56,In_135);
xnor U1154 (N_1154,In_522,In_93);
or U1155 (N_1155,In_244,In_442);
or U1156 (N_1156,In_324,In_925);
nand U1157 (N_1157,In_141,In_654);
and U1158 (N_1158,In_949,In_400);
nor U1159 (N_1159,In_263,In_679);
nor U1160 (N_1160,In_200,In_704);
nand U1161 (N_1161,In_542,In_701);
or U1162 (N_1162,In_857,In_897);
or U1163 (N_1163,In_607,In_281);
xor U1164 (N_1164,In_369,In_906);
and U1165 (N_1165,In_494,In_419);
xor U1166 (N_1166,In_594,In_617);
xnor U1167 (N_1167,In_925,In_962);
xnor U1168 (N_1168,In_73,In_787);
nand U1169 (N_1169,In_977,In_882);
or U1170 (N_1170,In_597,In_868);
xor U1171 (N_1171,In_407,In_982);
and U1172 (N_1172,In_497,In_3);
or U1173 (N_1173,In_275,In_782);
xnor U1174 (N_1174,In_446,In_932);
nor U1175 (N_1175,In_738,In_930);
xnor U1176 (N_1176,In_610,In_977);
and U1177 (N_1177,In_305,In_835);
nor U1178 (N_1178,In_375,In_141);
xor U1179 (N_1179,In_819,In_711);
or U1180 (N_1180,In_468,In_501);
or U1181 (N_1181,In_873,In_933);
nand U1182 (N_1182,In_403,In_123);
and U1183 (N_1183,In_164,In_904);
or U1184 (N_1184,In_44,In_0);
nand U1185 (N_1185,In_44,In_315);
xor U1186 (N_1186,In_411,In_413);
xor U1187 (N_1187,In_23,In_930);
and U1188 (N_1188,In_203,In_461);
xnor U1189 (N_1189,In_455,In_474);
or U1190 (N_1190,In_910,In_921);
nor U1191 (N_1191,In_441,In_288);
or U1192 (N_1192,In_20,In_53);
and U1193 (N_1193,In_679,In_884);
xnor U1194 (N_1194,In_939,In_290);
and U1195 (N_1195,In_519,In_466);
and U1196 (N_1196,In_24,In_846);
xor U1197 (N_1197,In_107,In_476);
xnor U1198 (N_1198,In_208,In_852);
nor U1199 (N_1199,In_772,In_266);
nor U1200 (N_1200,In_312,In_328);
or U1201 (N_1201,In_328,In_613);
xnor U1202 (N_1202,In_924,In_894);
nor U1203 (N_1203,In_80,In_508);
nand U1204 (N_1204,In_779,In_949);
and U1205 (N_1205,In_688,In_610);
or U1206 (N_1206,In_17,In_477);
xnor U1207 (N_1207,In_752,In_517);
nand U1208 (N_1208,In_802,In_997);
nand U1209 (N_1209,In_744,In_863);
xnor U1210 (N_1210,In_650,In_222);
nand U1211 (N_1211,In_748,In_624);
xnor U1212 (N_1212,In_189,In_764);
nand U1213 (N_1213,In_772,In_556);
or U1214 (N_1214,In_61,In_711);
and U1215 (N_1215,In_884,In_109);
xnor U1216 (N_1216,In_555,In_154);
or U1217 (N_1217,In_388,In_356);
nor U1218 (N_1218,In_586,In_288);
and U1219 (N_1219,In_168,In_230);
and U1220 (N_1220,In_260,In_583);
nor U1221 (N_1221,In_448,In_929);
nand U1222 (N_1222,In_585,In_922);
or U1223 (N_1223,In_840,In_190);
nor U1224 (N_1224,In_774,In_537);
nand U1225 (N_1225,In_907,In_850);
xor U1226 (N_1226,In_126,In_333);
xor U1227 (N_1227,In_959,In_978);
xnor U1228 (N_1228,In_487,In_629);
nand U1229 (N_1229,In_472,In_13);
xnor U1230 (N_1230,In_57,In_413);
nand U1231 (N_1231,In_495,In_900);
nor U1232 (N_1232,In_128,In_392);
nand U1233 (N_1233,In_320,In_175);
and U1234 (N_1234,In_60,In_654);
nand U1235 (N_1235,In_584,In_810);
nor U1236 (N_1236,In_682,In_642);
xnor U1237 (N_1237,In_799,In_715);
and U1238 (N_1238,In_868,In_255);
nor U1239 (N_1239,In_679,In_398);
and U1240 (N_1240,In_316,In_923);
or U1241 (N_1241,In_172,In_495);
nor U1242 (N_1242,In_71,In_579);
and U1243 (N_1243,In_456,In_719);
and U1244 (N_1244,In_72,In_540);
nor U1245 (N_1245,In_20,In_31);
and U1246 (N_1246,In_578,In_784);
nor U1247 (N_1247,In_159,In_655);
or U1248 (N_1248,In_890,In_649);
nor U1249 (N_1249,In_824,In_108);
xnor U1250 (N_1250,In_284,In_519);
and U1251 (N_1251,In_241,In_217);
xor U1252 (N_1252,In_784,In_430);
xor U1253 (N_1253,In_373,In_35);
xor U1254 (N_1254,In_585,In_419);
and U1255 (N_1255,In_209,In_974);
and U1256 (N_1256,In_679,In_616);
or U1257 (N_1257,In_705,In_187);
xor U1258 (N_1258,In_928,In_67);
nor U1259 (N_1259,In_565,In_480);
nand U1260 (N_1260,In_270,In_889);
xnor U1261 (N_1261,In_803,In_454);
nand U1262 (N_1262,In_772,In_192);
or U1263 (N_1263,In_87,In_872);
nand U1264 (N_1264,In_232,In_789);
nor U1265 (N_1265,In_153,In_21);
or U1266 (N_1266,In_200,In_455);
nor U1267 (N_1267,In_792,In_28);
and U1268 (N_1268,In_141,In_358);
xor U1269 (N_1269,In_39,In_655);
nor U1270 (N_1270,In_525,In_669);
or U1271 (N_1271,In_782,In_710);
nand U1272 (N_1272,In_992,In_364);
xnor U1273 (N_1273,In_664,In_395);
nor U1274 (N_1274,In_362,In_472);
or U1275 (N_1275,In_600,In_154);
nand U1276 (N_1276,In_486,In_379);
or U1277 (N_1277,In_919,In_298);
and U1278 (N_1278,In_520,In_67);
or U1279 (N_1279,In_345,In_597);
and U1280 (N_1280,In_622,In_868);
nand U1281 (N_1281,In_89,In_859);
nand U1282 (N_1282,In_349,In_155);
xnor U1283 (N_1283,In_468,In_936);
or U1284 (N_1284,In_6,In_209);
and U1285 (N_1285,In_571,In_478);
nand U1286 (N_1286,In_252,In_224);
xnor U1287 (N_1287,In_685,In_871);
nand U1288 (N_1288,In_3,In_825);
xor U1289 (N_1289,In_149,In_950);
nand U1290 (N_1290,In_895,In_291);
nor U1291 (N_1291,In_825,In_926);
xor U1292 (N_1292,In_997,In_319);
xor U1293 (N_1293,In_160,In_134);
and U1294 (N_1294,In_719,In_19);
xnor U1295 (N_1295,In_933,In_174);
nor U1296 (N_1296,In_118,In_130);
or U1297 (N_1297,In_936,In_482);
and U1298 (N_1298,In_460,In_51);
or U1299 (N_1299,In_584,In_165);
or U1300 (N_1300,In_172,In_33);
nand U1301 (N_1301,In_968,In_822);
and U1302 (N_1302,In_548,In_502);
nor U1303 (N_1303,In_174,In_861);
and U1304 (N_1304,In_240,In_640);
nor U1305 (N_1305,In_198,In_428);
xor U1306 (N_1306,In_19,In_925);
xor U1307 (N_1307,In_355,In_50);
or U1308 (N_1308,In_883,In_29);
nand U1309 (N_1309,In_361,In_557);
xor U1310 (N_1310,In_80,In_193);
or U1311 (N_1311,In_986,In_72);
and U1312 (N_1312,In_496,In_908);
nand U1313 (N_1313,In_466,In_82);
nor U1314 (N_1314,In_705,In_661);
and U1315 (N_1315,In_371,In_676);
nand U1316 (N_1316,In_646,In_306);
nand U1317 (N_1317,In_698,In_674);
xnor U1318 (N_1318,In_936,In_610);
nand U1319 (N_1319,In_537,In_702);
or U1320 (N_1320,In_686,In_771);
nand U1321 (N_1321,In_538,In_10);
and U1322 (N_1322,In_202,In_742);
nor U1323 (N_1323,In_537,In_403);
xor U1324 (N_1324,In_401,In_745);
xnor U1325 (N_1325,In_493,In_463);
or U1326 (N_1326,In_434,In_405);
nor U1327 (N_1327,In_42,In_125);
nor U1328 (N_1328,In_75,In_701);
xor U1329 (N_1329,In_557,In_756);
nand U1330 (N_1330,In_141,In_229);
nand U1331 (N_1331,In_343,In_366);
nor U1332 (N_1332,In_945,In_668);
and U1333 (N_1333,In_331,In_957);
nor U1334 (N_1334,In_877,In_875);
xnor U1335 (N_1335,In_260,In_575);
or U1336 (N_1336,In_680,In_254);
or U1337 (N_1337,In_538,In_580);
or U1338 (N_1338,In_528,In_214);
nor U1339 (N_1339,In_933,In_134);
or U1340 (N_1340,In_51,In_679);
and U1341 (N_1341,In_760,In_544);
or U1342 (N_1342,In_254,In_317);
and U1343 (N_1343,In_261,In_366);
nand U1344 (N_1344,In_648,In_880);
or U1345 (N_1345,In_102,In_385);
nand U1346 (N_1346,In_343,In_625);
nor U1347 (N_1347,In_256,In_48);
xnor U1348 (N_1348,In_933,In_478);
and U1349 (N_1349,In_610,In_793);
xor U1350 (N_1350,In_643,In_621);
nand U1351 (N_1351,In_974,In_255);
and U1352 (N_1352,In_897,In_894);
or U1353 (N_1353,In_327,In_275);
xnor U1354 (N_1354,In_232,In_282);
or U1355 (N_1355,In_595,In_17);
or U1356 (N_1356,In_703,In_322);
or U1357 (N_1357,In_28,In_382);
xnor U1358 (N_1358,In_546,In_971);
or U1359 (N_1359,In_336,In_419);
nand U1360 (N_1360,In_337,In_888);
xor U1361 (N_1361,In_485,In_7);
or U1362 (N_1362,In_221,In_89);
nor U1363 (N_1363,In_81,In_920);
and U1364 (N_1364,In_295,In_159);
nor U1365 (N_1365,In_909,In_627);
nor U1366 (N_1366,In_618,In_326);
xnor U1367 (N_1367,In_413,In_343);
and U1368 (N_1368,In_617,In_627);
nand U1369 (N_1369,In_319,In_921);
nor U1370 (N_1370,In_772,In_873);
and U1371 (N_1371,In_49,In_284);
nor U1372 (N_1372,In_24,In_116);
nor U1373 (N_1373,In_759,In_233);
xor U1374 (N_1374,In_857,In_902);
nand U1375 (N_1375,In_943,In_316);
xor U1376 (N_1376,In_212,In_163);
nand U1377 (N_1377,In_556,In_449);
or U1378 (N_1378,In_871,In_631);
nand U1379 (N_1379,In_958,In_622);
and U1380 (N_1380,In_927,In_946);
or U1381 (N_1381,In_614,In_630);
xor U1382 (N_1382,In_692,In_16);
or U1383 (N_1383,In_888,In_270);
nor U1384 (N_1384,In_348,In_40);
nor U1385 (N_1385,In_670,In_952);
and U1386 (N_1386,In_232,In_964);
or U1387 (N_1387,In_933,In_997);
and U1388 (N_1388,In_519,In_319);
xnor U1389 (N_1389,In_22,In_875);
nand U1390 (N_1390,In_33,In_404);
or U1391 (N_1391,In_496,In_838);
and U1392 (N_1392,In_35,In_166);
nand U1393 (N_1393,In_491,In_730);
nand U1394 (N_1394,In_139,In_602);
or U1395 (N_1395,In_611,In_621);
or U1396 (N_1396,In_83,In_785);
and U1397 (N_1397,In_343,In_870);
or U1398 (N_1398,In_345,In_526);
nand U1399 (N_1399,In_655,In_827);
nand U1400 (N_1400,In_539,In_320);
and U1401 (N_1401,In_386,In_521);
xor U1402 (N_1402,In_234,In_862);
nand U1403 (N_1403,In_355,In_322);
nor U1404 (N_1404,In_159,In_247);
and U1405 (N_1405,In_26,In_25);
nand U1406 (N_1406,In_596,In_59);
or U1407 (N_1407,In_631,In_386);
xnor U1408 (N_1408,In_96,In_922);
and U1409 (N_1409,In_769,In_339);
nor U1410 (N_1410,In_947,In_392);
or U1411 (N_1411,In_920,In_379);
nand U1412 (N_1412,In_609,In_478);
nand U1413 (N_1413,In_569,In_99);
and U1414 (N_1414,In_511,In_637);
or U1415 (N_1415,In_629,In_985);
or U1416 (N_1416,In_665,In_946);
nand U1417 (N_1417,In_419,In_724);
and U1418 (N_1418,In_659,In_30);
and U1419 (N_1419,In_536,In_560);
and U1420 (N_1420,In_282,In_3);
xor U1421 (N_1421,In_706,In_210);
or U1422 (N_1422,In_532,In_848);
xor U1423 (N_1423,In_561,In_176);
xor U1424 (N_1424,In_585,In_662);
or U1425 (N_1425,In_601,In_362);
nand U1426 (N_1426,In_198,In_330);
or U1427 (N_1427,In_282,In_186);
xnor U1428 (N_1428,In_25,In_894);
nor U1429 (N_1429,In_725,In_646);
nor U1430 (N_1430,In_855,In_496);
and U1431 (N_1431,In_737,In_839);
or U1432 (N_1432,In_307,In_878);
nand U1433 (N_1433,In_655,In_286);
nor U1434 (N_1434,In_288,In_40);
or U1435 (N_1435,In_818,In_102);
nor U1436 (N_1436,In_808,In_311);
or U1437 (N_1437,In_337,In_386);
xnor U1438 (N_1438,In_275,In_278);
or U1439 (N_1439,In_299,In_641);
nor U1440 (N_1440,In_191,In_224);
nor U1441 (N_1441,In_604,In_461);
nor U1442 (N_1442,In_344,In_89);
and U1443 (N_1443,In_16,In_770);
and U1444 (N_1444,In_604,In_376);
nor U1445 (N_1445,In_939,In_546);
xor U1446 (N_1446,In_673,In_62);
xnor U1447 (N_1447,In_824,In_755);
or U1448 (N_1448,In_630,In_821);
nor U1449 (N_1449,In_151,In_140);
nor U1450 (N_1450,In_340,In_841);
or U1451 (N_1451,In_525,In_9);
and U1452 (N_1452,In_42,In_247);
or U1453 (N_1453,In_821,In_950);
xor U1454 (N_1454,In_108,In_266);
nand U1455 (N_1455,In_398,In_252);
nand U1456 (N_1456,In_661,In_485);
nand U1457 (N_1457,In_333,In_553);
and U1458 (N_1458,In_885,In_628);
xnor U1459 (N_1459,In_601,In_179);
nor U1460 (N_1460,In_697,In_84);
nor U1461 (N_1461,In_58,In_985);
xor U1462 (N_1462,In_72,In_450);
nor U1463 (N_1463,In_157,In_695);
nand U1464 (N_1464,In_519,In_412);
and U1465 (N_1465,In_624,In_93);
or U1466 (N_1466,In_200,In_319);
and U1467 (N_1467,In_777,In_313);
xnor U1468 (N_1468,In_665,In_404);
nand U1469 (N_1469,In_589,In_685);
nor U1470 (N_1470,In_126,In_712);
and U1471 (N_1471,In_512,In_57);
nor U1472 (N_1472,In_539,In_461);
nand U1473 (N_1473,In_442,In_986);
or U1474 (N_1474,In_547,In_531);
or U1475 (N_1475,In_85,In_157);
or U1476 (N_1476,In_334,In_418);
xnor U1477 (N_1477,In_487,In_13);
nand U1478 (N_1478,In_992,In_994);
or U1479 (N_1479,In_2,In_220);
and U1480 (N_1480,In_961,In_315);
nand U1481 (N_1481,In_5,In_979);
xor U1482 (N_1482,In_131,In_229);
xnor U1483 (N_1483,In_802,In_29);
nor U1484 (N_1484,In_790,In_281);
xor U1485 (N_1485,In_876,In_736);
xor U1486 (N_1486,In_745,In_583);
xor U1487 (N_1487,In_701,In_896);
or U1488 (N_1488,In_412,In_8);
and U1489 (N_1489,In_640,In_692);
and U1490 (N_1490,In_899,In_779);
nand U1491 (N_1491,In_725,In_336);
or U1492 (N_1492,In_883,In_446);
and U1493 (N_1493,In_588,In_950);
xnor U1494 (N_1494,In_42,In_649);
and U1495 (N_1495,In_26,In_744);
nand U1496 (N_1496,In_269,In_319);
and U1497 (N_1497,In_842,In_449);
xnor U1498 (N_1498,In_454,In_328);
xor U1499 (N_1499,In_35,In_913);
or U1500 (N_1500,In_883,In_244);
nand U1501 (N_1501,In_135,In_62);
nand U1502 (N_1502,In_947,In_628);
xor U1503 (N_1503,In_812,In_846);
and U1504 (N_1504,In_132,In_988);
nor U1505 (N_1505,In_564,In_335);
nand U1506 (N_1506,In_989,In_563);
nand U1507 (N_1507,In_776,In_790);
and U1508 (N_1508,In_617,In_79);
nand U1509 (N_1509,In_823,In_714);
xnor U1510 (N_1510,In_306,In_437);
xnor U1511 (N_1511,In_508,In_35);
or U1512 (N_1512,In_582,In_486);
xor U1513 (N_1513,In_395,In_858);
and U1514 (N_1514,In_466,In_795);
nand U1515 (N_1515,In_787,In_288);
and U1516 (N_1516,In_993,In_321);
nand U1517 (N_1517,In_472,In_742);
and U1518 (N_1518,In_885,In_679);
and U1519 (N_1519,In_952,In_696);
nand U1520 (N_1520,In_75,In_8);
nand U1521 (N_1521,In_535,In_53);
nor U1522 (N_1522,In_44,In_155);
xor U1523 (N_1523,In_816,In_274);
nor U1524 (N_1524,In_157,In_949);
nand U1525 (N_1525,In_71,In_900);
and U1526 (N_1526,In_265,In_205);
and U1527 (N_1527,In_848,In_33);
nand U1528 (N_1528,In_943,In_726);
nor U1529 (N_1529,In_908,In_499);
and U1530 (N_1530,In_663,In_470);
nor U1531 (N_1531,In_257,In_819);
or U1532 (N_1532,In_814,In_373);
or U1533 (N_1533,In_344,In_973);
xnor U1534 (N_1534,In_852,In_199);
nand U1535 (N_1535,In_682,In_572);
xor U1536 (N_1536,In_219,In_733);
or U1537 (N_1537,In_796,In_707);
xor U1538 (N_1538,In_970,In_52);
xor U1539 (N_1539,In_64,In_325);
or U1540 (N_1540,In_87,In_566);
nand U1541 (N_1541,In_895,In_64);
or U1542 (N_1542,In_682,In_472);
or U1543 (N_1543,In_314,In_100);
or U1544 (N_1544,In_940,In_16);
and U1545 (N_1545,In_156,In_408);
xor U1546 (N_1546,In_479,In_984);
xor U1547 (N_1547,In_628,In_267);
or U1548 (N_1548,In_892,In_302);
nand U1549 (N_1549,In_886,In_649);
xnor U1550 (N_1550,In_304,In_93);
and U1551 (N_1551,In_523,In_341);
nor U1552 (N_1552,In_560,In_878);
xnor U1553 (N_1553,In_815,In_505);
nor U1554 (N_1554,In_452,In_773);
nand U1555 (N_1555,In_264,In_126);
nand U1556 (N_1556,In_164,In_839);
nor U1557 (N_1557,In_852,In_469);
and U1558 (N_1558,In_905,In_158);
or U1559 (N_1559,In_885,In_962);
and U1560 (N_1560,In_977,In_8);
xor U1561 (N_1561,In_354,In_52);
nand U1562 (N_1562,In_885,In_751);
nand U1563 (N_1563,In_964,In_316);
and U1564 (N_1564,In_3,In_314);
nor U1565 (N_1565,In_469,In_139);
nor U1566 (N_1566,In_0,In_482);
xor U1567 (N_1567,In_200,In_262);
xnor U1568 (N_1568,In_477,In_656);
xor U1569 (N_1569,In_468,In_199);
or U1570 (N_1570,In_923,In_68);
and U1571 (N_1571,In_37,In_825);
xnor U1572 (N_1572,In_553,In_810);
or U1573 (N_1573,In_593,In_10);
xnor U1574 (N_1574,In_181,In_225);
or U1575 (N_1575,In_276,In_777);
and U1576 (N_1576,In_216,In_170);
or U1577 (N_1577,In_502,In_501);
or U1578 (N_1578,In_453,In_948);
and U1579 (N_1579,In_677,In_582);
or U1580 (N_1580,In_478,In_286);
or U1581 (N_1581,In_92,In_556);
nand U1582 (N_1582,In_904,In_609);
and U1583 (N_1583,In_747,In_911);
nand U1584 (N_1584,In_562,In_843);
nand U1585 (N_1585,In_534,In_85);
nand U1586 (N_1586,In_835,In_946);
and U1587 (N_1587,In_190,In_451);
nand U1588 (N_1588,In_484,In_553);
xor U1589 (N_1589,In_869,In_640);
nor U1590 (N_1590,In_282,In_204);
xnor U1591 (N_1591,In_866,In_125);
nand U1592 (N_1592,In_9,In_238);
nor U1593 (N_1593,In_755,In_276);
and U1594 (N_1594,In_512,In_422);
nand U1595 (N_1595,In_349,In_579);
nand U1596 (N_1596,In_241,In_188);
or U1597 (N_1597,In_853,In_360);
and U1598 (N_1598,In_73,In_169);
xnor U1599 (N_1599,In_350,In_419);
nor U1600 (N_1600,In_605,In_165);
xnor U1601 (N_1601,In_69,In_396);
xor U1602 (N_1602,In_412,In_912);
and U1603 (N_1603,In_339,In_809);
nor U1604 (N_1604,In_137,In_888);
xnor U1605 (N_1605,In_322,In_379);
nand U1606 (N_1606,In_810,In_139);
xor U1607 (N_1607,In_973,In_408);
and U1608 (N_1608,In_686,In_110);
nor U1609 (N_1609,In_851,In_411);
and U1610 (N_1610,In_651,In_389);
and U1611 (N_1611,In_576,In_105);
and U1612 (N_1612,In_100,In_991);
xnor U1613 (N_1613,In_146,In_121);
nand U1614 (N_1614,In_477,In_950);
nand U1615 (N_1615,In_989,In_524);
and U1616 (N_1616,In_679,In_918);
xnor U1617 (N_1617,In_439,In_358);
xor U1618 (N_1618,In_391,In_976);
and U1619 (N_1619,In_144,In_136);
xor U1620 (N_1620,In_814,In_974);
nor U1621 (N_1621,In_613,In_472);
and U1622 (N_1622,In_491,In_329);
nor U1623 (N_1623,In_281,In_47);
and U1624 (N_1624,In_828,In_376);
or U1625 (N_1625,In_208,In_939);
or U1626 (N_1626,In_266,In_761);
nand U1627 (N_1627,In_724,In_130);
nand U1628 (N_1628,In_757,In_526);
xor U1629 (N_1629,In_35,In_132);
and U1630 (N_1630,In_696,In_341);
nor U1631 (N_1631,In_291,In_607);
xnor U1632 (N_1632,In_353,In_638);
nand U1633 (N_1633,In_754,In_500);
and U1634 (N_1634,In_756,In_672);
and U1635 (N_1635,In_183,In_264);
or U1636 (N_1636,In_711,In_847);
xor U1637 (N_1637,In_887,In_168);
xnor U1638 (N_1638,In_224,In_202);
nand U1639 (N_1639,In_164,In_479);
or U1640 (N_1640,In_849,In_885);
or U1641 (N_1641,In_856,In_59);
and U1642 (N_1642,In_992,In_588);
nand U1643 (N_1643,In_149,In_917);
or U1644 (N_1644,In_805,In_727);
xnor U1645 (N_1645,In_269,In_205);
nor U1646 (N_1646,In_410,In_8);
xnor U1647 (N_1647,In_530,In_79);
or U1648 (N_1648,In_760,In_739);
or U1649 (N_1649,In_305,In_726);
nand U1650 (N_1650,In_446,In_247);
or U1651 (N_1651,In_127,In_871);
nor U1652 (N_1652,In_627,In_514);
and U1653 (N_1653,In_323,In_72);
and U1654 (N_1654,In_526,In_669);
xor U1655 (N_1655,In_36,In_562);
xnor U1656 (N_1656,In_196,In_9);
nor U1657 (N_1657,In_524,In_370);
and U1658 (N_1658,In_655,In_673);
nand U1659 (N_1659,In_231,In_194);
nor U1660 (N_1660,In_831,In_156);
or U1661 (N_1661,In_990,In_878);
and U1662 (N_1662,In_930,In_237);
or U1663 (N_1663,In_819,In_363);
nand U1664 (N_1664,In_232,In_775);
nand U1665 (N_1665,In_456,In_782);
nor U1666 (N_1666,In_741,In_150);
and U1667 (N_1667,In_523,In_383);
and U1668 (N_1668,In_477,In_748);
nand U1669 (N_1669,In_303,In_60);
and U1670 (N_1670,In_833,In_581);
nand U1671 (N_1671,In_969,In_933);
nand U1672 (N_1672,In_689,In_780);
or U1673 (N_1673,In_762,In_440);
xor U1674 (N_1674,In_48,In_132);
nand U1675 (N_1675,In_96,In_155);
or U1676 (N_1676,In_602,In_815);
or U1677 (N_1677,In_876,In_734);
nand U1678 (N_1678,In_976,In_185);
xnor U1679 (N_1679,In_718,In_838);
or U1680 (N_1680,In_58,In_3);
or U1681 (N_1681,In_157,In_206);
and U1682 (N_1682,In_242,In_738);
nor U1683 (N_1683,In_138,In_496);
and U1684 (N_1684,In_336,In_715);
xor U1685 (N_1685,In_357,In_738);
or U1686 (N_1686,In_752,In_187);
nor U1687 (N_1687,In_531,In_339);
and U1688 (N_1688,In_942,In_57);
and U1689 (N_1689,In_27,In_864);
xor U1690 (N_1690,In_521,In_472);
xnor U1691 (N_1691,In_67,In_624);
and U1692 (N_1692,In_661,In_242);
nand U1693 (N_1693,In_290,In_573);
nand U1694 (N_1694,In_276,In_875);
and U1695 (N_1695,In_558,In_160);
nand U1696 (N_1696,In_190,In_184);
nand U1697 (N_1697,In_155,In_838);
or U1698 (N_1698,In_142,In_897);
nor U1699 (N_1699,In_52,In_919);
xor U1700 (N_1700,In_861,In_301);
nor U1701 (N_1701,In_803,In_891);
nand U1702 (N_1702,In_681,In_319);
and U1703 (N_1703,In_678,In_643);
or U1704 (N_1704,In_968,In_442);
nor U1705 (N_1705,In_341,In_120);
or U1706 (N_1706,In_810,In_970);
and U1707 (N_1707,In_108,In_445);
nor U1708 (N_1708,In_238,In_336);
nor U1709 (N_1709,In_538,In_859);
and U1710 (N_1710,In_467,In_324);
and U1711 (N_1711,In_595,In_764);
xor U1712 (N_1712,In_258,In_219);
and U1713 (N_1713,In_516,In_301);
or U1714 (N_1714,In_739,In_239);
nor U1715 (N_1715,In_721,In_404);
nand U1716 (N_1716,In_603,In_278);
and U1717 (N_1717,In_578,In_695);
and U1718 (N_1718,In_806,In_255);
nor U1719 (N_1719,In_695,In_110);
or U1720 (N_1720,In_339,In_759);
and U1721 (N_1721,In_710,In_270);
and U1722 (N_1722,In_216,In_854);
or U1723 (N_1723,In_710,In_622);
xor U1724 (N_1724,In_782,In_114);
xor U1725 (N_1725,In_852,In_957);
nor U1726 (N_1726,In_638,In_531);
and U1727 (N_1727,In_301,In_155);
nand U1728 (N_1728,In_862,In_716);
nor U1729 (N_1729,In_730,In_973);
nor U1730 (N_1730,In_879,In_339);
and U1731 (N_1731,In_880,In_388);
nor U1732 (N_1732,In_775,In_719);
xnor U1733 (N_1733,In_40,In_677);
xor U1734 (N_1734,In_155,In_716);
or U1735 (N_1735,In_189,In_505);
xnor U1736 (N_1736,In_496,In_489);
xnor U1737 (N_1737,In_986,In_953);
or U1738 (N_1738,In_246,In_500);
nand U1739 (N_1739,In_874,In_829);
xor U1740 (N_1740,In_692,In_505);
or U1741 (N_1741,In_885,In_371);
nor U1742 (N_1742,In_119,In_610);
xor U1743 (N_1743,In_653,In_281);
nor U1744 (N_1744,In_463,In_426);
nor U1745 (N_1745,In_291,In_717);
nand U1746 (N_1746,In_525,In_998);
and U1747 (N_1747,In_736,In_521);
or U1748 (N_1748,In_973,In_909);
or U1749 (N_1749,In_514,In_403);
xnor U1750 (N_1750,In_940,In_972);
nand U1751 (N_1751,In_702,In_708);
or U1752 (N_1752,In_543,In_860);
xnor U1753 (N_1753,In_944,In_527);
xor U1754 (N_1754,In_655,In_415);
nand U1755 (N_1755,In_324,In_927);
xor U1756 (N_1756,In_778,In_428);
xor U1757 (N_1757,In_521,In_238);
nand U1758 (N_1758,In_370,In_182);
xnor U1759 (N_1759,In_913,In_995);
xnor U1760 (N_1760,In_272,In_771);
and U1761 (N_1761,In_929,In_257);
or U1762 (N_1762,In_416,In_258);
and U1763 (N_1763,In_524,In_215);
and U1764 (N_1764,In_730,In_143);
and U1765 (N_1765,In_951,In_366);
nand U1766 (N_1766,In_553,In_873);
and U1767 (N_1767,In_384,In_64);
and U1768 (N_1768,In_451,In_170);
or U1769 (N_1769,In_263,In_168);
and U1770 (N_1770,In_515,In_290);
xor U1771 (N_1771,In_10,In_508);
nand U1772 (N_1772,In_84,In_530);
nand U1773 (N_1773,In_891,In_763);
and U1774 (N_1774,In_222,In_924);
and U1775 (N_1775,In_817,In_328);
xnor U1776 (N_1776,In_951,In_987);
nand U1777 (N_1777,In_145,In_334);
or U1778 (N_1778,In_837,In_784);
or U1779 (N_1779,In_82,In_123);
nor U1780 (N_1780,In_702,In_977);
or U1781 (N_1781,In_495,In_989);
or U1782 (N_1782,In_609,In_906);
nor U1783 (N_1783,In_927,In_516);
xnor U1784 (N_1784,In_103,In_946);
and U1785 (N_1785,In_407,In_562);
or U1786 (N_1786,In_362,In_441);
nand U1787 (N_1787,In_197,In_706);
nand U1788 (N_1788,In_249,In_752);
nand U1789 (N_1789,In_534,In_591);
xor U1790 (N_1790,In_505,In_805);
nand U1791 (N_1791,In_197,In_54);
or U1792 (N_1792,In_299,In_153);
nand U1793 (N_1793,In_880,In_653);
and U1794 (N_1794,In_545,In_199);
or U1795 (N_1795,In_525,In_650);
xor U1796 (N_1796,In_398,In_218);
xor U1797 (N_1797,In_285,In_717);
nor U1798 (N_1798,In_266,In_100);
nor U1799 (N_1799,In_371,In_443);
or U1800 (N_1800,In_438,In_88);
nand U1801 (N_1801,In_97,In_935);
and U1802 (N_1802,In_21,In_898);
xor U1803 (N_1803,In_23,In_948);
and U1804 (N_1804,In_300,In_520);
nor U1805 (N_1805,In_755,In_778);
or U1806 (N_1806,In_426,In_737);
and U1807 (N_1807,In_475,In_910);
or U1808 (N_1808,In_9,In_306);
nor U1809 (N_1809,In_764,In_707);
nand U1810 (N_1810,In_816,In_708);
nor U1811 (N_1811,In_420,In_226);
or U1812 (N_1812,In_916,In_976);
nor U1813 (N_1813,In_341,In_160);
xor U1814 (N_1814,In_452,In_69);
nor U1815 (N_1815,In_417,In_641);
and U1816 (N_1816,In_836,In_728);
xor U1817 (N_1817,In_359,In_681);
and U1818 (N_1818,In_812,In_153);
nand U1819 (N_1819,In_24,In_748);
nor U1820 (N_1820,In_371,In_515);
nor U1821 (N_1821,In_538,In_575);
nand U1822 (N_1822,In_467,In_506);
and U1823 (N_1823,In_107,In_374);
nor U1824 (N_1824,In_951,In_763);
nor U1825 (N_1825,In_741,In_304);
xor U1826 (N_1826,In_958,In_750);
and U1827 (N_1827,In_70,In_253);
nor U1828 (N_1828,In_941,In_828);
and U1829 (N_1829,In_86,In_655);
xor U1830 (N_1830,In_690,In_54);
and U1831 (N_1831,In_647,In_551);
nor U1832 (N_1832,In_918,In_884);
or U1833 (N_1833,In_671,In_281);
nand U1834 (N_1834,In_86,In_617);
or U1835 (N_1835,In_27,In_792);
nor U1836 (N_1836,In_389,In_299);
nand U1837 (N_1837,In_11,In_150);
xnor U1838 (N_1838,In_626,In_476);
and U1839 (N_1839,In_550,In_245);
and U1840 (N_1840,In_744,In_543);
or U1841 (N_1841,In_461,In_99);
nand U1842 (N_1842,In_232,In_107);
or U1843 (N_1843,In_289,In_76);
and U1844 (N_1844,In_847,In_121);
or U1845 (N_1845,In_78,In_35);
or U1846 (N_1846,In_384,In_24);
xor U1847 (N_1847,In_502,In_213);
or U1848 (N_1848,In_775,In_432);
nor U1849 (N_1849,In_263,In_865);
xnor U1850 (N_1850,In_916,In_974);
and U1851 (N_1851,In_19,In_275);
xnor U1852 (N_1852,In_593,In_211);
xor U1853 (N_1853,In_118,In_856);
nor U1854 (N_1854,In_238,In_29);
nor U1855 (N_1855,In_972,In_841);
nand U1856 (N_1856,In_196,In_609);
or U1857 (N_1857,In_673,In_402);
nor U1858 (N_1858,In_21,In_551);
xor U1859 (N_1859,In_436,In_219);
nor U1860 (N_1860,In_167,In_58);
and U1861 (N_1861,In_852,In_283);
nor U1862 (N_1862,In_440,In_654);
and U1863 (N_1863,In_563,In_340);
and U1864 (N_1864,In_698,In_564);
nand U1865 (N_1865,In_850,In_784);
nand U1866 (N_1866,In_564,In_507);
nor U1867 (N_1867,In_558,In_542);
or U1868 (N_1868,In_197,In_748);
nor U1869 (N_1869,In_846,In_100);
or U1870 (N_1870,In_849,In_720);
or U1871 (N_1871,In_493,In_980);
nand U1872 (N_1872,In_990,In_332);
or U1873 (N_1873,In_293,In_649);
nand U1874 (N_1874,In_708,In_70);
nor U1875 (N_1875,In_334,In_721);
nor U1876 (N_1876,In_544,In_614);
nand U1877 (N_1877,In_258,In_108);
xnor U1878 (N_1878,In_545,In_736);
or U1879 (N_1879,In_431,In_257);
nand U1880 (N_1880,In_61,In_621);
and U1881 (N_1881,In_803,In_374);
and U1882 (N_1882,In_182,In_715);
or U1883 (N_1883,In_498,In_520);
nor U1884 (N_1884,In_894,In_259);
or U1885 (N_1885,In_726,In_831);
nor U1886 (N_1886,In_866,In_661);
nor U1887 (N_1887,In_187,In_90);
or U1888 (N_1888,In_291,In_682);
nand U1889 (N_1889,In_546,In_60);
nand U1890 (N_1890,In_488,In_804);
or U1891 (N_1891,In_128,In_498);
nand U1892 (N_1892,In_571,In_991);
nand U1893 (N_1893,In_400,In_881);
nand U1894 (N_1894,In_795,In_781);
and U1895 (N_1895,In_189,In_715);
nand U1896 (N_1896,In_94,In_905);
and U1897 (N_1897,In_427,In_746);
xnor U1898 (N_1898,In_357,In_900);
or U1899 (N_1899,In_416,In_573);
xnor U1900 (N_1900,In_101,In_755);
xor U1901 (N_1901,In_895,In_722);
xor U1902 (N_1902,In_57,In_163);
and U1903 (N_1903,In_73,In_647);
nor U1904 (N_1904,In_479,In_668);
or U1905 (N_1905,In_103,In_24);
xnor U1906 (N_1906,In_874,In_117);
or U1907 (N_1907,In_661,In_528);
and U1908 (N_1908,In_555,In_157);
nand U1909 (N_1909,In_631,In_169);
or U1910 (N_1910,In_260,In_674);
or U1911 (N_1911,In_48,In_39);
xnor U1912 (N_1912,In_506,In_854);
or U1913 (N_1913,In_1,In_906);
and U1914 (N_1914,In_557,In_865);
xnor U1915 (N_1915,In_545,In_385);
nand U1916 (N_1916,In_207,In_974);
or U1917 (N_1917,In_333,In_455);
xor U1918 (N_1918,In_393,In_735);
nand U1919 (N_1919,In_167,In_322);
xor U1920 (N_1920,In_209,In_634);
and U1921 (N_1921,In_439,In_606);
or U1922 (N_1922,In_266,In_197);
and U1923 (N_1923,In_512,In_153);
nand U1924 (N_1924,In_534,In_74);
xnor U1925 (N_1925,In_405,In_117);
or U1926 (N_1926,In_857,In_886);
and U1927 (N_1927,In_376,In_583);
or U1928 (N_1928,In_754,In_254);
nor U1929 (N_1929,In_770,In_972);
and U1930 (N_1930,In_97,In_180);
and U1931 (N_1931,In_700,In_64);
nand U1932 (N_1932,In_27,In_413);
or U1933 (N_1933,In_44,In_926);
or U1934 (N_1934,In_638,In_298);
nor U1935 (N_1935,In_516,In_822);
xnor U1936 (N_1936,In_117,In_30);
nor U1937 (N_1937,In_165,In_806);
or U1938 (N_1938,In_295,In_27);
and U1939 (N_1939,In_343,In_875);
and U1940 (N_1940,In_537,In_222);
nor U1941 (N_1941,In_154,In_617);
nor U1942 (N_1942,In_455,In_975);
nand U1943 (N_1943,In_376,In_174);
nand U1944 (N_1944,In_901,In_598);
nand U1945 (N_1945,In_870,In_926);
nand U1946 (N_1946,In_639,In_439);
xnor U1947 (N_1947,In_432,In_592);
xnor U1948 (N_1948,In_347,In_659);
nand U1949 (N_1949,In_153,In_568);
nand U1950 (N_1950,In_834,In_873);
nand U1951 (N_1951,In_456,In_538);
and U1952 (N_1952,In_380,In_464);
nor U1953 (N_1953,In_22,In_849);
or U1954 (N_1954,In_946,In_672);
and U1955 (N_1955,In_560,In_702);
nor U1956 (N_1956,In_255,In_114);
nor U1957 (N_1957,In_337,In_112);
nor U1958 (N_1958,In_39,In_574);
nand U1959 (N_1959,In_993,In_442);
xor U1960 (N_1960,In_93,In_854);
or U1961 (N_1961,In_456,In_540);
and U1962 (N_1962,In_174,In_135);
xor U1963 (N_1963,In_711,In_740);
and U1964 (N_1964,In_493,In_430);
nor U1965 (N_1965,In_312,In_442);
nand U1966 (N_1966,In_312,In_356);
xor U1967 (N_1967,In_687,In_521);
nand U1968 (N_1968,In_175,In_676);
nand U1969 (N_1969,In_15,In_183);
and U1970 (N_1970,In_764,In_746);
nand U1971 (N_1971,In_853,In_476);
nor U1972 (N_1972,In_724,In_367);
nor U1973 (N_1973,In_959,In_919);
and U1974 (N_1974,In_537,In_551);
xnor U1975 (N_1975,In_133,In_675);
or U1976 (N_1976,In_441,In_980);
nor U1977 (N_1977,In_738,In_909);
nor U1978 (N_1978,In_785,In_556);
nor U1979 (N_1979,In_39,In_816);
and U1980 (N_1980,In_761,In_817);
and U1981 (N_1981,In_671,In_562);
and U1982 (N_1982,In_383,In_483);
and U1983 (N_1983,In_685,In_24);
nor U1984 (N_1984,In_946,In_948);
nand U1985 (N_1985,In_882,In_514);
nor U1986 (N_1986,In_153,In_136);
nor U1987 (N_1987,In_945,In_705);
or U1988 (N_1988,In_409,In_933);
xor U1989 (N_1989,In_981,In_167);
nor U1990 (N_1990,In_984,In_227);
or U1991 (N_1991,In_500,In_881);
and U1992 (N_1992,In_989,In_793);
nand U1993 (N_1993,In_463,In_406);
nand U1994 (N_1994,In_353,In_963);
or U1995 (N_1995,In_728,In_923);
nand U1996 (N_1996,In_464,In_738);
or U1997 (N_1997,In_217,In_243);
nor U1998 (N_1998,In_506,In_511);
or U1999 (N_1999,In_854,In_893);
nand U2000 (N_2000,In_958,In_938);
xor U2001 (N_2001,In_328,In_660);
nand U2002 (N_2002,In_300,In_173);
and U2003 (N_2003,In_659,In_804);
xor U2004 (N_2004,In_1,In_171);
nand U2005 (N_2005,In_235,In_57);
nor U2006 (N_2006,In_663,In_396);
nor U2007 (N_2007,In_444,In_837);
nand U2008 (N_2008,In_768,In_650);
or U2009 (N_2009,In_473,In_485);
or U2010 (N_2010,In_857,In_105);
nand U2011 (N_2011,In_875,In_954);
nand U2012 (N_2012,In_840,In_708);
nor U2013 (N_2013,In_927,In_335);
nor U2014 (N_2014,In_169,In_78);
or U2015 (N_2015,In_9,In_237);
or U2016 (N_2016,In_533,In_172);
xor U2017 (N_2017,In_853,In_393);
nand U2018 (N_2018,In_966,In_270);
or U2019 (N_2019,In_986,In_852);
xnor U2020 (N_2020,In_393,In_540);
xor U2021 (N_2021,In_182,In_5);
or U2022 (N_2022,In_728,In_705);
and U2023 (N_2023,In_335,In_256);
nand U2024 (N_2024,In_13,In_681);
xnor U2025 (N_2025,In_568,In_612);
or U2026 (N_2026,In_933,In_507);
nor U2027 (N_2027,In_943,In_733);
nor U2028 (N_2028,In_395,In_790);
or U2029 (N_2029,In_157,In_795);
xnor U2030 (N_2030,In_701,In_855);
nand U2031 (N_2031,In_937,In_282);
nand U2032 (N_2032,In_600,In_686);
nand U2033 (N_2033,In_658,In_319);
and U2034 (N_2034,In_439,In_411);
or U2035 (N_2035,In_93,In_791);
nand U2036 (N_2036,In_105,In_498);
nor U2037 (N_2037,In_633,In_158);
and U2038 (N_2038,In_822,In_44);
and U2039 (N_2039,In_302,In_965);
nor U2040 (N_2040,In_425,In_275);
nor U2041 (N_2041,In_200,In_804);
or U2042 (N_2042,In_791,In_519);
nand U2043 (N_2043,In_508,In_613);
and U2044 (N_2044,In_453,In_528);
xnor U2045 (N_2045,In_782,In_801);
and U2046 (N_2046,In_875,In_401);
and U2047 (N_2047,In_373,In_72);
nor U2048 (N_2048,In_908,In_775);
or U2049 (N_2049,In_980,In_76);
or U2050 (N_2050,In_778,In_677);
and U2051 (N_2051,In_364,In_349);
nand U2052 (N_2052,In_390,In_307);
xnor U2053 (N_2053,In_947,In_129);
nor U2054 (N_2054,In_574,In_848);
nor U2055 (N_2055,In_955,In_674);
xor U2056 (N_2056,In_772,In_304);
or U2057 (N_2057,In_500,In_223);
nand U2058 (N_2058,In_643,In_566);
xor U2059 (N_2059,In_201,In_382);
xnor U2060 (N_2060,In_952,In_778);
and U2061 (N_2061,In_631,In_934);
xor U2062 (N_2062,In_302,In_267);
xnor U2063 (N_2063,In_269,In_80);
and U2064 (N_2064,In_704,In_671);
xor U2065 (N_2065,In_505,In_133);
nand U2066 (N_2066,In_608,In_337);
or U2067 (N_2067,In_983,In_978);
or U2068 (N_2068,In_192,In_972);
xnor U2069 (N_2069,In_234,In_155);
nand U2070 (N_2070,In_744,In_891);
or U2071 (N_2071,In_877,In_836);
xnor U2072 (N_2072,In_738,In_920);
nor U2073 (N_2073,In_488,In_997);
nor U2074 (N_2074,In_868,In_19);
nor U2075 (N_2075,In_246,In_174);
nor U2076 (N_2076,In_796,In_56);
and U2077 (N_2077,In_868,In_875);
or U2078 (N_2078,In_529,In_66);
nor U2079 (N_2079,In_615,In_323);
xnor U2080 (N_2080,In_989,In_231);
nand U2081 (N_2081,In_613,In_937);
nor U2082 (N_2082,In_667,In_419);
or U2083 (N_2083,In_52,In_206);
or U2084 (N_2084,In_710,In_606);
or U2085 (N_2085,In_478,In_205);
and U2086 (N_2086,In_52,In_31);
and U2087 (N_2087,In_494,In_434);
nand U2088 (N_2088,In_783,In_843);
xor U2089 (N_2089,In_579,In_13);
or U2090 (N_2090,In_242,In_676);
nor U2091 (N_2091,In_754,In_681);
and U2092 (N_2092,In_187,In_452);
nand U2093 (N_2093,In_86,In_481);
nor U2094 (N_2094,In_688,In_525);
or U2095 (N_2095,In_491,In_892);
or U2096 (N_2096,In_0,In_364);
nand U2097 (N_2097,In_710,In_427);
xor U2098 (N_2098,In_403,In_636);
nor U2099 (N_2099,In_119,In_696);
or U2100 (N_2100,In_362,In_745);
nand U2101 (N_2101,In_142,In_421);
and U2102 (N_2102,In_344,In_331);
xnor U2103 (N_2103,In_148,In_263);
nor U2104 (N_2104,In_769,In_164);
xnor U2105 (N_2105,In_842,In_130);
and U2106 (N_2106,In_16,In_202);
and U2107 (N_2107,In_430,In_861);
or U2108 (N_2108,In_100,In_498);
and U2109 (N_2109,In_126,In_356);
and U2110 (N_2110,In_356,In_205);
xnor U2111 (N_2111,In_864,In_42);
xor U2112 (N_2112,In_317,In_160);
nor U2113 (N_2113,In_589,In_386);
xor U2114 (N_2114,In_139,In_672);
nand U2115 (N_2115,In_693,In_621);
or U2116 (N_2116,In_957,In_134);
and U2117 (N_2117,In_732,In_713);
nand U2118 (N_2118,In_645,In_422);
nor U2119 (N_2119,In_698,In_766);
nor U2120 (N_2120,In_98,In_809);
and U2121 (N_2121,In_939,In_476);
and U2122 (N_2122,In_73,In_249);
nor U2123 (N_2123,In_433,In_446);
and U2124 (N_2124,In_782,In_975);
xor U2125 (N_2125,In_912,In_943);
nand U2126 (N_2126,In_125,In_423);
nor U2127 (N_2127,In_793,In_105);
or U2128 (N_2128,In_672,In_233);
and U2129 (N_2129,In_623,In_122);
and U2130 (N_2130,In_88,In_314);
nand U2131 (N_2131,In_581,In_699);
nor U2132 (N_2132,In_314,In_417);
and U2133 (N_2133,In_529,In_174);
nand U2134 (N_2134,In_531,In_383);
xnor U2135 (N_2135,In_42,In_260);
nor U2136 (N_2136,In_893,In_624);
or U2137 (N_2137,In_288,In_992);
and U2138 (N_2138,In_887,In_988);
or U2139 (N_2139,In_648,In_696);
nand U2140 (N_2140,In_271,In_967);
and U2141 (N_2141,In_693,In_630);
xnor U2142 (N_2142,In_214,In_542);
and U2143 (N_2143,In_601,In_954);
or U2144 (N_2144,In_915,In_934);
nor U2145 (N_2145,In_770,In_234);
or U2146 (N_2146,In_686,In_769);
or U2147 (N_2147,In_838,In_922);
xnor U2148 (N_2148,In_898,In_367);
nand U2149 (N_2149,In_767,In_938);
or U2150 (N_2150,In_819,In_322);
or U2151 (N_2151,In_296,In_473);
and U2152 (N_2152,In_809,In_369);
nor U2153 (N_2153,In_270,In_605);
nor U2154 (N_2154,In_796,In_106);
nand U2155 (N_2155,In_327,In_886);
xor U2156 (N_2156,In_973,In_48);
nor U2157 (N_2157,In_670,In_685);
or U2158 (N_2158,In_729,In_627);
xnor U2159 (N_2159,In_926,In_146);
or U2160 (N_2160,In_227,In_268);
nor U2161 (N_2161,In_220,In_149);
nand U2162 (N_2162,In_475,In_241);
and U2163 (N_2163,In_443,In_573);
nand U2164 (N_2164,In_695,In_231);
nor U2165 (N_2165,In_118,In_667);
or U2166 (N_2166,In_637,In_629);
nand U2167 (N_2167,In_355,In_726);
xor U2168 (N_2168,In_82,In_792);
xnor U2169 (N_2169,In_447,In_126);
xnor U2170 (N_2170,In_63,In_183);
nand U2171 (N_2171,In_141,In_722);
and U2172 (N_2172,In_309,In_652);
nor U2173 (N_2173,In_213,In_35);
or U2174 (N_2174,In_93,In_249);
nand U2175 (N_2175,In_501,In_897);
and U2176 (N_2176,In_699,In_973);
nand U2177 (N_2177,In_163,In_156);
and U2178 (N_2178,In_166,In_633);
nand U2179 (N_2179,In_11,In_825);
nand U2180 (N_2180,In_236,In_950);
nand U2181 (N_2181,In_333,In_63);
and U2182 (N_2182,In_806,In_468);
nand U2183 (N_2183,In_189,In_557);
xor U2184 (N_2184,In_896,In_76);
xor U2185 (N_2185,In_79,In_697);
xnor U2186 (N_2186,In_136,In_528);
nor U2187 (N_2187,In_664,In_920);
nor U2188 (N_2188,In_771,In_912);
and U2189 (N_2189,In_497,In_43);
nand U2190 (N_2190,In_657,In_268);
nor U2191 (N_2191,In_74,In_710);
and U2192 (N_2192,In_998,In_630);
or U2193 (N_2193,In_503,In_13);
xnor U2194 (N_2194,In_726,In_576);
nor U2195 (N_2195,In_477,In_555);
or U2196 (N_2196,In_606,In_642);
and U2197 (N_2197,In_714,In_981);
xor U2198 (N_2198,In_928,In_939);
nand U2199 (N_2199,In_462,In_898);
xor U2200 (N_2200,In_484,In_297);
nor U2201 (N_2201,In_539,In_710);
nand U2202 (N_2202,In_690,In_688);
or U2203 (N_2203,In_401,In_793);
nor U2204 (N_2204,In_598,In_146);
xnor U2205 (N_2205,In_299,In_231);
nand U2206 (N_2206,In_207,In_59);
nand U2207 (N_2207,In_75,In_758);
xnor U2208 (N_2208,In_71,In_487);
or U2209 (N_2209,In_647,In_710);
and U2210 (N_2210,In_836,In_927);
xnor U2211 (N_2211,In_26,In_881);
xnor U2212 (N_2212,In_670,In_216);
and U2213 (N_2213,In_867,In_405);
nand U2214 (N_2214,In_927,In_910);
xor U2215 (N_2215,In_772,In_258);
nor U2216 (N_2216,In_757,In_760);
nand U2217 (N_2217,In_858,In_642);
or U2218 (N_2218,In_583,In_162);
nor U2219 (N_2219,In_871,In_710);
nor U2220 (N_2220,In_969,In_741);
or U2221 (N_2221,In_435,In_789);
nor U2222 (N_2222,In_480,In_539);
xor U2223 (N_2223,In_13,In_188);
xor U2224 (N_2224,In_244,In_183);
or U2225 (N_2225,In_365,In_118);
xor U2226 (N_2226,In_900,In_694);
xnor U2227 (N_2227,In_619,In_410);
and U2228 (N_2228,In_676,In_419);
or U2229 (N_2229,In_570,In_92);
nor U2230 (N_2230,In_774,In_885);
or U2231 (N_2231,In_52,In_4);
nor U2232 (N_2232,In_39,In_824);
nor U2233 (N_2233,In_953,In_952);
nor U2234 (N_2234,In_420,In_465);
nor U2235 (N_2235,In_846,In_888);
xor U2236 (N_2236,In_908,In_180);
and U2237 (N_2237,In_289,In_293);
and U2238 (N_2238,In_62,In_703);
or U2239 (N_2239,In_208,In_967);
nor U2240 (N_2240,In_271,In_102);
nor U2241 (N_2241,In_346,In_4);
or U2242 (N_2242,In_195,In_204);
or U2243 (N_2243,In_313,In_217);
nand U2244 (N_2244,In_428,In_280);
nand U2245 (N_2245,In_591,In_536);
or U2246 (N_2246,In_365,In_844);
and U2247 (N_2247,In_288,In_869);
nand U2248 (N_2248,In_721,In_471);
and U2249 (N_2249,In_330,In_876);
nand U2250 (N_2250,In_630,In_84);
and U2251 (N_2251,In_128,In_348);
xor U2252 (N_2252,In_312,In_570);
or U2253 (N_2253,In_957,In_658);
or U2254 (N_2254,In_364,In_400);
and U2255 (N_2255,In_750,In_155);
and U2256 (N_2256,In_652,In_920);
nor U2257 (N_2257,In_408,In_327);
or U2258 (N_2258,In_456,In_229);
nor U2259 (N_2259,In_237,In_614);
nor U2260 (N_2260,In_760,In_15);
and U2261 (N_2261,In_601,In_396);
xor U2262 (N_2262,In_444,In_581);
xor U2263 (N_2263,In_541,In_583);
and U2264 (N_2264,In_458,In_460);
and U2265 (N_2265,In_999,In_116);
nand U2266 (N_2266,In_428,In_997);
xor U2267 (N_2267,In_889,In_132);
xnor U2268 (N_2268,In_114,In_115);
or U2269 (N_2269,In_97,In_762);
or U2270 (N_2270,In_638,In_951);
and U2271 (N_2271,In_730,In_878);
or U2272 (N_2272,In_930,In_205);
xnor U2273 (N_2273,In_761,In_400);
xnor U2274 (N_2274,In_957,In_247);
xor U2275 (N_2275,In_974,In_704);
xnor U2276 (N_2276,In_143,In_422);
or U2277 (N_2277,In_826,In_435);
nor U2278 (N_2278,In_462,In_423);
or U2279 (N_2279,In_32,In_944);
nand U2280 (N_2280,In_282,In_563);
and U2281 (N_2281,In_780,In_665);
and U2282 (N_2282,In_756,In_201);
or U2283 (N_2283,In_699,In_462);
nor U2284 (N_2284,In_334,In_336);
or U2285 (N_2285,In_65,In_362);
or U2286 (N_2286,In_750,In_454);
nor U2287 (N_2287,In_3,In_828);
nand U2288 (N_2288,In_603,In_122);
xor U2289 (N_2289,In_27,In_811);
nor U2290 (N_2290,In_777,In_631);
or U2291 (N_2291,In_12,In_427);
nand U2292 (N_2292,In_38,In_925);
or U2293 (N_2293,In_413,In_443);
or U2294 (N_2294,In_781,In_98);
xnor U2295 (N_2295,In_185,In_177);
nor U2296 (N_2296,In_872,In_688);
xnor U2297 (N_2297,In_241,In_247);
or U2298 (N_2298,In_471,In_773);
nand U2299 (N_2299,In_147,In_33);
nor U2300 (N_2300,In_10,In_315);
or U2301 (N_2301,In_570,In_358);
and U2302 (N_2302,In_65,In_90);
nand U2303 (N_2303,In_665,In_497);
nor U2304 (N_2304,In_705,In_773);
and U2305 (N_2305,In_431,In_565);
or U2306 (N_2306,In_875,In_58);
or U2307 (N_2307,In_82,In_153);
or U2308 (N_2308,In_346,In_345);
or U2309 (N_2309,In_80,In_39);
or U2310 (N_2310,In_462,In_341);
xor U2311 (N_2311,In_499,In_856);
and U2312 (N_2312,In_451,In_212);
nand U2313 (N_2313,In_87,In_757);
and U2314 (N_2314,In_64,In_983);
xor U2315 (N_2315,In_801,In_123);
xnor U2316 (N_2316,In_353,In_913);
nor U2317 (N_2317,In_705,In_153);
nor U2318 (N_2318,In_545,In_12);
nand U2319 (N_2319,In_815,In_48);
nand U2320 (N_2320,In_369,In_901);
nor U2321 (N_2321,In_97,In_12);
nor U2322 (N_2322,In_807,In_459);
xnor U2323 (N_2323,In_309,In_798);
nor U2324 (N_2324,In_411,In_936);
and U2325 (N_2325,In_233,In_585);
xnor U2326 (N_2326,In_757,In_240);
nand U2327 (N_2327,In_754,In_262);
or U2328 (N_2328,In_486,In_395);
nor U2329 (N_2329,In_785,In_449);
and U2330 (N_2330,In_39,In_958);
or U2331 (N_2331,In_231,In_98);
nand U2332 (N_2332,In_378,In_869);
or U2333 (N_2333,In_782,In_119);
xnor U2334 (N_2334,In_799,In_217);
and U2335 (N_2335,In_874,In_584);
or U2336 (N_2336,In_538,In_88);
nand U2337 (N_2337,In_506,In_926);
nor U2338 (N_2338,In_359,In_943);
nand U2339 (N_2339,In_118,In_884);
and U2340 (N_2340,In_346,In_959);
nand U2341 (N_2341,In_226,In_579);
nor U2342 (N_2342,In_872,In_270);
nor U2343 (N_2343,In_228,In_213);
xor U2344 (N_2344,In_916,In_19);
and U2345 (N_2345,In_917,In_154);
nand U2346 (N_2346,In_234,In_697);
nor U2347 (N_2347,In_383,In_224);
nor U2348 (N_2348,In_50,In_138);
nor U2349 (N_2349,In_160,In_29);
or U2350 (N_2350,In_501,In_58);
xor U2351 (N_2351,In_478,In_128);
nor U2352 (N_2352,In_555,In_212);
or U2353 (N_2353,In_67,In_565);
nand U2354 (N_2354,In_919,In_584);
nor U2355 (N_2355,In_448,In_459);
nand U2356 (N_2356,In_174,In_606);
nor U2357 (N_2357,In_201,In_180);
or U2358 (N_2358,In_434,In_661);
xnor U2359 (N_2359,In_82,In_239);
or U2360 (N_2360,In_754,In_107);
nor U2361 (N_2361,In_906,In_558);
or U2362 (N_2362,In_920,In_455);
and U2363 (N_2363,In_290,In_165);
or U2364 (N_2364,In_788,In_796);
nor U2365 (N_2365,In_887,In_265);
and U2366 (N_2366,In_145,In_829);
nand U2367 (N_2367,In_867,In_653);
xor U2368 (N_2368,In_413,In_150);
xnor U2369 (N_2369,In_181,In_5);
xor U2370 (N_2370,In_42,In_408);
xnor U2371 (N_2371,In_571,In_438);
nand U2372 (N_2372,In_738,In_470);
or U2373 (N_2373,In_212,In_274);
and U2374 (N_2374,In_753,In_275);
xnor U2375 (N_2375,In_690,In_465);
nor U2376 (N_2376,In_875,In_244);
nor U2377 (N_2377,In_498,In_167);
or U2378 (N_2378,In_13,In_73);
xor U2379 (N_2379,In_873,In_580);
nand U2380 (N_2380,In_883,In_305);
nor U2381 (N_2381,In_652,In_315);
or U2382 (N_2382,In_542,In_863);
nand U2383 (N_2383,In_535,In_309);
and U2384 (N_2384,In_544,In_540);
xnor U2385 (N_2385,In_675,In_793);
and U2386 (N_2386,In_163,In_43);
xnor U2387 (N_2387,In_931,In_451);
nand U2388 (N_2388,In_985,In_953);
nor U2389 (N_2389,In_607,In_980);
and U2390 (N_2390,In_961,In_800);
nor U2391 (N_2391,In_895,In_593);
nor U2392 (N_2392,In_489,In_889);
xor U2393 (N_2393,In_940,In_917);
nand U2394 (N_2394,In_601,In_678);
or U2395 (N_2395,In_624,In_281);
nor U2396 (N_2396,In_394,In_649);
or U2397 (N_2397,In_953,In_77);
or U2398 (N_2398,In_235,In_813);
and U2399 (N_2399,In_323,In_447);
or U2400 (N_2400,In_93,In_76);
nor U2401 (N_2401,In_357,In_13);
xor U2402 (N_2402,In_648,In_232);
xnor U2403 (N_2403,In_977,In_880);
and U2404 (N_2404,In_192,In_758);
nand U2405 (N_2405,In_916,In_9);
nand U2406 (N_2406,In_534,In_95);
xnor U2407 (N_2407,In_239,In_84);
nand U2408 (N_2408,In_639,In_549);
or U2409 (N_2409,In_34,In_525);
nand U2410 (N_2410,In_678,In_991);
and U2411 (N_2411,In_867,In_120);
nor U2412 (N_2412,In_683,In_255);
or U2413 (N_2413,In_567,In_23);
and U2414 (N_2414,In_863,In_184);
or U2415 (N_2415,In_432,In_126);
nand U2416 (N_2416,In_157,In_415);
nand U2417 (N_2417,In_332,In_639);
nor U2418 (N_2418,In_870,In_987);
and U2419 (N_2419,In_745,In_430);
or U2420 (N_2420,In_291,In_702);
xor U2421 (N_2421,In_359,In_85);
xor U2422 (N_2422,In_653,In_735);
nand U2423 (N_2423,In_431,In_145);
xnor U2424 (N_2424,In_315,In_305);
xnor U2425 (N_2425,In_736,In_665);
nand U2426 (N_2426,In_831,In_263);
and U2427 (N_2427,In_189,In_369);
nand U2428 (N_2428,In_105,In_827);
and U2429 (N_2429,In_76,In_21);
xnor U2430 (N_2430,In_289,In_36);
nor U2431 (N_2431,In_286,In_310);
nor U2432 (N_2432,In_74,In_1);
nor U2433 (N_2433,In_641,In_808);
xor U2434 (N_2434,In_963,In_363);
nand U2435 (N_2435,In_370,In_998);
or U2436 (N_2436,In_210,In_472);
and U2437 (N_2437,In_88,In_32);
or U2438 (N_2438,In_725,In_754);
xor U2439 (N_2439,In_497,In_692);
xnor U2440 (N_2440,In_222,In_934);
xnor U2441 (N_2441,In_89,In_504);
nand U2442 (N_2442,In_565,In_950);
and U2443 (N_2443,In_647,In_277);
nor U2444 (N_2444,In_862,In_803);
nor U2445 (N_2445,In_602,In_56);
nand U2446 (N_2446,In_998,In_727);
nor U2447 (N_2447,In_327,In_181);
nand U2448 (N_2448,In_293,In_724);
or U2449 (N_2449,In_339,In_669);
and U2450 (N_2450,In_415,In_22);
nand U2451 (N_2451,In_778,In_767);
and U2452 (N_2452,In_477,In_182);
nor U2453 (N_2453,In_495,In_267);
or U2454 (N_2454,In_194,In_456);
nand U2455 (N_2455,In_724,In_618);
xor U2456 (N_2456,In_55,In_775);
nand U2457 (N_2457,In_323,In_837);
nand U2458 (N_2458,In_525,In_476);
nor U2459 (N_2459,In_636,In_919);
or U2460 (N_2460,In_161,In_844);
xor U2461 (N_2461,In_351,In_738);
xnor U2462 (N_2462,In_300,In_736);
nor U2463 (N_2463,In_200,In_336);
nand U2464 (N_2464,In_395,In_39);
xor U2465 (N_2465,In_87,In_466);
and U2466 (N_2466,In_824,In_315);
nor U2467 (N_2467,In_770,In_693);
or U2468 (N_2468,In_464,In_403);
or U2469 (N_2469,In_909,In_521);
xnor U2470 (N_2470,In_392,In_868);
or U2471 (N_2471,In_838,In_175);
and U2472 (N_2472,In_244,In_265);
nand U2473 (N_2473,In_312,In_6);
or U2474 (N_2474,In_509,In_964);
nand U2475 (N_2475,In_790,In_69);
or U2476 (N_2476,In_29,In_231);
or U2477 (N_2477,In_11,In_1);
xor U2478 (N_2478,In_780,In_401);
and U2479 (N_2479,In_528,In_107);
nor U2480 (N_2480,In_338,In_442);
nand U2481 (N_2481,In_390,In_585);
and U2482 (N_2482,In_895,In_485);
xor U2483 (N_2483,In_907,In_255);
nand U2484 (N_2484,In_326,In_76);
or U2485 (N_2485,In_28,In_191);
xor U2486 (N_2486,In_806,In_192);
or U2487 (N_2487,In_755,In_836);
nor U2488 (N_2488,In_494,In_139);
nor U2489 (N_2489,In_673,In_394);
or U2490 (N_2490,In_456,In_978);
nand U2491 (N_2491,In_633,In_615);
nor U2492 (N_2492,In_540,In_814);
xnor U2493 (N_2493,In_800,In_137);
xor U2494 (N_2494,In_399,In_201);
nand U2495 (N_2495,In_324,In_242);
or U2496 (N_2496,In_269,In_245);
nand U2497 (N_2497,In_276,In_582);
nor U2498 (N_2498,In_363,In_10);
xor U2499 (N_2499,In_485,In_588);
and U2500 (N_2500,N_2392,N_2177);
xnor U2501 (N_2501,N_790,N_1902);
xor U2502 (N_2502,N_2132,N_816);
or U2503 (N_2503,N_2418,N_1438);
xnor U2504 (N_2504,N_2310,N_1005);
and U2505 (N_2505,N_985,N_1255);
or U2506 (N_2506,N_1466,N_109);
and U2507 (N_2507,N_1998,N_1298);
and U2508 (N_2508,N_2184,N_1317);
and U2509 (N_2509,N_2147,N_2465);
nor U2510 (N_2510,N_2094,N_1692);
or U2511 (N_2511,N_2356,N_2098);
xnor U2512 (N_2512,N_1111,N_389);
or U2513 (N_2513,N_212,N_2081);
nor U2514 (N_2514,N_2220,N_2163);
and U2515 (N_2515,N_2388,N_882);
xor U2516 (N_2516,N_805,N_891);
xnor U2517 (N_2517,N_1425,N_1731);
or U2518 (N_2518,N_2330,N_0);
nor U2519 (N_2519,N_1453,N_436);
nand U2520 (N_2520,N_784,N_183);
xnor U2521 (N_2521,N_388,N_564);
xor U2522 (N_2522,N_1730,N_1521);
nor U2523 (N_2523,N_258,N_2375);
and U2524 (N_2524,N_1419,N_370);
or U2525 (N_2525,N_544,N_1959);
nand U2526 (N_2526,N_959,N_1756);
xnor U2527 (N_2527,N_1660,N_938);
or U2528 (N_2528,N_1485,N_992);
nor U2529 (N_2529,N_2275,N_1577);
and U2530 (N_2530,N_1527,N_2001);
xor U2531 (N_2531,N_1397,N_1482);
xnor U2532 (N_2532,N_1178,N_1934);
nor U2533 (N_2533,N_2076,N_2011);
nand U2534 (N_2534,N_1162,N_1243);
nand U2535 (N_2535,N_2302,N_511);
nand U2536 (N_2536,N_344,N_2316);
nor U2537 (N_2537,N_1291,N_2119);
nor U2538 (N_2538,N_1191,N_310);
and U2539 (N_2539,N_1781,N_1832);
or U2540 (N_2540,N_507,N_1018);
nand U2541 (N_2541,N_1327,N_1738);
nand U2542 (N_2542,N_291,N_802);
nand U2543 (N_2543,N_1887,N_2495);
and U2544 (N_2544,N_557,N_456);
xnor U2545 (N_2545,N_2442,N_2372);
xor U2546 (N_2546,N_1290,N_692);
xor U2547 (N_2547,N_115,N_725);
xor U2548 (N_2548,N_253,N_1475);
or U2549 (N_2549,N_948,N_1764);
or U2550 (N_2550,N_1450,N_1461);
or U2551 (N_2551,N_2291,N_1341);
nand U2552 (N_2552,N_1365,N_2438);
and U2553 (N_2553,N_1121,N_201);
and U2554 (N_2554,N_155,N_1616);
and U2555 (N_2555,N_1233,N_2385);
or U2556 (N_2556,N_1356,N_974);
xor U2557 (N_2557,N_2183,N_811);
nor U2558 (N_2558,N_2016,N_1359);
or U2559 (N_2559,N_2037,N_2355);
nand U2560 (N_2560,N_1463,N_1498);
xor U2561 (N_2561,N_2050,N_1938);
xnor U2562 (N_2562,N_2022,N_1589);
nor U2563 (N_2563,N_2267,N_425);
nor U2564 (N_2564,N_395,N_14);
nor U2565 (N_2565,N_1287,N_1911);
nor U2566 (N_2566,N_903,N_92);
nand U2567 (N_2567,N_2,N_625);
xor U2568 (N_2568,N_2226,N_2155);
or U2569 (N_2569,N_412,N_1247);
nor U2570 (N_2570,N_1590,N_2391);
or U2571 (N_2571,N_662,N_1802);
and U2572 (N_2572,N_398,N_772);
xnor U2573 (N_2573,N_1280,N_1770);
nor U2574 (N_2574,N_208,N_1686);
nor U2575 (N_2575,N_660,N_821);
and U2576 (N_2576,N_2031,N_1912);
xnor U2577 (N_2577,N_993,N_1156);
nor U2578 (N_2578,N_1544,N_367);
and U2579 (N_2579,N_2073,N_2100);
nand U2580 (N_2580,N_2018,N_1715);
nand U2581 (N_2581,N_1351,N_2317);
or U2582 (N_2582,N_1542,N_2200);
nand U2583 (N_2583,N_1908,N_1434);
or U2584 (N_2584,N_747,N_267);
and U2585 (N_2585,N_1098,N_1701);
xor U2586 (N_2586,N_1609,N_1622);
nand U2587 (N_2587,N_171,N_1009);
and U2588 (N_2588,N_1193,N_2087);
nand U2589 (N_2589,N_1946,N_1285);
xnor U2590 (N_2590,N_2093,N_1670);
nand U2591 (N_2591,N_304,N_1693);
and U2592 (N_2592,N_2494,N_1313);
nand U2593 (N_2593,N_755,N_1188);
nand U2594 (N_2594,N_1654,N_926);
xnor U2595 (N_2595,N_1179,N_676);
nand U2596 (N_2596,N_200,N_2111);
or U2597 (N_2597,N_1500,N_1245);
xnor U2598 (N_2598,N_1765,N_943);
and U2599 (N_2599,N_2270,N_257);
and U2600 (N_2600,N_1321,N_1926);
nor U2601 (N_2601,N_2125,N_1709);
or U2602 (N_2602,N_309,N_423);
or U2603 (N_2603,N_1920,N_1848);
and U2604 (N_2604,N_2199,N_333);
nand U2605 (N_2605,N_490,N_2015);
xor U2606 (N_2606,N_441,N_2334);
nand U2607 (N_2607,N_1746,N_1751);
xnor U2608 (N_2608,N_1889,N_1456);
xnor U2609 (N_2609,N_2107,N_1608);
or U2610 (N_2610,N_1969,N_347);
xnor U2611 (N_2611,N_247,N_1256);
and U2612 (N_2612,N_1523,N_1155);
and U2613 (N_2613,N_1673,N_1295);
xnor U2614 (N_2614,N_1535,N_1905);
nand U2615 (N_2615,N_470,N_236);
xor U2616 (N_2616,N_443,N_764);
and U2617 (N_2617,N_1424,N_2000);
xnor U2618 (N_2618,N_1587,N_2411);
nand U2619 (N_2619,N_1963,N_2196);
nand U2620 (N_2620,N_102,N_1449);
and U2621 (N_2621,N_1548,N_1723);
nor U2622 (N_2622,N_1404,N_2029);
nor U2623 (N_2623,N_941,N_2437);
or U2624 (N_2624,N_1480,N_1226);
nand U2625 (N_2625,N_553,N_2403);
nand U2626 (N_2626,N_1329,N_1965);
and U2627 (N_2627,N_2381,N_2401);
xor U2628 (N_2628,N_1993,N_1552);
nor U2629 (N_2629,N_763,N_1238);
nand U2630 (N_2630,N_2292,N_1721);
nand U2631 (N_2631,N_1279,N_1985);
and U2632 (N_2632,N_2272,N_2445);
nand U2633 (N_2633,N_513,N_193);
or U2634 (N_2634,N_1232,N_2090);
and U2635 (N_2635,N_972,N_1271);
nand U2636 (N_2636,N_1075,N_2305);
and U2637 (N_2637,N_2467,N_906);
nor U2638 (N_2638,N_775,N_1016);
nor U2639 (N_2639,N_778,N_1072);
xor U2640 (N_2640,N_1991,N_793);
and U2641 (N_2641,N_588,N_1793);
and U2642 (N_2642,N_2422,N_1070);
xor U2643 (N_2643,N_34,N_604);
nand U2644 (N_2644,N_1652,N_420);
or U2645 (N_2645,N_2407,N_1145);
xor U2646 (N_2646,N_113,N_1275);
or U2647 (N_2647,N_1180,N_1602);
and U2648 (N_2648,N_220,N_1357);
xor U2649 (N_2649,N_1923,N_1235);
xnor U2650 (N_2650,N_2065,N_1406);
or U2651 (N_2651,N_1541,N_917);
or U2652 (N_2652,N_1545,N_721);
xor U2653 (N_2653,N_1936,N_242);
nand U2654 (N_2654,N_2352,N_1328);
and U2655 (N_2655,N_2239,N_1713);
and U2656 (N_2656,N_1251,N_332);
nand U2657 (N_2657,N_1213,N_1375);
xor U2658 (N_2658,N_738,N_830);
nor U2659 (N_2659,N_1845,N_342);
or U2660 (N_2660,N_2099,N_1760);
xnor U2661 (N_2661,N_2363,N_2209);
or U2662 (N_2662,N_780,N_581);
nand U2663 (N_2663,N_524,N_2473);
xor U2664 (N_2664,N_639,N_103);
xnor U2665 (N_2665,N_3,N_1631);
nor U2666 (N_2666,N_1809,N_96);
xnor U2667 (N_2667,N_1847,N_1925);
xnor U2668 (N_2668,N_2179,N_1392);
or U2669 (N_2669,N_1276,N_2289);
nor U2670 (N_2670,N_1166,N_814);
nor U2671 (N_2671,N_495,N_2146);
nand U2672 (N_2672,N_213,N_1972);
xnor U2673 (N_2673,N_1083,N_890);
nand U2674 (N_2674,N_1000,N_2215);
or U2675 (N_2675,N_1398,N_506);
and U2676 (N_2676,N_1400,N_1019);
xnor U2677 (N_2677,N_679,N_1868);
or U2678 (N_2678,N_1761,N_1859);
or U2679 (N_2679,N_1687,N_230);
nor U2680 (N_2680,N_1600,N_1244);
nand U2681 (N_2681,N_187,N_925);
nand U2682 (N_2682,N_1223,N_1669);
xnor U2683 (N_2683,N_1754,N_669);
xor U2684 (N_2684,N_789,N_1879);
xnor U2685 (N_2685,N_1896,N_274);
xor U2686 (N_2686,N_1851,N_149);
nand U2687 (N_2687,N_769,N_1067);
xnor U2688 (N_2688,N_2410,N_5);
and U2689 (N_2689,N_1464,N_476);
nand U2690 (N_2690,N_1039,N_2482);
nand U2691 (N_2691,N_1488,N_964);
or U2692 (N_2692,N_2216,N_1592);
and U2693 (N_2693,N_602,N_1659);
and U2694 (N_2694,N_130,N_2026);
and U2695 (N_2695,N_259,N_2131);
and U2696 (N_2696,N_2174,N_411);
or U2697 (N_2697,N_1837,N_1818);
or U2698 (N_2698,N_1913,N_1556);
nand U2699 (N_2699,N_2472,N_991);
nand U2700 (N_2700,N_978,N_836);
nand U2701 (N_2701,N_633,N_792);
nor U2702 (N_2702,N_2181,N_808);
xor U2703 (N_2703,N_1508,N_1065);
nand U2704 (N_2704,N_1811,N_1248);
nor U2705 (N_2705,N_1787,N_1735);
nor U2706 (N_2706,N_1575,N_1873);
xnor U2707 (N_2707,N_2338,N_391);
xnor U2708 (N_2708,N_63,N_431);
nand U2709 (N_2709,N_225,N_451);
xor U2710 (N_2710,N_2164,N_17);
and U2711 (N_2711,N_1778,N_89);
nand U2712 (N_2712,N_2396,N_466);
nand U2713 (N_2713,N_718,N_1200);
nand U2714 (N_2714,N_1705,N_1246);
nand U2715 (N_2715,N_1827,N_413);
nor U2716 (N_2716,N_2167,N_1635);
nand U2717 (N_2717,N_859,N_2151);
xnor U2718 (N_2718,N_1459,N_1994);
nand U2719 (N_2719,N_1511,N_1046);
and U2720 (N_2720,N_1289,N_947);
nor U2721 (N_2721,N_1333,N_416);
xor U2722 (N_2722,N_1330,N_678);
nand U2723 (N_2723,N_138,N_1990);
nor U2724 (N_2724,N_1307,N_1355);
or U2725 (N_2725,N_605,N_2325);
xnor U2726 (N_2726,N_1992,N_781);
xnor U2727 (N_2727,N_167,N_1784);
nor U2728 (N_2728,N_417,N_742);
nor U2729 (N_2729,N_1060,N_1797);
and U2730 (N_2730,N_1995,N_1101);
or U2731 (N_2731,N_783,N_786);
or U2732 (N_2732,N_701,N_643);
and U2733 (N_2733,N_592,N_372);
xnor U2734 (N_2734,N_2150,N_1826);
and U2735 (N_2735,N_1426,N_1838);
and U2736 (N_2736,N_361,N_462);
nor U2737 (N_2737,N_1305,N_1619);
or U2738 (N_2738,N_1109,N_782);
xnor U2739 (N_2739,N_1,N_57);
or U2740 (N_2740,N_2428,N_1953);
and U2741 (N_2741,N_627,N_321);
or U2742 (N_2742,N_1979,N_862);
nor U2743 (N_2743,N_1052,N_1566);
nand U2744 (N_2744,N_2489,N_2149);
and U2745 (N_2745,N_2053,N_32);
and U2746 (N_2746,N_1804,N_170);
nand U2747 (N_2747,N_735,N_1565);
xnor U2748 (N_2748,N_145,N_350);
or U2749 (N_2749,N_734,N_572);
xnor U2750 (N_2750,N_1047,N_2319);
or U2751 (N_2751,N_2227,N_912);
nor U2752 (N_2752,N_410,N_1496);
and U2753 (N_2753,N_706,N_1173);
nand U2754 (N_2754,N_424,N_895);
or U2755 (N_2755,N_1624,N_573);
nand U2756 (N_2756,N_336,N_883);
nor U2757 (N_2757,N_897,N_1216);
or U2758 (N_2758,N_1401,N_2326);
nand U2759 (N_2759,N_1961,N_2478);
nor U2760 (N_2760,N_2176,N_488);
or U2761 (N_2761,N_2153,N_2349);
xnor U2762 (N_2762,N_1739,N_571);
and U2763 (N_2763,N_824,N_2331);
or U2764 (N_2764,N_2068,N_2004);
or U2765 (N_2765,N_8,N_2408);
nand U2766 (N_2766,N_329,N_2205);
xor U2767 (N_2767,N_2148,N_500);
and U2768 (N_2768,N_238,N_1741);
or U2769 (N_2769,N_642,N_1894);
xnor U2770 (N_2770,N_91,N_1656);
nand U2771 (N_2771,N_1583,N_319);
nor U2772 (N_2772,N_2033,N_41);
or U2773 (N_2773,N_2002,N_1205);
xnor U2774 (N_2774,N_714,N_1788);
nand U2775 (N_2775,N_2013,N_826);
and U2776 (N_2776,N_303,N_1691);
nand U2777 (N_2777,N_42,N_1407);
nor U2778 (N_2778,N_708,N_1817);
and U2779 (N_2779,N_2373,N_1884);
nor U2780 (N_2780,N_1020,N_671);
nor U2781 (N_2781,N_7,N_2282);
and U2782 (N_2782,N_736,N_920);
xor U2783 (N_2783,N_324,N_260);
nand U2784 (N_2784,N_2058,N_630);
nor U2785 (N_2785,N_371,N_737);
nand U2786 (N_2786,N_1803,N_554);
nand U2787 (N_2787,N_522,N_2371);
and U2788 (N_2788,N_2389,N_1582);
and U2789 (N_2789,N_1630,N_1444);
xor U2790 (N_2790,N_810,N_983);
xor U2791 (N_2791,N_527,N_1588);
and U2792 (N_2792,N_1664,N_120);
or U2793 (N_2793,N_760,N_2452);
and U2794 (N_2794,N_1984,N_503);
or U2795 (N_2795,N_1895,N_716);
xor U2796 (N_2796,N_1212,N_1732);
nor U2797 (N_2797,N_2429,N_555);
nor U2798 (N_2798,N_163,N_1906);
nand U2799 (N_2799,N_244,N_1505);
and U2800 (N_2800,N_1006,N_1015);
and U2801 (N_2801,N_1300,N_1642);
xor U2802 (N_2802,N_2402,N_1627);
nor U2803 (N_2803,N_1085,N_868);
nor U2804 (N_2804,N_954,N_93);
xnor U2805 (N_2805,N_1674,N_1152);
or U2806 (N_2806,N_2221,N_1331);
nor U2807 (N_2807,N_695,N_2191);
and U2808 (N_2808,N_966,N_1337);
nand U2809 (N_2809,N_128,N_2064);
nand U2810 (N_2810,N_1144,N_2104);
or U2811 (N_2811,N_2036,N_1265);
xor U2812 (N_2812,N_2406,N_942);
or U2813 (N_2813,N_803,N_795);
nor U2814 (N_2814,N_2170,N_2214);
and U2815 (N_2815,N_2311,N_381);
nor U2816 (N_2816,N_1737,N_741);
or U2817 (N_2817,N_1209,N_953);
xnor U2818 (N_2818,N_415,N_1682);
nand U2819 (N_2819,N_224,N_2010);
nor U2820 (N_2820,N_796,N_794);
xor U2821 (N_2821,N_287,N_2337);
nor U2822 (N_2822,N_1951,N_901);
nand U2823 (N_2823,N_1639,N_1530);
xnor U2824 (N_2824,N_2252,N_1146);
xor U2825 (N_2825,N_2212,N_730);
xnor U2826 (N_2826,N_2161,N_1258);
nor U2827 (N_2827,N_2458,N_117);
and U2828 (N_2828,N_222,N_1286);
xor U2829 (N_2829,N_66,N_647);
or U2830 (N_2830,N_1512,N_996);
or U2831 (N_2831,N_1763,N_894);
xor U2832 (N_2832,N_1448,N_1745);
nand U2833 (N_2833,N_1315,N_1550);
nor U2834 (N_2834,N_1880,N_1843);
or U2835 (N_2835,N_585,N_450);
and U2836 (N_2836,N_2320,N_663);
or U2837 (N_2837,N_72,N_1376);
or U2838 (N_2838,N_526,N_1395);
xnor U2839 (N_2839,N_378,N_1753);
xor U2840 (N_2840,N_1503,N_528);
and U2841 (N_2841,N_1458,N_2039);
nor U2842 (N_2842,N_1888,N_819);
nand U2843 (N_2843,N_865,N_1377);
or U2844 (N_2844,N_2229,N_85);
or U2845 (N_2845,N_297,N_237);
nor U2846 (N_2846,N_1573,N_904);
or U2847 (N_2847,N_746,N_1293);
or U2848 (N_2848,N_429,N_1164);
xnor U2849 (N_2849,N_1568,N_1270);
xor U2850 (N_2850,N_1743,N_1092);
nor U2851 (N_2851,N_2218,N_2069);
or U2852 (N_2852,N_1822,N_1358);
nor U2853 (N_2853,N_841,N_520);
and U2854 (N_2854,N_469,N_231);
and U2855 (N_2855,N_1779,N_586);
nor U2856 (N_2856,N_1928,N_1860);
or U2857 (N_2857,N_552,N_221);
xnor U2858 (N_2858,N_2444,N_448);
or U2859 (N_2859,N_1528,N_1679);
xnor U2860 (N_2860,N_1266,N_1833);
xor U2861 (N_2861,N_86,N_1176);
nor U2862 (N_2862,N_539,N_768);
xor U2863 (N_2863,N_1441,N_1457);
or U2864 (N_2864,N_376,N_2457);
or U2865 (N_2865,N_1495,N_141);
or U2866 (N_2866,N_628,N_1231);
xor U2867 (N_2867,N_2051,N_409);
or U2868 (N_2868,N_1727,N_493);
and U2869 (N_2869,N_1640,N_675);
nor U2870 (N_2870,N_1011,N_1201);
or U2871 (N_2871,N_617,N_2443);
and U2872 (N_2872,N_649,N_1489);
and U2873 (N_2873,N_1935,N_860);
xnor U2874 (N_2874,N_1432,N_1104);
nand U2875 (N_2875,N_1857,N_1914);
nor U2876 (N_2876,N_1783,N_2260);
nor U2877 (N_2877,N_1308,N_1676);
and U2878 (N_2878,N_1237,N_2084);
xnor U2879 (N_2879,N_2180,N_1350);
xor U2880 (N_2880,N_1522,N_1777);
nor U2881 (N_2881,N_1825,N_889);
nand U2882 (N_2882,N_22,N_2066);
or U2883 (N_2883,N_589,N_638);
xor U2884 (N_2884,N_843,N_1097);
and U2885 (N_2885,N_807,N_1875);
nand U2886 (N_2886,N_2424,N_584);
nor U2887 (N_2887,N_1971,N_1830);
nand U2888 (N_2888,N_1491,N_918);
or U2889 (N_2889,N_644,N_1786);
xor U2890 (N_2890,N_998,N_261);
or U2891 (N_2891,N_2460,N_1117);
nand U2892 (N_2892,N_272,N_2007);
nand U2893 (N_2893,N_2106,N_2294);
or U2894 (N_2894,N_24,N_1263);
xor U2895 (N_2895,N_2236,N_1282);
xnor U2896 (N_2896,N_1499,N_1975);
nand U2897 (N_2897,N_76,N_1253);
and U2898 (N_2898,N_1428,N_101);
nor U2899 (N_2899,N_965,N_1980);
xor U2900 (N_2900,N_538,N_933);
and U2901 (N_2901,N_1562,N_1613);
or U2902 (N_2902,N_54,N_26);
nor U2903 (N_2903,N_958,N_1623);
nor U2904 (N_2904,N_1274,N_2485);
and U2905 (N_2905,N_2207,N_2312);
or U2906 (N_2906,N_1234,N_375);
and U2907 (N_2907,N_1882,N_1941);
nor U2908 (N_2908,N_635,N_1211);
nand U2909 (N_2909,N_767,N_131);
nand U2910 (N_2910,N_922,N_2397);
nor U2911 (N_2911,N_67,N_2012);
xnor U2912 (N_2912,N_2258,N_2251);
nor U2913 (N_2913,N_366,N_1675);
and U2914 (N_2914,N_1782,N_570);
and U2915 (N_2915,N_1116,N_278);
and U2916 (N_2916,N_419,N_1045);
nor U2917 (N_2917,N_1267,N_80);
or U2918 (N_2918,N_368,N_726);
or U2919 (N_2919,N_981,N_2486);
or U2920 (N_2920,N_1034,N_1454);
or U2921 (N_2921,N_2208,N_2343);
xor U2922 (N_2922,N_1921,N_1372);
or U2923 (N_2923,N_1586,N_2059);
nand U2924 (N_2924,N_1944,N_2096);
xor U2925 (N_2925,N_1447,N_1703);
or U2926 (N_2926,N_1199,N_2024);
nand U2927 (N_2927,N_558,N_2113);
xnor U2928 (N_2928,N_655,N_1771);
and U2929 (N_2929,N_2194,N_1148);
nand U2930 (N_2930,N_2361,N_282);
nor U2931 (N_2931,N_2290,N_1048);
nand U2932 (N_2932,N_2233,N_219);
xnor U2933 (N_2933,N_1143,N_2123);
nand U2934 (N_2934,N_1384,N_1943);
nand U2935 (N_2935,N_2195,N_2197);
and U2936 (N_2936,N_911,N_1219);
and U2937 (N_2937,N_902,N_313);
or U2938 (N_2938,N_1643,N_254);
xnor U2939 (N_2939,N_1036,N_1641);
nor U2940 (N_2940,N_861,N_940);
nor U2941 (N_2941,N_353,N_1136);
nor U2942 (N_2942,N_1264,N_1089);
or U2943 (N_2943,N_1574,N_1685);
nor U2944 (N_2944,N_2217,N_1997);
nand U2945 (N_2945,N_1629,N_835);
or U2946 (N_2946,N_1494,N_334);
xnor U2947 (N_2947,N_1846,N_479);
nand U2948 (N_2948,N_1755,N_2359);
xor U2949 (N_2949,N_1471,N_809);
or U2950 (N_2950,N_2285,N_1854);
nor U2951 (N_2951,N_609,N_2379);
nand U2952 (N_2952,N_1138,N_1335);
nor U2953 (N_2953,N_1649,N_480);
or U2954 (N_2954,N_140,N_369);
xnor U2955 (N_2955,N_330,N_1093);
or U2956 (N_2956,N_1555,N_1645);
or U2957 (N_2957,N_1031,N_825);
or U2958 (N_2958,N_2109,N_2206);
nand U2959 (N_2959,N_1347,N_2415);
nor U2960 (N_2960,N_473,N_1340);
or U2961 (N_2961,N_1318,N_1957);
and U2962 (N_2962,N_641,N_615);
nand U2963 (N_2963,N_1988,N_48);
nor U2964 (N_2964,N_1815,N_530);
and U2965 (N_2965,N_1222,N_1954);
nand U2966 (N_2966,N_399,N_548);
or U2967 (N_2967,N_502,N_2431);
nand U2968 (N_2968,N_787,N_2336);
xnor U2969 (N_2969,N_65,N_1470);
xnor U2970 (N_2970,N_345,N_2187);
or U2971 (N_2971,N_1752,N_1174);
nand U2972 (N_2972,N_1572,N_1414);
or U2973 (N_2973,N_1462,N_2126);
and U2974 (N_2974,N_1418,N_428);
and U2975 (N_2975,N_945,N_464);
nor U2976 (N_2976,N_1017,N_540);
xnor U2977 (N_2977,N_2230,N_968);
nand U2978 (N_2978,N_1538,N_2315);
and U2979 (N_2979,N_771,N_1968);
nand U2980 (N_2980,N_50,N_59);
nor U2981 (N_2981,N_1103,N_1452);
nor U2982 (N_2982,N_887,N_1862);
nand U2983 (N_2983,N_1949,N_1539);
nor U2984 (N_2984,N_249,N_886);
or U2985 (N_2985,N_2287,N_1547);
and U2986 (N_2986,N_1805,N_1427);
xor U2987 (N_2987,N_724,N_999);
nor U2988 (N_2988,N_1194,N_1405);
or U2989 (N_2989,N_2169,N_1551);
nor U2990 (N_2990,N_266,N_543);
nor U2991 (N_2991,N_1310,N_1273);
and U2992 (N_2992,N_400,N_40);
or U2993 (N_2993,N_2116,N_294);
nand U2994 (N_2994,N_900,N_2426);
or U2995 (N_2995,N_636,N_2383);
nand U2996 (N_2996,N_1747,N_1278);
or U2997 (N_2997,N_850,N_600);
or U2998 (N_2998,N_1068,N_152);
xor U2999 (N_2999,N_132,N_1607);
nor U3000 (N_3000,N_1728,N_2095);
xor U3001 (N_3001,N_1885,N_610);
xor U3002 (N_3002,N_1362,N_957);
nand U3003 (N_3003,N_2466,N_256);
nor U3004 (N_3004,N_295,N_1982);
and U3005 (N_3005,N_1468,N_190);
nand U3006 (N_3006,N_2284,N_181);
xor U3007 (N_3007,N_380,N_2256);
or U3008 (N_3008,N_1014,N_2387);
or U3009 (N_3009,N_2470,N_732);
nand U3010 (N_3010,N_2313,N_1973);
nor U3011 (N_3011,N_439,N_892);
and U3012 (N_3012,N_74,N_1767);
nand U3013 (N_3013,N_289,N_1576);
nand U3014 (N_3014,N_444,N_1254);
nand U3015 (N_3015,N_2082,N_1531);
xnor U3016 (N_3016,N_845,N_56);
and U3017 (N_3017,N_1662,N_1718);
or U3018 (N_3018,N_967,N_563);
xor U3019 (N_3019,N_743,N_280);
or U3020 (N_3020,N_1634,N_250);
nor U3021 (N_3021,N_853,N_1716);
xnor U3022 (N_3022,N_2052,N_263);
nand U3023 (N_3023,N_1867,N_1169);
xor U3024 (N_3024,N_1187,N_637);
and U3025 (N_3025,N_1455,N_129);
xor U3026 (N_3026,N_913,N_1192);
and U3027 (N_3027,N_1239,N_1986);
nand U3028 (N_3028,N_1049,N_952);
nor U3029 (N_3029,N_39,N_688);
xnor U3030 (N_3030,N_2300,N_1033);
xor U3031 (N_3031,N_616,N_657);
xor U3032 (N_3032,N_82,N_2297);
or U3033 (N_3033,N_1106,N_1021);
xor U3034 (N_3034,N_1338,N_1465);
nor U3035 (N_3035,N_147,N_893);
xor U3036 (N_3036,N_2398,N_880);
and U3037 (N_3037,N_2061,N_707);
xor U3038 (N_3038,N_2014,N_1689);
nand U3039 (N_3039,N_2464,N_2158);
xnor U3040 (N_3040,N_1283,N_1821);
and U3041 (N_3041,N_1385,N_1740);
nand U3042 (N_3042,N_1240,N_1605);
and U3043 (N_3043,N_335,N_2144);
and U3044 (N_3044,N_119,N_2261);
nand U3045 (N_3045,N_2089,N_229);
or U3046 (N_3046,N_986,N_1323);
xnor U3047 (N_3047,N_112,N_848);
or U3048 (N_3048,N_594,N_750);
nor U3049 (N_3049,N_2419,N_1064);
xnor U3050 (N_3050,N_1115,N_1473);
nor U3051 (N_3051,N_189,N_460);
xor U3052 (N_3052,N_316,N_1836);
and U3053 (N_3053,N_317,N_651);
and U3054 (N_3054,N_9,N_124);
xor U3055 (N_3055,N_677,N_652);
xnor U3056 (N_3056,N_467,N_1415);
xnor U3057 (N_3057,N_844,N_545);
and U3058 (N_3058,N_2264,N_1750);
and U3059 (N_3059,N_1378,N_608);
and U3060 (N_3060,N_1729,N_1559);
and U3061 (N_3061,N_2461,N_449);
and U3062 (N_3062,N_90,N_2423);
nand U3063 (N_3063,N_800,N_1697);
or U3064 (N_3064,N_596,N_2474);
and U3065 (N_3065,N_1325,N_10);
and U3066 (N_3066,N_1696,N_1549);
nand U3067 (N_3067,N_1008,N_1416);
xnor U3068 (N_3068,N_1976,N_1610);
xnor U3069 (N_3069,N_2450,N_745);
nand U3070 (N_3070,N_123,N_1241);
and U3071 (N_3071,N_2340,N_1757);
nand U3072 (N_3072,N_1869,N_618);
nand U3073 (N_3073,N_207,N_1534);
and U3074 (N_3074,N_1858,N_1185);
and U3075 (N_3075,N_2362,N_1661);
nand U3076 (N_3076,N_833,N_1647);
nor U3077 (N_3077,N_52,N_2265);
nand U3078 (N_3078,N_1436,N_515);
nor U3079 (N_3079,N_2273,N_1038);
nor U3080 (N_3080,N_990,N_1677);
xor U3081 (N_3081,N_173,N_762);
xnor U3082 (N_3082,N_709,N_2222);
xnor U3083 (N_3083,N_246,N_318);
xnor U3084 (N_3084,N_1962,N_574);
or U3085 (N_3085,N_693,N_2257);
nor U3086 (N_3086,N_601,N_1883);
nor U3087 (N_3087,N_1369,N_1134);
and U3088 (N_3088,N_427,N_351);
or U3089 (N_3089,N_1850,N_1195);
and U3090 (N_3090,N_937,N_568);
nand U3091 (N_3091,N_1370,N_534);
xnor U3092 (N_3092,N_806,N_1277);
nor U3093 (N_3093,N_1563,N_118);
nand U3094 (N_3094,N_1903,N_1123);
and U3095 (N_3095,N_1671,N_1981);
nand U3096 (N_3096,N_1349,N_178);
nand U3097 (N_3097,N_97,N_2101);
nor U3098 (N_3098,N_1073,N_37);
and U3099 (N_3099,N_1655,N_1525);
nor U3100 (N_3100,N_1950,N_856);
nand U3101 (N_3101,N_414,N_1734);
and U3102 (N_3102,N_1524,N_536);
xnor U3103 (N_3103,N_1120,N_352);
nand U3104 (N_3104,N_1214,N_285);
or U3105 (N_3105,N_683,N_2455);
xnor U3106 (N_3106,N_6,N_1774);
xnor U3107 (N_3107,N_988,N_23);
or U3108 (N_3108,N_740,N_531);
nand U3109 (N_3109,N_2414,N_2203);
and U3110 (N_3110,N_2369,N_1520);
nand U3111 (N_3111,N_79,N_2143);
nand U3112 (N_3112,N_1632,N_2323);
nand U3113 (N_3113,N_1636,N_2333);
nand U3114 (N_3114,N_1110,N_134);
nand U3115 (N_3115,N_2157,N_1557);
xor U3116 (N_3116,N_1382,N_694);
and U3117 (N_3117,N_982,N_1403);
xor U3118 (N_3118,N_433,N_1813);
nor U3119 (N_3119,N_239,N_1390);
nor U3120 (N_3120,N_1167,N_1603);
nor U3121 (N_3121,N_1284,N_106);
or U3122 (N_3122,N_277,N_951);
nand U3123 (N_3123,N_857,N_1132);
and U3124 (N_3124,N_1054,N_2145);
and U3125 (N_3125,N_265,N_2479);
nand U3126 (N_3126,N_384,N_1844);
xor U3127 (N_3127,N_148,N_949);
and U3128 (N_3128,N_761,N_1644);
nor U3129 (N_3129,N_2025,N_607);
nand U3130 (N_3130,N_872,N_235);
nor U3131 (N_3131,N_226,N_2171);
xor U3132 (N_3132,N_1128,N_1561);
nand U3133 (N_3133,N_1720,N_2380);
xor U3134 (N_3134,N_98,N_874);
nand U3135 (N_3135,N_930,N_2045);
and U3136 (N_3136,N_139,N_923);
and U3137 (N_3137,N_497,N_1684);
nand U3138 (N_3138,N_465,N_1081);
or U3139 (N_3139,N_1227,N_161);
and U3140 (N_3140,N_325,N_1102);
or U3141 (N_3141,N_1824,N_1484);
or U3142 (N_3142,N_855,N_1726);
xnor U3143 (N_3143,N_1526,N_1901);
and U3144 (N_3144,N_2224,N_797);
nand U3145 (N_3145,N_47,N_2308);
nand U3146 (N_3146,N_2085,N_394);
nand U3147 (N_3147,N_829,N_2298);
nand U3148 (N_3148,N_1129,N_1748);
and U3149 (N_3149,N_1059,N_1864);
nand U3150 (N_3150,N_185,N_1137);
or U3151 (N_3151,N_1828,N_2348);
xor U3152 (N_3152,N_1126,N_1190);
xor U3153 (N_3153,N_455,N_1956);
xor U3154 (N_3154,N_2344,N_315);
xor U3155 (N_3155,N_211,N_1433);
or U3156 (N_3156,N_137,N_879);
and U3157 (N_3157,N_135,N_590);
nand U3158 (N_3158,N_1898,N_1853);
xor U3159 (N_3159,N_1744,N_2054);
nand U3160 (N_3160,N_2077,N_1028);
nor U3161 (N_3161,N_1929,N_2390);
and U3162 (N_3162,N_935,N_517);
nor U3163 (N_3163,N_1210,N_595);
and U3164 (N_3164,N_1628,N_1163);
and U3165 (N_3165,N_1578,N_2112);
and U3166 (N_3166,N_2159,N_1989);
or U3167 (N_3167,N_2043,N_1373);
nor U3168 (N_3168,N_842,N_405);
xor U3169 (N_3169,N_95,N_871);
nor U3170 (N_3170,N_668,N_2262);
nand U3171 (N_3171,N_426,N_125);
nand U3172 (N_3172,N_1421,N_1157);
and U3173 (N_3173,N_1236,N_228);
or U3174 (N_3174,N_1648,N_1829);
nor U3175 (N_3175,N_2374,N_2456);
nand U3176 (N_3176,N_1681,N_1082);
and U3177 (N_3177,N_1366,N_622);
nand U3178 (N_3178,N_1509,N_1814);
xor U3179 (N_3179,N_1303,N_656);
xor U3180 (N_3180,N_99,N_562);
or U3181 (N_3181,N_179,N_909);
and U3182 (N_3182,N_127,N_53);
or U3183 (N_3183,N_1225,N_442);
nor U3184 (N_3184,N_188,N_2046);
nand U3185 (N_3185,N_1127,N_1074);
nand U3186 (N_3186,N_111,N_348);
and U3187 (N_3187,N_341,N_1706);
nor U3188 (N_3188,N_1301,N_508);
nor U3189 (N_3189,N_1667,N_1791);
xor U3190 (N_3190,N_751,N_1442);
nor U3191 (N_3191,N_1119,N_723);
nor U3192 (N_3192,N_77,N_440);
nand U3193 (N_3193,N_195,N_1798);
nor U3194 (N_3194,N_1353,N_980);
nand U3195 (N_3195,N_489,N_496);
and U3196 (N_3196,N_687,N_1050);
nor U3197 (N_3197,N_1861,N_1261);
and U3198 (N_3198,N_2483,N_204);
and U3199 (N_3199,N_2488,N_2420);
nand U3200 (N_3200,N_598,N_583);
nor U3201 (N_3201,N_354,N_1474);
nand U3202 (N_3202,N_924,N_1876);
xnor U3203 (N_3203,N_1023,N_899);
nor U3204 (N_3204,N_1493,N_2080);
xnor U3205 (N_3205,N_1977,N_1711);
and U3206 (N_3206,N_2162,N_1759);
or U3207 (N_3207,N_1890,N_884);
nand U3208 (N_3208,N_363,N_180);
nor U3209 (N_3209,N_963,N_597);
or U3210 (N_3210,N_1823,N_477);
xor U3211 (N_3211,N_1483,N_905);
and U3212 (N_3212,N_241,N_1773);
nor U3213 (N_3213,N_1948,N_907);
or U3214 (N_3214,N_2127,N_2417);
nand U3215 (N_3215,N_2188,N_727);
nor U3216 (N_3216,N_302,N_827);
nand U3217 (N_3217,N_2321,N_214);
nor U3218 (N_3218,N_2288,N_1596);
and U3219 (N_3219,N_51,N_1177);
xnor U3220 (N_3220,N_365,N_1029);
nor U3221 (N_3221,N_1408,N_27);
nor U3222 (N_3222,N_2044,N_2324);
xnor U3223 (N_3223,N_1057,N_1186);
and U3224 (N_3224,N_160,N_2210);
nand U3225 (N_3225,N_215,N_1601);
nor U3226 (N_3226,N_1865,N_2243);
nand U3227 (N_3227,N_2286,N_1099);
xor U3228 (N_3228,N_704,N_753);
nand U3229 (N_3229,N_471,N_358);
nand U3230 (N_3230,N_1996,N_1035);
or U3231 (N_3231,N_1695,N_1259);
or U3232 (N_3232,N_2254,N_29);
and U3233 (N_3233,N_613,N_1516);
nor U3234 (N_3234,N_312,N_1160);
or U3235 (N_3235,N_2314,N_1165);
nor U3236 (N_3236,N_1095,N_1217);
nor U3237 (N_3237,N_665,N_1379);
or U3238 (N_3238,N_541,N_346);
nor U3239 (N_3239,N_151,N_243);
and U3240 (N_3240,N_485,N_576);
nand U3241 (N_3241,N_1532,N_21);
nor U3242 (N_3242,N_1699,N_1013);
nand U3243 (N_3243,N_197,N_2079);
xnor U3244 (N_3244,N_744,N_1297);
nor U3245 (N_3245,N_176,N_801);
or U3246 (N_3246,N_1620,N_2360);
and U3247 (N_3247,N_1514,N_108);
or U3248 (N_3248,N_1877,N_15);
xnor U3249 (N_3249,N_2427,N_1387);
nor U3250 (N_3250,N_614,N_248);
or U3251 (N_3251,N_698,N_301);
nand U3252 (N_3252,N_849,N_184);
xnor U3253 (N_3253,N_2142,N_1820);
xor U3254 (N_3254,N_1063,N_1388);
and U3255 (N_3255,N_205,N_1633);
xor U3256 (N_3256,N_1812,N_798);
and U3257 (N_3257,N_1422,N_1409);
xor U3258 (N_3258,N_929,N_110);
nand U3259 (N_3259,N_928,N_418);
or U3260 (N_3260,N_715,N_519);
nor U3261 (N_3261,N_1257,N_2165);
xor U3262 (N_3262,N_910,N_30);
nand U3263 (N_3263,N_578,N_159);
or U3264 (N_3264,N_2060,N_2134);
nor U3265 (N_3265,N_681,N_646);
nor U3266 (N_3266,N_1306,N_2232);
nand U3267 (N_3267,N_1168,N_2366);
nand U3268 (N_3268,N_712,N_196);
xor U3269 (N_3269,N_1700,N_397);
or U3270 (N_3270,N_1983,N_1540);
xor U3271 (N_3271,N_2436,N_1182);
nor U3272 (N_3272,N_623,N_1053);
nand U3273 (N_3273,N_1736,N_2354);
and U3274 (N_3274,N_995,N_1776);
or U3275 (N_3275,N_168,N_722);
and U3276 (N_3276,N_624,N_817);
or U3277 (N_3277,N_1124,N_2259);
xnor U3278 (N_3278,N_175,N_1076);
nor U3279 (N_3279,N_518,N_1688);
and U3280 (N_3280,N_1581,N_1130);
nor U3281 (N_3281,N_756,N_1606);
and U3282 (N_3282,N_603,N_973);
or U3283 (N_3283,N_1202,N_934);
nor U3284 (N_3284,N_474,N_2347);
xnor U3285 (N_3285,N_1105,N_1909);
nor U3286 (N_3286,N_1113,N_645);
and U3287 (N_3287,N_640,N_35);
or U3288 (N_3288,N_46,N_521);
and U3289 (N_3289,N_2190,N_1789);
nand U3290 (N_3290,N_1924,N_2129);
or U3291 (N_3291,N_1855,N_2481);
nor U3292 (N_3292,N_1964,N_1999);
or U3293 (N_3293,N_2299,N_1871);
or U3294 (N_3294,N_719,N_2156);
nand U3295 (N_3295,N_191,N_1108);
nor U3296 (N_3296,N_682,N_2462);
nor U3297 (N_3297,N_283,N_2204);
xnor U3298 (N_3298,N_505,N_542);
xnor U3299 (N_3299,N_2141,N_691);
xor U3300 (N_3300,N_360,N_25);
nand U3301 (N_3301,N_1611,N_1380);
and U3302 (N_3302,N_1580,N_2042);
or U3303 (N_3303,N_1086,N_2496);
and U3304 (N_3304,N_403,N_1796);
nor U3305 (N_3305,N_322,N_1412);
or U3306 (N_3306,N_281,N_1204);
nand U3307 (N_3307,N_591,N_2395);
nand U3308 (N_3308,N_2400,N_216);
nor U3309 (N_3309,N_2223,N_1170);
or U3310 (N_3310,N_1560,N_664);
xor U3311 (N_3311,N_1863,N_186);
or U3312 (N_3312,N_2476,N_387);
and U3313 (N_3313,N_472,N_1507);
nor U3314 (N_3314,N_206,N_1849);
and U3315 (N_3315,N_1348,N_1917);
or U3316 (N_3316,N_2468,N_2178);
and U3317 (N_3317,N_2103,N_2182);
and U3318 (N_3318,N_1090,N_339);
xor U3319 (N_3319,N_1658,N_1252);
nand U3320 (N_3320,N_308,N_537);
or U3321 (N_3321,N_1140,N_1970);
nor U3322 (N_3322,N_2449,N_1389);
and U3323 (N_3323,N_2448,N_1037);
nor U3324 (N_3324,N_1816,N_1125);
and U3325 (N_3325,N_1852,N_696);
and U3326 (N_3326,N_1078,N_494);
nand U3327 (N_3327,N_136,N_13);
nand U3328 (N_3328,N_950,N_839);
nor U3329 (N_3329,N_1663,N_1292);
nand U3330 (N_3330,N_2432,N_2160);
nor U3331 (N_3331,N_567,N_2038);
or U3332 (N_3332,N_832,N_486);
or U3333 (N_3333,N_927,N_2049);
nor U3334 (N_3334,N_379,N_1025);
xor U3335 (N_3335,N_620,N_2279);
and U3336 (N_3336,N_2353,N_2110);
nor U3337 (N_3337,N_2020,N_1374);
and U3338 (N_3338,N_914,N_1342);
and U3339 (N_3339,N_820,N_759);
or U3340 (N_3340,N_314,N_2271);
and U3341 (N_3341,N_818,N_1069);
nand U3342 (N_3342,N_104,N_1584);
nand U3343 (N_3343,N_2028,N_1175);
nand U3344 (N_3344,N_579,N_1717);
xor U3345 (N_3345,N_699,N_516);
and U3346 (N_3346,N_463,N_498);
and U3347 (N_3347,N_355,N_58);
and U3348 (N_3348,N_2122,N_2115);
and U3349 (N_3349,N_977,N_2309);
xnor U3350 (N_3350,N_711,N_153);
and U3351 (N_3351,N_976,N_2459);
nor U3352 (N_3352,N_252,N_2192);
nor U3353 (N_3353,N_1653,N_105);
or U3354 (N_3354,N_1502,N_16);
xor U3355 (N_3355,N_1363,N_612);
or U3356 (N_3356,N_1332,N_1044);
xor U3357 (N_3357,N_858,N_1615);
nand U3358 (N_3358,N_1451,N_1003);
and U3359 (N_3359,N_632,N_1710);
xnor U3360 (N_3360,N_837,N_932);
nor U3361 (N_3361,N_1383,N_1497);
and U3362 (N_3362,N_969,N_337);
nand U3363 (N_3363,N_94,N_1051);
xor U3364 (N_3364,N_2250,N_1872);
or U3365 (N_3365,N_1056,N_279);
and U3366 (N_3366,N_1543,N_1371);
nor U3367 (N_3367,N_1215,N_1437);
and U3368 (N_3368,N_1490,N_1554);
or U3369 (N_3369,N_2339,N_626);
and U3370 (N_3370,N_271,N_1614);
nand U3371 (N_3371,N_2041,N_788);
nor U3372 (N_3372,N_1041,N_1595);
nand U3373 (N_3373,N_1874,N_1001);
and U3374 (N_3374,N_1435,N_580);
nor U3375 (N_3375,N_765,N_587);
xor U3376 (N_3376,N_1360,N_1091);
nor U3377 (N_3377,N_2047,N_2211);
xnor U3378 (N_3378,N_2399,N_1571);
nand U3379 (N_3379,N_2097,N_754);
xor U3380 (N_3380,N_28,N_78);
nor U3381 (N_3381,N_2056,N_1396);
and U3382 (N_3382,N_2421,N_1907);
xor U3383 (N_3383,N_1203,N_2128);
and U3384 (N_3384,N_169,N_1479);
xor U3385 (N_3385,N_2276,N_1312);
and U3386 (N_3386,N_915,N_846);
xnor U3387 (N_3387,N_840,N_1446);
nand U3388 (N_3388,N_2023,N_1032);
xnor U3389 (N_3389,N_866,N_1766);
nand U3390 (N_3390,N_961,N_499);
nand U3391 (N_3391,N_1646,N_18);
nand U3392 (N_3392,N_2244,N_1808);
nand U3393 (N_3393,N_777,N_1423);
xor U3394 (N_3394,N_1100,N_1792);
or U3395 (N_3395,N_1221,N_1043);
or U3396 (N_3396,N_2055,N_1481);
and U3397 (N_3397,N_1087,N_828);
nor U3398 (N_3398,N_84,N_1900);
nor U3399 (N_3399,N_1391,N_1891);
and U3400 (N_3400,N_2283,N_203);
nand U3401 (N_3401,N_232,N_1733);
xor U3402 (N_3402,N_838,N_2017);
xnor U3403 (N_3403,N_2152,N_245);
xnor U3404 (N_3404,N_606,N_69);
or U3405 (N_3405,N_733,N_491);
xnor U3406 (N_3406,N_2480,N_327);
or U3407 (N_3407,N_1460,N_550);
xor U3408 (N_3408,N_2434,N_392);
nand U3409 (N_3409,N_1229,N_1506);
or U3410 (N_3410,N_2202,N_1309);
nand U3411 (N_3411,N_1842,N_752);
xor U3412 (N_3412,N_2034,N_199);
or U3413 (N_3413,N_88,N_1725);
nor U3414 (N_3414,N_2172,N_2075);
nor U3415 (N_3415,N_2019,N_1618);
nand U3416 (N_3416,N_1042,N_697);
nand U3417 (N_3417,N_2307,N_1260);
nor U3418 (N_3418,N_1945,N_2498);
or U3419 (N_3419,N_2035,N_434);
nor U3420 (N_3420,N_703,N_2409);
nand U3421 (N_3421,N_916,N_275);
nor U3422 (N_3422,N_1026,N_75);
xnor U3423 (N_3423,N_661,N_813);
nand U3424 (N_3424,N_487,N_770);
nand U3425 (N_3425,N_1445,N_182);
nand U3426 (N_3426,N_408,N_1055);
xnor U3427 (N_3427,N_956,N_1893);
and U3428 (N_3428,N_822,N_1558);
nand U3429 (N_3429,N_1207,N_869);
nand U3430 (N_3430,N_523,N_437);
xnor U3431 (N_3431,N_1302,N_1402);
or U3432 (N_3432,N_1918,N_299);
xnor U3433 (N_3433,N_1149,N_2306);
nor U3434 (N_3434,N_1564,N_532);
xor U3435 (N_3435,N_1153,N_264);
nand U3436 (N_3436,N_2382,N_673);
and U3437 (N_3437,N_989,N_1336);
and U3438 (N_3438,N_551,N_1381);
or U3439 (N_3439,N_43,N_684);
and U3440 (N_3440,N_338,N_2439);
nor U3441 (N_3441,N_919,N_1262);
nand U3442 (N_3442,N_457,N_728);
xnor U3443 (N_3443,N_1147,N_1904);
xor U3444 (N_3444,N_227,N_1916);
and U3445 (N_3445,N_458,N_2062);
or U3446 (N_3446,N_944,N_2130);
nor U3447 (N_3447,N_2358,N_2370);
nand U3448 (N_3448,N_1058,N_270);
nor U3449 (N_3449,N_667,N_328);
or U3450 (N_3450,N_446,N_1932);
or U3451 (N_3451,N_1518,N_717);
or U3452 (N_3452,N_144,N_223);
and U3453 (N_3453,N_2083,N_867);
and U3454 (N_3454,N_4,N_2228);
and U3455 (N_3455,N_382,N_1161);
nand U3456 (N_3456,N_2124,N_877);
nand U3457 (N_3457,N_481,N_2088);
xor U3458 (N_3458,N_1533,N_2303);
or U3459 (N_3459,N_38,N_1840);
nand U3460 (N_3460,N_611,N_1346);
nand U3461 (N_3461,N_68,N_2102);
or U3462 (N_3462,N_172,N_406);
nor U3463 (N_3463,N_2241,N_2138);
nand U3464 (N_3464,N_1344,N_2240);
nor U3465 (N_3465,N_1966,N_1299);
and U3466 (N_3466,N_1413,N_1919);
or U3467 (N_3467,N_1785,N_157);
or U3468 (N_3468,N_1319,N_560);
nor U3469 (N_3469,N_2114,N_1197);
or U3470 (N_3470,N_2248,N_19);
xnor U3471 (N_3471,N_2057,N_1394);
nor U3472 (N_3472,N_49,N_685);
xor U3473 (N_3473,N_422,N_1933);
nor U3474 (N_3474,N_979,N_1931);
nand U3475 (N_3475,N_1604,N_2277);
xor U3476 (N_3476,N_621,N_1158);
or U3477 (N_3477,N_2329,N_1004);
nor U3478 (N_3478,N_2201,N_1316);
nand U3479 (N_3479,N_774,N_1151);
xnor U3480 (N_3480,N_61,N_1841);
xnor U3481 (N_3481,N_1769,N_320);
nand U3482 (N_3482,N_1599,N_298);
and U3483 (N_3483,N_121,N_373);
nor U3484 (N_3484,N_834,N_1139);
xor U3485 (N_3485,N_2118,N_2376);
and U3486 (N_3486,N_1537,N_785);
and U3487 (N_3487,N_2186,N_2268);
nor U3488 (N_3488,N_323,N_1268);
xnor U3489 (N_3489,N_1570,N_1061);
or U3490 (N_3490,N_290,N_804);
nor U3491 (N_3491,N_1242,N_896);
xnor U3492 (N_3492,N_156,N_83);
nor U3493 (N_3493,N_158,N_2193);
xnor U3494 (N_3494,N_357,N_815);
or U3495 (N_3495,N_1910,N_251);
nand U3496 (N_3496,N_1122,N_533);
xnor U3497 (N_3497,N_452,N_217);
or U3498 (N_3498,N_1135,N_492);
xnor U3499 (N_3499,N_1492,N_1749);
nor U3500 (N_3500,N_2030,N_799);
nor U3501 (N_3501,N_1915,N_2499);
nor U3502 (N_3502,N_565,N_689);
nand U3503 (N_3503,N_1079,N_1930);
nor U3504 (N_3504,N_453,N_2246);
or U3505 (N_3505,N_852,N_881);
xor U3506 (N_3506,N_107,N_1007);
xnor U3507 (N_3507,N_1010,N_1417);
xnor U3508 (N_3508,N_62,N_2365);
or U3509 (N_3509,N_2351,N_1440);
and U3510 (N_3510,N_401,N_878);
nand U3511 (N_3511,N_2281,N_1198);
nand U3512 (N_3512,N_569,N_1598);
xor U3513 (N_3513,N_430,N_773);
and U3514 (N_3514,N_2447,N_1694);
and U3515 (N_3515,N_2105,N_482);
or U3516 (N_3516,N_1077,N_1856);
nand U3517 (N_3517,N_2117,N_1208);
xor U3518 (N_3518,N_60,N_177);
nor U3519 (N_3519,N_791,N_908);
xor U3520 (N_3520,N_1886,N_1002);
nor U3521 (N_3521,N_1183,N_1978);
or U3522 (N_3522,N_650,N_987);
nand U3523 (N_3523,N_356,N_1927);
nor U3524 (N_3524,N_936,N_1593);
xnor U3525 (N_3525,N_386,N_2231);
nor U3526 (N_3526,N_2198,N_1393);
xnor U3527 (N_3527,N_2341,N_2463);
or U3528 (N_3528,N_2247,N_1768);
nor U3529 (N_3529,N_939,N_1626);
and U3530 (N_3530,N_2108,N_70);
xor U3531 (N_3531,N_1794,N_619);
nor U3532 (N_3532,N_2249,N_970);
nand U3533 (N_3533,N_729,N_194);
nor U3534 (N_3534,N_1591,N_1469);
and U3535 (N_3535,N_1314,N_1172);
xor U3536 (N_3536,N_209,N_2446);
nand U3537 (N_3537,N_1133,N_1708);
xnor U3538 (N_3538,N_383,N_478);
nor U3539 (N_3539,N_700,N_269);
nor U3540 (N_3540,N_396,N_2067);
and U3541 (N_3541,N_2490,N_1683);
nand U3542 (N_3542,N_1690,N_2021);
nor U3543 (N_3543,N_854,N_1892);
nor U3544 (N_3544,N_2213,N_340);
or U3545 (N_3545,N_2377,N_2032);
xnor U3546 (N_3546,N_1801,N_293);
and U3547 (N_3547,N_1141,N_1040);
xnor U3548 (N_3548,N_461,N_2412);
nand U3549 (N_3549,N_1831,N_2295);
nand U3550 (N_3550,N_1780,N_306);
and U3551 (N_3551,N_2413,N_1281);
nand U3552 (N_3552,N_1411,N_1368);
or U3553 (N_3553,N_1218,N_1810);
xnor U3554 (N_3554,N_64,N_1958);
xor U3555 (N_3555,N_1594,N_165);
nand U3556 (N_3556,N_2274,N_233);
and U3557 (N_3557,N_2245,N_1224);
nand U3558 (N_3558,N_1567,N_192);
nor U3559 (N_3559,N_670,N_1352);
xor U3560 (N_3560,N_1476,N_2121);
or U3561 (N_3561,N_674,N_1478);
and U3562 (N_3562,N_404,N_1296);
and U3563 (N_3563,N_2135,N_876);
and U3564 (N_3564,N_1107,N_1772);
nor U3565 (N_3565,N_705,N_2074);
xnor U3566 (N_3566,N_1477,N_766);
xor U3567 (N_3567,N_1439,N_2430);
and U3568 (N_3568,N_307,N_504);
or U3569 (N_3569,N_654,N_1519);
or U3570 (N_3570,N_1758,N_1637);
nor U3571 (N_3571,N_702,N_2454);
xor U3572 (N_3572,N_779,N_1467);
xnor U3573 (N_3573,N_87,N_11);
nor U3574 (N_3574,N_1897,N_459);
xnor U3575 (N_3575,N_898,N_2350);
or U3576 (N_3576,N_2235,N_1184);
xor U3577 (N_3577,N_690,N_1621);
xnor U3578 (N_3578,N_2040,N_1343);
xor U3579 (N_3579,N_162,N_71);
nor U3580 (N_3580,N_407,N_1536);
xor U3581 (N_3581,N_2440,N_292);
or U3582 (N_3582,N_435,N_343);
or U3583 (N_3583,N_1878,N_1799);
nor U3584 (N_3584,N_198,N_1112);
nand U3585 (N_3585,N_873,N_823);
nand U3586 (N_3586,N_2367,N_971);
nor U3587 (N_3587,N_1702,N_133);
xor U3588 (N_3588,N_2491,N_851);
nor U3589 (N_3589,N_1947,N_2253);
nor U3590 (N_3590,N_1651,N_2492);
and U3591 (N_3591,N_311,N_126);
or U3592 (N_3592,N_2425,N_331);
and U3593 (N_3593,N_1881,N_2139);
and U3594 (N_3594,N_1150,N_1553);
or U3595 (N_3595,N_2168,N_475);
xor U3596 (N_3596,N_202,N_1866);
or U3597 (N_3597,N_1612,N_273);
nor U3598 (N_3598,N_1326,N_1722);
nand U3599 (N_3599,N_599,N_885);
and U3600 (N_3600,N_1668,N_863);
nand U3601 (N_3601,N_81,N_1939);
nand U3602 (N_3602,N_1529,N_1952);
nand U3603 (N_3603,N_2048,N_210);
and U3604 (N_3604,N_2497,N_2005);
nor U3605 (N_3605,N_1940,N_1546);
nor U3606 (N_3606,N_1806,N_1206);
nor U3607 (N_3607,N_2342,N_847);
or U3608 (N_3608,N_812,N_326);
and U3609 (N_3609,N_2234,N_1272);
or U3610 (N_3610,N_1579,N_305);
or U3611 (N_3611,N_2322,N_1597);
nand U3612 (N_3612,N_1672,N_1294);
or U3613 (N_3613,N_1942,N_234);
xor U3614 (N_3614,N_1322,N_875);
nor U3615 (N_3615,N_1839,N_577);
nand U3616 (N_3616,N_561,N_1486);
and U3617 (N_3617,N_154,N_1960);
and U3618 (N_3618,N_509,N_240);
or U3619 (N_3619,N_984,N_2238);
nand U3620 (N_3620,N_2304,N_1118);
xor U3621 (N_3621,N_1334,N_1650);
xor U3622 (N_3622,N_1250,N_629);
and U3623 (N_3623,N_1719,N_286);
and U3624 (N_3624,N_1987,N_2009);
xnor U3625 (N_3625,N_377,N_2405);
and U3626 (N_3626,N_2255,N_997);
xor U3627 (N_3627,N_514,N_2140);
or U3628 (N_3628,N_2175,N_1171);
and U3629 (N_3629,N_648,N_1835);
nand U3630 (N_3630,N_2451,N_483);
nor U3631 (N_3631,N_2293,N_142);
nor U3632 (N_3632,N_2364,N_262);
nand U3633 (N_3633,N_1024,N_2493);
nor U3634 (N_3634,N_864,N_921);
or U3635 (N_3635,N_1386,N_1795);
and U3636 (N_3636,N_1420,N_2378);
nor U3637 (N_3637,N_2484,N_1154);
and U3638 (N_3638,N_1707,N_2296);
nor U3639 (N_3639,N_164,N_1181);
nor U3640 (N_3640,N_1030,N_631);
xnor U3641 (N_3641,N_1320,N_390);
nor U3642 (N_3642,N_1665,N_1304);
and U3643 (N_3643,N_2185,N_359);
and U3644 (N_3644,N_1159,N_143);
or U3645 (N_3645,N_2433,N_559);
nand U3646 (N_3646,N_2269,N_374);
and U3647 (N_3647,N_659,N_55);
or U3648 (N_3648,N_122,N_634);
xnor U3649 (N_3649,N_955,N_2219);
and U3650 (N_3650,N_1955,N_447);
or U3651 (N_3651,N_1027,N_1084);
or U3652 (N_3652,N_2477,N_2475);
nand U3653 (N_3653,N_2120,N_1196);
and U3654 (N_3654,N_547,N_2263);
nand U3655 (N_3655,N_349,N_2063);
or U3656 (N_3656,N_484,N_1472);
xnor U3657 (N_3657,N_501,N_146);
and U3658 (N_3658,N_962,N_680);
xnor U3659 (N_3659,N_2453,N_2368);
xnor U3660 (N_3660,N_739,N_2136);
and U3661 (N_3661,N_1339,N_1220);
or U3662 (N_3662,N_1870,N_1698);
nand U3663 (N_3663,N_1066,N_758);
nand U3664 (N_3664,N_946,N_1142);
and U3665 (N_3665,N_2173,N_454);
nand U3666 (N_3666,N_1269,N_1487);
xor U3667 (N_3667,N_510,N_1410);
or U3668 (N_3668,N_31,N_1617);
and U3669 (N_3669,N_114,N_2280);
and U3670 (N_3670,N_73,N_1585);
or U3671 (N_3671,N_2225,N_421);
xor U3672 (N_3672,N_1742,N_549);
xnor U3673 (N_3673,N_2345,N_749);
and U3674 (N_3674,N_1361,N_2086);
xnor U3675 (N_3675,N_1114,N_1345);
and U3676 (N_3676,N_1680,N_566);
or U3677 (N_3677,N_2166,N_525);
nand U3678 (N_3678,N_672,N_2189);
and U3679 (N_3679,N_296,N_2346);
or U3680 (N_3680,N_748,N_1657);
nor U3681 (N_3681,N_174,N_535);
xor U3682 (N_3682,N_33,N_1513);
xnor U3683 (N_3683,N_445,N_218);
nor U3684 (N_3684,N_116,N_100);
and U3685 (N_3685,N_1922,N_2242);
nand U3686 (N_3686,N_1311,N_529);
or U3687 (N_3687,N_276,N_1807);
and U3688 (N_3688,N_1288,N_385);
nand U3689 (N_3689,N_1775,N_1012);
or U3690 (N_3690,N_2327,N_2154);
nor U3691 (N_3691,N_1501,N_1094);
and U3692 (N_3692,N_994,N_45);
nor U3693 (N_3693,N_1678,N_438);
nand U3694 (N_3694,N_2357,N_2393);
xor U3695 (N_3695,N_1666,N_255);
xor U3696 (N_3696,N_44,N_1569);
or U3697 (N_3697,N_1510,N_1515);
or U3698 (N_3698,N_468,N_362);
nor U3699 (N_3699,N_512,N_1088);
nor U3700 (N_3700,N_1096,N_2091);
or U3701 (N_3701,N_166,N_2328);
nor U3702 (N_3702,N_2384,N_2237);
nand U3703 (N_3703,N_1022,N_1704);
or U3704 (N_3704,N_2441,N_2078);
and U3705 (N_3705,N_2301,N_20);
nand U3706 (N_3706,N_1230,N_1625);
xor U3707 (N_3707,N_2133,N_870);
xor U3708 (N_3708,N_1071,N_1638);
or U3709 (N_3709,N_288,N_402);
and U3710 (N_3710,N_658,N_300);
nand U3711 (N_3711,N_1399,N_831);
nor U3712 (N_3712,N_2266,N_1324);
or U3713 (N_3713,N_2003,N_1367);
or U3714 (N_3714,N_1517,N_1800);
and U3715 (N_3715,N_582,N_150);
or U3716 (N_3716,N_2471,N_2137);
nand U3717 (N_3717,N_36,N_1364);
and U3718 (N_3718,N_546,N_975);
and U3719 (N_3719,N_575,N_1819);
or U3720 (N_3720,N_2027,N_1443);
and U3721 (N_3721,N_393,N_1967);
nor U3722 (N_3722,N_2332,N_1724);
xor U3723 (N_3723,N_432,N_713);
or U3724 (N_3724,N_1504,N_12);
and U3725 (N_3725,N_1131,N_666);
nor U3726 (N_3726,N_2092,N_888);
nand U3727 (N_3727,N_757,N_2335);
nand U3728 (N_3728,N_593,N_731);
nor U3729 (N_3729,N_1431,N_1790);
or U3730 (N_3730,N_284,N_2469);
xor U3731 (N_3731,N_710,N_2435);
or U3732 (N_3732,N_1974,N_2386);
xnor U3733 (N_3733,N_2072,N_1834);
nor U3734 (N_3734,N_1714,N_1062);
xor U3735 (N_3735,N_1228,N_364);
xnor U3736 (N_3736,N_268,N_776);
and U3737 (N_3737,N_931,N_2394);
or U3738 (N_3738,N_2487,N_1430);
and U3739 (N_3739,N_1354,N_1899);
nor U3740 (N_3740,N_2070,N_1249);
nor U3741 (N_3741,N_2318,N_653);
and U3742 (N_3742,N_1762,N_1937);
nor U3743 (N_3743,N_960,N_2404);
or U3744 (N_3744,N_2008,N_2006);
or U3745 (N_3745,N_720,N_556);
nand U3746 (N_3746,N_1712,N_2278);
xor U3747 (N_3747,N_1080,N_1189);
or U3748 (N_3748,N_686,N_2416);
and U3749 (N_3749,N_1429,N_2071);
nor U3750 (N_3750,N_850,N_2052);
or U3751 (N_3751,N_802,N_1685);
xnor U3752 (N_3752,N_2206,N_1115);
nand U3753 (N_3753,N_645,N_417);
nand U3754 (N_3754,N_1059,N_2212);
and U3755 (N_3755,N_89,N_1320);
or U3756 (N_3756,N_1390,N_1755);
nand U3757 (N_3757,N_2348,N_647);
and U3758 (N_3758,N_2162,N_297);
nand U3759 (N_3759,N_743,N_675);
and U3760 (N_3760,N_1912,N_1994);
xor U3761 (N_3761,N_955,N_1213);
nor U3762 (N_3762,N_1396,N_902);
xor U3763 (N_3763,N_762,N_1985);
nand U3764 (N_3764,N_2330,N_636);
nor U3765 (N_3765,N_100,N_661);
nand U3766 (N_3766,N_2283,N_122);
xnor U3767 (N_3767,N_1462,N_1232);
nand U3768 (N_3768,N_2335,N_1061);
or U3769 (N_3769,N_2258,N_2363);
xor U3770 (N_3770,N_646,N_344);
or U3771 (N_3771,N_496,N_248);
and U3772 (N_3772,N_1311,N_1505);
nor U3773 (N_3773,N_2208,N_506);
nor U3774 (N_3774,N_1484,N_94);
xor U3775 (N_3775,N_890,N_1107);
nor U3776 (N_3776,N_2300,N_2228);
and U3777 (N_3777,N_2209,N_1355);
nand U3778 (N_3778,N_400,N_1640);
or U3779 (N_3779,N_2186,N_1843);
nand U3780 (N_3780,N_163,N_162);
xor U3781 (N_3781,N_1497,N_1423);
xor U3782 (N_3782,N_1346,N_1058);
nand U3783 (N_3783,N_330,N_634);
nor U3784 (N_3784,N_791,N_1163);
xnor U3785 (N_3785,N_1479,N_2218);
and U3786 (N_3786,N_1206,N_282);
nand U3787 (N_3787,N_27,N_2340);
or U3788 (N_3788,N_277,N_1078);
or U3789 (N_3789,N_2377,N_1953);
xnor U3790 (N_3790,N_479,N_106);
nor U3791 (N_3791,N_490,N_75);
or U3792 (N_3792,N_605,N_1787);
or U3793 (N_3793,N_103,N_823);
and U3794 (N_3794,N_1655,N_2033);
and U3795 (N_3795,N_1030,N_1756);
or U3796 (N_3796,N_917,N_2251);
or U3797 (N_3797,N_453,N_240);
nor U3798 (N_3798,N_1351,N_1850);
and U3799 (N_3799,N_952,N_2008);
nand U3800 (N_3800,N_1102,N_1066);
nand U3801 (N_3801,N_185,N_2185);
nor U3802 (N_3802,N_2107,N_1322);
and U3803 (N_3803,N_1442,N_1018);
xor U3804 (N_3804,N_1669,N_2323);
and U3805 (N_3805,N_663,N_1154);
nand U3806 (N_3806,N_559,N_249);
nand U3807 (N_3807,N_111,N_1652);
and U3808 (N_3808,N_1542,N_898);
nand U3809 (N_3809,N_1515,N_866);
xnor U3810 (N_3810,N_1059,N_2226);
nand U3811 (N_3811,N_623,N_2048);
nand U3812 (N_3812,N_1104,N_516);
and U3813 (N_3813,N_1075,N_2165);
nor U3814 (N_3814,N_583,N_2499);
or U3815 (N_3815,N_2098,N_502);
nor U3816 (N_3816,N_781,N_1924);
and U3817 (N_3817,N_1918,N_1214);
xnor U3818 (N_3818,N_802,N_859);
or U3819 (N_3819,N_74,N_1513);
xor U3820 (N_3820,N_1274,N_545);
xnor U3821 (N_3821,N_2303,N_2121);
nand U3822 (N_3822,N_2092,N_1098);
nand U3823 (N_3823,N_2028,N_1216);
nor U3824 (N_3824,N_1386,N_2126);
nand U3825 (N_3825,N_1546,N_1806);
nand U3826 (N_3826,N_2217,N_2400);
and U3827 (N_3827,N_967,N_1192);
and U3828 (N_3828,N_2350,N_138);
nor U3829 (N_3829,N_654,N_1859);
and U3830 (N_3830,N_1165,N_1336);
nor U3831 (N_3831,N_549,N_2322);
and U3832 (N_3832,N_1909,N_2425);
or U3833 (N_3833,N_2117,N_1648);
xnor U3834 (N_3834,N_682,N_1610);
nor U3835 (N_3835,N_804,N_1338);
nand U3836 (N_3836,N_1095,N_101);
nor U3837 (N_3837,N_49,N_1572);
nand U3838 (N_3838,N_1363,N_573);
or U3839 (N_3839,N_1734,N_2236);
xor U3840 (N_3840,N_2133,N_2026);
nand U3841 (N_3841,N_1023,N_774);
xor U3842 (N_3842,N_733,N_791);
and U3843 (N_3843,N_1976,N_2448);
nor U3844 (N_3844,N_1219,N_130);
or U3845 (N_3845,N_2080,N_76);
and U3846 (N_3846,N_540,N_1820);
or U3847 (N_3847,N_2046,N_1717);
xnor U3848 (N_3848,N_1912,N_1294);
xor U3849 (N_3849,N_355,N_1333);
or U3850 (N_3850,N_2306,N_1156);
and U3851 (N_3851,N_1764,N_393);
nand U3852 (N_3852,N_1272,N_1694);
xor U3853 (N_3853,N_1476,N_1645);
or U3854 (N_3854,N_1638,N_1742);
nor U3855 (N_3855,N_2357,N_2030);
nor U3856 (N_3856,N_1955,N_2042);
nand U3857 (N_3857,N_1712,N_1924);
and U3858 (N_3858,N_1973,N_920);
nor U3859 (N_3859,N_2255,N_664);
nand U3860 (N_3860,N_519,N_1397);
xor U3861 (N_3861,N_483,N_1131);
xor U3862 (N_3862,N_1245,N_338);
or U3863 (N_3863,N_2403,N_2371);
or U3864 (N_3864,N_974,N_821);
xor U3865 (N_3865,N_1975,N_971);
nor U3866 (N_3866,N_59,N_519);
or U3867 (N_3867,N_1017,N_193);
nand U3868 (N_3868,N_1741,N_785);
and U3869 (N_3869,N_2318,N_2139);
xnor U3870 (N_3870,N_984,N_175);
nand U3871 (N_3871,N_2182,N_667);
xnor U3872 (N_3872,N_1468,N_383);
and U3873 (N_3873,N_1248,N_1405);
or U3874 (N_3874,N_2496,N_1066);
and U3875 (N_3875,N_1891,N_500);
xor U3876 (N_3876,N_2228,N_39);
nor U3877 (N_3877,N_1266,N_754);
nand U3878 (N_3878,N_736,N_840);
and U3879 (N_3879,N_581,N_397);
nor U3880 (N_3880,N_1084,N_465);
xnor U3881 (N_3881,N_1846,N_2468);
nor U3882 (N_3882,N_127,N_1470);
xor U3883 (N_3883,N_930,N_1094);
xnor U3884 (N_3884,N_1818,N_154);
nor U3885 (N_3885,N_222,N_287);
and U3886 (N_3886,N_2348,N_60);
xor U3887 (N_3887,N_1241,N_814);
nor U3888 (N_3888,N_73,N_817);
nor U3889 (N_3889,N_1923,N_113);
or U3890 (N_3890,N_443,N_1914);
and U3891 (N_3891,N_1162,N_1904);
or U3892 (N_3892,N_1240,N_1102);
nand U3893 (N_3893,N_654,N_357);
nand U3894 (N_3894,N_1754,N_1163);
xor U3895 (N_3895,N_1310,N_291);
and U3896 (N_3896,N_1193,N_1492);
and U3897 (N_3897,N_275,N_303);
nand U3898 (N_3898,N_1710,N_379);
or U3899 (N_3899,N_647,N_756);
nor U3900 (N_3900,N_1683,N_2314);
nand U3901 (N_3901,N_90,N_506);
or U3902 (N_3902,N_56,N_1423);
xor U3903 (N_3903,N_2125,N_875);
or U3904 (N_3904,N_124,N_1145);
nand U3905 (N_3905,N_116,N_1296);
or U3906 (N_3906,N_2314,N_2368);
xnor U3907 (N_3907,N_1479,N_2014);
nand U3908 (N_3908,N_2022,N_1960);
nor U3909 (N_3909,N_2333,N_365);
nor U3910 (N_3910,N_886,N_2211);
xor U3911 (N_3911,N_987,N_401);
nand U3912 (N_3912,N_1006,N_2028);
nand U3913 (N_3913,N_102,N_160);
nor U3914 (N_3914,N_2150,N_615);
or U3915 (N_3915,N_1254,N_682);
and U3916 (N_3916,N_1170,N_1956);
xor U3917 (N_3917,N_589,N_928);
or U3918 (N_3918,N_1780,N_1976);
and U3919 (N_3919,N_2135,N_403);
nand U3920 (N_3920,N_718,N_1403);
and U3921 (N_3921,N_906,N_472);
xor U3922 (N_3922,N_1993,N_157);
xnor U3923 (N_3923,N_124,N_1800);
xor U3924 (N_3924,N_2001,N_2468);
xnor U3925 (N_3925,N_1253,N_1849);
or U3926 (N_3926,N_2013,N_1006);
or U3927 (N_3927,N_738,N_1412);
nor U3928 (N_3928,N_1944,N_2208);
or U3929 (N_3929,N_527,N_2231);
or U3930 (N_3930,N_943,N_181);
and U3931 (N_3931,N_681,N_1396);
nand U3932 (N_3932,N_55,N_150);
nand U3933 (N_3933,N_524,N_693);
xnor U3934 (N_3934,N_187,N_107);
xnor U3935 (N_3935,N_1893,N_607);
and U3936 (N_3936,N_2239,N_1621);
or U3937 (N_3937,N_1904,N_795);
nor U3938 (N_3938,N_1662,N_788);
xor U3939 (N_3939,N_1478,N_1985);
xor U3940 (N_3940,N_915,N_686);
nand U3941 (N_3941,N_2078,N_1966);
and U3942 (N_3942,N_32,N_2428);
and U3943 (N_3943,N_1601,N_2423);
xor U3944 (N_3944,N_444,N_256);
xor U3945 (N_3945,N_553,N_876);
xnor U3946 (N_3946,N_1046,N_1099);
xnor U3947 (N_3947,N_877,N_2210);
xor U3948 (N_3948,N_1833,N_125);
and U3949 (N_3949,N_1309,N_287);
or U3950 (N_3950,N_2156,N_1346);
and U3951 (N_3951,N_323,N_1449);
nor U3952 (N_3952,N_353,N_609);
nand U3953 (N_3953,N_91,N_1526);
xnor U3954 (N_3954,N_2364,N_2020);
or U3955 (N_3955,N_689,N_210);
nand U3956 (N_3956,N_954,N_271);
nand U3957 (N_3957,N_1092,N_1378);
or U3958 (N_3958,N_1934,N_203);
nand U3959 (N_3959,N_692,N_2204);
xnor U3960 (N_3960,N_227,N_1505);
xnor U3961 (N_3961,N_1901,N_1797);
nand U3962 (N_3962,N_203,N_1104);
or U3963 (N_3963,N_1878,N_1537);
nand U3964 (N_3964,N_754,N_1843);
xnor U3965 (N_3965,N_1839,N_887);
nand U3966 (N_3966,N_760,N_1431);
and U3967 (N_3967,N_1144,N_705);
nand U3968 (N_3968,N_2373,N_219);
or U3969 (N_3969,N_30,N_1987);
and U3970 (N_3970,N_726,N_794);
or U3971 (N_3971,N_695,N_375);
and U3972 (N_3972,N_940,N_1988);
or U3973 (N_3973,N_1006,N_1556);
or U3974 (N_3974,N_431,N_1519);
or U3975 (N_3975,N_1818,N_671);
xor U3976 (N_3976,N_307,N_2314);
or U3977 (N_3977,N_567,N_1047);
nor U3978 (N_3978,N_1523,N_491);
or U3979 (N_3979,N_525,N_1559);
nor U3980 (N_3980,N_507,N_1022);
nor U3981 (N_3981,N_50,N_2170);
and U3982 (N_3982,N_1446,N_393);
xor U3983 (N_3983,N_2066,N_887);
nor U3984 (N_3984,N_2182,N_1570);
and U3985 (N_3985,N_949,N_438);
or U3986 (N_3986,N_760,N_2476);
and U3987 (N_3987,N_1331,N_1760);
nand U3988 (N_3988,N_250,N_1914);
or U3989 (N_3989,N_687,N_1402);
nor U3990 (N_3990,N_437,N_427);
xor U3991 (N_3991,N_2045,N_1347);
nor U3992 (N_3992,N_1902,N_69);
or U3993 (N_3993,N_2153,N_15);
and U3994 (N_3994,N_1296,N_1694);
or U3995 (N_3995,N_1330,N_2065);
nand U3996 (N_3996,N_246,N_1886);
xnor U3997 (N_3997,N_855,N_987);
nor U3998 (N_3998,N_1782,N_277);
nor U3999 (N_3999,N_654,N_1073);
and U4000 (N_4000,N_398,N_1744);
xnor U4001 (N_4001,N_1389,N_139);
nand U4002 (N_4002,N_875,N_2178);
and U4003 (N_4003,N_1745,N_2058);
xnor U4004 (N_4004,N_575,N_854);
and U4005 (N_4005,N_1724,N_694);
nand U4006 (N_4006,N_291,N_657);
xnor U4007 (N_4007,N_1318,N_141);
or U4008 (N_4008,N_2076,N_626);
nand U4009 (N_4009,N_418,N_1478);
nand U4010 (N_4010,N_623,N_262);
nand U4011 (N_4011,N_1077,N_1882);
nor U4012 (N_4012,N_823,N_945);
nand U4013 (N_4013,N_2064,N_350);
nand U4014 (N_4014,N_1726,N_463);
xor U4015 (N_4015,N_2117,N_814);
nor U4016 (N_4016,N_708,N_2151);
nand U4017 (N_4017,N_1297,N_760);
nor U4018 (N_4018,N_926,N_1791);
nor U4019 (N_4019,N_1793,N_384);
and U4020 (N_4020,N_197,N_2134);
xnor U4021 (N_4021,N_1503,N_511);
nand U4022 (N_4022,N_1474,N_1472);
nor U4023 (N_4023,N_2113,N_1770);
or U4024 (N_4024,N_748,N_2478);
xor U4025 (N_4025,N_1797,N_154);
and U4026 (N_4026,N_826,N_679);
xnor U4027 (N_4027,N_372,N_2384);
nand U4028 (N_4028,N_1376,N_2);
nand U4029 (N_4029,N_393,N_350);
or U4030 (N_4030,N_2450,N_584);
nand U4031 (N_4031,N_2110,N_75);
xor U4032 (N_4032,N_1410,N_2396);
nor U4033 (N_4033,N_2366,N_1029);
and U4034 (N_4034,N_184,N_584);
xor U4035 (N_4035,N_1266,N_128);
and U4036 (N_4036,N_398,N_118);
xor U4037 (N_4037,N_587,N_1509);
and U4038 (N_4038,N_2406,N_1530);
nand U4039 (N_4039,N_1501,N_1662);
and U4040 (N_4040,N_78,N_1090);
xor U4041 (N_4041,N_2299,N_2224);
xor U4042 (N_4042,N_741,N_553);
or U4043 (N_4043,N_1701,N_293);
and U4044 (N_4044,N_2202,N_1317);
and U4045 (N_4045,N_240,N_187);
nor U4046 (N_4046,N_11,N_1901);
or U4047 (N_4047,N_2369,N_1187);
and U4048 (N_4048,N_2050,N_746);
nand U4049 (N_4049,N_1727,N_628);
nand U4050 (N_4050,N_1207,N_1771);
xor U4051 (N_4051,N_2219,N_2334);
xor U4052 (N_4052,N_1297,N_2273);
nand U4053 (N_4053,N_1818,N_2097);
or U4054 (N_4054,N_2028,N_208);
and U4055 (N_4055,N_952,N_624);
nor U4056 (N_4056,N_997,N_182);
nand U4057 (N_4057,N_661,N_1109);
xnor U4058 (N_4058,N_240,N_271);
nand U4059 (N_4059,N_2093,N_981);
nand U4060 (N_4060,N_104,N_1473);
xnor U4061 (N_4061,N_969,N_645);
nand U4062 (N_4062,N_656,N_139);
nor U4063 (N_4063,N_19,N_821);
nor U4064 (N_4064,N_1330,N_1430);
xor U4065 (N_4065,N_1155,N_1088);
and U4066 (N_4066,N_1418,N_570);
xnor U4067 (N_4067,N_1185,N_1593);
or U4068 (N_4068,N_1620,N_1273);
xor U4069 (N_4069,N_1455,N_142);
xor U4070 (N_4070,N_1322,N_1937);
and U4071 (N_4071,N_766,N_1891);
or U4072 (N_4072,N_1423,N_1200);
nor U4073 (N_4073,N_102,N_1269);
nand U4074 (N_4074,N_200,N_1392);
nand U4075 (N_4075,N_1845,N_1726);
nor U4076 (N_4076,N_1911,N_893);
or U4077 (N_4077,N_331,N_492);
and U4078 (N_4078,N_618,N_674);
or U4079 (N_4079,N_1798,N_1728);
nand U4080 (N_4080,N_710,N_1420);
nor U4081 (N_4081,N_531,N_1234);
nor U4082 (N_4082,N_1641,N_213);
nand U4083 (N_4083,N_1100,N_707);
nand U4084 (N_4084,N_2111,N_2407);
and U4085 (N_4085,N_2291,N_2369);
and U4086 (N_4086,N_397,N_1435);
xor U4087 (N_4087,N_948,N_1248);
xnor U4088 (N_4088,N_665,N_908);
nand U4089 (N_4089,N_139,N_944);
xnor U4090 (N_4090,N_42,N_1917);
and U4091 (N_4091,N_1520,N_1393);
xor U4092 (N_4092,N_15,N_1941);
or U4093 (N_4093,N_650,N_362);
nand U4094 (N_4094,N_930,N_865);
or U4095 (N_4095,N_1954,N_193);
xor U4096 (N_4096,N_1224,N_541);
nand U4097 (N_4097,N_92,N_974);
and U4098 (N_4098,N_713,N_1495);
xor U4099 (N_4099,N_1078,N_1951);
xnor U4100 (N_4100,N_1606,N_1198);
nand U4101 (N_4101,N_1066,N_1912);
nor U4102 (N_4102,N_1656,N_243);
xnor U4103 (N_4103,N_886,N_834);
nand U4104 (N_4104,N_1971,N_2186);
xnor U4105 (N_4105,N_1692,N_2433);
nand U4106 (N_4106,N_622,N_1970);
nand U4107 (N_4107,N_1968,N_845);
and U4108 (N_4108,N_1261,N_841);
nor U4109 (N_4109,N_1357,N_2107);
nand U4110 (N_4110,N_1420,N_897);
or U4111 (N_4111,N_511,N_497);
and U4112 (N_4112,N_491,N_1314);
and U4113 (N_4113,N_1359,N_2170);
nor U4114 (N_4114,N_1632,N_2111);
nor U4115 (N_4115,N_2282,N_1722);
xnor U4116 (N_4116,N_2210,N_1394);
nand U4117 (N_4117,N_256,N_285);
or U4118 (N_4118,N_1701,N_385);
nand U4119 (N_4119,N_1679,N_140);
xnor U4120 (N_4120,N_1306,N_1337);
and U4121 (N_4121,N_432,N_512);
or U4122 (N_4122,N_1164,N_1682);
and U4123 (N_4123,N_2355,N_623);
or U4124 (N_4124,N_185,N_2174);
or U4125 (N_4125,N_1055,N_521);
or U4126 (N_4126,N_2325,N_646);
or U4127 (N_4127,N_1322,N_189);
or U4128 (N_4128,N_2168,N_101);
or U4129 (N_4129,N_1583,N_2328);
nor U4130 (N_4130,N_2383,N_30);
xnor U4131 (N_4131,N_1363,N_1745);
and U4132 (N_4132,N_3,N_1685);
xnor U4133 (N_4133,N_935,N_1234);
xnor U4134 (N_4134,N_948,N_1813);
xnor U4135 (N_4135,N_2041,N_166);
or U4136 (N_4136,N_431,N_1357);
xnor U4137 (N_4137,N_67,N_1704);
or U4138 (N_4138,N_2004,N_948);
xnor U4139 (N_4139,N_2141,N_2172);
nor U4140 (N_4140,N_1272,N_412);
or U4141 (N_4141,N_803,N_738);
and U4142 (N_4142,N_888,N_2252);
xnor U4143 (N_4143,N_2125,N_194);
nor U4144 (N_4144,N_566,N_2182);
or U4145 (N_4145,N_2443,N_1669);
nor U4146 (N_4146,N_2042,N_207);
and U4147 (N_4147,N_460,N_1794);
xor U4148 (N_4148,N_461,N_1068);
nor U4149 (N_4149,N_1409,N_1490);
and U4150 (N_4150,N_1939,N_1082);
and U4151 (N_4151,N_1912,N_1910);
xnor U4152 (N_4152,N_722,N_1606);
nand U4153 (N_4153,N_2460,N_1782);
nand U4154 (N_4154,N_1921,N_1695);
nor U4155 (N_4155,N_121,N_462);
xnor U4156 (N_4156,N_832,N_2256);
xnor U4157 (N_4157,N_1838,N_1772);
nand U4158 (N_4158,N_2266,N_1695);
xor U4159 (N_4159,N_2473,N_671);
and U4160 (N_4160,N_1753,N_263);
nor U4161 (N_4161,N_67,N_651);
or U4162 (N_4162,N_684,N_1294);
or U4163 (N_4163,N_1396,N_2256);
and U4164 (N_4164,N_2233,N_853);
nor U4165 (N_4165,N_223,N_2347);
xor U4166 (N_4166,N_209,N_1424);
nor U4167 (N_4167,N_875,N_590);
xor U4168 (N_4168,N_1907,N_1946);
nor U4169 (N_4169,N_1392,N_201);
nand U4170 (N_4170,N_1639,N_1745);
and U4171 (N_4171,N_185,N_2325);
and U4172 (N_4172,N_521,N_1058);
nor U4173 (N_4173,N_37,N_256);
nand U4174 (N_4174,N_980,N_1096);
or U4175 (N_4175,N_238,N_1327);
nor U4176 (N_4176,N_667,N_2132);
nor U4177 (N_4177,N_1467,N_756);
and U4178 (N_4178,N_1481,N_1908);
nor U4179 (N_4179,N_1301,N_2311);
nand U4180 (N_4180,N_983,N_1909);
nor U4181 (N_4181,N_2161,N_1768);
nor U4182 (N_4182,N_517,N_406);
nor U4183 (N_4183,N_820,N_1657);
nor U4184 (N_4184,N_1889,N_2140);
nand U4185 (N_4185,N_732,N_44);
nand U4186 (N_4186,N_2451,N_1082);
and U4187 (N_4187,N_503,N_444);
nor U4188 (N_4188,N_323,N_1130);
nor U4189 (N_4189,N_1930,N_1344);
nand U4190 (N_4190,N_1530,N_1809);
and U4191 (N_4191,N_670,N_2477);
or U4192 (N_4192,N_452,N_2181);
and U4193 (N_4193,N_1602,N_913);
and U4194 (N_4194,N_1376,N_2257);
nor U4195 (N_4195,N_1772,N_340);
nor U4196 (N_4196,N_822,N_627);
nor U4197 (N_4197,N_1698,N_730);
nand U4198 (N_4198,N_861,N_331);
or U4199 (N_4199,N_605,N_1327);
and U4200 (N_4200,N_810,N_930);
and U4201 (N_4201,N_2056,N_1691);
and U4202 (N_4202,N_2008,N_364);
nand U4203 (N_4203,N_2051,N_2399);
and U4204 (N_4204,N_38,N_747);
nand U4205 (N_4205,N_2327,N_1512);
or U4206 (N_4206,N_788,N_2388);
nor U4207 (N_4207,N_704,N_1866);
and U4208 (N_4208,N_701,N_1243);
xnor U4209 (N_4209,N_1306,N_1827);
nor U4210 (N_4210,N_1242,N_1660);
or U4211 (N_4211,N_1665,N_926);
and U4212 (N_4212,N_1413,N_1334);
xor U4213 (N_4213,N_2434,N_2124);
xor U4214 (N_4214,N_2465,N_837);
nor U4215 (N_4215,N_1124,N_1563);
xnor U4216 (N_4216,N_203,N_15);
xnor U4217 (N_4217,N_1614,N_898);
or U4218 (N_4218,N_2208,N_633);
xor U4219 (N_4219,N_1194,N_14);
or U4220 (N_4220,N_1326,N_266);
nor U4221 (N_4221,N_1638,N_1450);
or U4222 (N_4222,N_182,N_251);
and U4223 (N_4223,N_569,N_384);
nor U4224 (N_4224,N_2488,N_2038);
xor U4225 (N_4225,N_1311,N_450);
xor U4226 (N_4226,N_2324,N_1838);
nor U4227 (N_4227,N_1611,N_314);
nor U4228 (N_4228,N_2493,N_559);
xor U4229 (N_4229,N_193,N_1636);
or U4230 (N_4230,N_905,N_2149);
and U4231 (N_4231,N_2495,N_694);
nor U4232 (N_4232,N_1819,N_1491);
nor U4233 (N_4233,N_565,N_937);
and U4234 (N_4234,N_1463,N_2446);
nor U4235 (N_4235,N_1256,N_872);
xnor U4236 (N_4236,N_844,N_224);
nor U4237 (N_4237,N_2314,N_2029);
nand U4238 (N_4238,N_491,N_82);
nand U4239 (N_4239,N_677,N_1137);
or U4240 (N_4240,N_1958,N_1528);
nand U4241 (N_4241,N_1691,N_2224);
nand U4242 (N_4242,N_668,N_848);
nand U4243 (N_4243,N_1390,N_1927);
and U4244 (N_4244,N_1366,N_1154);
nand U4245 (N_4245,N_1091,N_493);
nor U4246 (N_4246,N_704,N_1156);
nand U4247 (N_4247,N_766,N_2474);
or U4248 (N_4248,N_521,N_1689);
nand U4249 (N_4249,N_173,N_1110);
nand U4250 (N_4250,N_1702,N_2);
and U4251 (N_4251,N_252,N_1057);
nor U4252 (N_4252,N_111,N_1992);
or U4253 (N_4253,N_589,N_220);
nand U4254 (N_4254,N_1030,N_56);
and U4255 (N_4255,N_1055,N_60);
nor U4256 (N_4256,N_894,N_1920);
nand U4257 (N_4257,N_1191,N_2244);
or U4258 (N_4258,N_1566,N_1636);
nor U4259 (N_4259,N_1021,N_1560);
xnor U4260 (N_4260,N_861,N_922);
or U4261 (N_4261,N_136,N_951);
nand U4262 (N_4262,N_1271,N_210);
nand U4263 (N_4263,N_826,N_1167);
or U4264 (N_4264,N_1676,N_2418);
or U4265 (N_4265,N_1654,N_88);
nand U4266 (N_4266,N_651,N_1313);
nand U4267 (N_4267,N_1075,N_375);
nor U4268 (N_4268,N_253,N_2472);
and U4269 (N_4269,N_236,N_1704);
or U4270 (N_4270,N_1370,N_1540);
and U4271 (N_4271,N_981,N_2051);
or U4272 (N_4272,N_1935,N_2369);
or U4273 (N_4273,N_778,N_326);
nor U4274 (N_4274,N_500,N_1112);
or U4275 (N_4275,N_2214,N_2421);
xor U4276 (N_4276,N_873,N_1198);
nand U4277 (N_4277,N_599,N_2007);
nand U4278 (N_4278,N_213,N_2158);
and U4279 (N_4279,N_1609,N_1899);
and U4280 (N_4280,N_572,N_206);
or U4281 (N_4281,N_2457,N_2160);
and U4282 (N_4282,N_822,N_425);
nor U4283 (N_4283,N_1238,N_451);
or U4284 (N_4284,N_199,N_1850);
xor U4285 (N_4285,N_804,N_1253);
xor U4286 (N_4286,N_628,N_301);
or U4287 (N_4287,N_1171,N_1565);
and U4288 (N_4288,N_1819,N_1889);
xor U4289 (N_4289,N_1545,N_2170);
and U4290 (N_4290,N_1709,N_752);
and U4291 (N_4291,N_1956,N_2159);
and U4292 (N_4292,N_1409,N_1880);
and U4293 (N_4293,N_1989,N_1726);
or U4294 (N_4294,N_1710,N_928);
nor U4295 (N_4295,N_2252,N_1909);
or U4296 (N_4296,N_1901,N_1583);
and U4297 (N_4297,N_2469,N_523);
or U4298 (N_4298,N_2375,N_1105);
and U4299 (N_4299,N_416,N_798);
and U4300 (N_4300,N_2033,N_1659);
xnor U4301 (N_4301,N_1003,N_476);
nand U4302 (N_4302,N_1166,N_1334);
and U4303 (N_4303,N_235,N_1570);
nor U4304 (N_4304,N_1228,N_1154);
or U4305 (N_4305,N_2388,N_642);
or U4306 (N_4306,N_1864,N_1019);
nand U4307 (N_4307,N_1959,N_2424);
nor U4308 (N_4308,N_2152,N_2025);
or U4309 (N_4309,N_1287,N_1434);
nand U4310 (N_4310,N_2178,N_1505);
nor U4311 (N_4311,N_1806,N_2493);
nand U4312 (N_4312,N_2305,N_1368);
xor U4313 (N_4313,N_931,N_1007);
xnor U4314 (N_4314,N_2097,N_453);
xnor U4315 (N_4315,N_204,N_601);
or U4316 (N_4316,N_409,N_1836);
nand U4317 (N_4317,N_2111,N_1744);
or U4318 (N_4318,N_402,N_435);
nor U4319 (N_4319,N_1799,N_1333);
and U4320 (N_4320,N_855,N_1541);
nor U4321 (N_4321,N_1400,N_704);
and U4322 (N_4322,N_145,N_1907);
nand U4323 (N_4323,N_2440,N_1062);
nand U4324 (N_4324,N_121,N_2152);
nand U4325 (N_4325,N_2132,N_2216);
nor U4326 (N_4326,N_1759,N_1812);
nand U4327 (N_4327,N_48,N_1796);
and U4328 (N_4328,N_116,N_1370);
xnor U4329 (N_4329,N_61,N_1583);
nand U4330 (N_4330,N_1361,N_1310);
xnor U4331 (N_4331,N_710,N_1509);
xor U4332 (N_4332,N_1514,N_2416);
or U4333 (N_4333,N_1781,N_1216);
nor U4334 (N_4334,N_252,N_734);
or U4335 (N_4335,N_1136,N_194);
nand U4336 (N_4336,N_493,N_62);
nand U4337 (N_4337,N_1547,N_353);
and U4338 (N_4338,N_404,N_288);
xnor U4339 (N_4339,N_813,N_1035);
xnor U4340 (N_4340,N_374,N_2121);
xor U4341 (N_4341,N_2202,N_380);
or U4342 (N_4342,N_2108,N_1108);
or U4343 (N_4343,N_1014,N_1168);
or U4344 (N_4344,N_2397,N_2190);
xnor U4345 (N_4345,N_1709,N_1351);
nor U4346 (N_4346,N_688,N_2250);
nor U4347 (N_4347,N_509,N_2215);
or U4348 (N_4348,N_817,N_2380);
xor U4349 (N_4349,N_1622,N_1873);
nand U4350 (N_4350,N_936,N_1067);
or U4351 (N_4351,N_482,N_1566);
nand U4352 (N_4352,N_452,N_191);
and U4353 (N_4353,N_1938,N_185);
xnor U4354 (N_4354,N_1022,N_324);
xnor U4355 (N_4355,N_2454,N_85);
nand U4356 (N_4356,N_66,N_273);
or U4357 (N_4357,N_1793,N_988);
nor U4358 (N_4358,N_705,N_1737);
nor U4359 (N_4359,N_2273,N_479);
or U4360 (N_4360,N_1931,N_2485);
nor U4361 (N_4361,N_2094,N_1907);
nor U4362 (N_4362,N_2266,N_2344);
nor U4363 (N_4363,N_154,N_159);
or U4364 (N_4364,N_1264,N_1951);
nor U4365 (N_4365,N_1860,N_1348);
or U4366 (N_4366,N_1648,N_805);
nand U4367 (N_4367,N_1416,N_448);
or U4368 (N_4368,N_1784,N_2196);
nand U4369 (N_4369,N_2043,N_2421);
and U4370 (N_4370,N_897,N_261);
and U4371 (N_4371,N_2470,N_540);
and U4372 (N_4372,N_2050,N_6);
nand U4373 (N_4373,N_466,N_2078);
nor U4374 (N_4374,N_1901,N_966);
and U4375 (N_4375,N_1261,N_2293);
nor U4376 (N_4376,N_407,N_2061);
or U4377 (N_4377,N_759,N_938);
xor U4378 (N_4378,N_2116,N_897);
xor U4379 (N_4379,N_122,N_2244);
or U4380 (N_4380,N_829,N_389);
xor U4381 (N_4381,N_423,N_1938);
and U4382 (N_4382,N_1712,N_1611);
and U4383 (N_4383,N_923,N_1567);
and U4384 (N_4384,N_284,N_503);
xor U4385 (N_4385,N_720,N_2163);
nand U4386 (N_4386,N_1832,N_987);
nor U4387 (N_4387,N_1190,N_652);
or U4388 (N_4388,N_2351,N_1519);
and U4389 (N_4389,N_2008,N_1635);
and U4390 (N_4390,N_970,N_1808);
or U4391 (N_4391,N_1104,N_1218);
nor U4392 (N_4392,N_1612,N_499);
and U4393 (N_4393,N_1726,N_2449);
or U4394 (N_4394,N_6,N_1035);
nand U4395 (N_4395,N_277,N_2024);
xor U4396 (N_4396,N_1107,N_2117);
nor U4397 (N_4397,N_630,N_52);
nand U4398 (N_4398,N_490,N_1498);
nor U4399 (N_4399,N_210,N_109);
nor U4400 (N_4400,N_1888,N_1884);
nand U4401 (N_4401,N_873,N_1586);
and U4402 (N_4402,N_447,N_968);
nand U4403 (N_4403,N_2034,N_2118);
nand U4404 (N_4404,N_1820,N_2030);
and U4405 (N_4405,N_2281,N_2463);
xor U4406 (N_4406,N_1541,N_987);
nor U4407 (N_4407,N_530,N_2181);
nor U4408 (N_4408,N_1500,N_2160);
or U4409 (N_4409,N_1390,N_699);
nor U4410 (N_4410,N_927,N_111);
or U4411 (N_4411,N_1608,N_489);
nand U4412 (N_4412,N_1839,N_1213);
and U4413 (N_4413,N_2058,N_875);
and U4414 (N_4414,N_1565,N_143);
and U4415 (N_4415,N_1802,N_346);
or U4416 (N_4416,N_1681,N_1186);
xor U4417 (N_4417,N_815,N_2268);
nand U4418 (N_4418,N_1122,N_1148);
xnor U4419 (N_4419,N_608,N_2489);
xnor U4420 (N_4420,N_748,N_1121);
xnor U4421 (N_4421,N_1302,N_2419);
and U4422 (N_4422,N_957,N_259);
nor U4423 (N_4423,N_2465,N_1527);
or U4424 (N_4424,N_1557,N_2093);
nand U4425 (N_4425,N_790,N_2418);
nand U4426 (N_4426,N_204,N_18);
nor U4427 (N_4427,N_931,N_1175);
nand U4428 (N_4428,N_1623,N_1129);
nor U4429 (N_4429,N_137,N_798);
xnor U4430 (N_4430,N_885,N_670);
or U4431 (N_4431,N_2104,N_886);
and U4432 (N_4432,N_1159,N_1431);
nand U4433 (N_4433,N_2117,N_146);
nor U4434 (N_4434,N_2151,N_793);
xor U4435 (N_4435,N_137,N_1191);
nand U4436 (N_4436,N_593,N_1056);
xor U4437 (N_4437,N_259,N_1579);
xnor U4438 (N_4438,N_1462,N_1150);
nand U4439 (N_4439,N_1252,N_2028);
and U4440 (N_4440,N_1985,N_697);
and U4441 (N_4441,N_442,N_376);
or U4442 (N_4442,N_7,N_1898);
xor U4443 (N_4443,N_516,N_2272);
or U4444 (N_4444,N_1402,N_865);
nor U4445 (N_4445,N_244,N_778);
or U4446 (N_4446,N_2129,N_683);
nand U4447 (N_4447,N_436,N_942);
nand U4448 (N_4448,N_1726,N_455);
xnor U4449 (N_4449,N_269,N_987);
nand U4450 (N_4450,N_242,N_1081);
nor U4451 (N_4451,N_1144,N_1110);
or U4452 (N_4452,N_2409,N_255);
or U4453 (N_4453,N_2432,N_1925);
or U4454 (N_4454,N_2215,N_1741);
xor U4455 (N_4455,N_630,N_857);
and U4456 (N_4456,N_1490,N_1474);
nand U4457 (N_4457,N_1119,N_1946);
and U4458 (N_4458,N_2385,N_2272);
nand U4459 (N_4459,N_1498,N_1547);
and U4460 (N_4460,N_639,N_847);
nor U4461 (N_4461,N_1996,N_1710);
nand U4462 (N_4462,N_1121,N_712);
xnor U4463 (N_4463,N_1234,N_648);
nand U4464 (N_4464,N_505,N_774);
nor U4465 (N_4465,N_2147,N_2464);
xor U4466 (N_4466,N_2192,N_699);
nand U4467 (N_4467,N_2238,N_186);
or U4468 (N_4468,N_2402,N_1484);
nand U4469 (N_4469,N_1995,N_1893);
xnor U4470 (N_4470,N_689,N_1);
and U4471 (N_4471,N_1546,N_2437);
nor U4472 (N_4472,N_1565,N_87);
and U4473 (N_4473,N_1313,N_392);
xnor U4474 (N_4474,N_1340,N_223);
and U4475 (N_4475,N_166,N_1424);
and U4476 (N_4476,N_1510,N_2291);
nor U4477 (N_4477,N_530,N_324);
nor U4478 (N_4478,N_239,N_2280);
and U4479 (N_4479,N_783,N_2375);
xor U4480 (N_4480,N_691,N_100);
xnor U4481 (N_4481,N_105,N_2379);
and U4482 (N_4482,N_1738,N_488);
nor U4483 (N_4483,N_661,N_348);
nand U4484 (N_4484,N_484,N_591);
xor U4485 (N_4485,N_1566,N_2467);
or U4486 (N_4486,N_2033,N_1322);
and U4487 (N_4487,N_465,N_1997);
xnor U4488 (N_4488,N_2036,N_1599);
or U4489 (N_4489,N_940,N_2160);
and U4490 (N_4490,N_503,N_1191);
and U4491 (N_4491,N_229,N_1257);
and U4492 (N_4492,N_1421,N_381);
nand U4493 (N_4493,N_956,N_230);
nor U4494 (N_4494,N_1886,N_282);
or U4495 (N_4495,N_2048,N_2363);
xnor U4496 (N_4496,N_1327,N_1640);
nor U4497 (N_4497,N_211,N_1418);
xnor U4498 (N_4498,N_1883,N_723);
or U4499 (N_4499,N_461,N_427);
nand U4500 (N_4500,N_1653,N_50);
nor U4501 (N_4501,N_2405,N_86);
nor U4502 (N_4502,N_2229,N_1299);
xor U4503 (N_4503,N_2243,N_220);
or U4504 (N_4504,N_104,N_1649);
or U4505 (N_4505,N_2454,N_386);
and U4506 (N_4506,N_1213,N_1107);
and U4507 (N_4507,N_1572,N_1307);
nor U4508 (N_4508,N_1569,N_251);
or U4509 (N_4509,N_352,N_214);
xnor U4510 (N_4510,N_1363,N_2185);
or U4511 (N_4511,N_1509,N_2465);
and U4512 (N_4512,N_1153,N_697);
and U4513 (N_4513,N_2306,N_1547);
xor U4514 (N_4514,N_856,N_2485);
nand U4515 (N_4515,N_1600,N_826);
xnor U4516 (N_4516,N_699,N_2464);
xnor U4517 (N_4517,N_991,N_378);
or U4518 (N_4518,N_1878,N_1706);
nor U4519 (N_4519,N_1456,N_680);
or U4520 (N_4520,N_1358,N_1349);
nand U4521 (N_4521,N_576,N_632);
nand U4522 (N_4522,N_1914,N_1181);
or U4523 (N_4523,N_2412,N_1265);
nand U4524 (N_4524,N_1328,N_2161);
xor U4525 (N_4525,N_983,N_757);
xor U4526 (N_4526,N_531,N_1161);
nand U4527 (N_4527,N_1487,N_346);
or U4528 (N_4528,N_690,N_290);
and U4529 (N_4529,N_1873,N_453);
nor U4530 (N_4530,N_1923,N_1765);
and U4531 (N_4531,N_1498,N_1831);
xnor U4532 (N_4532,N_1146,N_2362);
nand U4533 (N_4533,N_652,N_38);
or U4534 (N_4534,N_1405,N_2473);
nor U4535 (N_4535,N_712,N_2256);
and U4536 (N_4536,N_2285,N_907);
and U4537 (N_4537,N_370,N_474);
or U4538 (N_4538,N_1839,N_989);
or U4539 (N_4539,N_2465,N_2209);
xor U4540 (N_4540,N_719,N_1763);
nor U4541 (N_4541,N_1697,N_893);
nor U4542 (N_4542,N_603,N_1218);
and U4543 (N_4543,N_194,N_1186);
nor U4544 (N_4544,N_1404,N_1907);
nor U4545 (N_4545,N_2292,N_930);
or U4546 (N_4546,N_1803,N_1316);
nor U4547 (N_4547,N_24,N_1958);
or U4548 (N_4548,N_1987,N_1947);
xnor U4549 (N_4549,N_2497,N_2342);
and U4550 (N_4550,N_225,N_604);
xnor U4551 (N_4551,N_1396,N_2231);
nand U4552 (N_4552,N_508,N_2044);
nand U4553 (N_4553,N_511,N_1679);
nand U4554 (N_4554,N_62,N_1734);
xor U4555 (N_4555,N_1010,N_1337);
nand U4556 (N_4556,N_370,N_1366);
nor U4557 (N_4557,N_673,N_1003);
or U4558 (N_4558,N_2177,N_1877);
nand U4559 (N_4559,N_952,N_385);
and U4560 (N_4560,N_1907,N_1087);
nor U4561 (N_4561,N_2001,N_610);
or U4562 (N_4562,N_1,N_1482);
nand U4563 (N_4563,N_218,N_408);
xor U4564 (N_4564,N_1582,N_1850);
xnor U4565 (N_4565,N_2304,N_1631);
or U4566 (N_4566,N_1545,N_2215);
xor U4567 (N_4567,N_25,N_1303);
or U4568 (N_4568,N_1495,N_39);
nor U4569 (N_4569,N_339,N_1522);
and U4570 (N_4570,N_2214,N_1164);
or U4571 (N_4571,N_2263,N_2425);
nand U4572 (N_4572,N_2492,N_245);
xor U4573 (N_4573,N_783,N_298);
nand U4574 (N_4574,N_1089,N_2201);
nor U4575 (N_4575,N_1792,N_498);
nand U4576 (N_4576,N_663,N_2439);
nand U4577 (N_4577,N_1974,N_801);
nand U4578 (N_4578,N_2094,N_1086);
nor U4579 (N_4579,N_1663,N_2159);
nor U4580 (N_4580,N_1396,N_10);
nand U4581 (N_4581,N_2054,N_217);
and U4582 (N_4582,N_2258,N_1722);
or U4583 (N_4583,N_905,N_1080);
xor U4584 (N_4584,N_800,N_755);
and U4585 (N_4585,N_140,N_2143);
or U4586 (N_4586,N_686,N_751);
xor U4587 (N_4587,N_569,N_2261);
nand U4588 (N_4588,N_460,N_1003);
nand U4589 (N_4589,N_467,N_596);
and U4590 (N_4590,N_1101,N_1464);
and U4591 (N_4591,N_5,N_248);
or U4592 (N_4592,N_2238,N_1643);
nand U4593 (N_4593,N_549,N_2199);
or U4594 (N_4594,N_17,N_8);
and U4595 (N_4595,N_1665,N_1492);
nor U4596 (N_4596,N_614,N_1488);
xor U4597 (N_4597,N_1704,N_775);
and U4598 (N_4598,N_1361,N_364);
xor U4599 (N_4599,N_1887,N_784);
or U4600 (N_4600,N_2014,N_761);
nand U4601 (N_4601,N_720,N_565);
nand U4602 (N_4602,N_199,N_2096);
nor U4603 (N_4603,N_1901,N_1213);
and U4604 (N_4604,N_187,N_1480);
and U4605 (N_4605,N_1087,N_276);
and U4606 (N_4606,N_2396,N_598);
nand U4607 (N_4607,N_1033,N_1691);
and U4608 (N_4608,N_2351,N_2133);
or U4609 (N_4609,N_1566,N_1827);
or U4610 (N_4610,N_217,N_27);
or U4611 (N_4611,N_6,N_2023);
nor U4612 (N_4612,N_1687,N_457);
and U4613 (N_4613,N_939,N_1678);
and U4614 (N_4614,N_1131,N_2341);
or U4615 (N_4615,N_2214,N_2257);
or U4616 (N_4616,N_1577,N_1173);
and U4617 (N_4617,N_1889,N_2205);
xor U4618 (N_4618,N_1017,N_1406);
xnor U4619 (N_4619,N_1473,N_208);
xor U4620 (N_4620,N_2014,N_857);
nand U4621 (N_4621,N_1332,N_1698);
nor U4622 (N_4622,N_1281,N_1404);
nand U4623 (N_4623,N_1198,N_298);
nor U4624 (N_4624,N_2499,N_395);
nor U4625 (N_4625,N_2413,N_621);
xor U4626 (N_4626,N_160,N_701);
or U4627 (N_4627,N_1422,N_1538);
nor U4628 (N_4628,N_156,N_1031);
xnor U4629 (N_4629,N_34,N_981);
nand U4630 (N_4630,N_1545,N_1506);
or U4631 (N_4631,N_1140,N_764);
nand U4632 (N_4632,N_965,N_583);
and U4633 (N_4633,N_1918,N_1386);
nand U4634 (N_4634,N_145,N_711);
or U4635 (N_4635,N_1530,N_2391);
xor U4636 (N_4636,N_2108,N_1382);
nand U4637 (N_4637,N_2356,N_566);
nand U4638 (N_4638,N_387,N_26);
and U4639 (N_4639,N_1537,N_511);
and U4640 (N_4640,N_1816,N_2410);
and U4641 (N_4641,N_1816,N_1036);
nand U4642 (N_4642,N_2423,N_415);
and U4643 (N_4643,N_992,N_1610);
nor U4644 (N_4644,N_972,N_2364);
or U4645 (N_4645,N_974,N_2285);
or U4646 (N_4646,N_1316,N_1477);
xor U4647 (N_4647,N_789,N_1727);
xor U4648 (N_4648,N_149,N_1184);
xnor U4649 (N_4649,N_624,N_250);
and U4650 (N_4650,N_2127,N_264);
and U4651 (N_4651,N_1957,N_1694);
nand U4652 (N_4652,N_331,N_633);
xnor U4653 (N_4653,N_1555,N_1374);
and U4654 (N_4654,N_1471,N_1747);
or U4655 (N_4655,N_1895,N_347);
nor U4656 (N_4656,N_1250,N_1849);
nand U4657 (N_4657,N_1357,N_1522);
nor U4658 (N_4658,N_546,N_1698);
nor U4659 (N_4659,N_63,N_122);
xor U4660 (N_4660,N_962,N_2176);
xnor U4661 (N_4661,N_891,N_998);
xor U4662 (N_4662,N_1879,N_2020);
nor U4663 (N_4663,N_364,N_233);
nor U4664 (N_4664,N_568,N_2082);
or U4665 (N_4665,N_2486,N_1413);
nor U4666 (N_4666,N_1243,N_2019);
xnor U4667 (N_4667,N_1815,N_837);
or U4668 (N_4668,N_683,N_2051);
xor U4669 (N_4669,N_1900,N_147);
and U4670 (N_4670,N_266,N_1580);
nor U4671 (N_4671,N_1937,N_671);
nor U4672 (N_4672,N_1537,N_1273);
nor U4673 (N_4673,N_1235,N_94);
or U4674 (N_4674,N_238,N_2025);
nand U4675 (N_4675,N_1257,N_1985);
nor U4676 (N_4676,N_1113,N_159);
nor U4677 (N_4677,N_1875,N_994);
nand U4678 (N_4678,N_1110,N_99);
and U4679 (N_4679,N_1795,N_728);
nand U4680 (N_4680,N_1952,N_1811);
nand U4681 (N_4681,N_546,N_1014);
xor U4682 (N_4682,N_2359,N_797);
nand U4683 (N_4683,N_2428,N_2081);
or U4684 (N_4684,N_1909,N_1648);
xor U4685 (N_4685,N_2180,N_403);
nor U4686 (N_4686,N_1028,N_951);
nand U4687 (N_4687,N_148,N_1202);
nand U4688 (N_4688,N_1310,N_2463);
and U4689 (N_4689,N_1276,N_1515);
or U4690 (N_4690,N_1583,N_1945);
nor U4691 (N_4691,N_731,N_213);
xnor U4692 (N_4692,N_1200,N_350);
nor U4693 (N_4693,N_1742,N_1868);
nor U4694 (N_4694,N_2346,N_1314);
nor U4695 (N_4695,N_125,N_755);
xnor U4696 (N_4696,N_1871,N_95);
nor U4697 (N_4697,N_405,N_2152);
or U4698 (N_4698,N_1860,N_562);
or U4699 (N_4699,N_2392,N_7);
or U4700 (N_4700,N_513,N_1894);
nand U4701 (N_4701,N_672,N_405);
nor U4702 (N_4702,N_1975,N_1824);
or U4703 (N_4703,N_1390,N_2344);
nor U4704 (N_4704,N_2074,N_1612);
or U4705 (N_4705,N_384,N_1587);
and U4706 (N_4706,N_1844,N_977);
xor U4707 (N_4707,N_2143,N_434);
and U4708 (N_4708,N_1612,N_110);
and U4709 (N_4709,N_1317,N_2116);
nand U4710 (N_4710,N_365,N_1124);
nand U4711 (N_4711,N_2025,N_2304);
or U4712 (N_4712,N_431,N_2487);
nand U4713 (N_4713,N_1483,N_470);
xor U4714 (N_4714,N_1389,N_2353);
nor U4715 (N_4715,N_307,N_2092);
nor U4716 (N_4716,N_1569,N_1159);
xnor U4717 (N_4717,N_1900,N_1294);
and U4718 (N_4718,N_56,N_2287);
xor U4719 (N_4719,N_1422,N_567);
nor U4720 (N_4720,N_563,N_931);
and U4721 (N_4721,N_126,N_479);
and U4722 (N_4722,N_140,N_277);
or U4723 (N_4723,N_687,N_2451);
nand U4724 (N_4724,N_1705,N_445);
xnor U4725 (N_4725,N_909,N_351);
nand U4726 (N_4726,N_1961,N_1043);
nand U4727 (N_4727,N_686,N_209);
xor U4728 (N_4728,N_1916,N_1786);
nor U4729 (N_4729,N_709,N_2346);
nand U4730 (N_4730,N_2244,N_2218);
xor U4731 (N_4731,N_1759,N_1343);
nand U4732 (N_4732,N_1895,N_1217);
or U4733 (N_4733,N_1006,N_1898);
nand U4734 (N_4734,N_499,N_1957);
or U4735 (N_4735,N_379,N_1001);
xor U4736 (N_4736,N_1897,N_1433);
nand U4737 (N_4737,N_422,N_33);
nand U4738 (N_4738,N_2288,N_1881);
nand U4739 (N_4739,N_1268,N_383);
nand U4740 (N_4740,N_54,N_241);
xor U4741 (N_4741,N_1470,N_467);
and U4742 (N_4742,N_1480,N_1255);
and U4743 (N_4743,N_1263,N_313);
or U4744 (N_4744,N_2285,N_176);
xor U4745 (N_4745,N_1665,N_1708);
or U4746 (N_4746,N_1874,N_1586);
xnor U4747 (N_4747,N_586,N_1538);
or U4748 (N_4748,N_363,N_1470);
nand U4749 (N_4749,N_885,N_234);
nor U4750 (N_4750,N_501,N_373);
nand U4751 (N_4751,N_1497,N_1549);
or U4752 (N_4752,N_1000,N_1062);
or U4753 (N_4753,N_211,N_1036);
nand U4754 (N_4754,N_825,N_941);
nor U4755 (N_4755,N_77,N_2329);
nor U4756 (N_4756,N_804,N_1982);
nor U4757 (N_4757,N_2487,N_814);
xor U4758 (N_4758,N_1772,N_1677);
nand U4759 (N_4759,N_2316,N_2260);
and U4760 (N_4760,N_1629,N_1207);
nand U4761 (N_4761,N_639,N_1411);
nand U4762 (N_4762,N_240,N_892);
nor U4763 (N_4763,N_1288,N_786);
nand U4764 (N_4764,N_2104,N_2315);
or U4765 (N_4765,N_1018,N_2192);
or U4766 (N_4766,N_1837,N_1624);
nand U4767 (N_4767,N_522,N_2252);
xor U4768 (N_4768,N_1376,N_2465);
nand U4769 (N_4769,N_197,N_2415);
xor U4770 (N_4770,N_1429,N_887);
nand U4771 (N_4771,N_1952,N_950);
and U4772 (N_4772,N_1114,N_197);
nand U4773 (N_4773,N_1566,N_512);
nand U4774 (N_4774,N_1134,N_830);
xnor U4775 (N_4775,N_2269,N_2225);
and U4776 (N_4776,N_1464,N_98);
and U4777 (N_4777,N_1673,N_1038);
and U4778 (N_4778,N_1393,N_2448);
nand U4779 (N_4779,N_429,N_2439);
nor U4780 (N_4780,N_1331,N_999);
xor U4781 (N_4781,N_928,N_1346);
or U4782 (N_4782,N_627,N_1228);
nor U4783 (N_4783,N_2032,N_1407);
or U4784 (N_4784,N_1713,N_2487);
xnor U4785 (N_4785,N_1491,N_1975);
or U4786 (N_4786,N_2432,N_1421);
nor U4787 (N_4787,N_458,N_914);
or U4788 (N_4788,N_109,N_1910);
and U4789 (N_4789,N_2046,N_2445);
or U4790 (N_4790,N_1818,N_1982);
xnor U4791 (N_4791,N_203,N_2472);
nor U4792 (N_4792,N_606,N_1502);
or U4793 (N_4793,N_2248,N_2258);
xor U4794 (N_4794,N_1465,N_1047);
nand U4795 (N_4795,N_525,N_2491);
nor U4796 (N_4796,N_129,N_1534);
xnor U4797 (N_4797,N_173,N_1231);
or U4798 (N_4798,N_198,N_2011);
or U4799 (N_4799,N_1218,N_1936);
or U4800 (N_4800,N_1754,N_224);
nand U4801 (N_4801,N_143,N_653);
or U4802 (N_4802,N_1368,N_2130);
nor U4803 (N_4803,N_998,N_488);
and U4804 (N_4804,N_2179,N_1796);
nor U4805 (N_4805,N_2256,N_1156);
xnor U4806 (N_4806,N_11,N_1091);
nand U4807 (N_4807,N_1555,N_394);
and U4808 (N_4808,N_171,N_2215);
xor U4809 (N_4809,N_2375,N_181);
nor U4810 (N_4810,N_2358,N_1593);
xor U4811 (N_4811,N_2394,N_1467);
nand U4812 (N_4812,N_1422,N_2081);
or U4813 (N_4813,N_1899,N_450);
or U4814 (N_4814,N_1402,N_260);
and U4815 (N_4815,N_1120,N_2324);
nand U4816 (N_4816,N_1039,N_498);
or U4817 (N_4817,N_2318,N_956);
nand U4818 (N_4818,N_2174,N_1230);
nor U4819 (N_4819,N_433,N_1624);
nor U4820 (N_4820,N_2190,N_2300);
or U4821 (N_4821,N_383,N_1050);
and U4822 (N_4822,N_611,N_1179);
or U4823 (N_4823,N_723,N_261);
nor U4824 (N_4824,N_2015,N_1536);
and U4825 (N_4825,N_2087,N_2025);
nor U4826 (N_4826,N_354,N_730);
and U4827 (N_4827,N_676,N_1108);
nand U4828 (N_4828,N_1452,N_1168);
or U4829 (N_4829,N_143,N_103);
and U4830 (N_4830,N_2362,N_1878);
and U4831 (N_4831,N_1543,N_258);
and U4832 (N_4832,N_1178,N_1880);
nand U4833 (N_4833,N_715,N_1566);
nor U4834 (N_4834,N_1553,N_896);
and U4835 (N_4835,N_274,N_1773);
nand U4836 (N_4836,N_242,N_1636);
or U4837 (N_4837,N_985,N_56);
nor U4838 (N_4838,N_2061,N_1807);
nor U4839 (N_4839,N_1174,N_1309);
or U4840 (N_4840,N_2216,N_289);
nand U4841 (N_4841,N_211,N_2078);
nand U4842 (N_4842,N_2309,N_2354);
and U4843 (N_4843,N_2065,N_1973);
xor U4844 (N_4844,N_967,N_400);
nand U4845 (N_4845,N_1802,N_1461);
xnor U4846 (N_4846,N_453,N_1154);
xnor U4847 (N_4847,N_161,N_762);
nor U4848 (N_4848,N_221,N_1774);
nor U4849 (N_4849,N_1399,N_1905);
nand U4850 (N_4850,N_1382,N_1140);
or U4851 (N_4851,N_1101,N_706);
xor U4852 (N_4852,N_975,N_1997);
xnor U4853 (N_4853,N_509,N_70);
xor U4854 (N_4854,N_1425,N_987);
or U4855 (N_4855,N_759,N_1370);
nor U4856 (N_4856,N_1184,N_1781);
or U4857 (N_4857,N_469,N_1650);
and U4858 (N_4858,N_466,N_1932);
nor U4859 (N_4859,N_2295,N_1275);
or U4860 (N_4860,N_1068,N_2139);
nor U4861 (N_4861,N_653,N_1675);
nor U4862 (N_4862,N_888,N_1308);
nor U4863 (N_4863,N_206,N_2123);
or U4864 (N_4864,N_2313,N_8);
xor U4865 (N_4865,N_200,N_509);
nor U4866 (N_4866,N_2016,N_584);
nand U4867 (N_4867,N_900,N_1313);
xor U4868 (N_4868,N_2486,N_1893);
nor U4869 (N_4869,N_532,N_369);
nor U4870 (N_4870,N_191,N_1110);
or U4871 (N_4871,N_2296,N_1581);
and U4872 (N_4872,N_1357,N_970);
xor U4873 (N_4873,N_1048,N_93);
nand U4874 (N_4874,N_1035,N_1005);
nor U4875 (N_4875,N_207,N_1444);
and U4876 (N_4876,N_610,N_1123);
or U4877 (N_4877,N_1962,N_2190);
nand U4878 (N_4878,N_312,N_1435);
nand U4879 (N_4879,N_266,N_403);
and U4880 (N_4880,N_418,N_1827);
nand U4881 (N_4881,N_1407,N_262);
nor U4882 (N_4882,N_821,N_2370);
nor U4883 (N_4883,N_643,N_521);
xnor U4884 (N_4884,N_1387,N_250);
and U4885 (N_4885,N_1263,N_129);
xnor U4886 (N_4886,N_2108,N_1806);
nor U4887 (N_4887,N_2180,N_1395);
xor U4888 (N_4888,N_2284,N_589);
nand U4889 (N_4889,N_317,N_1986);
nor U4890 (N_4890,N_1810,N_484);
nor U4891 (N_4891,N_965,N_1699);
or U4892 (N_4892,N_2084,N_1995);
nor U4893 (N_4893,N_1320,N_2235);
and U4894 (N_4894,N_161,N_918);
nor U4895 (N_4895,N_2115,N_404);
xor U4896 (N_4896,N_1484,N_1364);
xnor U4897 (N_4897,N_22,N_2119);
or U4898 (N_4898,N_494,N_1376);
nor U4899 (N_4899,N_846,N_2126);
nor U4900 (N_4900,N_25,N_2247);
nand U4901 (N_4901,N_2385,N_805);
xnor U4902 (N_4902,N_997,N_1996);
or U4903 (N_4903,N_1466,N_1278);
xnor U4904 (N_4904,N_1125,N_2390);
or U4905 (N_4905,N_2074,N_1428);
nand U4906 (N_4906,N_578,N_1150);
nand U4907 (N_4907,N_228,N_1114);
xnor U4908 (N_4908,N_4,N_1405);
and U4909 (N_4909,N_34,N_1413);
and U4910 (N_4910,N_408,N_2477);
or U4911 (N_4911,N_1254,N_2077);
and U4912 (N_4912,N_2190,N_1223);
nand U4913 (N_4913,N_1524,N_2085);
nand U4914 (N_4914,N_683,N_2066);
nand U4915 (N_4915,N_2034,N_1677);
nand U4916 (N_4916,N_199,N_337);
nor U4917 (N_4917,N_1016,N_1018);
or U4918 (N_4918,N_152,N_1491);
or U4919 (N_4919,N_1723,N_1081);
nor U4920 (N_4920,N_275,N_1126);
nor U4921 (N_4921,N_2284,N_853);
nand U4922 (N_4922,N_796,N_669);
xor U4923 (N_4923,N_1974,N_277);
nand U4924 (N_4924,N_1852,N_1611);
or U4925 (N_4925,N_2181,N_1355);
nor U4926 (N_4926,N_2189,N_233);
and U4927 (N_4927,N_1929,N_1842);
xnor U4928 (N_4928,N_834,N_1958);
or U4929 (N_4929,N_22,N_1562);
or U4930 (N_4930,N_542,N_1039);
or U4931 (N_4931,N_2447,N_1453);
xor U4932 (N_4932,N_2124,N_226);
and U4933 (N_4933,N_651,N_1854);
xor U4934 (N_4934,N_1060,N_1387);
xor U4935 (N_4935,N_218,N_1665);
nand U4936 (N_4936,N_1203,N_2292);
xnor U4937 (N_4937,N_1223,N_152);
nand U4938 (N_4938,N_1228,N_1725);
xor U4939 (N_4939,N_1484,N_1709);
and U4940 (N_4940,N_716,N_1667);
nor U4941 (N_4941,N_1982,N_322);
xnor U4942 (N_4942,N_2100,N_322);
xor U4943 (N_4943,N_1255,N_235);
and U4944 (N_4944,N_1365,N_587);
nand U4945 (N_4945,N_1219,N_2461);
nor U4946 (N_4946,N_1011,N_17);
nand U4947 (N_4947,N_709,N_697);
nand U4948 (N_4948,N_1504,N_1814);
xnor U4949 (N_4949,N_1092,N_2052);
or U4950 (N_4950,N_122,N_1994);
nor U4951 (N_4951,N_165,N_2223);
nor U4952 (N_4952,N_1007,N_763);
or U4953 (N_4953,N_595,N_2081);
and U4954 (N_4954,N_1903,N_582);
nand U4955 (N_4955,N_150,N_1240);
nor U4956 (N_4956,N_622,N_2166);
and U4957 (N_4957,N_1249,N_1866);
nand U4958 (N_4958,N_1302,N_1635);
and U4959 (N_4959,N_2477,N_1635);
or U4960 (N_4960,N_922,N_299);
nor U4961 (N_4961,N_465,N_521);
nand U4962 (N_4962,N_490,N_2390);
nor U4963 (N_4963,N_2498,N_756);
xor U4964 (N_4964,N_1761,N_1234);
nand U4965 (N_4965,N_1398,N_1088);
or U4966 (N_4966,N_2468,N_1327);
or U4967 (N_4967,N_1559,N_259);
or U4968 (N_4968,N_424,N_313);
and U4969 (N_4969,N_2311,N_1499);
nand U4970 (N_4970,N_1880,N_1265);
nor U4971 (N_4971,N_2498,N_1201);
or U4972 (N_4972,N_1447,N_1541);
xnor U4973 (N_4973,N_702,N_1994);
or U4974 (N_4974,N_1144,N_1646);
or U4975 (N_4975,N_2142,N_553);
xnor U4976 (N_4976,N_2461,N_1);
or U4977 (N_4977,N_2302,N_450);
or U4978 (N_4978,N_896,N_2210);
and U4979 (N_4979,N_2273,N_2090);
nor U4980 (N_4980,N_921,N_805);
nor U4981 (N_4981,N_1977,N_81);
nand U4982 (N_4982,N_210,N_2477);
xnor U4983 (N_4983,N_1013,N_913);
and U4984 (N_4984,N_1230,N_698);
or U4985 (N_4985,N_1791,N_2068);
nor U4986 (N_4986,N_997,N_1402);
nor U4987 (N_4987,N_10,N_1678);
nand U4988 (N_4988,N_787,N_515);
and U4989 (N_4989,N_2357,N_1783);
xnor U4990 (N_4990,N_805,N_326);
and U4991 (N_4991,N_188,N_1096);
or U4992 (N_4992,N_1275,N_969);
and U4993 (N_4993,N_1670,N_2078);
and U4994 (N_4994,N_2476,N_644);
or U4995 (N_4995,N_1259,N_2395);
or U4996 (N_4996,N_1288,N_935);
nand U4997 (N_4997,N_1010,N_1639);
or U4998 (N_4998,N_2038,N_1789);
nand U4999 (N_4999,N_28,N_981);
xnor U5000 (N_5000,N_3844,N_4722);
nor U5001 (N_5001,N_3052,N_2847);
nand U5002 (N_5002,N_3022,N_4709);
and U5003 (N_5003,N_4477,N_4531);
or U5004 (N_5004,N_2964,N_3036);
xor U5005 (N_5005,N_3965,N_4365);
xor U5006 (N_5006,N_4987,N_4756);
and U5007 (N_5007,N_3862,N_3067);
or U5008 (N_5008,N_4530,N_2939);
or U5009 (N_5009,N_3251,N_4809);
or U5010 (N_5010,N_3684,N_2543);
nand U5011 (N_5011,N_4579,N_3248);
xor U5012 (N_5012,N_3742,N_4986);
xor U5013 (N_5013,N_4710,N_3352);
nand U5014 (N_5014,N_3317,N_4187);
and U5015 (N_5015,N_4868,N_3370);
xnor U5016 (N_5016,N_4397,N_3705);
and U5017 (N_5017,N_3641,N_4604);
xor U5018 (N_5018,N_4570,N_4832);
nor U5019 (N_5019,N_4626,N_3518);
xnor U5020 (N_5020,N_2871,N_4129);
nor U5021 (N_5021,N_2639,N_4552);
nand U5022 (N_5022,N_2647,N_2644);
nor U5023 (N_5023,N_4931,N_3607);
xnor U5024 (N_5024,N_4482,N_3743);
xor U5025 (N_5025,N_3362,N_3791);
nand U5026 (N_5026,N_4313,N_3861);
nor U5027 (N_5027,N_4914,N_2777);
nand U5028 (N_5028,N_3343,N_2584);
or U5029 (N_5029,N_4069,N_4301);
nor U5030 (N_5030,N_2548,N_3212);
nand U5031 (N_5031,N_3000,N_3615);
nor U5032 (N_5032,N_2841,N_4864);
nand U5033 (N_5033,N_4408,N_3787);
xor U5034 (N_5034,N_3383,N_4022);
nor U5035 (N_5035,N_3957,N_4012);
nand U5036 (N_5036,N_4291,N_4984);
and U5037 (N_5037,N_2505,N_3735);
xor U5038 (N_5038,N_4102,N_3007);
or U5039 (N_5039,N_4370,N_3860);
nor U5040 (N_5040,N_4594,N_3297);
or U5041 (N_5041,N_4638,N_3775);
xnor U5042 (N_5042,N_2982,N_4972);
nand U5043 (N_5043,N_3665,N_2558);
nand U5044 (N_5044,N_4259,N_3407);
or U5045 (N_5045,N_4352,N_4598);
xnor U5046 (N_5046,N_3188,N_4556);
or U5047 (N_5047,N_4091,N_3652);
and U5048 (N_5048,N_3525,N_4215);
xnor U5049 (N_5049,N_2627,N_4835);
xor U5050 (N_5050,N_4608,N_3601);
xor U5051 (N_5051,N_4532,N_3654);
and U5052 (N_5052,N_2878,N_3139);
nor U5053 (N_5053,N_2973,N_4305);
xor U5054 (N_5054,N_2530,N_3121);
nand U5055 (N_5055,N_3475,N_3260);
nor U5056 (N_5056,N_3392,N_4980);
nor U5057 (N_5057,N_3995,N_2771);
and U5058 (N_5058,N_3226,N_4618);
and U5059 (N_5059,N_3398,N_3667);
nand U5060 (N_5060,N_3024,N_4188);
nand U5061 (N_5061,N_3659,N_4077);
xor U5062 (N_5062,N_4386,N_4090);
nand U5063 (N_5063,N_4228,N_3267);
and U5064 (N_5064,N_3298,N_2793);
and U5065 (N_5065,N_3907,N_3394);
xnor U5066 (N_5066,N_4302,N_4669);
xnor U5067 (N_5067,N_4210,N_4330);
nor U5068 (N_5068,N_4032,N_4013);
or U5069 (N_5069,N_3959,N_4031);
xor U5070 (N_5070,N_3470,N_2708);
nor U5071 (N_5071,N_2974,N_4534);
xor U5072 (N_5072,N_3945,N_3540);
nand U5073 (N_5073,N_3090,N_4250);
nor U5074 (N_5074,N_4150,N_2534);
nor U5075 (N_5075,N_4285,N_2523);
xnor U5076 (N_5076,N_4272,N_4586);
nor U5077 (N_5077,N_2821,N_4391);
and U5078 (N_5078,N_3771,N_4175);
and U5079 (N_5079,N_3115,N_2660);
nor U5080 (N_5080,N_3837,N_3277);
nor U5081 (N_5081,N_4645,N_4702);
and U5082 (N_5082,N_4019,N_3127);
or U5083 (N_5083,N_2870,N_3678);
nand U5084 (N_5084,N_2780,N_4548);
nand U5085 (N_5085,N_3094,N_3190);
xnor U5086 (N_5086,N_3523,N_2752);
xor U5087 (N_5087,N_3363,N_2633);
or U5088 (N_5088,N_4288,N_4425);
and U5089 (N_5089,N_3335,N_3967);
nand U5090 (N_5090,N_3295,N_3627);
or U5091 (N_5091,N_2667,N_3878);
or U5092 (N_5092,N_3016,N_3818);
or U5093 (N_5093,N_2642,N_3309);
nand U5094 (N_5094,N_2938,N_4078);
and U5095 (N_5095,N_2989,N_4520);
and U5096 (N_5096,N_3199,N_4494);
nor U5097 (N_5097,N_3790,N_2672);
nand U5098 (N_5098,N_4575,N_4084);
nand U5099 (N_5099,N_2836,N_3749);
and U5100 (N_5100,N_2865,N_4427);
and U5101 (N_5101,N_3417,N_4344);
nand U5102 (N_5102,N_4171,N_4884);
nand U5103 (N_5103,N_4178,N_4642);
xor U5104 (N_5104,N_2719,N_3713);
and U5105 (N_5105,N_4267,N_4071);
and U5106 (N_5106,N_4591,N_4599);
nor U5107 (N_5107,N_4453,N_4802);
and U5108 (N_5108,N_3934,N_3474);
nor U5109 (N_5109,N_2741,N_3689);
xnor U5110 (N_5110,N_2869,N_2852);
nor U5111 (N_5111,N_2882,N_4717);
and U5112 (N_5112,N_2967,N_3874);
nand U5113 (N_5113,N_4002,N_3425);
xnor U5114 (N_5114,N_3906,N_3402);
nand U5115 (N_5115,N_4103,N_3597);
nor U5116 (N_5116,N_2541,N_2568);
nor U5117 (N_5117,N_3501,N_3221);
and U5118 (N_5118,N_4533,N_4962);
or U5119 (N_5119,N_2735,N_2886);
nand U5120 (N_5120,N_2892,N_3952);
xnor U5121 (N_5121,N_4118,N_3073);
or U5122 (N_5122,N_4023,N_3924);
or U5123 (N_5123,N_4412,N_4966);
nand U5124 (N_5124,N_4863,N_4158);
and U5125 (N_5125,N_3881,N_3421);
nor U5126 (N_5126,N_4108,N_3648);
xnor U5127 (N_5127,N_3733,N_3761);
xor U5128 (N_5128,N_2794,N_4892);
nand U5129 (N_5129,N_4908,N_3804);
nor U5130 (N_5130,N_2962,N_3633);
nand U5131 (N_5131,N_4004,N_2686);
xor U5132 (N_5132,N_3075,N_3657);
and U5133 (N_5133,N_4172,N_3991);
xnor U5134 (N_5134,N_3023,N_4732);
nor U5135 (N_5135,N_4311,N_3429);
nand U5136 (N_5136,N_4678,N_2928);
nand U5137 (N_5137,N_4212,N_2643);
or U5138 (N_5138,N_3005,N_4481);
xnor U5139 (N_5139,N_4584,N_3579);
nor U5140 (N_5140,N_2858,N_4195);
nand U5141 (N_5141,N_4409,N_4848);
xor U5142 (N_5142,N_4493,N_4491);
xor U5143 (N_5143,N_4997,N_4774);
nor U5144 (N_5144,N_3949,N_4364);
nand U5145 (N_5145,N_2900,N_4658);
and U5146 (N_5146,N_4429,N_4968);
xnor U5147 (N_5147,N_3119,N_3836);
or U5148 (N_5148,N_3511,N_4255);
nor U5149 (N_5149,N_3165,N_3574);
xnor U5150 (N_5150,N_2727,N_4615);
xnor U5151 (N_5151,N_4437,N_4508);
nand U5152 (N_5152,N_3027,N_2760);
xor U5153 (N_5153,N_4055,N_4740);
nand U5154 (N_5154,N_3903,N_2833);
nand U5155 (N_5155,N_2898,N_4010);
xnor U5156 (N_5156,N_4148,N_2818);
nor U5157 (N_5157,N_3400,N_4219);
xor U5158 (N_5158,N_2516,N_3688);
or U5159 (N_5159,N_4231,N_4957);
and U5160 (N_5160,N_4241,N_4325);
and U5161 (N_5161,N_4112,N_2823);
or U5162 (N_5162,N_4001,N_3643);
nor U5163 (N_5163,N_4380,N_3189);
or U5164 (N_5164,N_2612,N_4300);
or U5165 (N_5165,N_3292,N_4782);
xor U5166 (N_5166,N_2744,N_3035);
xnor U5167 (N_5167,N_4203,N_3063);
or U5168 (N_5168,N_3435,N_4839);
nand U5169 (N_5169,N_4478,N_4003);
xor U5170 (N_5170,N_3405,N_3500);
and U5171 (N_5171,N_2810,N_3453);
xnor U5172 (N_5172,N_4253,N_4788);
nand U5173 (N_5173,N_4854,N_2528);
nor U5174 (N_5174,N_4866,N_2976);
xor U5175 (N_5175,N_4298,N_3782);
or U5176 (N_5176,N_3240,N_4655);
nand U5177 (N_5177,N_4257,N_4544);
nor U5178 (N_5178,N_4551,N_2932);
nand U5179 (N_5179,N_3484,N_4217);
nor U5180 (N_5180,N_4878,N_3043);
xor U5181 (N_5181,N_4941,N_2956);
xnor U5182 (N_5182,N_4064,N_3593);
nand U5183 (N_5183,N_3046,N_4160);
nor U5184 (N_5184,N_4211,N_3485);
and U5185 (N_5185,N_3290,N_4152);
or U5186 (N_5186,N_2666,N_2677);
nand U5187 (N_5187,N_4665,N_2840);
or U5188 (N_5188,N_2606,N_4454);
or U5189 (N_5189,N_3055,N_3704);
or U5190 (N_5190,N_4484,N_2656);
nor U5191 (N_5191,N_3029,N_4214);
xor U5192 (N_5192,N_4810,N_4817);
nor U5193 (N_5193,N_3465,N_3553);
and U5194 (N_5194,N_3685,N_4492);
and U5195 (N_5195,N_3296,N_2637);
and U5196 (N_5196,N_4773,N_3451);
nor U5197 (N_5197,N_2628,N_4335);
xnor U5198 (N_5198,N_3589,N_2854);
nand U5199 (N_5199,N_4646,N_2990);
nor U5200 (N_5200,N_4673,N_2876);
nand U5201 (N_5201,N_3674,N_2911);
nor U5202 (N_5202,N_3867,N_3011);
nand U5203 (N_5203,N_3032,N_2873);
nor U5204 (N_5204,N_3707,N_3879);
nor U5205 (N_5205,N_3087,N_2707);
nor U5206 (N_5206,N_2802,N_4679);
nand U5207 (N_5207,N_4037,N_4222);
nand U5208 (N_5208,N_4807,N_4590);
or U5209 (N_5209,N_4097,N_4252);
or U5210 (N_5210,N_2631,N_3992);
nand U5211 (N_5211,N_3929,N_4913);
nor U5212 (N_5212,N_2515,N_3580);
nor U5213 (N_5213,N_3457,N_2908);
xor U5214 (N_5214,N_4657,N_2977);
or U5215 (N_5215,N_4474,N_3626);
nor U5216 (N_5216,N_2703,N_2893);
nand U5217 (N_5217,N_3086,N_4336);
nand U5218 (N_5218,N_4342,N_3192);
and U5219 (N_5219,N_4648,N_2683);
nand U5220 (N_5220,N_4902,N_3964);
nor U5221 (N_5221,N_4943,N_4378);
xnor U5222 (N_5222,N_3859,N_3077);
xor U5223 (N_5223,N_4053,N_3134);
nor U5224 (N_5224,N_3618,N_3231);
nor U5225 (N_5225,N_4956,N_3869);
nor U5226 (N_5226,N_3532,N_3610);
nand U5227 (N_5227,N_3699,N_3026);
nand U5228 (N_5228,N_4280,N_2694);
nand U5229 (N_5229,N_2815,N_3373);
and U5230 (N_5230,N_2776,N_3458);
nor U5231 (N_5231,N_4376,N_4169);
or U5232 (N_5232,N_3410,N_4467);
and U5233 (N_5233,N_4528,N_2618);
nor U5234 (N_5234,N_4396,N_4703);
and U5235 (N_5235,N_3198,N_4511);
nor U5236 (N_5236,N_2577,N_4200);
xor U5237 (N_5237,N_4652,N_2540);
nor U5238 (N_5238,N_4597,N_3592);
nand U5239 (N_5239,N_2593,N_3197);
nor U5240 (N_5240,N_2688,N_3954);
nor U5241 (N_5241,N_3731,N_3507);
nand U5242 (N_5242,N_3760,N_3960);
xor U5243 (N_5243,N_3982,N_2894);
nand U5244 (N_5244,N_3703,N_3060);
nor U5245 (N_5245,N_3681,N_2529);
nand U5246 (N_5246,N_4881,N_2806);
xor U5247 (N_5247,N_3926,N_3477);
and U5248 (N_5248,N_2653,N_3160);
nand U5249 (N_5249,N_3176,N_3441);
xnor U5250 (N_5250,N_3680,N_2713);
and U5251 (N_5251,N_3144,N_3279);
or U5252 (N_5252,N_2906,N_4547);
or U5253 (N_5253,N_4821,N_3191);
and U5254 (N_5254,N_3811,N_4106);
nand U5255 (N_5255,N_4994,N_3019);
and U5256 (N_5256,N_4314,N_3084);
nand U5257 (N_5257,N_3423,N_2917);
and U5258 (N_5258,N_3840,N_3196);
or U5259 (N_5259,N_2872,N_2820);
and U5260 (N_5260,N_4310,N_3637);
and U5261 (N_5261,N_3428,N_3272);
and U5262 (N_5262,N_2947,N_3720);
nand U5263 (N_5263,N_4056,N_3533);
xor U5264 (N_5264,N_2550,N_2759);
or U5265 (N_5265,N_4517,N_2738);
and U5266 (N_5266,N_4974,N_3630);
nand U5267 (N_5267,N_4113,N_4826);
and U5268 (N_5268,N_3440,N_4025);
or U5269 (N_5269,N_3670,N_4727);
nand U5270 (N_5270,N_4576,N_3033);
nor U5271 (N_5271,N_3752,N_4524);
or U5272 (N_5272,N_3105,N_3694);
xnor U5273 (N_5273,N_2599,N_2791);
and U5274 (N_5274,N_4050,N_3017);
nor U5275 (N_5275,N_2680,N_3085);
and U5276 (N_5276,N_3223,N_3909);
nor U5277 (N_5277,N_2909,N_2749);
nand U5278 (N_5278,N_4070,N_4621);
and U5279 (N_5279,N_3936,N_2664);
nand U5280 (N_5280,N_4379,N_3885);
or U5281 (N_5281,N_2920,N_4539);
nor U5282 (N_5282,N_2551,N_2895);
and U5283 (N_5283,N_4742,N_4185);
or U5284 (N_5284,N_3541,N_3057);
nor U5285 (N_5285,N_4096,N_2506);
nor U5286 (N_5286,N_3535,N_3767);
xor U5287 (N_5287,N_4345,N_3640);
nor U5288 (N_5288,N_3820,N_4985);
nor U5289 (N_5289,N_4327,N_4698);
nand U5290 (N_5290,N_4855,N_4093);
nand U5291 (N_5291,N_3464,N_3166);
xor U5292 (N_5292,N_2996,N_4582);
or U5293 (N_5293,N_3389,N_3887);
nor U5294 (N_5294,N_3886,N_4546);
nor U5295 (N_5295,N_4704,N_2681);
or U5296 (N_5296,N_2740,N_4205);
xor U5297 (N_5297,N_4906,N_3283);
or U5298 (N_5298,N_2991,N_3696);
xnor U5299 (N_5299,N_4870,N_3275);
xor U5300 (N_5300,N_4443,N_3985);
or U5301 (N_5301,N_3493,N_4201);
and U5302 (N_5302,N_4929,N_4693);
nor U5303 (N_5303,N_4353,N_4033);
or U5304 (N_5304,N_4394,N_2696);
and U5305 (N_5305,N_4795,N_3956);
xor U5306 (N_5306,N_4134,N_4476);
or U5307 (N_5307,N_2959,N_3690);
and U5308 (N_5308,N_4721,N_3664);
xor U5309 (N_5309,N_3567,N_4079);
or U5310 (N_5310,N_4373,N_3675);
or U5311 (N_5311,N_3255,N_2834);
nor U5312 (N_5312,N_4877,N_3237);
nor U5313 (N_5313,N_3986,N_3408);
nor U5314 (N_5314,N_2769,N_4293);
nor U5315 (N_5315,N_3012,N_4390);
nand U5316 (N_5316,N_3941,N_4781);
xnor U5317 (N_5317,N_3118,N_3088);
and U5318 (N_5318,N_2746,N_2508);
nor U5319 (N_5319,N_4262,N_3774);
xor U5320 (N_5320,N_3506,N_4515);
or U5321 (N_5321,N_4587,N_3576);
and U5322 (N_5322,N_3748,N_4016);
and U5323 (N_5323,N_3286,N_3747);
nor U5324 (N_5324,N_3289,N_3328);
or U5325 (N_5325,N_2571,N_4470);
nor U5326 (N_5326,N_3128,N_4082);
nor U5327 (N_5327,N_4741,N_3508);
and U5328 (N_5328,N_3209,N_4653);
and U5329 (N_5329,N_2921,N_4447);
nand U5330 (N_5330,N_3438,N_4871);
xor U5331 (N_5331,N_3487,N_4921);
and U5332 (N_5332,N_3801,N_4209);
or U5333 (N_5333,N_4975,N_4847);
xnor U5334 (N_5334,N_3683,N_2957);
nor U5335 (N_5335,N_4923,N_3009);
or U5336 (N_5336,N_3071,N_3880);
or U5337 (N_5337,N_3824,N_4486);
and U5338 (N_5338,N_4705,N_3828);
or U5339 (N_5339,N_3386,N_4308);
nor U5340 (N_5340,N_4242,N_2965);
or U5341 (N_5341,N_4748,N_3489);
nand U5342 (N_5342,N_2796,N_2961);
nor U5343 (N_5343,N_3725,N_3452);
nor U5344 (N_5344,N_4076,N_4468);
nand U5345 (N_5345,N_4808,N_3799);
nor U5346 (N_5346,N_2545,N_3499);
nor U5347 (N_5347,N_3053,N_3894);
nand U5348 (N_5348,N_3572,N_3854);
nand U5349 (N_5349,N_2723,N_4979);
or U5350 (N_5350,N_4651,N_3534);
nor U5351 (N_5351,N_3602,N_3174);
xnor U5352 (N_5352,N_3536,N_2718);
xnor U5353 (N_5353,N_3235,N_3242);
or U5354 (N_5354,N_3784,N_3315);
xnor U5355 (N_5355,N_4020,N_3645);
and U5356 (N_5356,N_4989,N_4284);
nor U5357 (N_5357,N_2853,N_3763);
nand U5358 (N_5358,N_4101,N_4747);
nand U5359 (N_5359,N_4874,N_3401);
xor U5360 (N_5360,N_2654,N_3314);
nand U5361 (N_5361,N_3687,N_4928);
nand U5362 (N_5362,N_3180,N_3918);
nor U5363 (N_5363,N_3716,N_4950);
nor U5364 (N_5364,N_3708,N_3783);
xnor U5365 (N_5365,N_4382,N_3418);
or U5366 (N_5366,N_4662,N_4132);
and U5367 (N_5367,N_4690,N_3575);
nor U5368 (N_5368,N_3817,N_3167);
nor U5369 (N_5369,N_3301,N_4912);
nor U5370 (N_5370,N_3133,N_4700);
nand U5371 (N_5371,N_4381,N_3395);
and U5372 (N_5372,N_4851,N_4512);
nand U5373 (N_5373,N_4945,N_3455);
xor U5374 (N_5374,N_3900,N_4857);
and U5375 (N_5375,N_2502,N_3809);
and U5376 (N_5376,N_2819,N_4341);
xor U5377 (N_5377,N_4392,N_4724);
nand U5378 (N_5378,N_2679,N_2665);
and U5379 (N_5379,N_2983,N_3920);
nor U5380 (N_5380,N_4971,N_4068);
xnor U5381 (N_5381,N_3510,N_3320);
xor U5382 (N_5382,N_3996,N_2509);
nand U5383 (N_5383,N_2620,N_4860);
xnor U5384 (N_5384,N_2586,N_4766);
nand U5385 (N_5385,N_4790,N_3365);
and U5386 (N_5386,N_3195,N_3944);
or U5387 (N_5387,N_3061,N_3788);
or U5388 (N_5388,N_4299,N_4525);
xnor U5389 (N_5389,N_3310,N_4909);
xnor U5390 (N_5390,N_3066,N_4123);
or U5391 (N_5391,N_3529,N_4918);
xor U5392 (N_5392,N_2557,N_4716);
and U5393 (N_5393,N_3897,N_3514);
or U5394 (N_5394,N_2765,N_3110);
nand U5395 (N_5395,N_2597,N_2874);
nor U5396 (N_5396,N_4339,N_2658);
and U5397 (N_5397,N_3865,N_2531);
nand U5398 (N_5398,N_2995,N_3276);
and U5399 (N_5399,N_3014,N_3230);
nor U5400 (N_5400,N_3293,N_2607);
and U5401 (N_5401,N_2579,N_3182);
nand U5402 (N_5402,N_3300,N_4824);
nor U5403 (N_5403,N_2555,N_4351);
and U5404 (N_5404,N_4736,N_4347);
xor U5405 (N_5405,N_4779,N_2725);
or U5406 (N_5406,N_4089,N_4996);
and U5407 (N_5407,N_4275,N_4085);
and U5408 (N_5408,N_2942,N_3851);
nor U5409 (N_5409,N_3768,N_3064);
or U5410 (N_5410,N_4269,N_2785);
nor U5411 (N_5411,N_3635,N_2927);
nor U5412 (N_5412,N_4497,N_4930);
nor U5413 (N_5413,N_3983,N_4965);
or U5414 (N_5414,N_3222,N_2783);
and U5415 (N_5415,N_4751,N_3349);
and U5416 (N_5416,N_3476,N_3562);
or U5417 (N_5417,N_2668,N_4009);
xor U5418 (N_5418,N_3414,N_3432);
or U5419 (N_5419,N_2797,N_3411);
xor U5420 (N_5420,N_3561,N_3096);
nand U5421 (N_5421,N_3829,N_4501);
xor U5422 (N_5422,N_4977,N_3265);
nand U5423 (N_5423,N_3693,N_4610);
nor U5424 (N_5424,N_3107,N_2972);
nand U5425 (N_5425,N_4925,N_4042);
xor U5426 (N_5426,N_4014,N_2559);
xor U5427 (N_5427,N_2649,N_4385);
nor U5428 (N_5428,N_3890,N_2761);
and U5429 (N_5429,N_3156,N_4561);
nor U5430 (N_5430,N_3148,N_3179);
nand U5431 (N_5431,N_2650,N_4852);
or U5432 (N_5432,N_4159,N_3051);
xnor U5433 (N_5433,N_4260,N_3917);
nand U5434 (N_5434,N_4235,N_4565);
xnor U5435 (N_5435,N_4762,N_2803);
nor U5436 (N_5436,N_3905,N_4282);
or U5437 (N_5437,N_4448,N_4630);
or U5438 (N_5438,N_3138,N_3596);
or U5439 (N_5439,N_3792,N_4639);
nor U5440 (N_5440,N_4733,N_4937);
and U5441 (N_5441,N_4641,N_4328);
or U5442 (N_5442,N_3726,N_3651);
nand U5443 (N_5443,N_3578,N_3661);
nor U5444 (N_5444,N_3856,N_3157);
and U5445 (N_5445,N_4503,N_3263);
or U5446 (N_5446,N_3910,N_2601);
xor U5447 (N_5447,N_4073,N_2661);
and U5448 (N_5448,N_4221,N_3072);
xnor U5449 (N_5449,N_4601,N_4208);
nand U5450 (N_5450,N_3672,N_4225);
xor U5451 (N_5451,N_3981,N_2788);
and U5452 (N_5452,N_4027,N_4567);
xnor U5453 (N_5453,N_3439,N_4283);
nand U5454 (N_5454,N_2883,N_2844);
and U5455 (N_5455,N_2764,N_3236);
nand U5456 (N_5456,N_4580,N_3698);
and U5457 (N_5457,N_4940,N_4605);
and U5458 (N_5458,N_4899,N_3473);
xor U5459 (N_5459,N_4463,N_4677);
nor U5460 (N_5460,N_2945,N_2602);
xnor U5461 (N_5461,N_3587,N_4263);
nand U5462 (N_5462,N_2801,N_2901);
nand U5463 (N_5463,N_3388,N_3241);
nand U5464 (N_5464,N_4768,N_2630);
xor U5465 (N_5465,N_3340,N_3614);
and U5466 (N_5466,N_3099,N_2697);
or U5467 (N_5467,N_4746,N_4624);
xor U5468 (N_5468,N_2678,N_4088);
xor U5469 (N_5469,N_2565,N_2918);
and U5470 (N_5470,N_2503,N_3980);
or U5471 (N_5471,N_3264,N_4656);
nand U5472 (N_5472,N_3495,N_3010);
or U5473 (N_5473,N_2774,N_4338);
xor U5474 (N_5474,N_4227,N_3660);
or U5475 (N_5475,N_2889,N_4264);
nand U5476 (N_5476,N_4021,N_4086);
nor U5477 (N_5477,N_4276,N_2808);
and U5478 (N_5478,N_4369,N_4048);
nor U5479 (N_5479,N_4969,N_3204);
and U5480 (N_5480,N_4880,N_2993);
xnor U5481 (N_5481,N_4018,N_3599);
xor U5482 (N_5482,N_3268,N_3445);
nand U5483 (N_5483,N_4933,N_4504);
or U5484 (N_5484,N_3346,N_3316);
nor U5485 (N_5485,N_4804,N_2507);
nand U5486 (N_5486,N_3126,N_3409);
nand U5487 (N_5487,N_3835,N_4745);
or U5488 (N_5488,N_2714,N_4991);
nor U5489 (N_5489,N_3039,N_3323);
nor U5490 (N_5490,N_3249,N_2888);
nor U5491 (N_5491,N_4220,N_4560);
xor U5492 (N_5492,N_2553,N_4720);
xor U5493 (N_5493,N_3858,N_3978);
and U5494 (N_5494,N_3530,N_2722);
and U5495 (N_5495,N_3162,N_3712);
xor U5496 (N_5496,N_4008,N_3412);
or U5497 (N_5497,N_3962,N_3082);
or U5498 (N_5498,N_3243,N_4238);
nor U5499 (N_5499,N_4674,N_4963);
nand U5500 (N_5500,N_4758,N_3617);
or U5501 (N_5501,N_3246,N_4387);
or U5502 (N_5502,N_2574,N_4041);
xnor U5503 (N_5503,N_3478,N_4566);
or U5504 (N_5504,N_4793,N_4803);
and U5505 (N_5505,N_4876,N_4417);
nor U5506 (N_5506,N_4792,N_3140);
nor U5507 (N_5507,N_3915,N_4932);
or U5508 (N_5508,N_2645,N_4654);
and U5509 (N_5509,N_4649,N_2615);
or U5510 (N_5510,N_4738,N_4559);
and U5511 (N_5511,N_3278,N_3252);
or U5512 (N_5512,N_3989,N_4697);
and U5513 (N_5513,N_4323,N_4182);
nand U5514 (N_5514,N_3103,N_4265);
or U5515 (N_5515,N_2638,N_3914);
nand U5516 (N_5516,N_4435,N_3717);
nor U5517 (N_5517,N_4815,N_4038);
or U5518 (N_5518,N_2795,N_2899);
nand U5519 (N_5519,N_2655,N_4872);
nor U5520 (N_5520,N_4249,N_2712);
or U5521 (N_5521,N_2971,N_4357);
nor U5522 (N_5522,N_3390,N_4204);
nor U5523 (N_5523,N_4413,N_3427);
or U5524 (N_5524,N_3522,N_3422);
or U5525 (N_5525,N_3330,N_3822);
nor U5526 (N_5526,N_4127,N_3169);
nor U5527 (N_5527,N_3494,N_3564);
xor U5528 (N_5528,N_3932,N_4754);
or U5529 (N_5529,N_2610,N_4192);
nand U5530 (N_5530,N_3244,N_4891);
xnor U5531 (N_5531,N_3324,N_4753);
xnor U5532 (N_5532,N_2813,N_3814);
nor U5533 (N_5533,N_2671,N_4767);
nand U5534 (N_5534,N_3955,N_3083);
and U5535 (N_5535,N_4680,N_2952);
nand U5536 (N_5536,N_4224,N_4549);
nand U5537 (N_5537,N_3838,N_3294);
or U5538 (N_5538,N_4812,N_2941);
xnor U5539 (N_5539,N_3546,N_3449);
nand U5540 (N_5540,N_3342,N_4361);
and U5541 (N_5541,N_4954,N_4777);
xor U5542 (N_5542,N_4853,N_4051);
nand U5543 (N_5543,N_3504,N_3582);
or U5544 (N_5544,N_2994,N_2781);
and U5545 (N_5545,N_2809,N_4814);
and U5546 (N_5546,N_4251,N_3644);
xor U5547 (N_5547,N_4279,N_3808);
nand U5548 (N_5548,N_3786,N_4240);
xnor U5549 (N_5549,N_4449,N_3623);
xor U5550 (N_5550,N_3888,N_3381);
and U5551 (N_5551,N_3111,N_4946);
xnor U5552 (N_5552,N_3512,N_4322);
or U5553 (N_5553,N_2913,N_2689);
xor U5554 (N_5554,N_4569,N_2617);
xnor U5555 (N_5555,N_3415,N_2979);
nor U5556 (N_5556,N_4516,N_2835);
or U5557 (N_5557,N_3348,N_4540);
and U5558 (N_5558,N_3399,N_4978);
xnor U5559 (N_5559,N_2673,N_3892);
xor U5560 (N_5560,N_4469,N_3045);
nand U5561 (N_5561,N_4480,N_4244);
and U5562 (N_5562,N_2662,N_3737);
and U5563 (N_5563,N_3498,N_3555);
or U5564 (N_5564,N_3318,N_3701);
and U5565 (N_5565,N_3563,N_2830);
or U5566 (N_5566,N_2817,N_2739);
and U5567 (N_5567,N_4439,N_4695);
nor U5568 (N_5568,N_3895,N_2953);
or U5569 (N_5569,N_4156,N_3686);
and U5570 (N_5570,N_3754,N_3379);
or U5571 (N_5571,N_4355,N_4760);
and U5572 (N_5572,N_3911,N_4407);
xnor U5573 (N_5573,N_3622,N_4065);
or U5574 (N_5574,N_3143,N_4634);
xor U5575 (N_5575,N_2582,N_3702);
or U5576 (N_5576,N_4568,N_4755);
nand U5577 (N_5577,N_3729,N_3842);
nor U5578 (N_5578,N_3406,N_2903);
nand U5579 (N_5579,N_4672,N_4131);
or U5580 (N_5580,N_2792,N_4348);
or U5581 (N_5581,N_3668,N_3603);
nor U5582 (N_5582,N_3021,N_3117);
nor U5583 (N_5583,N_4947,N_2598);
and U5584 (N_5584,N_4360,N_2915);
and U5585 (N_5585,N_3795,N_3606);
nand U5586 (N_5586,N_4109,N_2619);
xnor U5587 (N_5587,N_4723,N_4699);
nand U5588 (N_5588,N_3527,N_4428);
xnor U5589 (N_5589,N_4995,N_3149);
or U5590 (N_5590,N_4136,N_4865);
and U5591 (N_5591,N_2837,N_3345);
xor U5592 (N_5592,N_3004,N_4592);
nand U5593 (N_5593,N_3825,N_3727);
xnor U5594 (N_5594,N_4562,N_2682);
xnor U5595 (N_5595,N_3155,N_4418);
or U5596 (N_5596,N_4434,N_4199);
nor U5597 (N_5597,N_3649,N_4887);
nor U5598 (N_5598,N_3079,N_4890);
and U5599 (N_5599,N_2698,N_4161);
nor U5600 (N_5600,N_4910,N_2850);
nor U5601 (N_5601,N_2500,N_4837);
and U5602 (N_5602,N_3256,N_4938);
xnor U5603 (N_5603,N_3031,N_4411);
nor U5604 (N_5604,N_4862,N_4976);
nor U5605 (N_5605,N_2726,N_4828);
and U5606 (N_5606,N_3028,N_4170);
xnor U5607 (N_5607,N_4318,N_4692);
or U5608 (N_5608,N_4867,N_3030);
or U5609 (N_5609,N_3319,N_3376);
and U5610 (N_5610,N_4554,N_4149);
or U5611 (N_5611,N_4521,N_4684);
nor U5612 (N_5612,N_3939,N_2730);
and U5613 (N_5613,N_4885,N_4233);
xnor U5614 (N_5614,N_3184,N_3805);
nand U5615 (N_5615,N_3104,N_2949);
xnor U5616 (N_5616,N_3454,N_3848);
xor U5617 (N_5617,N_2860,N_2904);
nand U5618 (N_5618,N_4181,N_2925);
xor U5619 (N_5619,N_4708,N_3745);
or U5620 (N_5620,N_4664,N_3170);
nor U5621 (N_5621,N_4799,N_4207);
nand U5622 (N_5622,N_4595,N_3247);
nor U5623 (N_5623,N_3830,N_3908);
and U5624 (N_5624,N_4627,N_2826);
nand U5625 (N_5625,N_4295,N_3718);
and U5626 (N_5626,N_4218,N_2849);
nand U5627 (N_5627,N_3671,N_3719);
xor U5628 (N_5628,N_2861,N_4153);
nor U5629 (N_5629,N_3513,N_3145);
nand U5630 (N_5630,N_4354,N_4660);
and U5631 (N_5631,N_3647,N_2828);
xor U5632 (N_5632,N_3308,N_2720);
xor U5633 (N_5633,N_4459,N_3437);
or U5634 (N_5634,N_4216,N_4307);
xor U5635 (N_5635,N_4286,N_4663);
and U5636 (N_5636,N_3872,N_4829);
xor U5637 (N_5637,N_2825,N_2690);
and U5638 (N_5638,N_3516,N_4505);
xnor U5639 (N_5639,N_4197,N_4919);
or U5640 (N_5640,N_2581,N_4557);
nand U5641 (N_5641,N_3779,N_3738);
xor U5642 (N_5642,N_3459,N_4952);
and U5643 (N_5643,N_4063,N_3547);
xor U5644 (N_5644,N_3695,N_3491);
nor U5645 (N_5645,N_4206,N_2799);
or U5646 (N_5646,N_4422,N_3583);
nor U5647 (N_5647,N_3385,N_4744);
xor U5648 (N_5648,N_4545,N_4377);
nand U5649 (N_5649,N_2798,N_2859);
xnor U5650 (N_5650,N_4588,N_2621);
nor U5651 (N_5651,N_3595,N_4317);
and U5652 (N_5652,N_4800,N_4772);
nand U5653 (N_5653,N_2884,N_2547);
nor U5654 (N_5654,N_3434,N_2659);
nor U5655 (N_5655,N_4460,N_3311);
or U5656 (N_5656,N_2561,N_4479);
or U5657 (N_5657,N_2919,N_3544);
xor U5658 (N_5658,N_4958,N_3109);
and U5659 (N_5659,N_3839,N_3150);
or U5660 (N_5660,N_4312,N_3360);
xnor U5661 (N_5661,N_4990,N_3785);
xor U5662 (N_5662,N_3832,N_2511);
xnor U5663 (N_5663,N_4362,N_3325);
nor U5664 (N_5664,N_3173,N_4104);
and U5665 (N_5665,N_4403,N_3101);
nand U5666 (N_5666,N_4761,N_3923);
and U5667 (N_5667,N_3520,N_2526);
or U5668 (N_5668,N_3001,N_3662);
nand U5669 (N_5669,N_3653,N_4500);
or U5670 (N_5670,N_3789,N_2951);
nand U5671 (N_5671,N_2814,N_3769);
and U5672 (N_5672,N_3517,N_3969);
or U5673 (N_5673,N_3928,N_2552);
xnor U5674 (N_5674,N_4006,N_3539);
nor U5675 (N_5675,N_4951,N_3628);
and U5676 (N_5676,N_2839,N_2657);
xor U5677 (N_5677,N_2734,N_2695);
and U5678 (N_5678,N_3568,N_4915);
xnor U5679 (N_5679,N_4110,N_4162);
nor U5680 (N_5680,N_3519,N_4405);
nor U5681 (N_5681,N_4689,N_2922);
and U5682 (N_5682,N_2881,N_3129);
nor U5683 (N_5683,N_4518,N_3632);
and U5684 (N_5684,N_4813,N_3676);
or U5685 (N_5685,N_2514,N_3081);
and U5686 (N_5686,N_4239,N_3624);
or U5687 (N_5687,N_4072,N_3673);
xnor U5688 (N_5688,N_3321,N_3152);
nand U5689 (N_5689,N_3545,N_4400);
nand U5690 (N_5690,N_3431,N_2867);
and U5691 (N_5691,N_3068,N_2916);
and U5692 (N_5692,N_3261,N_2729);
or U5693 (N_5693,N_2804,N_2702);
xnor U5694 (N_5694,N_3163,N_4332);
xnor U5695 (N_5695,N_3058,N_4596);
nand U5696 (N_5696,N_2778,N_3443);
nor U5697 (N_5697,N_3875,N_2575);
xor U5698 (N_5698,N_2950,N_4273);
xor U5699 (N_5699,N_4398,N_2757);
xnor U5700 (N_5700,N_4879,N_2848);
or U5701 (N_5701,N_4416,N_2933);
nor U5702 (N_5702,N_3334,N_2533);
xnor U5703 (N_5703,N_3559,N_3354);
and U5704 (N_5704,N_3285,N_2902);
or U5705 (N_5705,N_4838,N_3227);
and U5706 (N_5706,N_3629,N_4270);
xor U5707 (N_5707,N_3382,N_4246);
nand U5708 (N_5708,N_3958,N_3159);
nand U5709 (N_5709,N_3691,N_3393);
or U5710 (N_5710,N_3515,N_3313);
and U5711 (N_5711,N_2758,N_4640);
nand U5712 (N_5712,N_4294,N_4043);
xnor U5713 (N_5713,N_2674,N_3542);
and U5714 (N_5714,N_4527,N_4436);
xnor U5715 (N_5715,N_3403,N_4180);
nand U5716 (N_5716,N_3044,N_3966);
and U5717 (N_5717,N_3819,N_3669);
nand U5718 (N_5718,N_3446,N_3259);
nor U5719 (N_5719,N_2544,N_3091);
nand U5720 (N_5720,N_4691,N_4074);
and U5721 (N_5721,N_4374,N_2685);
and U5722 (N_5722,N_3776,N_2701);
xor U5723 (N_5723,N_3217,N_2742);
nand U5724 (N_5724,N_3714,N_4523);
nor U5725 (N_5725,N_4564,N_3375);
or U5726 (N_5726,N_2747,N_3764);
or U5727 (N_5727,N_4289,N_3942);
nor U5728 (N_5728,N_2652,N_2585);
nand U5729 (N_5729,N_2984,N_3736);
and U5730 (N_5730,N_2699,N_4128);
xor U5731 (N_5731,N_3481,N_2963);
and U5732 (N_5732,N_2613,N_4775);
nand U5733 (N_5733,N_4124,N_3883);
or U5734 (N_5734,N_3979,N_2980);
or U5735 (N_5735,N_2700,N_3214);
xor U5736 (N_5736,N_4898,N_4278);
xnor U5737 (N_5737,N_2724,N_3078);
xnor U5738 (N_5738,N_2562,N_4230);
or U5739 (N_5739,N_4039,N_4581);
nand U5740 (N_5740,N_3469,N_3270);
xor U5741 (N_5741,N_4026,N_4366);
or U5742 (N_5742,N_4035,N_2969);
and U5743 (N_5743,N_2556,N_2968);
nor U5744 (N_5744,N_4901,N_3374);
xor U5745 (N_5745,N_4707,N_3076);
nand U5746 (N_5746,N_3232,N_3999);
nor U5747 (N_5747,N_3153,N_4442);
or U5748 (N_5748,N_3852,N_3552);
nand U5749 (N_5749,N_4138,N_4126);
nor U5750 (N_5750,N_3739,N_3397);
nor U5751 (N_5751,N_4513,N_4682);
and U5752 (N_5752,N_3927,N_2768);
or U5753 (N_5753,N_3003,N_2706);
xnor U5754 (N_5754,N_3609,N_2524);
and U5755 (N_5755,N_3537,N_4542);
xor U5756 (N_5756,N_4731,N_4713);
nor U5757 (N_5757,N_2709,N_4798);
and U5758 (N_5758,N_4472,N_2546);
nand U5759 (N_5759,N_2717,N_4119);
or U5760 (N_5760,N_4805,N_3639);
xnor U5761 (N_5761,N_2880,N_3050);
xnor U5762 (N_5762,N_3147,N_2912);
xnor U5763 (N_5763,N_4541,N_4819);
nor U5764 (N_5764,N_3178,N_4927);
nor U5765 (N_5765,N_4894,N_3070);
or U5766 (N_5766,N_3864,N_4553);
nor U5767 (N_5767,N_2751,N_3245);
nand U5768 (N_5768,N_4420,N_3413);
xnor U5769 (N_5769,N_3141,N_2590);
and U5770 (N_5770,N_4236,N_3492);
or U5771 (N_5771,N_4406,N_2907);
nor U5772 (N_5772,N_3740,N_3447);
and U5773 (N_5773,N_3975,N_2538);
and U5774 (N_5774,N_3218,N_4701);
or U5775 (N_5775,N_3074,N_4749);
and U5776 (N_5776,N_3585,N_3538);
nand U5777 (N_5777,N_3976,N_4506);
and U5778 (N_5778,N_3573,N_4452);
nand U5779 (N_5779,N_3646,N_4315);
or U5780 (N_5780,N_4047,N_4917);
xor U5781 (N_5781,N_4526,N_4959);
nor U5782 (N_5782,N_3531,N_3937);
nand U5783 (N_5783,N_3893,N_2772);
xor U5784 (N_5784,N_3377,N_3116);
xnor U5785 (N_5785,N_3993,N_4060);
and U5786 (N_5786,N_4688,N_4942);
nand U5787 (N_5787,N_3420,N_3018);
or U5788 (N_5788,N_3131,N_3560);
or U5789 (N_5789,N_4237,N_4735);
and U5790 (N_5790,N_4087,N_4607);
and U5791 (N_5791,N_4636,N_3097);
or U5792 (N_5792,N_4498,N_4611);
xnor U5793 (N_5793,N_3366,N_4686);
xnor U5794 (N_5794,N_4816,N_3876);
nor U5795 (N_5795,N_2522,N_4823);
nor U5796 (N_5796,N_4712,N_3821);
nand U5797 (N_5797,N_4784,N_4536);
or U5798 (N_5798,N_4743,N_4223);
nor U5799 (N_5799,N_4840,N_3436);
nor U5800 (N_5800,N_3488,N_4811);
or U5801 (N_5801,N_3168,N_3971);
and U5802 (N_5802,N_4757,N_4137);
xnor U5803 (N_5803,N_4146,N_3773);
or U5804 (N_5804,N_4765,N_3800);
nand U5805 (N_5805,N_3734,N_4797);
xor U5806 (N_5806,N_3600,N_3306);
xnor U5807 (N_5807,N_3896,N_3479);
and U5808 (N_5808,N_4430,N_4316);
and U5809 (N_5809,N_4613,N_4629);
or U5810 (N_5810,N_4644,N_4488);
nand U5811 (N_5811,N_2624,N_4174);
xnor U5812 (N_5812,N_2525,N_3793);
nor U5813 (N_5813,N_3238,N_4122);
or U5814 (N_5814,N_4176,N_4130);
and U5815 (N_5815,N_3898,N_4147);
xor U5816 (N_5816,N_3666,N_3947);
or U5817 (N_5817,N_3521,N_3813);
and U5818 (N_5818,N_3746,N_2632);
nor U5819 (N_5819,N_3305,N_3450);
nor U5820 (N_5820,N_4970,N_4842);
nand U5821 (N_5821,N_3047,N_2827);
and U5822 (N_5822,N_3847,N_4786);
xor U5823 (N_5823,N_3391,N_2504);
and U5824 (N_5824,N_4261,N_3815);
xor U5825 (N_5825,N_3997,N_2779);
xor U5826 (N_5826,N_4949,N_4165);
nor U5827 (N_5827,N_3200,N_3584);
xor U5828 (N_5828,N_3177,N_2591);
and U5829 (N_5829,N_3744,N_3151);
or U5830 (N_5830,N_2934,N_4719);
and U5831 (N_5831,N_2966,N_4920);
xor U5832 (N_5832,N_3333,N_4993);
or U5833 (N_5833,N_3557,N_3984);
and U5834 (N_5834,N_3480,N_3211);
and U5835 (N_5835,N_4558,N_3855);
or U5836 (N_5836,N_2930,N_2864);
or U5837 (N_5837,N_4393,N_4334);
and U5838 (N_5838,N_4081,N_3326);
xnor U5839 (N_5839,N_3619,N_4167);
and U5840 (N_5840,N_4953,N_3095);
nor U5841 (N_5841,N_3302,N_4499);
or U5842 (N_5842,N_3591,N_4245);
xnor U5843 (N_5843,N_4806,N_2831);
or U5844 (N_5844,N_4936,N_4168);
xor U5845 (N_5845,N_2782,N_4818);
or U5846 (N_5846,N_4830,N_2510);
xnor U5847 (N_5847,N_3943,N_2535);
nand U5848 (N_5848,N_4603,N_4066);
nor U5849 (N_5849,N_3990,N_2676);
xnor U5850 (N_5850,N_4116,N_4046);
and U5851 (N_5851,N_4157,N_3797);
xor U5852 (N_5852,N_2675,N_3120);
nor U5853 (N_5853,N_3757,N_3581);
nor U5854 (N_5854,N_3798,N_4706);
and U5855 (N_5855,N_2756,N_2773);
xor U5856 (N_5856,N_2816,N_4896);
xnor U5857 (N_5857,N_3625,N_4198);
and U5858 (N_5858,N_3037,N_4141);
and U5859 (N_5859,N_2986,N_3806);
nand U5860 (N_5860,N_3948,N_4384);
nor U5861 (N_5861,N_3902,N_3951);
and U5862 (N_5862,N_4028,N_4256);
nor U5863 (N_5863,N_2992,N_4875);
nor U5864 (N_5864,N_3631,N_2716);
and U5865 (N_5865,N_4905,N_4831);
or U5866 (N_5866,N_3758,N_4186);
or U5867 (N_5867,N_4297,N_3216);
nand U5868 (N_5868,N_3503,N_3380);
nand U5869 (N_5869,N_4529,N_4189);
nor U5870 (N_5870,N_3106,N_2517);
nand U5871 (N_5871,N_3146,N_3466);
nand U5872 (N_5872,N_4040,N_4924);
or U5873 (N_5873,N_4457,N_2542);
or U5874 (N_5874,N_3765,N_2669);
xnor U5875 (N_5875,N_4683,N_4350);
nor U5876 (N_5876,N_4602,N_4058);
xor U5877 (N_5877,N_3974,N_2935);
or U5878 (N_5878,N_4730,N_4888);
nor U5879 (N_5879,N_4320,N_2611);
xnor U5880 (N_5880,N_4117,N_4992);
xor U5881 (N_5881,N_2897,N_3723);
nand U5882 (N_5882,N_4173,N_2891);
or U5883 (N_5883,N_2924,N_3008);
nand U5884 (N_5884,N_4363,N_4234);
nor U5885 (N_5885,N_2731,N_3338);
xor U5886 (N_5886,N_4099,N_2651);
nand U5887 (N_5887,N_2885,N_4319);
and U5888 (N_5888,N_3598,N_4631);
nor U5889 (N_5889,N_4739,N_3807);
and U5890 (N_5890,N_2887,N_3502);
nand U5891 (N_5891,N_2634,N_4401);
nand U5892 (N_5892,N_2829,N_3715);
nand U5893 (N_5893,N_2616,N_3239);
nand U5894 (N_5894,N_2958,N_4166);
and U5895 (N_5895,N_2583,N_4955);
nand U5896 (N_5896,N_4495,N_3772);
or U5897 (N_5897,N_2875,N_4675);
xor U5898 (N_5898,N_3750,N_4681);
xnor U5899 (N_5899,N_2572,N_4671);
nor U5900 (N_5900,N_3636,N_4062);
xor U5901 (N_5901,N_4787,N_3677);
nor U5902 (N_5902,N_4822,N_3404);
nand U5903 (N_5903,N_3102,N_4052);
xnor U5904 (N_5904,N_4628,N_3638);
or U5905 (N_5905,N_3549,N_4143);
nand U5906 (N_5906,N_4154,N_4778);
and U5907 (N_5907,N_3040,N_3950);
xor U5908 (N_5908,N_2563,N_2587);
or U5909 (N_5909,N_2960,N_3841);
or U5910 (N_5910,N_3271,N_2929);
xnor U5911 (N_5911,N_3332,N_4593);
and U5912 (N_5912,N_2863,N_4226);
nand U5913 (N_5913,N_2931,N_2527);
xor U5914 (N_5914,N_2691,N_4292);
xor U5915 (N_5915,N_3312,N_4144);
and U5916 (N_5916,N_2603,N_2914);
nand U5917 (N_5917,N_4213,N_4092);
xor U5918 (N_5918,N_2580,N_3987);
and U5919 (N_5919,N_4612,N_4054);
nand U5920 (N_5920,N_4044,N_3006);
xor U5921 (N_5921,N_3843,N_3065);
xnor U5922 (N_5922,N_3353,N_4326);
nand U5923 (N_5923,N_2711,N_4535);
or U5924 (N_5924,N_4789,N_4858);
nand U5925 (N_5925,N_3322,N_4190);
and U5926 (N_5926,N_4659,N_4140);
xnor U5927 (N_5927,N_3274,N_4897);
nand U5928 (N_5928,N_4419,N_3853);
or U5929 (N_5929,N_3857,N_3015);
nor U5930 (N_5930,N_3961,N_3777);
nand U5931 (N_5931,N_3384,N_4485);
nor U5932 (N_5932,N_3273,N_4005);
nor U5933 (N_5933,N_4100,N_3972);
nor U5934 (N_5934,N_3780,N_4024);
xor U5935 (N_5935,N_3845,N_2770);
and U5936 (N_5936,N_3172,N_4661);
xnor U5937 (N_5937,N_4321,N_3925);
nor U5938 (N_5938,N_4343,N_4451);
or U5939 (N_5939,N_4349,N_3225);
xnor U5940 (N_5940,N_4011,N_4973);
or U5941 (N_5941,N_3548,N_3364);
and U5942 (N_5942,N_4183,N_4537);
and U5943 (N_5943,N_3114,N_4466);
nand U5944 (N_5944,N_4045,N_4676);
and U5945 (N_5945,N_3194,N_3280);
nor U5946 (N_5946,N_3953,N_4421);
nor U5947 (N_5947,N_4281,N_4000);
xnor U5948 (N_5948,N_3812,N_4886);
or U5949 (N_5949,N_4725,N_2705);
xnor U5950 (N_5950,N_4614,N_3863);
xor U5951 (N_5951,N_2721,N_3056);
and U5952 (N_5952,N_4563,N_4125);
xor U5953 (N_5953,N_3336,N_2857);
nor U5954 (N_5954,N_4836,N_3998);
or U5955 (N_5955,N_2737,N_3919);
and U5956 (N_5956,N_4944,N_3284);
or U5957 (N_5957,N_2812,N_3372);
nand U5958 (N_5958,N_4415,N_2910);
and U5959 (N_5959,N_4667,N_2736);
nor U5960 (N_5960,N_4825,N_4907);
xnor U5961 (N_5961,N_2824,N_3092);
xor U5962 (N_5962,N_3588,N_2753);
nand U5963 (N_5963,N_4988,N_4248);
xnor U5964 (N_5964,N_4922,N_3866);
or U5965 (N_5965,N_4633,N_3233);
or U5966 (N_5966,N_3543,N_2519);
xor U5967 (N_5967,N_2567,N_4934);
and U5968 (N_5968,N_4414,N_4635);
xnor U5969 (N_5969,N_3679,N_3616);
and U5970 (N_5970,N_3059,N_3655);
nand U5971 (N_5971,N_2588,N_2636);
and U5972 (N_5972,N_3164,N_4196);
and U5973 (N_5973,N_2978,N_3186);
nand U5974 (N_5974,N_4850,N_3282);
nand U5975 (N_5975,N_4059,N_2520);
or U5976 (N_5976,N_4893,N_4687);
xnor U5977 (N_5977,N_3554,N_4861);
nor U5978 (N_5978,N_4869,N_3213);
nand U5979 (N_5979,N_3724,N_2513);
nor U5980 (N_5980,N_3137,N_4450);
or U5981 (N_5981,N_4483,N_2943);
and U5982 (N_5982,N_4998,N_2625);
or U5983 (N_5983,N_3368,N_3889);
nor U5984 (N_5984,N_4737,N_3123);
nand U5985 (N_5985,N_3387,N_4948);
nand U5986 (N_5986,N_3658,N_4771);
xnor U5987 (N_5987,N_4522,N_2975);
xor U5988 (N_5988,N_4846,N_2501);
nand U5989 (N_5989,N_3329,N_3125);
and U5990 (N_5990,N_2838,N_3304);
or U5991 (N_5991,N_4844,N_3721);
nor U5992 (N_5992,N_3823,N_3916);
or U5993 (N_5993,N_4734,N_3416);
nor U5994 (N_5994,N_3281,N_4111);
and U5995 (N_5995,N_4367,N_4685);
xnor U5996 (N_5996,N_2748,N_3433);
nor U5997 (N_5997,N_4543,N_3621);
and U5998 (N_5998,N_2622,N_2937);
xnor U5999 (N_5999,N_3831,N_3396);
xnor U6000 (N_6000,N_4462,N_2570);
nor U6001 (N_6001,N_4960,N_2684);
nor U6002 (N_6002,N_4845,N_2614);
and U6003 (N_6003,N_2856,N_3357);
xor U6004 (N_6004,N_2896,N_4465);
and U6005 (N_6005,N_4801,N_4967);
xnor U6006 (N_6006,N_2784,N_2536);
nand U6007 (N_6007,N_3973,N_4752);
nor U6008 (N_6008,N_4356,N_4389);
nand U6009 (N_6009,N_4650,N_3471);
xnor U6010 (N_6010,N_4764,N_4151);
nor U6011 (N_6011,N_4358,N_3175);
nor U6012 (N_6012,N_4783,N_4461);
nor U6013 (N_6013,N_4647,N_3802);
and U6014 (N_6014,N_3253,N_4903);
xor U6015 (N_6015,N_2755,N_3034);
and U6016 (N_6016,N_2866,N_3940);
and U6017 (N_6017,N_2595,N_3054);
xnor U6018 (N_6018,N_2846,N_2998);
nor U6019 (N_6019,N_3577,N_2997);
nand U6020 (N_6020,N_3509,N_3307);
xnor U6021 (N_6021,N_3262,N_4796);
and U6022 (N_6022,N_4271,N_4632);
nand U6023 (N_6023,N_3870,N_2745);
or U6024 (N_6024,N_2560,N_4142);
xnor U6025 (N_6025,N_4287,N_4464);
or U6026 (N_6026,N_3634,N_3605);
and U6027 (N_6027,N_4668,N_4770);
nor U6028 (N_6028,N_2987,N_2868);
nand U6029 (N_6029,N_4961,N_3778);
and U6030 (N_6030,N_4637,N_2743);
nand U6031 (N_6031,N_2890,N_2518);
xnor U6032 (N_6032,N_4550,N_4135);
nor U6033 (N_6033,N_4115,N_2762);
or U6034 (N_6034,N_2767,N_4337);
and U6035 (N_6035,N_3303,N_3371);
xnor U6036 (N_6036,N_4194,N_3025);
or U6037 (N_6037,N_3565,N_4303);
nand U6038 (N_6038,N_3258,N_3755);
and U6039 (N_6039,N_4833,N_3350);
nand U6040 (N_6040,N_4371,N_3135);
or U6041 (N_6041,N_4114,N_4139);
nor U6042 (N_6042,N_4177,N_4456);
xor U6043 (N_6043,N_2789,N_4620);
nor U6044 (N_6044,N_3367,N_3611);
nor U6045 (N_6045,N_4426,N_2687);
nand U6046 (N_6046,N_3002,N_3124);
nor U6047 (N_6047,N_3781,N_4229);
and U6048 (N_6048,N_3287,N_4424);
xnor U6049 (N_6049,N_3692,N_2569);
or U6050 (N_6050,N_3891,N_3551);
nand U6051 (N_6051,N_4121,N_4105);
nand U6052 (N_6052,N_4820,N_4296);
and U6053 (N_6053,N_3706,N_3069);
nor U6054 (N_6054,N_4191,N_2640);
or U6055 (N_6055,N_3205,N_4049);
and U6056 (N_6056,N_3711,N_3827);
nor U6057 (N_6057,N_2862,N_4133);
or U6058 (N_6058,N_4431,N_3020);
nand U6059 (N_6059,N_4372,N_4164);
nand U6060 (N_6060,N_3193,N_4184);
and U6061 (N_6061,N_4904,N_4926);
nor U6062 (N_6062,N_3041,N_4395);
or U6063 (N_6063,N_3570,N_4882);
nor U6064 (N_6064,N_3710,N_4368);
and U6065 (N_6065,N_4057,N_3656);
nand U6066 (N_6066,N_3766,N_2750);
and U6067 (N_6067,N_3608,N_3331);
or U6068 (N_6068,N_3524,N_3472);
and U6069 (N_6069,N_3566,N_3207);
or U6070 (N_6070,N_4583,N_3486);
nor U6071 (N_6071,N_3871,N_3751);
xnor U6072 (N_6072,N_2822,N_3448);
and U6073 (N_6073,N_3796,N_3931);
and U6074 (N_6074,N_4939,N_2981);
and U6075 (N_6075,N_3700,N_4306);
or U6076 (N_6076,N_4776,N_2754);
or U6077 (N_6077,N_4007,N_3463);
nand U6078 (N_6078,N_3460,N_3161);
nand U6079 (N_6079,N_3327,N_4496);
and U6080 (N_6080,N_2554,N_3994);
nor U6081 (N_6081,N_4277,N_2646);
xor U6082 (N_6082,N_2605,N_4094);
nand U6083 (N_6083,N_2592,N_4841);
nand U6084 (N_6084,N_4538,N_4843);
or U6085 (N_6085,N_2532,N_2609);
nand U6086 (N_6086,N_3682,N_2641);
xor U6087 (N_6087,N_3663,N_4694);
xnor U6088 (N_6088,N_3100,N_3762);
and U6089 (N_6089,N_2843,N_4080);
xnor U6090 (N_6090,N_3080,N_3930);
xnor U6091 (N_6091,N_4856,N_4514);
and U6092 (N_6092,N_3921,N_3224);
and U6093 (N_6093,N_3569,N_3912);
or U6094 (N_6094,N_3132,N_2704);
or U6095 (N_6095,N_3849,N_4340);
nor U6096 (N_6096,N_3369,N_4555);
nand U6097 (N_6097,N_4791,N_4274);
nor U6098 (N_6098,N_3048,N_2905);
nand U6099 (N_6099,N_4475,N_4333);
nand U6100 (N_6100,N_2600,N_4359);
or U6101 (N_6101,N_4616,N_4509);
or U6102 (N_6102,N_2763,N_2710);
xor U6103 (N_6103,N_2940,N_3759);
nand U6104 (N_6104,N_4410,N_3254);
xor U6105 (N_6105,N_3185,N_4433);
or U6106 (N_6106,N_3351,N_4643);
or U6107 (N_6107,N_2608,N_3424);
xor U6108 (N_6108,N_4145,N_4440);
or U6109 (N_6109,N_4388,N_3013);
nor U6110 (N_6110,N_4600,N_3339);
xnor U6111 (N_6111,N_2589,N_2800);
nor U6112 (N_6112,N_3220,N_2549);
nor U6113 (N_6113,N_2936,N_3203);
nor U6114 (N_6114,N_4304,N_3130);
nor U6115 (N_6115,N_3229,N_3935);
and U6116 (N_6116,N_3266,N_4432);
nor U6117 (N_6117,N_4589,N_4983);
nor U6118 (N_6118,N_2955,N_4981);
xnor U6119 (N_6119,N_4729,N_4916);
nor U6120 (N_6120,N_3467,N_4623);
nor U6121 (N_6121,N_4446,N_2842);
and U6122 (N_6122,N_4346,N_3288);
and U6123 (N_6123,N_2732,N_3946);
and U6124 (N_6124,N_2596,N_2576);
or U6125 (N_6125,N_2629,N_3113);
nor U6126 (N_6126,N_3816,N_4324);
or U6127 (N_6127,N_3586,N_4696);
or U6128 (N_6128,N_2670,N_3210);
xor U6129 (N_6129,N_3722,N_4510);
xnor U6130 (N_6130,N_4029,N_3142);
or U6131 (N_6131,N_2926,N_3988);
or U6132 (N_6132,N_4849,N_4578);
nor U6133 (N_6133,N_3556,N_2766);
nand U6134 (N_6134,N_2648,N_4574);
and U6135 (N_6135,N_4243,N_3826);
nand U6136 (N_6136,N_3462,N_3709);
nand U6137 (N_6137,N_3968,N_4399);
nor U6138 (N_6138,N_3933,N_4711);
xor U6139 (N_6139,N_3899,N_3136);
xor U6140 (N_6140,N_4489,N_3356);
nor U6141 (N_6141,N_2728,N_3154);
and U6142 (N_6142,N_2985,N_2693);
or U6143 (N_6143,N_3257,N_3741);
xnor U6144 (N_6144,N_4179,N_2604);
and U6145 (N_6145,N_3430,N_4585);
nand U6146 (N_6146,N_3528,N_4769);
xnor U6147 (N_6147,N_3358,N_4606);
xor U6148 (N_6148,N_3468,N_3650);
or U6149 (N_6149,N_2537,N_3347);
xor U6150 (N_6150,N_3038,N_3850);
nand U6151 (N_6151,N_4718,N_3833);
or U6152 (N_6152,N_3234,N_3697);
xor U6153 (N_6153,N_4889,N_3970);
or U6154 (N_6154,N_3359,N_2879);
or U6155 (N_6155,N_4017,N_2811);
or U6156 (N_6156,N_2946,N_3112);
and U6157 (N_6157,N_4728,N_3206);
xnor U6158 (N_6158,N_2877,N_3496);
and U6159 (N_6159,N_3904,N_4402);
nor U6160 (N_6160,N_4193,N_4763);
or U6161 (N_6161,N_2845,N_2692);
xor U6162 (N_6162,N_3977,N_4015);
nand U6163 (N_6163,N_4095,N_4714);
nand U6164 (N_6164,N_3810,N_2923);
or U6165 (N_6165,N_4266,N_3834);
and U6166 (N_6166,N_3442,N_4107);
and U6167 (N_6167,N_4827,N_3482);
and U6168 (N_6168,N_4036,N_4726);
and U6169 (N_6169,N_3558,N_4573);
and U6170 (N_6170,N_2566,N_4155);
nor U6171 (N_6171,N_3049,N_4759);
or U6172 (N_6172,N_4622,N_2715);
or U6173 (N_6173,N_3215,N_4383);
and U6174 (N_6174,N_3594,N_4895);
nor U6175 (N_6175,N_3461,N_3612);
nor U6176 (N_6176,N_4487,N_2512);
and U6177 (N_6177,N_3098,N_3062);
nor U6178 (N_6178,N_4163,N_2805);
nand U6179 (N_6179,N_2573,N_3171);
nand U6180 (N_6180,N_2832,N_2999);
or U6181 (N_6181,N_4471,N_3426);
and U6182 (N_6182,N_4247,N_4859);
or U6183 (N_6183,N_2594,N_4502);
and U6184 (N_6184,N_3361,N_4404);
nand U6185 (N_6185,N_4794,N_2790);
nor U6186 (N_6186,N_2944,N_4780);
or U6187 (N_6187,N_4900,N_4666);
nand U6188 (N_6188,N_2855,N_3378);
and U6189 (N_6189,N_2663,N_3208);
nor U6190 (N_6190,N_4571,N_4445);
and U6191 (N_6191,N_4067,N_3642);
nand U6192 (N_6192,N_2970,N_3269);
xnor U6193 (N_6193,N_4098,N_3728);
xnor U6194 (N_6194,N_2786,N_3604);
nand U6195 (N_6195,N_4268,N_4572);
or U6196 (N_6196,N_4617,N_2635);
nand U6197 (N_6197,N_2954,N_4232);
nand U6198 (N_6198,N_3963,N_3042);
xor U6199 (N_6199,N_2988,N_3228);
xor U6200 (N_6200,N_4982,N_3730);
nand U6201 (N_6201,N_3882,N_2626);
nor U6202 (N_6202,N_4715,N_4911);
nor U6203 (N_6203,N_4441,N_3490);
and U6204 (N_6204,N_4075,N_4883);
nand U6205 (N_6205,N_3181,N_2807);
nor U6206 (N_6206,N_4455,N_3158);
and U6207 (N_6207,N_3770,N_4258);
or U6208 (N_6208,N_3341,N_3590);
xnor U6209 (N_6209,N_4619,N_3444);
nand U6210 (N_6210,N_4375,N_3355);
nand U6211 (N_6211,N_3913,N_4785);
nor U6212 (N_6212,N_4964,N_3550);
and U6213 (N_6213,N_4290,N_2733);
nand U6214 (N_6214,N_2851,N_3794);
nor U6215 (N_6215,N_4438,N_3922);
nand U6216 (N_6216,N_3344,N_3250);
and U6217 (N_6217,N_4444,N_2775);
nand U6218 (N_6218,N_3202,N_3884);
and U6219 (N_6219,N_4609,N_3620);
xor U6220 (N_6220,N_2623,N_3873);
or U6221 (N_6221,N_4309,N_4423);
nor U6222 (N_6222,N_3497,N_4999);
nor U6223 (N_6223,N_3183,N_3846);
nand U6224 (N_6224,N_3201,N_4061);
xnor U6225 (N_6225,N_4873,N_3187);
and U6226 (N_6226,N_3419,N_3337);
nand U6227 (N_6227,N_3868,N_4490);
or U6228 (N_6228,N_4202,N_4834);
and U6229 (N_6229,N_2787,N_4458);
and U6230 (N_6230,N_3219,N_3122);
nand U6231 (N_6231,N_3732,N_3093);
xnor U6232 (N_6232,N_3613,N_4670);
or U6233 (N_6233,N_2564,N_3299);
and U6234 (N_6234,N_4030,N_3456);
and U6235 (N_6235,N_4935,N_2539);
xor U6236 (N_6236,N_4120,N_3108);
or U6237 (N_6237,N_4519,N_3526);
nor U6238 (N_6238,N_2948,N_3803);
nor U6239 (N_6239,N_3877,N_4254);
nand U6240 (N_6240,N_2578,N_4083);
nor U6241 (N_6241,N_4329,N_3938);
nor U6242 (N_6242,N_4331,N_4473);
xor U6243 (N_6243,N_3089,N_3756);
nor U6244 (N_6244,N_4577,N_4625);
nand U6245 (N_6245,N_3291,N_3753);
xor U6246 (N_6246,N_2521,N_3505);
nand U6247 (N_6247,N_4507,N_3483);
or U6248 (N_6248,N_4034,N_3571);
nand U6249 (N_6249,N_4750,N_3901);
nand U6250 (N_6250,N_4698,N_3598);
and U6251 (N_6251,N_3751,N_2541);
and U6252 (N_6252,N_4083,N_4840);
or U6253 (N_6253,N_2810,N_4610);
xor U6254 (N_6254,N_2596,N_3826);
or U6255 (N_6255,N_4059,N_3866);
nand U6256 (N_6256,N_3404,N_2902);
xor U6257 (N_6257,N_3189,N_2594);
or U6258 (N_6258,N_2715,N_3101);
nor U6259 (N_6259,N_4526,N_2676);
xnor U6260 (N_6260,N_3085,N_3528);
nor U6261 (N_6261,N_3987,N_4148);
nand U6262 (N_6262,N_4159,N_2867);
and U6263 (N_6263,N_4132,N_3899);
nand U6264 (N_6264,N_3386,N_2542);
xnor U6265 (N_6265,N_4414,N_2853);
and U6266 (N_6266,N_3678,N_3875);
nand U6267 (N_6267,N_4047,N_4891);
or U6268 (N_6268,N_4049,N_3978);
and U6269 (N_6269,N_4157,N_4910);
or U6270 (N_6270,N_3864,N_3405);
xor U6271 (N_6271,N_4473,N_4303);
and U6272 (N_6272,N_3269,N_4385);
xnor U6273 (N_6273,N_3402,N_4560);
and U6274 (N_6274,N_2743,N_3391);
nor U6275 (N_6275,N_4908,N_3246);
and U6276 (N_6276,N_4666,N_3174);
xor U6277 (N_6277,N_3640,N_3243);
or U6278 (N_6278,N_4915,N_4951);
nand U6279 (N_6279,N_3128,N_3343);
nand U6280 (N_6280,N_4207,N_4425);
nand U6281 (N_6281,N_3250,N_3938);
nor U6282 (N_6282,N_3810,N_2917);
nand U6283 (N_6283,N_4884,N_3018);
nand U6284 (N_6284,N_3454,N_3701);
and U6285 (N_6285,N_4608,N_4853);
nor U6286 (N_6286,N_3822,N_4396);
nor U6287 (N_6287,N_3979,N_2533);
and U6288 (N_6288,N_3888,N_4003);
and U6289 (N_6289,N_3820,N_3304);
or U6290 (N_6290,N_4037,N_4300);
nand U6291 (N_6291,N_4094,N_4725);
and U6292 (N_6292,N_3723,N_4232);
and U6293 (N_6293,N_2963,N_3093);
nor U6294 (N_6294,N_3850,N_3753);
xor U6295 (N_6295,N_4676,N_4706);
xnor U6296 (N_6296,N_3377,N_4133);
or U6297 (N_6297,N_4439,N_4605);
or U6298 (N_6298,N_3135,N_2569);
and U6299 (N_6299,N_3088,N_4768);
nor U6300 (N_6300,N_3602,N_2983);
and U6301 (N_6301,N_3658,N_3322);
nor U6302 (N_6302,N_4325,N_3988);
nand U6303 (N_6303,N_3025,N_4763);
or U6304 (N_6304,N_4026,N_3757);
or U6305 (N_6305,N_2878,N_2632);
or U6306 (N_6306,N_2503,N_4342);
xor U6307 (N_6307,N_3406,N_4042);
nor U6308 (N_6308,N_4097,N_4249);
or U6309 (N_6309,N_3077,N_3461);
nand U6310 (N_6310,N_3665,N_3347);
xnor U6311 (N_6311,N_2767,N_3544);
nor U6312 (N_6312,N_3214,N_4741);
xor U6313 (N_6313,N_3292,N_3627);
or U6314 (N_6314,N_3341,N_4944);
xnor U6315 (N_6315,N_4826,N_4848);
or U6316 (N_6316,N_4665,N_4986);
nand U6317 (N_6317,N_3617,N_3142);
nor U6318 (N_6318,N_2508,N_3111);
or U6319 (N_6319,N_4063,N_3520);
nor U6320 (N_6320,N_2501,N_4552);
and U6321 (N_6321,N_3834,N_3999);
and U6322 (N_6322,N_3814,N_3551);
nor U6323 (N_6323,N_2697,N_4951);
nor U6324 (N_6324,N_3709,N_2762);
or U6325 (N_6325,N_3024,N_3583);
and U6326 (N_6326,N_2881,N_4385);
nand U6327 (N_6327,N_3243,N_3428);
and U6328 (N_6328,N_4392,N_4710);
and U6329 (N_6329,N_3215,N_4290);
and U6330 (N_6330,N_2971,N_4774);
and U6331 (N_6331,N_2557,N_4469);
and U6332 (N_6332,N_3842,N_3028);
and U6333 (N_6333,N_4615,N_4955);
xnor U6334 (N_6334,N_4570,N_3454);
nor U6335 (N_6335,N_2633,N_3834);
nor U6336 (N_6336,N_3823,N_4119);
xnor U6337 (N_6337,N_2803,N_3796);
xnor U6338 (N_6338,N_3787,N_4398);
nand U6339 (N_6339,N_4907,N_3341);
nor U6340 (N_6340,N_2731,N_3997);
nor U6341 (N_6341,N_3734,N_3265);
and U6342 (N_6342,N_4080,N_4680);
nor U6343 (N_6343,N_4027,N_4343);
nand U6344 (N_6344,N_3474,N_3283);
nor U6345 (N_6345,N_3623,N_3327);
xor U6346 (N_6346,N_3624,N_2725);
and U6347 (N_6347,N_3592,N_4325);
or U6348 (N_6348,N_4624,N_4551);
or U6349 (N_6349,N_4295,N_3111);
and U6350 (N_6350,N_4168,N_3727);
and U6351 (N_6351,N_3979,N_4581);
nand U6352 (N_6352,N_3474,N_4496);
nor U6353 (N_6353,N_2524,N_2886);
or U6354 (N_6354,N_4053,N_4990);
nor U6355 (N_6355,N_3909,N_3141);
nand U6356 (N_6356,N_3134,N_4708);
nand U6357 (N_6357,N_4128,N_4747);
nand U6358 (N_6358,N_4749,N_3969);
and U6359 (N_6359,N_2589,N_2919);
nor U6360 (N_6360,N_2787,N_4864);
nand U6361 (N_6361,N_3025,N_4307);
nand U6362 (N_6362,N_3551,N_4951);
nand U6363 (N_6363,N_3570,N_2731);
nor U6364 (N_6364,N_3388,N_3253);
and U6365 (N_6365,N_4295,N_3372);
and U6366 (N_6366,N_2824,N_3604);
nor U6367 (N_6367,N_4924,N_4372);
xor U6368 (N_6368,N_3029,N_4866);
nor U6369 (N_6369,N_2982,N_3597);
and U6370 (N_6370,N_4875,N_3506);
or U6371 (N_6371,N_3549,N_3149);
and U6372 (N_6372,N_4714,N_4613);
or U6373 (N_6373,N_3317,N_4960);
and U6374 (N_6374,N_3326,N_4014);
and U6375 (N_6375,N_3684,N_2756);
or U6376 (N_6376,N_4417,N_3484);
nor U6377 (N_6377,N_4461,N_4343);
nand U6378 (N_6378,N_3870,N_4857);
or U6379 (N_6379,N_4528,N_4216);
xnor U6380 (N_6380,N_4107,N_3128);
xor U6381 (N_6381,N_3187,N_3325);
or U6382 (N_6382,N_2703,N_3194);
or U6383 (N_6383,N_2581,N_3181);
or U6384 (N_6384,N_4238,N_3752);
nor U6385 (N_6385,N_3175,N_3511);
xor U6386 (N_6386,N_4695,N_3787);
nor U6387 (N_6387,N_3375,N_2844);
and U6388 (N_6388,N_2571,N_4089);
xor U6389 (N_6389,N_4699,N_3175);
and U6390 (N_6390,N_4704,N_2989);
or U6391 (N_6391,N_3168,N_3783);
xor U6392 (N_6392,N_4048,N_4228);
xor U6393 (N_6393,N_4079,N_2578);
nor U6394 (N_6394,N_2571,N_2894);
nor U6395 (N_6395,N_3550,N_4115);
xor U6396 (N_6396,N_3298,N_4109);
or U6397 (N_6397,N_2952,N_3005);
nor U6398 (N_6398,N_3699,N_4510);
and U6399 (N_6399,N_3951,N_3051);
or U6400 (N_6400,N_3000,N_4413);
xnor U6401 (N_6401,N_4977,N_4310);
xnor U6402 (N_6402,N_4784,N_2694);
nand U6403 (N_6403,N_2641,N_3505);
nand U6404 (N_6404,N_3505,N_4069);
and U6405 (N_6405,N_2720,N_4496);
xor U6406 (N_6406,N_4911,N_2658);
or U6407 (N_6407,N_4729,N_4663);
xor U6408 (N_6408,N_3711,N_2717);
nor U6409 (N_6409,N_4200,N_2727);
and U6410 (N_6410,N_2683,N_4895);
nand U6411 (N_6411,N_2655,N_4554);
nand U6412 (N_6412,N_4512,N_2667);
or U6413 (N_6413,N_4520,N_3385);
nor U6414 (N_6414,N_2767,N_3000);
and U6415 (N_6415,N_3598,N_3832);
and U6416 (N_6416,N_3010,N_2594);
nand U6417 (N_6417,N_3158,N_3597);
nor U6418 (N_6418,N_4828,N_3602);
or U6419 (N_6419,N_4823,N_3104);
nor U6420 (N_6420,N_2690,N_4948);
xnor U6421 (N_6421,N_4601,N_4031);
nand U6422 (N_6422,N_3938,N_2502);
nor U6423 (N_6423,N_2914,N_4197);
or U6424 (N_6424,N_2827,N_2989);
or U6425 (N_6425,N_3242,N_4652);
and U6426 (N_6426,N_4383,N_3223);
nor U6427 (N_6427,N_4806,N_2835);
or U6428 (N_6428,N_2739,N_4629);
nand U6429 (N_6429,N_2578,N_3518);
or U6430 (N_6430,N_3058,N_3571);
and U6431 (N_6431,N_3847,N_4892);
nor U6432 (N_6432,N_3502,N_2509);
and U6433 (N_6433,N_3575,N_3862);
and U6434 (N_6434,N_2544,N_3824);
and U6435 (N_6435,N_3767,N_2769);
or U6436 (N_6436,N_4204,N_2595);
and U6437 (N_6437,N_3440,N_3203);
nor U6438 (N_6438,N_4048,N_4575);
and U6439 (N_6439,N_4067,N_3483);
or U6440 (N_6440,N_3321,N_4540);
or U6441 (N_6441,N_3886,N_4001);
xnor U6442 (N_6442,N_3821,N_2779);
nor U6443 (N_6443,N_3378,N_2660);
nor U6444 (N_6444,N_2515,N_2706);
nor U6445 (N_6445,N_2775,N_3778);
or U6446 (N_6446,N_4340,N_3395);
nand U6447 (N_6447,N_2902,N_3124);
and U6448 (N_6448,N_3113,N_4973);
nand U6449 (N_6449,N_3766,N_4804);
or U6450 (N_6450,N_3535,N_3888);
and U6451 (N_6451,N_3853,N_3173);
or U6452 (N_6452,N_3969,N_4131);
xnor U6453 (N_6453,N_3083,N_4056);
nand U6454 (N_6454,N_3756,N_3368);
and U6455 (N_6455,N_2625,N_3573);
xnor U6456 (N_6456,N_2889,N_2621);
nor U6457 (N_6457,N_4740,N_3310);
nor U6458 (N_6458,N_3241,N_2853);
nand U6459 (N_6459,N_3816,N_4412);
or U6460 (N_6460,N_2504,N_3525);
nand U6461 (N_6461,N_3074,N_4109);
nor U6462 (N_6462,N_3671,N_3399);
xnor U6463 (N_6463,N_4643,N_4290);
and U6464 (N_6464,N_3457,N_3802);
or U6465 (N_6465,N_4232,N_3265);
nor U6466 (N_6466,N_3316,N_2771);
nand U6467 (N_6467,N_3205,N_4068);
nand U6468 (N_6468,N_3902,N_3449);
nor U6469 (N_6469,N_4497,N_4913);
nand U6470 (N_6470,N_3645,N_2685);
xnor U6471 (N_6471,N_4771,N_3242);
nor U6472 (N_6472,N_2579,N_3890);
and U6473 (N_6473,N_3334,N_4459);
nor U6474 (N_6474,N_4453,N_4472);
nand U6475 (N_6475,N_4048,N_3208);
xor U6476 (N_6476,N_4412,N_4942);
and U6477 (N_6477,N_2508,N_4299);
xor U6478 (N_6478,N_3223,N_4010);
and U6479 (N_6479,N_3141,N_4982);
xor U6480 (N_6480,N_2899,N_4126);
or U6481 (N_6481,N_3861,N_4045);
nor U6482 (N_6482,N_2517,N_4967);
nor U6483 (N_6483,N_3214,N_2561);
and U6484 (N_6484,N_2833,N_4609);
nor U6485 (N_6485,N_4255,N_2798);
nor U6486 (N_6486,N_3033,N_4951);
and U6487 (N_6487,N_2651,N_4320);
and U6488 (N_6488,N_4273,N_3368);
nand U6489 (N_6489,N_3734,N_4646);
xor U6490 (N_6490,N_4405,N_2912);
and U6491 (N_6491,N_2890,N_3151);
or U6492 (N_6492,N_2716,N_2806);
and U6493 (N_6493,N_4567,N_4993);
nand U6494 (N_6494,N_3903,N_3945);
nand U6495 (N_6495,N_4572,N_4614);
nand U6496 (N_6496,N_4725,N_4702);
nor U6497 (N_6497,N_3875,N_2853);
or U6498 (N_6498,N_2575,N_3839);
nand U6499 (N_6499,N_4707,N_4300);
xor U6500 (N_6500,N_3388,N_3841);
and U6501 (N_6501,N_2658,N_3777);
nand U6502 (N_6502,N_4764,N_4507);
xor U6503 (N_6503,N_3750,N_3421);
and U6504 (N_6504,N_4490,N_3245);
nor U6505 (N_6505,N_4610,N_3178);
and U6506 (N_6506,N_4936,N_2731);
or U6507 (N_6507,N_3883,N_2878);
and U6508 (N_6508,N_3884,N_4877);
nand U6509 (N_6509,N_3504,N_4718);
xor U6510 (N_6510,N_3258,N_3121);
xnor U6511 (N_6511,N_3606,N_4237);
and U6512 (N_6512,N_4154,N_4747);
xor U6513 (N_6513,N_4437,N_2676);
and U6514 (N_6514,N_4556,N_3139);
nor U6515 (N_6515,N_4629,N_3441);
nor U6516 (N_6516,N_2841,N_3628);
nor U6517 (N_6517,N_3339,N_3476);
and U6518 (N_6518,N_4331,N_3659);
nand U6519 (N_6519,N_3851,N_2611);
xnor U6520 (N_6520,N_3737,N_4334);
nor U6521 (N_6521,N_4002,N_3337);
xor U6522 (N_6522,N_3833,N_3507);
nand U6523 (N_6523,N_2782,N_2842);
nand U6524 (N_6524,N_2761,N_3041);
or U6525 (N_6525,N_3847,N_2890);
xor U6526 (N_6526,N_4394,N_2534);
xor U6527 (N_6527,N_3386,N_3748);
and U6528 (N_6528,N_2828,N_4500);
and U6529 (N_6529,N_4589,N_2666);
xor U6530 (N_6530,N_3918,N_4329);
or U6531 (N_6531,N_4580,N_4964);
xor U6532 (N_6532,N_2536,N_4026);
nand U6533 (N_6533,N_4859,N_3549);
nor U6534 (N_6534,N_2626,N_4677);
nand U6535 (N_6535,N_4208,N_2923);
or U6536 (N_6536,N_2516,N_4616);
nand U6537 (N_6537,N_4154,N_3288);
or U6538 (N_6538,N_4029,N_4986);
nor U6539 (N_6539,N_4188,N_4312);
or U6540 (N_6540,N_3660,N_3118);
or U6541 (N_6541,N_2966,N_4522);
nor U6542 (N_6542,N_2835,N_3381);
xnor U6543 (N_6543,N_4380,N_3392);
or U6544 (N_6544,N_2506,N_3701);
nor U6545 (N_6545,N_3844,N_4865);
and U6546 (N_6546,N_4939,N_2993);
nor U6547 (N_6547,N_2998,N_3477);
xor U6548 (N_6548,N_3755,N_4184);
nor U6549 (N_6549,N_4258,N_2924);
and U6550 (N_6550,N_2910,N_3868);
nand U6551 (N_6551,N_3819,N_2978);
or U6552 (N_6552,N_3949,N_2742);
xnor U6553 (N_6553,N_4279,N_3336);
nor U6554 (N_6554,N_3265,N_3065);
xnor U6555 (N_6555,N_4414,N_3568);
nor U6556 (N_6556,N_3635,N_2511);
or U6557 (N_6557,N_2842,N_3356);
and U6558 (N_6558,N_3205,N_4263);
xor U6559 (N_6559,N_3478,N_3723);
xnor U6560 (N_6560,N_3657,N_3375);
or U6561 (N_6561,N_3674,N_3787);
nor U6562 (N_6562,N_3861,N_2869);
nand U6563 (N_6563,N_4921,N_4772);
and U6564 (N_6564,N_3794,N_3426);
and U6565 (N_6565,N_4198,N_4440);
nor U6566 (N_6566,N_2505,N_4168);
and U6567 (N_6567,N_4869,N_3619);
xnor U6568 (N_6568,N_4986,N_4375);
nand U6569 (N_6569,N_3642,N_4687);
xor U6570 (N_6570,N_3223,N_4361);
nand U6571 (N_6571,N_3620,N_3430);
nor U6572 (N_6572,N_3477,N_4867);
nand U6573 (N_6573,N_4206,N_2638);
nand U6574 (N_6574,N_3151,N_3851);
nand U6575 (N_6575,N_4228,N_4974);
nor U6576 (N_6576,N_3377,N_3309);
xor U6577 (N_6577,N_3003,N_3486);
nor U6578 (N_6578,N_4194,N_4920);
or U6579 (N_6579,N_3055,N_4272);
nor U6580 (N_6580,N_4163,N_2537);
or U6581 (N_6581,N_4903,N_3616);
or U6582 (N_6582,N_4025,N_3534);
or U6583 (N_6583,N_3241,N_2904);
nor U6584 (N_6584,N_4511,N_4826);
xor U6585 (N_6585,N_4206,N_3243);
xor U6586 (N_6586,N_4119,N_4587);
and U6587 (N_6587,N_4813,N_2817);
xor U6588 (N_6588,N_3786,N_4671);
xnor U6589 (N_6589,N_2902,N_4445);
xnor U6590 (N_6590,N_4681,N_4926);
xnor U6591 (N_6591,N_3399,N_3036);
or U6592 (N_6592,N_4521,N_4626);
and U6593 (N_6593,N_3859,N_2739);
xnor U6594 (N_6594,N_3225,N_3932);
xor U6595 (N_6595,N_4221,N_3630);
nand U6596 (N_6596,N_4726,N_3607);
nor U6597 (N_6597,N_4837,N_4625);
and U6598 (N_6598,N_3872,N_3322);
nand U6599 (N_6599,N_2736,N_3554);
nand U6600 (N_6600,N_2955,N_3145);
or U6601 (N_6601,N_4021,N_2796);
xnor U6602 (N_6602,N_4196,N_4233);
nand U6603 (N_6603,N_2753,N_3733);
xor U6604 (N_6604,N_2743,N_4008);
xor U6605 (N_6605,N_2671,N_4313);
or U6606 (N_6606,N_2909,N_4609);
nand U6607 (N_6607,N_3566,N_2634);
or U6608 (N_6608,N_4279,N_3421);
nor U6609 (N_6609,N_4127,N_2566);
nand U6610 (N_6610,N_4430,N_3289);
and U6611 (N_6611,N_4860,N_3004);
nor U6612 (N_6612,N_4019,N_3484);
nor U6613 (N_6613,N_2556,N_4353);
xnor U6614 (N_6614,N_3565,N_3556);
and U6615 (N_6615,N_2885,N_3743);
xor U6616 (N_6616,N_4474,N_4114);
nand U6617 (N_6617,N_3428,N_3653);
and U6618 (N_6618,N_3420,N_2951);
xnor U6619 (N_6619,N_4391,N_3821);
xnor U6620 (N_6620,N_4749,N_2687);
nor U6621 (N_6621,N_3535,N_4570);
xnor U6622 (N_6622,N_3990,N_4351);
nand U6623 (N_6623,N_4724,N_2796);
xnor U6624 (N_6624,N_2587,N_4935);
xor U6625 (N_6625,N_2738,N_3163);
xnor U6626 (N_6626,N_4780,N_4242);
and U6627 (N_6627,N_3089,N_4360);
xor U6628 (N_6628,N_3933,N_4008);
and U6629 (N_6629,N_2843,N_3519);
nand U6630 (N_6630,N_4112,N_4256);
nor U6631 (N_6631,N_3215,N_2534);
and U6632 (N_6632,N_3046,N_3743);
nand U6633 (N_6633,N_3268,N_4764);
or U6634 (N_6634,N_3850,N_3048);
nor U6635 (N_6635,N_3965,N_3552);
and U6636 (N_6636,N_4173,N_3143);
xnor U6637 (N_6637,N_4660,N_4784);
or U6638 (N_6638,N_4115,N_3275);
or U6639 (N_6639,N_2870,N_2782);
nand U6640 (N_6640,N_4674,N_3683);
and U6641 (N_6641,N_4604,N_2898);
xnor U6642 (N_6642,N_2614,N_3631);
xnor U6643 (N_6643,N_3996,N_3478);
and U6644 (N_6644,N_2955,N_3653);
xor U6645 (N_6645,N_4356,N_4456);
nor U6646 (N_6646,N_3888,N_3053);
and U6647 (N_6647,N_3882,N_4203);
nand U6648 (N_6648,N_3783,N_2921);
nor U6649 (N_6649,N_3839,N_4582);
nand U6650 (N_6650,N_2883,N_4200);
xnor U6651 (N_6651,N_2623,N_4739);
nand U6652 (N_6652,N_4345,N_2777);
xor U6653 (N_6653,N_3046,N_4565);
xor U6654 (N_6654,N_3899,N_2994);
or U6655 (N_6655,N_4087,N_4262);
or U6656 (N_6656,N_3508,N_3135);
or U6657 (N_6657,N_3886,N_2862);
nand U6658 (N_6658,N_4540,N_4133);
xor U6659 (N_6659,N_3008,N_2539);
xor U6660 (N_6660,N_4299,N_3932);
xnor U6661 (N_6661,N_4348,N_4598);
nand U6662 (N_6662,N_3916,N_3865);
or U6663 (N_6663,N_3703,N_4342);
or U6664 (N_6664,N_3416,N_3842);
nand U6665 (N_6665,N_4017,N_3557);
xnor U6666 (N_6666,N_3554,N_4342);
or U6667 (N_6667,N_3056,N_4050);
nand U6668 (N_6668,N_3286,N_2680);
xor U6669 (N_6669,N_4990,N_4490);
nand U6670 (N_6670,N_4876,N_3346);
nor U6671 (N_6671,N_4129,N_3695);
or U6672 (N_6672,N_2988,N_4989);
xor U6673 (N_6673,N_3513,N_2676);
or U6674 (N_6674,N_2500,N_3949);
xnor U6675 (N_6675,N_3689,N_3978);
xor U6676 (N_6676,N_3311,N_3862);
xnor U6677 (N_6677,N_4262,N_2713);
xnor U6678 (N_6678,N_4687,N_4959);
nand U6679 (N_6679,N_2527,N_4574);
nand U6680 (N_6680,N_3342,N_3834);
or U6681 (N_6681,N_4827,N_3168);
xor U6682 (N_6682,N_4288,N_2812);
nor U6683 (N_6683,N_4157,N_4664);
and U6684 (N_6684,N_3353,N_3954);
nand U6685 (N_6685,N_2948,N_4182);
nor U6686 (N_6686,N_4072,N_4356);
xor U6687 (N_6687,N_4960,N_2610);
nand U6688 (N_6688,N_3729,N_4070);
nand U6689 (N_6689,N_2604,N_3491);
nor U6690 (N_6690,N_3776,N_4638);
nand U6691 (N_6691,N_3389,N_3856);
nor U6692 (N_6692,N_3101,N_3467);
nand U6693 (N_6693,N_2681,N_3179);
nand U6694 (N_6694,N_4875,N_3861);
nand U6695 (N_6695,N_3949,N_4636);
xnor U6696 (N_6696,N_4704,N_4273);
nand U6697 (N_6697,N_4435,N_2756);
xnor U6698 (N_6698,N_4863,N_3499);
and U6699 (N_6699,N_3187,N_4823);
xor U6700 (N_6700,N_3439,N_3353);
nand U6701 (N_6701,N_3152,N_4562);
nor U6702 (N_6702,N_3559,N_2896);
nor U6703 (N_6703,N_3796,N_4472);
or U6704 (N_6704,N_2650,N_2789);
nand U6705 (N_6705,N_4191,N_3840);
or U6706 (N_6706,N_4238,N_3036);
xor U6707 (N_6707,N_4303,N_4275);
or U6708 (N_6708,N_3873,N_4470);
and U6709 (N_6709,N_2520,N_4452);
and U6710 (N_6710,N_2766,N_3333);
nand U6711 (N_6711,N_3089,N_4871);
and U6712 (N_6712,N_2844,N_3973);
or U6713 (N_6713,N_4178,N_3915);
xnor U6714 (N_6714,N_2632,N_4412);
xor U6715 (N_6715,N_3878,N_3604);
nor U6716 (N_6716,N_3256,N_4470);
and U6717 (N_6717,N_4041,N_3701);
nor U6718 (N_6718,N_3339,N_4164);
and U6719 (N_6719,N_4907,N_4103);
xnor U6720 (N_6720,N_3314,N_3052);
xnor U6721 (N_6721,N_4135,N_4721);
nor U6722 (N_6722,N_4205,N_2705);
and U6723 (N_6723,N_4991,N_4116);
nand U6724 (N_6724,N_3329,N_3427);
nor U6725 (N_6725,N_4634,N_3573);
nor U6726 (N_6726,N_2753,N_4064);
nor U6727 (N_6727,N_3972,N_4930);
or U6728 (N_6728,N_4588,N_2704);
and U6729 (N_6729,N_3642,N_2755);
or U6730 (N_6730,N_3498,N_3789);
nand U6731 (N_6731,N_3584,N_3236);
or U6732 (N_6732,N_4680,N_2652);
or U6733 (N_6733,N_4504,N_4743);
xor U6734 (N_6734,N_3106,N_3585);
nor U6735 (N_6735,N_4627,N_2521);
or U6736 (N_6736,N_4845,N_2948);
xnor U6737 (N_6737,N_3421,N_3767);
nand U6738 (N_6738,N_4668,N_2595);
nor U6739 (N_6739,N_4866,N_3643);
xnor U6740 (N_6740,N_2735,N_3262);
nor U6741 (N_6741,N_3516,N_4750);
nor U6742 (N_6742,N_2865,N_4529);
or U6743 (N_6743,N_3690,N_3545);
or U6744 (N_6744,N_2910,N_2965);
or U6745 (N_6745,N_4118,N_4573);
nand U6746 (N_6746,N_3934,N_3166);
or U6747 (N_6747,N_3700,N_4252);
nor U6748 (N_6748,N_2687,N_2632);
xor U6749 (N_6749,N_3063,N_4600);
xnor U6750 (N_6750,N_4255,N_4329);
nor U6751 (N_6751,N_2967,N_3415);
and U6752 (N_6752,N_3910,N_2509);
nor U6753 (N_6753,N_3525,N_4089);
nor U6754 (N_6754,N_3324,N_3811);
nor U6755 (N_6755,N_4366,N_3431);
xnor U6756 (N_6756,N_2924,N_4012);
and U6757 (N_6757,N_4601,N_3087);
xor U6758 (N_6758,N_4265,N_2955);
nand U6759 (N_6759,N_4239,N_3310);
xor U6760 (N_6760,N_3451,N_4094);
nand U6761 (N_6761,N_4523,N_4513);
nand U6762 (N_6762,N_2998,N_3880);
xor U6763 (N_6763,N_2932,N_2608);
and U6764 (N_6764,N_2911,N_3382);
nand U6765 (N_6765,N_3198,N_2695);
nand U6766 (N_6766,N_3240,N_2793);
and U6767 (N_6767,N_3437,N_4204);
xnor U6768 (N_6768,N_3918,N_2969);
nor U6769 (N_6769,N_3488,N_4936);
nand U6770 (N_6770,N_4513,N_4790);
and U6771 (N_6771,N_4664,N_3943);
nor U6772 (N_6772,N_3140,N_2651);
nand U6773 (N_6773,N_4949,N_3141);
xor U6774 (N_6774,N_3701,N_4997);
xnor U6775 (N_6775,N_4168,N_3541);
nor U6776 (N_6776,N_3469,N_4463);
and U6777 (N_6777,N_3544,N_4749);
nor U6778 (N_6778,N_4982,N_4337);
nand U6779 (N_6779,N_2798,N_4269);
and U6780 (N_6780,N_3518,N_2562);
and U6781 (N_6781,N_3393,N_3093);
nor U6782 (N_6782,N_4437,N_3609);
and U6783 (N_6783,N_4919,N_3867);
or U6784 (N_6784,N_4519,N_4332);
xnor U6785 (N_6785,N_3607,N_3945);
nand U6786 (N_6786,N_2865,N_4265);
nand U6787 (N_6787,N_3131,N_2577);
xor U6788 (N_6788,N_3183,N_3589);
nor U6789 (N_6789,N_2819,N_3933);
and U6790 (N_6790,N_4109,N_4462);
nor U6791 (N_6791,N_4247,N_3194);
and U6792 (N_6792,N_2734,N_4993);
or U6793 (N_6793,N_3966,N_4542);
xnor U6794 (N_6794,N_2755,N_3496);
and U6795 (N_6795,N_4553,N_2742);
nand U6796 (N_6796,N_4569,N_4720);
nor U6797 (N_6797,N_2837,N_4296);
nor U6798 (N_6798,N_4159,N_3069);
nand U6799 (N_6799,N_4395,N_4997);
nand U6800 (N_6800,N_2618,N_3296);
nand U6801 (N_6801,N_3502,N_4697);
nor U6802 (N_6802,N_2696,N_2800);
nor U6803 (N_6803,N_4797,N_4603);
xnor U6804 (N_6804,N_2964,N_4531);
and U6805 (N_6805,N_3576,N_4381);
and U6806 (N_6806,N_3321,N_4720);
and U6807 (N_6807,N_3955,N_3261);
and U6808 (N_6808,N_4995,N_2559);
xnor U6809 (N_6809,N_2852,N_4330);
or U6810 (N_6810,N_4458,N_3471);
or U6811 (N_6811,N_2947,N_3470);
and U6812 (N_6812,N_4679,N_2660);
and U6813 (N_6813,N_2794,N_3848);
nor U6814 (N_6814,N_4158,N_4650);
or U6815 (N_6815,N_4158,N_2576);
nand U6816 (N_6816,N_4804,N_4560);
nor U6817 (N_6817,N_3507,N_4748);
or U6818 (N_6818,N_4231,N_3633);
xor U6819 (N_6819,N_3894,N_3103);
nand U6820 (N_6820,N_3415,N_4184);
or U6821 (N_6821,N_2776,N_4516);
nand U6822 (N_6822,N_2995,N_3392);
or U6823 (N_6823,N_2592,N_3213);
nor U6824 (N_6824,N_4015,N_2796);
and U6825 (N_6825,N_3542,N_3541);
nand U6826 (N_6826,N_3839,N_4246);
xnor U6827 (N_6827,N_2946,N_3913);
nor U6828 (N_6828,N_3513,N_3059);
and U6829 (N_6829,N_2511,N_4412);
xor U6830 (N_6830,N_4902,N_3615);
and U6831 (N_6831,N_3297,N_3925);
nor U6832 (N_6832,N_3623,N_2659);
and U6833 (N_6833,N_2761,N_3043);
nor U6834 (N_6834,N_2750,N_2518);
or U6835 (N_6835,N_3559,N_3568);
nand U6836 (N_6836,N_4189,N_4524);
nand U6837 (N_6837,N_4502,N_2702);
nor U6838 (N_6838,N_3504,N_3001);
xor U6839 (N_6839,N_2609,N_3934);
xor U6840 (N_6840,N_2977,N_2931);
nor U6841 (N_6841,N_4197,N_2720);
or U6842 (N_6842,N_2833,N_3792);
nand U6843 (N_6843,N_3257,N_4018);
and U6844 (N_6844,N_3820,N_3398);
nor U6845 (N_6845,N_4702,N_2959);
xor U6846 (N_6846,N_3968,N_4033);
xnor U6847 (N_6847,N_3147,N_4288);
nand U6848 (N_6848,N_3389,N_3392);
xor U6849 (N_6849,N_4318,N_3382);
and U6850 (N_6850,N_3329,N_3899);
and U6851 (N_6851,N_4741,N_4126);
or U6852 (N_6852,N_3384,N_3833);
xnor U6853 (N_6853,N_3863,N_3408);
nor U6854 (N_6854,N_2562,N_3406);
xnor U6855 (N_6855,N_2857,N_3084);
nand U6856 (N_6856,N_4300,N_4849);
nand U6857 (N_6857,N_4886,N_4304);
and U6858 (N_6858,N_4132,N_2916);
xnor U6859 (N_6859,N_2530,N_2917);
nand U6860 (N_6860,N_2954,N_3720);
or U6861 (N_6861,N_3030,N_3344);
nor U6862 (N_6862,N_3518,N_3493);
xnor U6863 (N_6863,N_4815,N_3514);
and U6864 (N_6864,N_3241,N_4526);
or U6865 (N_6865,N_2872,N_3245);
nand U6866 (N_6866,N_3001,N_4004);
nor U6867 (N_6867,N_3458,N_2615);
xor U6868 (N_6868,N_2961,N_4286);
nor U6869 (N_6869,N_4690,N_4613);
or U6870 (N_6870,N_2919,N_4771);
xor U6871 (N_6871,N_3368,N_3920);
xor U6872 (N_6872,N_3884,N_2541);
or U6873 (N_6873,N_4806,N_3195);
nor U6874 (N_6874,N_3655,N_4124);
and U6875 (N_6875,N_3031,N_4163);
and U6876 (N_6876,N_3013,N_2776);
or U6877 (N_6877,N_3273,N_4324);
nor U6878 (N_6878,N_3301,N_4169);
nor U6879 (N_6879,N_2780,N_4090);
nand U6880 (N_6880,N_3632,N_4710);
or U6881 (N_6881,N_3497,N_2794);
or U6882 (N_6882,N_3764,N_3110);
or U6883 (N_6883,N_2544,N_3198);
xor U6884 (N_6884,N_4510,N_3277);
nor U6885 (N_6885,N_4252,N_4777);
or U6886 (N_6886,N_3592,N_3684);
xnor U6887 (N_6887,N_4022,N_4890);
nand U6888 (N_6888,N_3400,N_3244);
or U6889 (N_6889,N_3763,N_3550);
or U6890 (N_6890,N_3844,N_2856);
and U6891 (N_6891,N_3865,N_3910);
and U6892 (N_6892,N_3596,N_3525);
nor U6893 (N_6893,N_4051,N_3416);
and U6894 (N_6894,N_3007,N_3381);
and U6895 (N_6895,N_3003,N_3242);
and U6896 (N_6896,N_4008,N_4323);
nand U6897 (N_6897,N_3666,N_4361);
and U6898 (N_6898,N_3711,N_4077);
nand U6899 (N_6899,N_4820,N_4750);
nand U6900 (N_6900,N_3572,N_3627);
and U6901 (N_6901,N_4941,N_3860);
and U6902 (N_6902,N_3244,N_3473);
or U6903 (N_6903,N_3749,N_2699);
xnor U6904 (N_6904,N_2642,N_2715);
xnor U6905 (N_6905,N_3632,N_4429);
and U6906 (N_6906,N_4179,N_2822);
xnor U6907 (N_6907,N_4281,N_3697);
nor U6908 (N_6908,N_3562,N_3153);
or U6909 (N_6909,N_4782,N_3596);
nor U6910 (N_6910,N_4876,N_4434);
nor U6911 (N_6911,N_4302,N_3514);
nor U6912 (N_6912,N_4565,N_4889);
and U6913 (N_6913,N_4792,N_4164);
nand U6914 (N_6914,N_4676,N_2823);
and U6915 (N_6915,N_4133,N_3732);
xor U6916 (N_6916,N_3814,N_4062);
nand U6917 (N_6917,N_3164,N_2876);
and U6918 (N_6918,N_4053,N_2775);
nand U6919 (N_6919,N_4181,N_3687);
and U6920 (N_6920,N_3971,N_4681);
nor U6921 (N_6921,N_3396,N_4169);
nand U6922 (N_6922,N_4431,N_3929);
xor U6923 (N_6923,N_2989,N_3946);
and U6924 (N_6924,N_4844,N_4389);
nand U6925 (N_6925,N_2619,N_4779);
nand U6926 (N_6926,N_4296,N_3420);
and U6927 (N_6927,N_4295,N_3308);
or U6928 (N_6928,N_2881,N_4573);
xnor U6929 (N_6929,N_2836,N_4139);
xor U6930 (N_6930,N_4383,N_4209);
and U6931 (N_6931,N_3603,N_4579);
and U6932 (N_6932,N_4839,N_3720);
or U6933 (N_6933,N_2554,N_3560);
and U6934 (N_6934,N_2517,N_4266);
nor U6935 (N_6935,N_4608,N_3670);
nand U6936 (N_6936,N_4320,N_4948);
nor U6937 (N_6937,N_3500,N_3133);
nor U6938 (N_6938,N_4669,N_4579);
nor U6939 (N_6939,N_3971,N_3002);
and U6940 (N_6940,N_4491,N_3108);
xor U6941 (N_6941,N_3087,N_3716);
nor U6942 (N_6942,N_4348,N_4034);
nand U6943 (N_6943,N_4040,N_3290);
or U6944 (N_6944,N_4981,N_2931);
nor U6945 (N_6945,N_3032,N_3545);
and U6946 (N_6946,N_4629,N_4491);
or U6947 (N_6947,N_4529,N_4616);
nor U6948 (N_6948,N_4858,N_3856);
or U6949 (N_6949,N_4326,N_2752);
nor U6950 (N_6950,N_2751,N_2505);
nand U6951 (N_6951,N_2574,N_4298);
xor U6952 (N_6952,N_4727,N_4450);
nor U6953 (N_6953,N_4870,N_4748);
nand U6954 (N_6954,N_2735,N_3933);
and U6955 (N_6955,N_3255,N_2894);
xnor U6956 (N_6956,N_2796,N_4249);
nand U6957 (N_6957,N_4989,N_3823);
or U6958 (N_6958,N_4894,N_2507);
xnor U6959 (N_6959,N_2632,N_3816);
and U6960 (N_6960,N_4380,N_4182);
or U6961 (N_6961,N_2697,N_2765);
nor U6962 (N_6962,N_4959,N_2915);
nor U6963 (N_6963,N_2587,N_3044);
or U6964 (N_6964,N_4235,N_4254);
nand U6965 (N_6965,N_4074,N_3727);
or U6966 (N_6966,N_3488,N_2513);
nor U6967 (N_6967,N_2665,N_3754);
xnor U6968 (N_6968,N_4718,N_3544);
xnor U6969 (N_6969,N_3895,N_2944);
and U6970 (N_6970,N_3172,N_3561);
nand U6971 (N_6971,N_4401,N_2979);
nor U6972 (N_6972,N_3204,N_3284);
nand U6973 (N_6973,N_3430,N_4596);
xnor U6974 (N_6974,N_4065,N_3853);
nand U6975 (N_6975,N_2650,N_4849);
and U6976 (N_6976,N_4827,N_4094);
nand U6977 (N_6977,N_4765,N_3461);
xnor U6978 (N_6978,N_4510,N_3554);
and U6979 (N_6979,N_2550,N_3463);
or U6980 (N_6980,N_4935,N_3105);
xor U6981 (N_6981,N_3483,N_4851);
and U6982 (N_6982,N_4932,N_2711);
xor U6983 (N_6983,N_3311,N_4623);
nor U6984 (N_6984,N_4183,N_4319);
nand U6985 (N_6985,N_3158,N_4528);
xnor U6986 (N_6986,N_4151,N_4277);
xor U6987 (N_6987,N_4457,N_3571);
or U6988 (N_6988,N_2970,N_2555);
nor U6989 (N_6989,N_4050,N_4206);
xnor U6990 (N_6990,N_2793,N_3033);
xnor U6991 (N_6991,N_4842,N_4195);
nor U6992 (N_6992,N_2997,N_3337);
nand U6993 (N_6993,N_2807,N_4754);
nand U6994 (N_6994,N_3961,N_4487);
xnor U6995 (N_6995,N_3066,N_2647);
xor U6996 (N_6996,N_4850,N_4035);
and U6997 (N_6997,N_3300,N_3523);
nand U6998 (N_6998,N_4631,N_2743);
nand U6999 (N_6999,N_3497,N_2970);
nor U7000 (N_7000,N_4131,N_4209);
nor U7001 (N_7001,N_4526,N_3065);
and U7002 (N_7002,N_4927,N_3138);
xor U7003 (N_7003,N_2945,N_3461);
and U7004 (N_7004,N_2544,N_4569);
xor U7005 (N_7005,N_4535,N_3565);
nand U7006 (N_7006,N_3821,N_3748);
xor U7007 (N_7007,N_4406,N_3569);
nand U7008 (N_7008,N_3615,N_3811);
or U7009 (N_7009,N_2944,N_3346);
and U7010 (N_7010,N_4069,N_4281);
and U7011 (N_7011,N_2830,N_3521);
nor U7012 (N_7012,N_2661,N_3779);
and U7013 (N_7013,N_4783,N_4099);
nand U7014 (N_7014,N_3324,N_2713);
xnor U7015 (N_7015,N_3734,N_3715);
nor U7016 (N_7016,N_3071,N_2536);
xor U7017 (N_7017,N_4449,N_4677);
and U7018 (N_7018,N_4159,N_3182);
nor U7019 (N_7019,N_3346,N_3918);
xor U7020 (N_7020,N_4966,N_3401);
or U7021 (N_7021,N_4086,N_4020);
nand U7022 (N_7022,N_3991,N_4485);
nand U7023 (N_7023,N_3884,N_4172);
xor U7024 (N_7024,N_3515,N_3653);
nor U7025 (N_7025,N_3941,N_3218);
and U7026 (N_7026,N_2615,N_2724);
nor U7027 (N_7027,N_3527,N_2865);
xnor U7028 (N_7028,N_4461,N_3766);
nand U7029 (N_7029,N_3534,N_3824);
nor U7030 (N_7030,N_4527,N_2560);
and U7031 (N_7031,N_2521,N_4305);
nor U7032 (N_7032,N_3813,N_3220);
and U7033 (N_7033,N_3651,N_4179);
xor U7034 (N_7034,N_3354,N_2921);
and U7035 (N_7035,N_3128,N_4983);
nand U7036 (N_7036,N_4277,N_4607);
xor U7037 (N_7037,N_4288,N_4330);
nor U7038 (N_7038,N_3134,N_3247);
nand U7039 (N_7039,N_2614,N_4227);
nand U7040 (N_7040,N_4101,N_4956);
nor U7041 (N_7041,N_4058,N_3104);
or U7042 (N_7042,N_4154,N_4806);
nand U7043 (N_7043,N_4746,N_4155);
or U7044 (N_7044,N_4281,N_3155);
and U7045 (N_7045,N_3689,N_3926);
and U7046 (N_7046,N_3805,N_3961);
xnor U7047 (N_7047,N_4107,N_4705);
nand U7048 (N_7048,N_2509,N_3401);
and U7049 (N_7049,N_4992,N_2766);
nor U7050 (N_7050,N_4915,N_4524);
and U7051 (N_7051,N_3658,N_4528);
or U7052 (N_7052,N_3204,N_4500);
or U7053 (N_7053,N_3683,N_3580);
nand U7054 (N_7054,N_4000,N_4245);
and U7055 (N_7055,N_4454,N_2531);
or U7056 (N_7056,N_4841,N_4589);
or U7057 (N_7057,N_4705,N_4185);
xor U7058 (N_7058,N_4553,N_4080);
xnor U7059 (N_7059,N_3327,N_3069);
nand U7060 (N_7060,N_3572,N_3879);
or U7061 (N_7061,N_4723,N_2551);
or U7062 (N_7062,N_3063,N_4993);
and U7063 (N_7063,N_4918,N_2943);
and U7064 (N_7064,N_4800,N_2926);
and U7065 (N_7065,N_3153,N_4599);
or U7066 (N_7066,N_3078,N_4797);
and U7067 (N_7067,N_2836,N_4068);
and U7068 (N_7068,N_3597,N_2505);
xnor U7069 (N_7069,N_4093,N_2901);
nand U7070 (N_7070,N_3189,N_3419);
and U7071 (N_7071,N_3459,N_2899);
and U7072 (N_7072,N_4877,N_3446);
xor U7073 (N_7073,N_3739,N_4431);
nor U7074 (N_7074,N_3169,N_3851);
or U7075 (N_7075,N_4035,N_4762);
or U7076 (N_7076,N_3120,N_3228);
xor U7077 (N_7077,N_3669,N_2629);
nor U7078 (N_7078,N_3620,N_3776);
nor U7079 (N_7079,N_4420,N_3426);
xnor U7080 (N_7080,N_2942,N_3394);
and U7081 (N_7081,N_3835,N_3075);
nand U7082 (N_7082,N_3662,N_3923);
or U7083 (N_7083,N_3707,N_4115);
xor U7084 (N_7084,N_2647,N_4539);
nand U7085 (N_7085,N_2913,N_3012);
nor U7086 (N_7086,N_4958,N_3865);
nand U7087 (N_7087,N_4647,N_4377);
and U7088 (N_7088,N_2523,N_3102);
xor U7089 (N_7089,N_3519,N_3184);
nor U7090 (N_7090,N_3412,N_4043);
or U7091 (N_7091,N_2921,N_3718);
nor U7092 (N_7092,N_3339,N_4808);
and U7093 (N_7093,N_3749,N_2840);
or U7094 (N_7094,N_3867,N_4182);
xor U7095 (N_7095,N_3247,N_3943);
nor U7096 (N_7096,N_2895,N_3237);
and U7097 (N_7097,N_4396,N_4562);
xor U7098 (N_7098,N_4768,N_4407);
and U7099 (N_7099,N_3775,N_2925);
nor U7100 (N_7100,N_3211,N_3946);
nand U7101 (N_7101,N_4939,N_4341);
xor U7102 (N_7102,N_3951,N_4130);
nand U7103 (N_7103,N_3637,N_3629);
nand U7104 (N_7104,N_3284,N_2730);
or U7105 (N_7105,N_4830,N_4381);
nor U7106 (N_7106,N_3972,N_4191);
nand U7107 (N_7107,N_3155,N_4082);
nor U7108 (N_7108,N_3928,N_4283);
nor U7109 (N_7109,N_4708,N_3207);
xor U7110 (N_7110,N_2760,N_3874);
or U7111 (N_7111,N_3809,N_4780);
nor U7112 (N_7112,N_3565,N_3122);
nand U7113 (N_7113,N_4235,N_4430);
xnor U7114 (N_7114,N_4785,N_3616);
xor U7115 (N_7115,N_2740,N_3445);
and U7116 (N_7116,N_4199,N_4208);
nor U7117 (N_7117,N_4949,N_4907);
nand U7118 (N_7118,N_4866,N_3355);
xnor U7119 (N_7119,N_3886,N_2922);
xor U7120 (N_7120,N_4256,N_3903);
or U7121 (N_7121,N_4528,N_3700);
nor U7122 (N_7122,N_4887,N_4684);
and U7123 (N_7123,N_4819,N_3501);
nor U7124 (N_7124,N_4806,N_2986);
xor U7125 (N_7125,N_2676,N_2514);
and U7126 (N_7126,N_3499,N_2694);
or U7127 (N_7127,N_3258,N_4003);
and U7128 (N_7128,N_2811,N_3747);
xnor U7129 (N_7129,N_2657,N_2697);
nand U7130 (N_7130,N_3847,N_4361);
or U7131 (N_7131,N_4451,N_4408);
nor U7132 (N_7132,N_2778,N_3044);
xor U7133 (N_7133,N_4275,N_3864);
nor U7134 (N_7134,N_4978,N_2798);
and U7135 (N_7135,N_4814,N_3762);
xnor U7136 (N_7136,N_4314,N_3240);
and U7137 (N_7137,N_4724,N_4160);
xnor U7138 (N_7138,N_4718,N_3620);
nor U7139 (N_7139,N_3334,N_3647);
nor U7140 (N_7140,N_4406,N_4346);
nor U7141 (N_7141,N_3883,N_4491);
nand U7142 (N_7142,N_3818,N_3999);
nor U7143 (N_7143,N_3739,N_3126);
nand U7144 (N_7144,N_4254,N_3444);
xnor U7145 (N_7145,N_3751,N_3847);
or U7146 (N_7146,N_3704,N_4931);
nor U7147 (N_7147,N_4278,N_4766);
nand U7148 (N_7148,N_2758,N_4629);
or U7149 (N_7149,N_4126,N_3204);
or U7150 (N_7150,N_4670,N_3028);
nand U7151 (N_7151,N_2757,N_2501);
nand U7152 (N_7152,N_3247,N_3256);
nand U7153 (N_7153,N_3251,N_3512);
or U7154 (N_7154,N_3925,N_4601);
nor U7155 (N_7155,N_4279,N_2717);
nor U7156 (N_7156,N_3087,N_4215);
or U7157 (N_7157,N_3060,N_3331);
nor U7158 (N_7158,N_3713,N_3652);
nor U7159 (N_7159,N_4136,N_3677);
xor U7160 (N_7160,N_4664,N_2586);
nor U7161 (N_7161,N_2719,N_3649);
nand U7162 (N_7162,N_4397,N_3599);
nor U7163 (N_7163,N_2814,N_3912);
nand U7164 (N_7164,N_3054,N_2798);
nand U7165 (N_7165,N_3316,N_2603);
or U7166 (N_7166,N_4584,N_3632);
nand U7167 (N_7167,N_3377,N_3128);
xor U7168 (N_7168,N_4206,N_2967);
nand U7169 (N_7169,N_3371,N_3259);
nor U7170 (N_7170,N_4250,N_4946);
xor U7171 (N_7171,N_3215,N_4061);
or U7172 (N_7172,N_3146,N_4618);
nand U7173 (N_7173,N_3215,N_3963);
nor U7174 (N_7174,N_3574,N_2827);
and U7175 (N_7175,N_3819,N_2715);
and U7176 (N_7176,N_4308,N_2842);
xnor U7177 (N_7177,N_3037,N_3227);
or U7178 (N_7178,N_3900,N_3514);
nor U7179 (N_7179,N_2871,N_2795);
xor U7180 (N_7180,N_4691,N_3050);
and U7181 (N_7181,N_3076,N_2577);
or U7182 (N_7182,N_3621,N_4610);
nand U7183 (N_7183,N_3536,N_3915);
nand U7184 (N_7184,N_4568,N_2906);
or U7185 (N_7185,N_2511,N_3618);
or U7186 (N_7186,N_4689,N_2517);
or U7187 (N_7187,N_4552,N_2858);
and U7188 (N_7188,N_4209,N_3638);
xor U7189 (N_7189,N_4850,N_2617);
or U7190 (N_7190,N_3167,N_2724);
nor U7191 (N_7191,N_3404,N_4496);
or U7192 (N_7192,N_2503,N_4167);
and U7193 (N_7193,N_4728,N_2651);
and U7194 (N_7194,N_3146,N_2550);
xor U7195 (N_7195,N_4757,N_3269);
nand U7196 (N_7196,N_4207,N_2762);
nor U7197 (N_7197,N_2529,N_3089);
xnor U7198 (N_7198,N_2576,N_2927);
or U7199 (N_7199,N_3756,N_2818);
nor U7200 (N_7200,N_4623,N_3186);
nor U7201 (N_7201,N_3785,N_3565);
nor U7202 (N_7202,N_4822,N_4171);
and U7203 (N_7203,N_4953,N_3477);
nand U7204 (N_7204,N_4684,N_4555);
nand U7205 (N_7205,N_3716,N_4238);
nor U7206 (N_7206,N_3618,N_4148);
or U7207 (N_7207,N_4825,N_4945);
and U7208 (N_7208,N_3153,N_4914);
xnor U7209 (N_7209,N_2824,N_4971);
and U7210 (N_7210,N_2873,N_2769);
xnor U7211 (N_7211,N_4511,N_2746);
nand U7212 (N_7212,N_2900,N_4053);
xor U7213 (N_7213,N_4676,N_3669);
nand U7214 (N_7214,N_2649,N_3030);
nor U7215 (N_7215,N_2865,N_3841);
and U7216 (N_7216,N_3631,N_2663);
xnor U7217 (N_7217,N_3766,N_4983);
xnor U7218 (N_7218,N_4315,N_4558);
nor U7219 (N_7219,N_2842,N_3432);
nand U7220 (N_7220,N_4232,N_3513);
xor U7221 (N_7221,N_4939,N_2577);
xnor U7222 (N_7222,N_4887,N_4302);
xor U7223 (N_7223,N_4212,N_3967);
or U7224 (N_7224,N_4737,N_3642);
and U7225 (N_7225,N_3295,N_3740);
and U7226 (N_7226,N_2702,N_3233);
and U7227 (N_7227,N_4974,N_2608);
nand U7228 (N_7228,N_4807,N_2735);
nand U7229 (N_7229,N_4005,N_4134);
or U7230 (N_7230,N_3969,N_3461);
and U7231 (N_7231,N_4665,N_4612);
and U7232 (N_7232,N_4081,N_4392);
nor U7233 (N_7233,N_4161,N_3408);
nand U7234 (N_7234,N_4183,N_3727);
and U7235 (N_7235,N_3836,N_3335);
and U7236 (N_7236,N_2902,N_3351);
xor U7237 (N_7237,N_3703,N_3011);
or U7238 (N_7238,N_4167,N_3735);
xnor U7239 (N_7239,N_3098,N_3533);
nor U7240 (N_7240,N_3575,N_3925);
nor U7241 (N_7241,N_4695,N_4656);
or U7242 (N_7242,N_3571,N_3741);
nand U7243 (N_7243,N_4111,N_3541);
nor U7244 (N_7244,N_3773,N_4344);
and U7245 (N_7245,N_3815,N_4070);
and U7246 (N_7246,N_4568,N_2758);
nor U7247 (N_7247,N_2733,N_2812);
xor U7248 (N_7248,N_4565,N_2978);
and U7249 (N_7249,N_4819,N_3866);
or U7250 (N_7250,N_4624,N_4716);
nand U7251 (N_7251,N_2562,N_3222);
or U7252 (N_7252,N_4387,N_2715);
xnor U7253 (N_7253,N_3461,N_4465);
and U7254 (N_7254,N_3165,N_3905);
nor U7255 (N_7255,N_4608,N_3243);
and U7256 (N_7256,N_3783,N_4838);
xor U7257 (N_7257,N_3324,N_2672);
xnor U7258 (N_7258,N_3178,N_2591);
nor U7259 (N_7259,N_4650,N_4717);
or U7260 (N_7260,N_2672,N_3445);
and U7261 (N_7261,N_3425,N_2611);
or U7262 (N_7262,N_4933,N_2548);
nor U7263 (N_7263,N_2588,N_3411);
or U7264 (N_7264,N_3497,N_3200);
xnor U7265 (N_7265,N_3846,N_4449);
and U7266 (N_7266,N_3672,N_4183);
nand U7267 (N_7267,N_2981,N_4764);
or U7268 (N_7268,N_3518,N_3755);
and U7269 (N_7269,N_3668,N_4876);
and U7270 (N_7270,N_4854,N_3690);
and U7271 (N_7271,N_3353,N_3274);
and U7272 (N_7272,N_4414,N_4415);
or U7273 (N_7273,N_2968,N_3682);
xor U7274 (N_7274,N_3388,N_2690);
and U7275 (N_7275,N_4608,N_3885);
and U7276 (N_7276,N_3359,N_3363);
xnor U7277 (N_7277,N_4665,N_2536);
nor U7278 (N_7278,N_4755,N_2711);
nand U7279 (N_7279,N_3695,N_3305);
and U7280 (N_7280,N_4698,N_4294);
or U7281 (N_7281,N_4053,N_2599);
nand U7282 (N_7282,N_3437,N_4833);
nand U7283 (N_7283,N_2609,N_2735);
nor U7284 (N_7284,N_3185,N_3439);
or U7285 (N_7285,N_2991,N_2890);
or U7286 (N_7286,N_2927,N_4902);
and U7287 (N_7287,N_4263,N_4985);
and U7288 (N_7288,N_4468,N_4319);
and U7289 (N_7289,N_2971,N_3519);
nand U7290 (N_7290,N_4736,N_3736);
and U7291 (N_7291,N_3804,N_2693);
or U7292 (N_7292,N_4141,N_3620);
xor U7293 (N_7293,N_3291,N_3992);
or U7294 (N_7294,N_3738,N_4489);
xnor U7295 (N_7295,N_4839,N_2860);
and U7296 (N_7296,N_3708,N_4730);
or U7297 (N_7297,N_4862,N_4329);
and U7298 (N_7298,N_3433,N_4954);
nand U7299 (N_7299,N_4904,N_3797);
xor U7300 (N_7300,N_3429,N_2981);
nand U7301 (N_7301,N_3740,N_3528);
nor U7302 (N_7302,N_4496,N_4399);
nor U7303 (N_7303,N_3558,N_3033);
nand U7304 (N_7304,N_2775,N_4302);
nand U7305 (N_7305,N_3398,N_4939);
nand U7306 (N_7306,N_4615,N_4399);
xor U7307 (N_7307,N_4797,N_3203);
nor U7308 (N_7308,N_4791,N_4764);
and U7309 (N_7309,N_3503,N_4592);
and U7310 (N_7310,N_2849,N_4581);
xnor U7311 (N_7311,N_3099,N_2523);
nor U7312 (N_7312,N_4093,N_4321);
and U7313 (N_7313,N_2708,N_3761);
xnor U7314 (N_7314,N_4701,N_4990);
and U7315 (N_7315,N_4133,N_3379);
or U7316 (N_7316,N_4889,N_3948);
and U7317 (N_7317,N_3465,N_4487);
xnor U7318 (N_7318,N_3529,N_4517);
or U7319 (N_7319,N_4369,N_3970);
or U7320 (N_7320,N_4348,N_4674);
xor U7321 (N_7321,N_3314,N_4502);
xnor U7322 (N_7322,N_3769,N_3671);
nor U7323 (N_7323,N_3155,N_2698);
or U7324 (N_7324,N_2967,N_4368);
nor U7325 (N_7325,N_3001,N_3527);
xnor U7326 (N_7326,N_4745,N_3459);
nor U7327 (N_7327,N_3903,N_3675);
or U7328 (N_7328,N_3447,N_4855);
nand U7329 (N_7329,N_2822,N_3145);
nor U7330 (N_7330,N_4010,N_3258);
and U7331 (N_7331,N_4367,N_4190);
xnor U7332 (N_7332,N_2751,N_2674);
nand U7333 (N_7333,N_4448,N_4395);
and U7334 (N_7334,N_3268,N_2625);
nor U7335 (N_7335,N_3014,N_3447);
nor U7336 (N_7336,N_4516,N_4446);
nor U7337 (N_7337,N_3583,N_4815);
nand U7338 (N_7338,N_2733,N_4993);
nor U7339 (N_7339,N_3699,N_3907);
nor U7340 (N_7340,N_2720,N_3545);
nand U7341 (N_7341,N_2542,N_2791);
or U7342 (N_7342,N_4355,N_2844);
nor U7343 (N_7343,N_3050,N_3499);
or U7344 (N_7344,N_3836,N_4929);
xor U7345 (N_7345,N_3424,N_3120);
xnor U7346 (N_7346,N_4798,N_4943);
and U7347 (N_7347,N_4773,N_2823);
nor U7348 (N_7348,N_2767,N_4194);
nand U7349 (N_7349,N_4030,N_3070);
nor U7350 (N_7350,N_3908,N_4615);
and U7351 (N_7351,N_3738,N_4281);
nor U7352 (N_7352,N_4819,N_2756);
nor U7353 (N_7353,N_4157,N_3673);
or U7354 (N_7354,N_3278,N_4316);
nor U7355 (N_7355,N_2794,N_2899);
and U7356 (N_7356,N_3254,N_3242);
and U7357 (N_7357,N_4860,N_4405);
nand U7358 (N_7358,N_4964,N_3457);
nand U7359 (N_7359,N_3581,N_4281);
or U7360 (N_7360,N_3399,N_3130);
and U7361 (N_7361,N_4130,N_4924);
or U7362 (N_7362,N_4684,N_4876);
or U7363 (N_7363,N_4743,N_4421);
nor U7364 (N_7364,N_4764,N_4740);
or U7365 (N_7365,N_4276,N_4804);
xor U7366 (N_7366,N_4297,N_3682);
nand U7367 (N_7367,N_4731,N_4617);
nor U7368 (N_7368,N_3652,N_2900);
nor U7369 (N_7369,N_4328,N_4589);
xor U7370 (N_7370,N_4865,N_4972);
or U7371 (N_7371,N_4319,N_3321);
nor U7372 (N_7372,N_4685,N_3722);
nand U7373 (N_7373,N_2507,N_4095);
nand U7374 (N_7374,N_4803,N_3794);
and U7375 (N_7375,N_2773,N_2594);
or U7376 (N_7376,N_3001,N_2585);
or U7377 (N_7377,N_3395,N_4571);
or U7378 (N_7378,N_4221,N_2603);
nor U7379 (N_7379,N_2709,N_2644);
and U7380 (N_7380,N_3312,N_2868);
nand U7381 (N_7381,N_3813,N_4083);
and U7382 (N_7382,N_4010,N_2866);
and U7383 (N_7383,N_3616,N_4993);
and U7384 (N_7384,N_3581,N_4684);
nor U7385 (N_7385,N_2705,N_4290);
nor U7386 (N_7386,N_4771,N_3001);
nor U7387 (N_7387,N_4889,N_3386);
or U7388 (N_7388,N_3360,N_4067);
xnor U7389 (N_7389,N_2737,N_4219);
nand U7390 (N_7390,N_4848,N_2746);
and U7391 (N_7391,N_4714,N_2921);
or U7392 (N_7392,N_2847,N_3954);
and U7393 (N_7393,N_2671,N_4677);
nand U7394 (N_7394,N_2512,N_4372);
or U7395 (N_7395,N_3641,N_3442);
or U7396 (N_7396,N_3214,N_4185);
and U7397 (N_7397,N_3398,N_2961);
nor U7398 (N_7398,N_4905,N_4126);
xnor U7399 (N_7399,N_3893,N_3268);
nor U7400 (N_7400,N_4111,N_2765);
nor U7401 (N_7401,N_3208,N_2592);
nand U7402 (N_7402,N_3584,N_3287);
xor U7403 (N_7403,N_4560,N_4095);
and U7404 (N_7404,N_3591,N_4276);
nand U7405 (N_7405,N_2527,N_4404);
or U7406 (N_7406,N_3184,N_3336);
nor U7407 (N_7407,N_4100,N_3826);
nand U7408 (N_7408,N_4398,N_3209);
nand U7409 (N_7409,N_3422,N_3880);
nand U7410 (N_7410,N_4282,N_4810);
xnor U7411 (N_7411,N_4063,N_3171);
nand U7412 (N_7412,N_3299,N_3988);
and U7413 (N_7413,N_3290,N_3805);
nand U7414 (N_7414,N_2718,N_3779);
and U7415 (N_7415,N_2748,N_2672);
nor U7416 (N_7416,N_2883,N_4919);
or U7417 (N_7417,N_2851,N_3606);
nand U7418 (N_7418,N_3828,N_3537);
nor U7419 (N_7419,N_3248,N_3932);
nor U7420 (N_7420,N_3222,N_4775);
and U7421 (N_7421,N_3843,N_2652);
and U7422 (N_7422,N_3340,N_2647);
and U7423 (N_7423,N_4734,N_3927);
nor U7424 (N_7424,N_3296,N_4813);
and U7425 (N_7425,N_3644,N_3523);
nand U7426 (N_7426,N_4882,N_4731);
nand U7427 (N_7427,N_3888,N_4824);
and U7428 (N_7428,N_3101,N_4342);
and U7429 (N_7429,N_3901,N_2512);
nor U7430 (N_7430,N_4464,N_4522);
nand U7431 (N_7431,N_2927,N_2506);
xor U7432 (N_7432,N_3926,N_3362);
or U7433 (N_7433,N_4647,N_4616);
nand U7434 (N_7434,N_3760,N_4442);
nand U7435 (N_7435,N_3371,N_3311);
nand U7436 (N_7436,N_3666,N_4749);
nand U7437 (N_7437,N_3526,N_2579);
nor U7438 (N_7438,N_4805,N_3777);
nor U7439 (N_7439,N_3951,N_3375);
xnor U7440 (N_7440,N_3494,N_3080);
and U7441 (N_7441,N_3986,N_4304);
nor U7442 (N_7442,N_2568,N_3908);
nor U7443 (N_7443,N_4136,N_4984);
nor U7444 (N_7444,N_3637,N_3245);
nand U7445 (N_7445,N_4031,N_3461);
or U7446 (N_7446,N_4485,N_3395);
xnor U7447 (N_7447,N_4395,N_3486);
nor U7448 (N_7448,N_2655,N_3140);
nand U7449 (N_7449,N_4702,N_3467);
or U7450 (N_7450,N_4327,N_4638);
xor U7451 (N_7451,N_4368,N_2673);
and U7452 (N_7452,N_4120,N_3654);
xor U7453 (N_7453,N_3327,N_3388);
or U7454 (N_7454,N_3331,N_3699);
and U7455 (N_7455,N_4437,N_2980);
or U7456 (N_7456,N_3252,N_3371);
and U7457 (N_7457,N_3728,N_3451);
or U7458 (N_7458,N_4265,N_4974);
and U7459 (N_7459,N_3030,N_3712);
nor U7460 (N_7460,N_2545,N_4419);
or U7461 (N_7461,N_2627,N_4038);
xor U7462 (N_7462,N_3571,N_4273);
nor U7463 (N_7463,N_2531,N_2676);
nor U7464 (N_7464,N_4797,N_3236);
nand U7465 (N_7465,N_4746,N_4866);
xor U7466 (N_7466,N_3150,N_3952);
nor U7467 (N_7467,N_3033,N_4444);
or U7468 (N_7468,N_2990,N_2614);
and U7469 (N_7469,N_4080,N_4513);
or U7470 (N_7470,N_2581,N_2995);
and U7471 (N_7471,N_3042,N_2910);
nor U7472 (N_7472,N_3342,N_4222);
nand U7473 (N_7473,N_3746,N_3922);
and U7474 (N_7474,N_4242,N_3305);
nor U7475 (N_7475,N_3037,N_3672);
xor U7476 (N_7476,N_4391,N_4056);
xnor U7477 (N_7477,N_3961,N_3552);
nor U7478 (N_7478,N_2789,N_4762);
or U7479 (N_7479,N_2895,N_3191);
nand U7480 (N_7480,N_3387,N_2888);
or U7481 (N_7481,N_4337,N_3345);
nand U7482 (N_7482,N_2752,N_3839);
nor U7483 (N_7483,N_3765,N_4425);
nand U7484 (N_7484,N_3229,N_2953);
nand U7485 (N_7485,N_3397,N_4121);
nor U7486 (N_7486,N_4246,N_4711);
or U7487 (N_7487,N_3485,N_3305);
nand U7488 (N_7488,N_2994,N_2982);
nor U7489 (N_7489,N_4111,N_4562);
xor U7490 (N_7490,N_4817,N_4287);
nor U7491 (N_7491,N_3274,N_2618);
or U7492 (N_7492,N_3888,N_2972);
and U7493 (N_7493,N_4537,N_4147);
or U7494 (N_7494,N_4291,N_4095);
xnor U7495 (N_7495,N_3484,N_3930);
xnor U7496 (N_7496,N_2588,N_3667);
and U7497 (N_7497,N_3944,N_2733);
nor U7498 (N_7498,N_3612,N_3559);
nand U7499 (N_7499,N_2857,N_3647);
nand U7500 (N_7500,N_6810,N_5673);
nor U7501 (N_7501,N_5569,N_7280);
or U7502 (N_7502,N_6325,N_5026);
and U7503 (N_7503,N_7407,N_5722);
nand U7504 (N_7504,N_5980,N_7394);
and U7505 (N_7505,N_6474,N_7140);
xor U7506 (N_7506,N_7341,N_6735);
xnor U7507 (N_7507,N_6676,N_7127);
and U7508 (N_7508,N_5140,N_6523);
or U7509 (N_7509,N_6637,N_5446);
xor U7510 (N_7510,N_7314,N_6576);
nand U7511 (N_7511,N_6538,N_5636);
nand U7512 (N_7512,N_6989,N_6135);
nand U7513 (N_7513,N_6387,N_5715);
xnor U7514 (N_7514,N_7091,N_6549);
nand U7515 (N_7515,N_6980,N_5575);
nand U7516 (N_7516,N_7068,N_6867);
xnor U7517 (N_7517,N_5764,N_6361);
and U7518 (N_7518,N_7219,N_5330);
nand U7519 (N_7519,N_5899,N_6636);
nand U7520 (N_7520,N_6746,N_6555);
xnor U7521 (N_7521,N_5107,N_5091);
nor U7522 (N_7522,N_5783,N_7398);
and U7523 (N_7523,N_6578,N_5061);
xor U7524 (N_7524,N_6440,N_6318);
and U7525 (N_7525,N_5676,N_5336);
and U7526 (N_7526,N_6109,N_6292);
or U7527 (N_7527,N_7387,N_5317);
nor U7528 (N_7528,N_5025,N_6048);
or U7529 (N_7529,N_7285,N_5931);
or U7530 (N_7530,N_7049,N_6221);
or U7531 (N_7531,N_6525,N_6872);
and U7532 (N_7532,N_5611,N_7082);
nor U7533 (N_7533,N_5641,N_5349);
nand U7534 (N_7534,N_5697,N_6967);
or U7535 (N_7535,N_6428,N_6897);
and U7536 (N_7536,N_5406,N_5017);
and U7537 (N_7537,N_5364,N_6561);
nand U7538 (N_7538,N_5370,N_6698);
or U7539 (N_7539,N_6899,N_6548);
xor U7540 (N_7540,N_5066,N_6353);
nor U7541 (N_7541,N_6700,N_5344);
or U7542 (N_7542,N_5958,N_5634);
nor U7543 (N_7543,N_5982,N_7184);
and U7544 (N_7544,N_6058,N_7443);
nand U7545 (N_7545,N_5795,N_5933);
nand U7546 (N_7546,N_7456,N_6130);
or U7547 (N_7547,N_6757,N_6365);
or U7548 (N_7548,N_7470,N_6328);
nor U7549 (N_7549,N_6175,N_5886);
nor U7550 (N_7550,N_6953,N_5721);
xor U7551 (N_7551,N_5667,N_5918);
xnor U7552 (N_7552,N_5837,N_6044);
or U7553 (N_7553,N_6028,N_5964);
and U7554 (N_7554,N_7332,N_5038);
or U7555 (N_7555,N_6189,N_5591);
xor U7556 (N_7556,N_6117,N_5099);
xor U7557 (N_7557,N_6783,N_5490);
or U7558 (N_7558,N_5741,N_6624);
and U7559 (N_7559,N_6139,N_6784);
nor U7560 (N_7560,N_6731,N_5503);
nand U7561 (N_7561,N_6808,N_5170);
or U7562 (N_7562,N_6707,N_5206);
or U7563 (N_7563,N_5421,N_5102);
and U7564 (N_7564,N_6644,N_6078);
or U7565 (N_7565,N_5515,N_5513);
or U7566 (N_7566,N_7324,N_7196);
xor U7567 (N_7567,N_6686,N_5160);
xnor U7568 (N_7568,N_7411,N_7263);
nand U7569 (N_7569,N_7180,N_5353);
nand U7570 (N_7570,N_5689,N_6488);
xnor U7571 (N_7571,N_5560,N_7273);
or U7572 (N_7572,N_5050,N_7118);
or U7573 (N_7573,N_6569,N_6478);
nor U7574 (N_7574,N_5435,N_5523);
nand U7575 (N_7575,N_6815,N_5376);
or U7576 (N_7576,N_5028,N_5031);
nand U7577 (N_7577,N_6640,N_7017);
or U7578 (N_7578,N_5557,N_5599);
and U7579 (N_7579,N_5529,N_7120);
nand U7580 (N_7580,N_5694,N_5766);
or U7581 (N_7581,N_7141,N_6678);
or U7582 (N_7582,N_7201,N_5022);
nor U7583 (N_7583,N_6094,N_6276);
xor U7584 (N_7584,N_6055,N_6579);
nand U7585 (N_7585,N_6209,N_7087);
xnor U7586 (N_7586,N_5105,N_5930);
and U7587 (N_7587,N_6881,N_7464);
xor U7588 (N_7588,N_5462,N_7230);
and U7589 (N_7589,N_5765,N_6661);
nand U7590 (N_7590,N_7137,N_5583);
nand U7591 (N_7591,N_6312,N_6880);
nand U7592 (N_7592,N_5302,N_5554);
nor U7593 (N_7593,N_7382,N_6616);
xnor U7594 (N_7594,N_6900,N_5112);
xnor U7595 (N_7595,N_5073,N_5094);
nand U7596 (N_7596,N_6649,N_5185);
and U7597 (N_7597,N_6740,N_6546);
nand U7598 (N_7598,N_6340,N_5171);
nor U7599 (N_7599,N_6412,N_6211);
xnor U7600 (N_7600,N_6539,N_7028);
or U7601 (N_7601,N_5922,N_6823);
and U7602 (N_7602,N_5772,N_5954);
nand U7603 (N_7603,N_6030,N_7298);
and U7604 (N_7604,N_5823,N_7401);
xnor U7605 (N_7605,N_7089,N_7156);
and U7606 (N_7606,N_5374,N_7154);
xnor U7607 (N_7607,N_6051,N_5324);
or U7608 (N_7608,N_5100,N_6775);
nor U7609 (N_7609,N_6876,N_7258);
and U7610 (N_7610,N_6862,N_7202);
and U7611 (N_7611,N_6490,N_5626);
and U7612 (N_7612,N_6970,N_5287);
nand U7613 (N_7613,N_6090,N_7211);
or U7614 (N_7614,N_5145,N_5834);
and U7615 (N_7615,N_6527,N_6992);
nor U7616 (N_7616,N_7374,N_5419);
xor U7617 (N_7617,N_6948,N_6036);
nand U7618 (N_7618,N_5769,N_7316);
nand U7619 (N_7619,N_5427,N_5447);
xor U7620 (N_7620,N_7397,N_5276);
nor U7621 (N_7621,N_6151,N_5904);
or U7622 (N_7622,N_7376,N_5104);
nand U7623 (N_7623,N_5985,N_5008);
nand U7624 (N_7624,N_6081,N_7418);
or U7625 (N_7625,N_5870,N_6057);
or U7626 (N_7626,N_7479,N_5361);
or U7627 (N_7627,N_6356,N_6766);
nor U7628 (N_7628,N_7060,N_6760);
or U7629 (N_7629,N_7023,N_6973);
or U7630 (N_7630,N_5572,N_6886);
and U7631 (N_7631,N_6242,N_6213);
xor U7632 (N_7632,N_6960,N_5144);
nor U7633 (N_7633,N_5563,N_6714);
and U7634 (N_7634,N_6289,N_6215);
or U7635 (N_7635,N_7168,N_6153);
and U7636 (N_7636,N_5113,N_6482);
and U7637 (N_7637,N_6080,N_6227);
nor U7638 (N_7638,N_7099,N_7182);
nor U7639 (N_7639,N_5776,N_6790);
or U7640 (N_7640,N_6988,N_6985);
or U7641 (N_7641,N_5372,N_6866);
or U7642 (N_7642,N_7132,N_7183);
or U7643 (N_7643,N_6912,N_5895);
nor U7644 (N_7644,N_5506,N_6835);
and U7645 (N_7645,N_7352,N_6099);
or U7646 (N_7646,N_7311,N_6620);
xor U7647 (N_7647,N_5040,N_7419);
nand U7648 (N_7648,N_6805,N_7152);
and U7649 (N_7649,N_5258,N_5822);
xnor U7650 (N_7650,N_7414,N_6662);
nor U7651 (N_7651,N_5928,N_6550);
xnor U7652 (N_7652,N_5936,N_5656);
and U7653 (N_7653,N_5538,N_5340);
xor U7654 (N_7654,N_5134,N_5248);
nand U7655 (N_7655,N_6019,N_5015);
and U7656 (N_7656,N_7482,N_6405);
nand U7657 (N_7657,N_6646,N_6319);
xnor U7658 (N_7658,N_5821,N_5130);
nand U7659 (N_7659,N_6481,N_7448);
xor U7660 (N_7660,N_6721,N_7425);
xor U7661 (N_7661,N_6503,N_6241);
and U7662 (N_7662,N_7042,N_5163);
and U7663 (N_7663,N_7217,N_5800);
or U7664 (N_7664,N_5357,N_5830);
nor U7665 (N_7665,N_5345,N_6379);
nor U7666 (N_7666,N_6495,N_5784);
xor U7667 (N_7667,N_5388,N_5927);
or U7668 (N_7668,N_6350,N_5897);
and U7669 (N_7669,N_7383,N_5207);
or U7670 (N_7670,N_5632,N_7244);
and U7671 (N_7671,N_5255,N_5054);
nor U7672 (N_7672,N_6982,N_6339);
nor U7673 (N_7673,N_6123,N_6670);
nand U7674 (N_7674,N_5643,N_7429);
or U7675 (N_7675,N_6372,N_5310);
xor U7676 (N_7676,N_7121,N_6655);
nand U7677 (N_7677,N_6699,N_6924);
xnor U7678 (N_7678,N_7377,N_7058);
nand U7679 (N_7679,N_6929,N_6791);
nand U7680 (N_7680,N_5670,N_5649);
nor U7681 (N_7681,N_7350,N_7021);
nor U7682 (N_7682,N_7150,N_6622);
nand U7683 (N_7683,N_6293,N_6895);
nand U7684 (N_7684,N_5901,N_7436);
or U7685 (N_7685,N_6060,N_5423);
and U7686 (N_7686,N_5270,N_7052);
nand U7687 (N_7687,N_7094,N_5177);
nor U7688 (N_7688,N_5346,N_5146);
nand U7689 (N_7689,N_6681,N_6724);
or U7690 (N_7690,N_5159,N_5035);
nand U7691 (N_7691,N_7103,N_7165);
xnor U7692 (N_7692,N_5459,N_5525);
nand U7693 (N_7693,N_6910,N_6770);
xnor U7694 (N_7694,N_5707,N_7148);
xnor U7695 (N_7695,N_6217,N_5612);
xor U7696 (N_7696,N_7432,N_7162);
nor U7697 (N_7697,N_5095,N_6723);
or U7698 (N_7698,N_5908,N_5751);
nand U7699 (N_7699,N_7122,N_6607);
nand U7700 (N_7700,N_7307,N_7193);
nand U7701 (N_7701,N_7435,N_5812);
or U7702 (N_7702,N_6146,N_7197);
xor U7703 (N_7703,N_6891,N_5963);
or U7704 (N_7704,N_7281,N_6034);
or U7705 (N_7705,N_6167,N_5978);
nor U7706 (N_7706,N_5037,N_6604);
or U7707 (N_7707,N_7430,N_6869);
xnor U7708 (N_7708,N_5023,N_6336);
and U7709 (N_7709,N_6961,N_7093);
nor U7710 (N_7710,N_5524,N_7223);
and U7711 (N_7711,N_6065,N_5631);
and U7712 (N_7712,N_5150,N_6235);
or U7713 (N_7713,N_7337,N_7255);
nand U7714 (N_7714,N_6863,N_5141);
nor U7715 (N_7715,N_6926,N_5905);
xor U7716 (N_7716,N_6202,N_5381);
xor U7717 (N_7717,N_6243,N_5466);
and U7718 (N_7718,N_6377,N_5979);
and U7719 (N_7719,N_5749,N_5573);
and U7720 (N_7720,N_6087,N_5412);
xnor U7721 (N_7721,N_6160,N_7266);
nor U7722 (N_7722,N_7359,N_7420);
nor U7723 (N_7723,N_5120,N_5483);
nand U7724 (N_7724,N_6608,N_5202);
and U7725 (N_7725,N_6126,N_6837);
and U7726 (N_7726,N_5881,N_6934);
nand U7727 (N_7727,N_7050,N_5385);
nor U7728 (N_7728,N_5789,N_5313);
and U7729 (N_7729,N_6291,N_6749);
and U7730 (N_7730,N_5970,N_6868);
and U7731 (N_7731,N_7416,N_7207);
xor U7732 (N_7732,N_5735,N_6422);
nand U7733 (N_7733,N_7031,N_5086);
xor U7734 (N_7734,N_6930,N_6816);
or U7735 (N_7735,N_6819,N_7145);
or U7736 (N_7736,N_5314,N_7380);
and U7737 (N_7737,N_6439,N_5977);
and U7738 (N_7738,N_5873,N_6432);
nor U7739 (N_7739,N_5407,N_6337);
nand U7740 (N_7740,N_6807,N_6609);
nor U7741 (N_7741,N_6580,N_6086);
and U7742 (N_7742,N_6246,N_5953);
or U7743 (N_7743,N_5659,N_5833);
nand U7744 (N_7744,N_5375,N_6716);
and U7745 (N_7745,N_7431,N_6203);
and U7746 (N_7746,N_6951,N_7423);
and U7747 (N_7747,N_7349,N_5685);
and U7748 (N_7748,N_6720,N_6529);
nor U7749 (N_7749,N_7488,N_6403);
nand U7750 (N_7750,N_5485,N_5175);
nor U7751 (N_7751,N_5846,N_5080);
nor U7752 (N_7752,N_7008,N_5477);
nor U7753 (N_7753,N_6586,N_6536);
nor U7754 (N_7754,N_6178,N_6210);
nand U7755 (N_7755,N_7262,N_6730);
nand U7756 (N_7756,N_6769,N_6093);
xor U7757 (N_7757,N_6185,N_5014);
nand U7758 (N_7758,N_6096,N_5530);
or U7759 (N_7759,N_6307,N_6205);
xnor U7760 (N_7760,N_6045,N_5840);
nand U7761 (N_7761,N_6346,N_5131);
or U7762 (N_7762,N_7185,N_6727);
nand U7763 (N_7763,N_7055,N_5859);
nor U7764 (N_7764,N_6174,N_6582);
and U7765 (N_7765,N_6861,N_7459);
xnor U7766 (N_7766,N_6062,N_5536);
nor U7767 (N_7767,N_6283,N_5642);
and U7768 (N_7768,N_6452,N_6925);
xnor U7769 (N_7769,N_5855,N_5083);
and U7770 (N_7770,N_5709,N_5938);
nor U7771 (N_7771,N_5590,N_5373);
nor U7772 (N_7772,N_5829,N_6966);
or U7773 (N_7773,N_5620,N_5706);
xor U7774 (N_7774,N_7417,N_5433);
nand U7775 (N_7775,N_5195,N_5574);
nand U7776 (N_7776,N_7097,N_5016);
xor U7777 (N_7777,N_5497,N_7059);
nand U7778 (N_7778,N_5587,N_5501);
or U7779 (N_7779,N_6944,N_7231);
and U7780 (N_7780,N_5075,N_7393);
and U7781 (N_7781,N_7327,N_6273);
nand U7782 (N_7782,N_5352,N_5168);
xor U7783 (N_7783,N_5174,N_6445);
and U7784 (N_7784,N_6437,N_5096);
nand U7785 (N_7785,N_7191,N_7075);
nand U7786 (N_7786,N_5799,N_7080);
nor U7787 (N_7787,N_6463,N_7354);
nor U7788 (N_7788,N_7379,N_7226);
nand U7789 (N_7789,N_6237,N_5369);
or U7790 (N_7790,N_6214,N_7335);
nand U7791 (N_7791,N_5615,N_6165);
nor U7792 (N_7792,N_6855,N_5520);
and U7793 (N_7793,N_5850,N_6554);
and U7794 (N_7794,N_5937,N_5084);
nand U7795 (N_7795,N_7428,N_7392);
nor U7796 (N_7796,N_6390,N_5186);
nor U7797 (N_7797,N_5955,N_6595);
and U7798 (N_7798,N_5624,N_7493);
and U7799 (N_7799,N_5147,N_6528);
nand U7800 (N_7800,N_6419,N_6804);
nor U7801 (N_7801,N_7025,N_5235);
or U7802 (N_7802,N_7063,N_6193);
xnor U7803 (N_7803,N_6026,N_6141);
nor U7804 (N_7804,N_6994,N_7071);
or U7805 (N_7805,N_6074,N_6476);
and U7806 (N_7806,N_5001,N_5883);
and U7807 (N_7807,N_6706,N_5814);
nand U7808 (N_7808,N_5902,N_5754);
and U7809 (N_7809,N_5876,N_7312);
or U7810 (N_7810,N_5924,N_6679);
xnor U7811 (N_7811,N_7339,N_5951);
xnor U7812 (N_7812,N_6313,N_5909);
nand U7813 (N_7813,N_7208,N_7013);
nand U7814 (N_7814,N_5728,N_5994);
and U7815 (N_7815,N_6611,N_6396);
or U7816 (N_7816,N_5380,N_6279);
nor U7817 (N_7817,N_5191,N_5565);
nand U7818 (N_7818,N_6230,N_6603);
and U7819 (N_7819,N_6460,N_7295);
xnor U7820 (N_7820,N_7471,N_6436);
nand U7821 (N_7821,N_6272,N_6562);
nor U7822 (N_7822,N_5420,N_5097);
xnor U7823 (N_7823,N_7302,N_6913);
xor U7824 (N_7824,N_5041,N_5085);
nor U7825 (N_7825,N_5956,N_5469);
nor U7826 (N_7826,N_7111,N_6635);
xor U7827 (N_7827,N_6471,N_6750);
or U7828 (N_7828,N_6623,N_5705);
or U7829 (N_7829,N_5440,N_5647);
xor U7830 (N_7830,N_5010,N_6889);
and U7831 (N_7831,N_5788,N_5323);
xor U7832 (N_7832,N_5786,N_6564);
xnor U7833 (N_7833,N_6035,N_5853);
xor U7834 (N_7834,N_5983,N_5959);
nand U7835 (N_7835,N_6475,N_7344);
xnor U7836 (N_7836,N_5939,N_7485);
or U7837 (N_7837,N_7402,N_7283);
nand U7838 (N_7838,N_5542,N_6504);
nand U7839 (N_7839,N_6169,N_6263);
nand U7840 (N_7840,N_6088,N_5465);
nor U7841 (N_7841,N_7495,N_5377);
or U7842 (N_7842,N_6903,N_5960);
xor U7843 (N_7843,N_5334,N_5681);
nand U7844 (N_7844,N_6306,N_6113);
or U7845 (N_7845,N_5657,N_6414);
nand U7846 (N_7846,N_5032,N_6752);
nand U7847 (N_7847,N_6887,N_6736);
and U7848 (N_7848,N_7483,N_6505);
nand U7849 (N_7849,N_5819,N_6589);
xor U7850 (N_7850,N_5582,N_5318);
or U7851 (N_7851,N_6812,N_6741);
nor U7852 (N_7852,N_5121,N_6309);
xnor U7853 (N_7853,N_5230,N_6726);
or U7854 (N_7854,N_7010,N_7198);
and U7855 (N_7855,N_5312,N_7444);
xnor U7856 (N_7856,N_6355,N_6249);
or U7857 (N_7857,N_5589,N_6000);
and U7858 (N_7858,N_5273,N_5940);
and U7859 (N_7859,N_6147,N_6570);
and U7860 (N_7860,N_6711,N_5730);
or U7861 (N_7861,N_6981,N_5247);
xor U7862 (N_7862,N_7427,N_5319);
nand U7863 (N_7863,N_5036,N_6118);
or U7864 (N_7864,N_7346,N_5482);
nor U7865 (N_7865,N_5126,N_7496);
and U7866 (N_7866,N_6575,N_6950);
nand U7867 (N_7867,N_6733,N_5006);
nand U7868 (N_7868,N_6168,N_5498);
and U7869 (N_7869,N_6500,N_5777);
or U7870 (N_7870,N_6932,N_5387);
xor U7871 (N_7871,N_6280,N_6373);
nor U7872 (N_7872,N_5478,N_6158);
nand U7873 (N_7873,N_7134,N_7454);
and U7874 (N_7874,N_6621,N_6535);
nand U7875 (N_7875,N_5935,N_6239);
or U7876 (N_7876,N_5556,N_6421);
or U7877 (N_7877,N_6702,N_6278);
nor U7878 (N_7878,N_5961,N_5226);
xnor U7879 (N_7879,N_5396,N_5910);
and U7880 (N_7880,N_6923,N_6516);
and U7881 (N_7881,N_5753,N_5617);
and U7882 (N_7882,N_6438,N_6545);
xnor U7883 (N_7883,N_5154,N_5791);
nor U7884 (N_7884,N_5947,N_5383);
and U7885 (N_7885,N_6795,N_7026);
xor U7886 (N_7886,N_5241,N_6049);
nor U7887 (N_7887,N_6761,N_5835);
nor U7888 (N_7888,N_5921,N_5005);
nor U7889 (N_7889,N_5212,N_7369);
nand U7890 (N_7890,N_5309,N_6255);
xnor U7891 (N_7891,N_6543,N_5680);
nand U7892 (N_7892,N_7250,N_6917);
or U7893 (N_7893,N_5790,N_5796);
xnor U7894 (N_7894,N_6378,N_6004);
or U7895 (N_7895,N_6745,N_5417);
or U7896 (N_7896,N_5359,N_5335);
and U7897 (N_7897,N_6494,N_6918);
xnor U7898 (N_7898,N_5729,N_5923);
and U7899 (N_7899,N_5217,N_6006);
nand U7900 (N_7900,N_5090,N_5687);
nand U7901 (N_7901,N_5962,N_5944);
nand U7902 (N_7902,N_6939,N_6898);
and U7903 (N_7903,N_5138,N_6018);
and U7904 (N_7904,N_7360,N_7037);
nor U7905 (N_7905,N_5699,N_5180);
xnor U7906 (N_7906,N_6778,N_5606);
nand U7907 (N_7907,N_7494,N_7351);
and U7908 (N_7908,N_7022,N_6825);
nor U7909 (N_7909,N_6888,N_5222);
or U7910 (N_7910,N_6864,N_7469);
nor U7911 (N_7911,N_5453,N_5432);
nand U7912 (N_7912,N_5744,N_5852);
xor U7913 (N_7913,N_7426,N_6433);
xor U7914 (N_7914,N_7294,N_7161);
and U7915 (N_7915,N_6739,N_6834);
nor U7916 (N_7916,N_5455,N_7203);
nand U7917 (N_7917,N_6393,N_6491);
nand U7918 (N_7918,N_7288,N_6371);
or U7919 (N_7919,N_5275,N_5629);
xor U7920 (N_7920,N_5691,N_7229);
nor U7921 (N_7921,N_5018,N_5069);
nor U7922 (N_7922,N_6773,N_5906);
and U7923 (N_7923,N_5547,N_6541);
nand U7924 (N_7924,N_7274,N_6056);
nor U7925 (N_7925,N_5300,N_7001);
xor U7926 (N_7926,N_6497,N_5434);
xnor U7927 (N_7927,N_5004,N_7319);
nand U7928 (N_7928,N_7254,N_6183);
xnor U7929 (N_7929,N_6010,N_5618);
and U7930 (N_7930,N_5172,N_7061);
nand U7931 (N_7931,N_6803,N_6493);
and U7932 (N_7932,N_6188,N_6369);
nand U7933 (N_7933,N_5968,N_5484);
and U7934 (N_7934,N_5243,N_5291);
and U7935 (N_7935,N_6231,N_5623);
xor U7936 (N_7936,N_6597,N_6376);
nand U7937 (N_7937,N_7460,N_6250);
xnor U7938 (N_7938,N_5062,N_6818);
nand U7939 (N_7939,N_5189,N_6492);
or U7940 (N_7940,N_6708,N_5761);
xnor U7941 (N_7941,N_6634,N_5945);
xor U7942 (N_7942,N_6968,N_6831);
or U7943 (N_7943,N_5165,N_6097);
or U7944 (N_7944,N_5675,N_7073);
xnor U7945 (N_7945,N_5898,N_7291);
and U7946 (N_7946,N_6942,N_6301);
nand U7947 (N_7947,N_6534,N_6284);
nand U7948 (N_7948,N_5133,N_6382);
nand U7949 (N_7949,N_7019,N_5651);
xor U7950 (N_7950,N_5739,N_6977);
nor U7951 (N_7951,N_6738,N_5566);
nor U7952 (N_7952,N_5668,N_7098);
xnor U7953 (N_7953,N_7345,N_5003);
xnor U7954 (N_7954,N_6201,N_6519);
nand U7955 (N_7955,N_7035,N_5841);
or U7956 (N_7956,N_7070,N_6271);
or U7957 (N_7957,N_7476,N_5253);
xnor U7958 (N_7958,N_6039,N_7085);
or U7959 (N_7959,N_7451,N_5662);
nor U7960 (N_7960,N_7498,N_6285);
or U7961 (N_7961,N_5495,N_6793);
or U7962 (N_7962,N_5584,N_7064);
or U7963 (N_7963,N_5362,N_7405);
xnor U7964 (N_7964,N_5757,N_5678);
nor U7965 (N_7965,N_6647,N_7278);
or U7966 (N_7966,N_7030,N_5998);
and U7967 (N_7967,N_6817,N_5518);
xor U7968 (N_7968,N_5449,N_6316);
and U7969 (N_7969,N_6384,N_6643);
xnor U7970 (N_7970,N_5225,N_5999);
nor U7971 (N_7971,N_5535,N_5868);
or U7972 (N_7972,N_5077,N_6565);
or U7973 (N_7973,N_5988,N_7433);
nand U7974 (N_7974,N_6177,N_5803);
nor U7975 (N_7975,N_6194,N_7391);
nand U7976 (N_7976,N_6061,N_6811);
nand U7977 (N_7977,N_5805,N_6509);
or U7978 (N_7978,N_6996,N_6479);
nand U7979 (N_7979,N_5162,N_7304);
xnor U7980 (N_7980,N_5622,N_6728);
and U7981 (N_7981,N_7367,N_5671);
or U7982 (N_7982,N_6990,N_6557);
or U7983 (N_7983,N_5747,N_7045);
nand U7984 (N_7984,N_6143,N_6986);
and U7985 (N_7985,N_5941,N_5250);
xnor U7986 (N_7986,N_7321,N_6764);
xnor U7987 (N_7987,N_7239,N_6873);
and U7988 (N_7988,N_6311,N_7357);
nand U7989 (N_7989,N_5932,N_5598);
xnor U7990 (N_7990,N_6959,N_6001);
and U7991 (N_7991,N_5211,N_6341);
xor U7992 (N_7992,N_6703,N_7331);
and U7993 (N_7993,N_6729,N_6386);
nor U7994 (N_7994,N_6751,N_7100);
xor U7995 (N_7995,N_6518,N_7300);
or U7996 (N_7996,N_6907,N_7264);
nand U7997 (N_7997,N_6206,N_6305);
xor U7998 (N_7998,N_6298,N_6134);
nand U7999 (N_7999,N_6652,N_6521);
nand U8000 (N_8000,N_5176,N_6780);
nand U8001 (N_8001,N_6625,N_5297);
and U8002 (N_8002,N_5282,N_7155);
nand U8003 (N_8003,N_5604,N_5745);
and U8004 (N_8004,N_5976,N_7039);
xor U8005 (N_8005,N_6105,N_6600);
nor U8006 (N_8006,N_5652,N_5700);
and U8007 (N_8007,N_5644,N_6448);
xnor U8008 (N_8008,N_6477,N_6840);
nand U8009 (N_8009,N_7490,N_7083);
and U8010 (N_8010,N_5608,N_5801);
xor U8011 (N_8011,N_6264,N_5781);
xnor U8012 (N_8012,N_6449,N_7396);
or U8013 (N_8013,N_7113,N_6208);
nor U8014 (N_8014,N_5480,N_5158);
nor U8015 (N_8015,N_6326,N_6672);
xor U8016 (N_8016,N_6122,N_7361);
nor U8017 (N_8017,N_7293,N_6904);
nand U8018 (N_8018,N_5078,N_6011);
xnor U8019 (N_8019,N_5065,N_7318);
nand U8020 (N_8020,N_6614,N_6645);
nand U8021 (N_8021,N_5301,N_6294);
nand U8022 (N_8022,N_6976,N_6330);
nand U8023 (N_8023,N_7408,N_5184);
xor U8024 (N_8024,N_5862,N_7313);
nor U8025 (N_8025,N_5737,N_7385);
nand U8026 (N_8026,N_5048,N_6259);
and U8027 (N_8027,N_5044,N_6940);
and U8028 (N_8028,N_6660,N_5021);
nand U8029 (N_8029,N_6234,N_6046);
nand U8030 (N_8030,N_6511,N_7124);
xnor U8031 (N_8031,N_6956,N_7389);
or U8032 (N_8032,N_7188,N_6483);
and U8033 (N_8033,N_6591,N_6995);
and U8034 (N_8034,N_6257,N_5129);
nor U8035 (N_8035,N_7114,N_7175);
xor U8036 (N_8036,N_7478,N_7186);
or U8037 (N_8037,N_5020,N_6027);
and U8038 (N_8038,N_5029,N_6446);
nand U8039 (N_8039,N_6743,N_5646);
xor U8040 (N_8040,N_6828,N_5267);
and U8041 (N_8041,N_5993,N_5592);
xor U8042 (N_8042,N_6725,N_5588);
nand U8043 (N_8043,N_6559,N_5391);
and U8044 (N_8044,N_5702,N_7149);
and U8045 (N_8045,N_5692,N_5292);
or U8046 (N_8046,N_7365,N_5467);
xor U8047 (N_8047,N_6719,N_7003);
and U8048 (N_8048,N_6410,N_5511);
nand U8049 (N_8049,N_6499,N_5718);
or U8050 (N_8050,N_7204,N_5546);
xor U8051 (N_8051,N_6400,N_5308);
and U8052 (N_8052,N_6532,N_6181);
nand U8053 (N_8053,N_6128,N_5414);
xor U8054 (N_8054,N_5277,N_7271);
xnor U8055 (N_8055,N_5279,N_7009);
or U8056 (N_8056,N_5024,N_7450);
or U8057 (N_8057,N_6091,N_7116);
and U8058 (N_8058,N_6347,N_5514);
or U8059 (N_8059,N_5502,N_5264);
or U8060 (N_8060,N_6732,N_7348);
and U8061 (N_8061,N_5354,N_6406);
nand U8062 (N_8062,N_6013,N_5000);
and U8063 (N_8063,N_5695,N_7218);
nor U8064 (N_8064,N_7437,N_6100);
and U8065 (N_8065,N_5393,N_5661);
or U8066 (N_8066,N_5194,N_7353);
xor U8067 (N_8067,N_5710,N_5303);
nor U8068 (N_8068,N_6965,N_5794);
nand U8069 (N_8069,N_5454,N_5068);
or U8070 (N_8070,N_7325,N_6915);
xnor U8071 (N_8071,N_7486,N_5328);
and U8072 (N_8072,N_6069,N_6526);
nor U8073 (N_8073,N_7153,N_5294);
nand U8074 (N_8074,N_7147,N_5060);
and U8075 (N_8075,N_6787,N_6360);
xor U8076 (N_8076,N_6870,N_5797);
xnor U8077 (N_8077,N_5223,N_6874);
or U8078 (N_8078,N_6852,N_6473);
nor U8079 (N_8079,N_7257,N_7163);
or U8080 (N_8080,N_6401,N_6157);
nand U8081 (N_8081,N_7347,N_6759);
nor U8082 (N_8082,N_6663,N_6882);
nand U8083 (N_8083,N_5155,N_7123);
nor U8084 (N_8084,N_6429,N_7115);
and U8085 (N_8085,N_6275,N_6149);
or U8086 (N_8086,N_6936,N_6848);
xor U8087 (N_8087,N_5252,N_5428);
or U8088 (N_8088,N_7146,N_5716);
nand U8089 (N_8089,N_5070,N_5768);
nand U8090 (N_8090,N_5128,N_7395);
and U8091 (N_8091,N_7276,N_5839);
or U8092 (N_8092,N_5600,N_6020);
nor U8093 (N_8093,N_6832,N_6824);
or U8094 (N_8094,N_5742,N_6423);
and U8095 (N_8095,N_6015,N_6763);
nor U8096 (N_8096,N_5915,N_5299);
nor U8097 (N_8097,N_5476,N_5079);
nor U8098 (N_8098,N_6332,N_7238);
or U8099 (N_8099,N_6674,N_5027);
nor U8100 (N_8100,N_5510,N_7403);
xnor U8101 (N_8101,N_5259,N_6974);
xnor U8102 (N_8102,N_6116,N_5925);
nand U8103 (N_8103,N_5343,N_5865);
nor U8104 (N_8104,N_6718,N_6033);
and U8105 (N_8105,N_5148,N_5663);
nor U8106 (N_8106,N_7381,N_6198);
nand U8107 (N_8107,N_6830,N_5266);
nand U8108 (N_8108,N_5750,N_5679);
xnor U8109 (N_8109,N_7102,N_7221);
nor U8110 (N_8110,N_6688,N_7260);
and U8111 (N_8111,N_7463,N_6082);
or U8112 (N_8112,N_6552,N_7249);
xnor U8113 (N_8113,N_6658,N_7272);
or U8114 (N_8114,N_5047,N_5851);
nor U8115 (N_8115,N_6002,N_6712);
xor U8116 (N_8116,N_6469,N_6821);
or U8117 (N_8117,N_5114,N_6754);
and U8118 (N_8118,N_5758,N_5395);
xnor U8119 (N_8119,N_7322,N_5603);
xor U8120 (N_8120,N_7170,N_6544);
nand U8121 (N_8121,N_5286,N_5012);
nor U8122 (N_8122,N_5288,N_7214);
or U8123 (N_8123,N_7029,N_5567);
nand U8124 (N_8124,N_5053,N_7400);
or U8125 (N_8125,N_5544,N_7067);
nor U8126 (N_8126,N_6651,N_6687);
and U8127 (N_8127,N_5055,N_6949);
or U8128 (N_8128,N_5143,N_6394);
and U8129 (N_8129,N_6098,N_7309);
or U8130 (N_8130,N_7461,N_5648);
or U8131 (N_8131,N_6262,N_6618);
nor U8132 (N_8132,N_7449,N_7240);
or U8133 (N_8133,N_6388,N_5703);
xnor U8134 (N_8134,N_6290,N_7047);
nor U8135 (N_8135,N_5725,N_6583);
or U8136 (N_8136,N_7477,N_7474);
nand U8137 (N_8137,N_5320,N_5293);
xor U8138 (N_8138,N_6779,N_5106);
nand U8139 (N_8139,N_5409,N_5281);
nor U8140 (N_8140,N_5949,N_7192);
and U8141 (N_8141,N_7235,N_7040);
nand U8142 (N_8142,N_6680,N_5785);
nand U8143 (N_8143,N_7412,N_5221);
or U8144 (N_8144,N_6121,N_5167);
nor U8145 (N_8145,N_5704,N_6850);
xor U8146 (N_8146,N_7489,N_6962);
xnor U8147 (N_8147,N_5063,N_6064);
and U8148 (N_8148,N_7421,N_5736);
xnor U8149 (N_8149,N_6331,N_5942);
xor U8150 (N_8150,N_7016,N_5806);
or U8151 (N_8151,N_6734,N_7406);
and U8152 (N_8152,N_6502,N_6125);
xor U8153 (N_8153,N_7078,N_5124);
and U8154 (N_8154,N_5879,N_5278);
nor U8155 (N_8155,N_5326,N_5316);
nand U8156 (N_8156,N_7452,N_6042);
nand U8157 (N_8157,N_6771,N_7119);
xnor U8158 (N_8158,N_6038,N_6434);
nand U8159 (N_8159,N_5386,N_5755);
nor U8160 (N_8160,N_5698,N_5553);
or U8161 (N_8161,N_7158,N_5492);
or U8162 (N_8162,N_7056,N_7259);
xnor U8163 (N_8163,N_5965,N_5531);
nor U8164 (N_8164,N_6150,N_6031);
nand U8165 (N_8165,N_6851,N_7181);
xor U8166 (N_8166,N_5204,N_6300);
nand U8167 (N_8167,N_6857,N_7173);
nor U8168 (N_8168,N_6798,N_6999);
nor U8169 (N_8169,N_5011,N_5110);
nor U8170 (N_8170,N_7005,N_5505);
nand U8171 (N_8171,N_5578,N_6173);
or U8172 (N_8172,N_6642,N_5550);
xor U8173 (N_8173,N_6207,N_5863);
nand U8174 (N_8174,N_5779,N_6144);
nand U8175 (N_8175,N_6127,N_6408);
and U8176 (N_8176,N_7326,N_6073);
nor U8177 (N_8177,N_5838,N_6137);
or U8178 (N_8178,N_5762,N_5613);
and U8179 (N_8179,N_5367,N_7057);
or U8180 (N_8180,N_6957,N_7242);
xor U8181 (N_8181,N_5660,N_6040);
nand U8182 (N_8182,N_5986,N_6024);
and U8183 (N_8183,N_5888,N_6129);
nor U8184 (N_8184,N_6180,N_6650);
xor U8185 (N_8185,N_6108,N_6596);
and U8186 (N_8186,N_6659,N_6520);
and U8187 (N_8187,N_6154,N_6767);
nand U8188 (N_8188,N_5161,N_5033);
and U8189 (N_8189,N_5782,N_6133);
xnor U8190 (N_8190,N_5152,N_5360);
xor U8191 (N_8191,N_5593,N_7105);
xnor U8192 (N_8192,N_5200,N_5237);
nor U8193 (N_8193,N_6717,N_5990);
or U8194 (N_8194,N_5997,N_6524);
nor U8195 (N_8195,N_5832,N_6963);
nand U8196 (N_8196,N_6162,N_6542);
xnor U8197 (N_8197,N_6050,N_6875);
and U8198 (N_8198,N_5139,N_7000);
and U8199 (N_8199,N_7222,N_7034);
nor U8200 (N_8200,N_6801,N_5664);
and U8201 (N_8201,N_6517,N_5082);
nor U8202 (N_8202,N_7006,N_7164);
and U8203 (N_8203,N_7292,N_7410);
and U8204 (N_8204,N_6451,N_6638);
nand U8205 (N_8205,N_5254,N_6954);
nor U8206 (N_8206,N_5576,N_7330);
and U8207 (N_8207,N_5734,N_5216);
nand U8208 (N_8208,N_6553,N_5724);
nand U8209 (N_8209,N_6315,N_6598);
xor U8210 (N_8210,N_6772,N_5770);
nor U8211 (N_8211,N_7342,N_7265);
nand U8212 (N_8212,N_5325,N_6792);
nor U8213 (N_8213,N_5464,N_6946);
xor U8214 (N_8214,N_5614,N_5410);
and U8215 (N_8215,N_5813,N_7143);
or U8216 (N_8216,N_5793,N_5625);
nand U8217 (N_8217,N_7328,N_6829);
nor U8218 (N_8218,N_6902,N_5871);
nand U8219 (N_8219,N_5713,N_6402);
or U8220 (N_8220,N_6814,N_6431);
nand U8221 (N_8221,N_5493,N_6588);
or U8222 (N_8222,N_6043,N_5802);
or U8223 (N_8223,N_6426,N_5701);
xnor U8224 (N_8224,N_6222,N_6813);
or U8225 (N_8225,N_5844,N_5450);
nor U8226 (N_8226,N_5552,N_7447);
xor U8227 (N_8227,N_5242,N_5992);
xnor U8228 (N_8228,N_7227,N_6470);
nand U8229 (N_8229,N_7305,N_5234);
or U8230 (N_8230,N_7036,N_7492);
xor U8231 (N_8231,N_7388,N_6119);
or U8232 (N_8232,N_7213,N_7054);
and U8233 (N_8233,N_5429,N_5122);
nor U8234 (N_8234,N_7236,N_6581);
and U8235 (N_8235,N_7135,N_6079);
nor U8236 (N_8236,N_5488,N_7362);
xor U8237 (N_8237,N_6344,N_6556);
nand U8238 (N_8238,N_5456,N_5817);
and U8239 (N_8239,N_6197,N_6204);
and U8240 (N_8240,N_5422,N_7364);
or U8241 (N_8241,N_5379,N_5290);
xor U8242 (N_8242,N_5125,N_6480);
nor U8243 (N_8243,N_7044,N_5169);
xnor U8244 (N_8244,N_5717,N_5153);
nand U8245 (N_8245,N_6958,N_6605);
xnor U8246 (N_8246,N_7333,N_6566);
nand U8247 (N_8247,N_6537,N_6694);
xnor U8248 (N_8248,N_6456,N_7445);
nor U8249 (N_8249,N_6357,N_6335);
nand U8250 (N_8250,N_6409,N_6395);
nand U8251 (N_8251,N_6756,N_6299);
xor U8252 (N_8252,N_6286,N_6114);
and U8253 (N_8253,N_5683,N_7225);
nor U8254 (N_8254,N_6427,N_6927);
or U8255 (N_8255,N_6496,N_6367);
or U8256 (N_8256,N_5262,N_5056);
nor U8257 (N_8257,N_6327,N_6964);
nor U8258 (N_8258,N_6744,N_7409);
nor U8259 (N_8259,N_7290,N_5411);
nor U8260 (N_8260,N_5405,N_6685);
nand U8261 (N_8261,N_6796,N_5307);
nand U8262 (N_8262,N_6997,N_6691);
xor U8263 (N_8263,N_6920,N_6314);
nor U8264 (N_8264,N_6176,N_6705);
xnor U8265 (N_8265,N_6103,N_5013);
nand U8266 (N_8266,N_5843,N_7439);
nand U8267 (N_8267,N_7109,N_7338);
or U8268 (N_8268,N_5969,N_6251);
and U8269 (N_8269,N_6606,N_6172);
and U8270 (N_8270,N_5682,N_6095);
nor U8271 (N_8271,N_6228,N_7171);
xor U8272 (N_8272,N_6224,N_7306);
nand U8273 (N_8273,N_5653,N_6602);
nor U8274 (N_8274,N_6709,N_7157);
and U8275 (N_8275,N_5869,N_5527);
nand U8276 (N_8276,N_6430,N_7199);
or U8277 (N_8277,N_6458,N_6673);
and U8278 (N_8278,N_6317,N_5943);
nand U8279 (N_8279,N_5321,N_7020);
or U8280 (N_8280,N_5798,N_6288);
nand U8281 (N_8281,N_5621,N_5472);
and U8282 (N_8282,N_7275,N_7261);
xnor U8283 (N_8283,N_5399,N_6668);
nor U8284 (N_8284,N_5586,N_5283);
or U8285 (N_8285,N_5981,N_6684);
nor U8286 (N_8286,N_5727,N_7267);
or U8287 (N_8287,N_6594,N_5763);
nor U8288 (N_8288,N_5526,N_6901);
and U8289 (N_8289,N_7210,N_6682);
nand U8290 (N_8290,N_7024,N_7032);
nor U8291 (N_8291,N_5496,N_5448);
nand U8292 (N_8292,N_6802,N_5007);
and U8293 (N_8293,N_6633,N_6037);
and U8294 (N_8294,N_6191,N_6363);
xnor U8295 (N_8295,N_7303,N_5348);
or U8296 (N_8296,N_6945,N_6742);
nor U8297 (N_8297,N_5305,N_5585);
nor U8298 (N_8298,N_6572,N_5076);
and U8299 (N_8299,N_7413,N_6383);
and U8300 (N_8300,N_5402,N_7117);
nor U8301 (N_8301,N_6653,N_6247);
or U8302 (N_8302,N_5489,N_5441);
nor U8303 (N_8303,N_7106,N_6059);
xnor U8304 (N_8304,N_6522,N_5355);
nand U8305 (N_8305,N_5991,N_5807);
nor U8306 (N_8306,N_6417,N_5109);
or U8307 (N_8307,N_7144,N_5596);
nor U8308 (N_8308,N_5712,N_7200);
and U8309 (N_8309,N_6392,N_6854);
nor U8310 (N_8310,N_5052,N_6689);
nand U8311 (N_8311,N_6845,N_6937);
or U8312 (N_8312,N_6136,N_6587);
nand U8313 (N_8313,N_6457,N_7475);
or U8314 (N_8314,N_6577,N_6233);
nor U8315 (N_8315,N_5342,N_6822);
and U8316 (N_8316,N_5088,N_5043);
or U8317 (N_8317,N_5665,N_6164);
nand U8318 (N_8318,N_7212,N_6182);
xor U8319 (N_8319,N_5347,N_5332);
or U8320 (N_8320,N_7216,N_5628);
or U8321 (N_8321,N_7015,N_7256);
nand U8322 (N_8322,N_6321,N_6485);
nor U8323 (N_8323,N_5119,N_7434);
xnor U8324 (N_8324,N_7138,N_7334);
nor U8325 (N_8325,N_5808,N_7172);
and U8326 (N_8326,N_6248,N_5828);
nor U8327 (N_8327,N_7497,N_5327);
or U8328 (N_8328,N_5605,N_6998);
xnor U8329 (N_8329,N_5210,N_6993);
xor U8330 (N_8330,N_7310,N_6590);
nor U8331 (N_8331,N_5508,N_6032);
and U8332 (N_8332,N_7027,N_5509);
nor U8333 (N_8333,N_5042,N_5192);
nor U8334 (N_8334,N_5975,N_5792);
and U8335 (N_8335,N_5948,N_7446);
nor U8336 (N_8336,N_5522,N_5394);
or U8337 (N_8337,N_6671,N_6800);
nor U8338 (N_8338,N_7375,N_6132);
xnor U8339 (N_8339,N_6758,N_5672);
xnor U8340 (N_8340,N_6334,N_7131);
and U8341 (N_8341,N_5461,N_5714);
nand U8342 (N_8342,N_7112,N_5401);
nand U8343 (N_8343,N_6931,N_6896);
or U8344 (N_8344,N_6935,N_7011);
nand U8345 (N_8345,N_6110,N_6484);
nor U8346 (N_8346,N_5289,N_6047);
xor U8347 (N_8347,N_6277,N_6017);
nand U8348 (N_8348,N_6601,N_5431);
nor U8349 (N_8349,N_5213,N_7195);
nor U8350 (N_8350,N_7299,N_7051);
or U8351 (N_8351,N_7234,N_5046);
and U8352 (N_8352,N_5571,N_6089);
or U8353 (N_8353,N_5356,N_6860);
and U8354 (N_8354,N_7069,N_5919);
nor U8355 (N_8355,N_5284,N_5306);
nor U8356 (N_8356,N_5397,N_5157);
xor U8357 (N_8357,N_7176,N_6381);
and U8358 (N_8358,N_6858,N_5438);
xor U8359 (N_8359,N_6398,N_5842);
nor U8360 (N_8360,N_5911,N_7142);
and U8361 (N_8361,N_6613,N_7232);
nand U8362 (N_8362,N_6461,N_5856);
nand U8363 (N_8363,N_6952,N_5220);
and U8364 (N_8364,N_6219,N_7241);
nand U8365 (N_8365,N_5836,N_5658);
and U8366 (N_8366,N_7296,N_5272);
xnor U8367 (N_8367,N_7269,N_5913);
nor U8368 (N_8368,N_6138,N_5098);
or U8369 (N_8369,N_5731,N_5568);
nor U8370 (N_8370,N_5481,N_5363);
or U8371 (N_8371,N_5890,N_5451);
and U8372 (N_8372,N_5579,N_5089);
xnor U8373 (N_8373,N_5627,N_6066);
or U8374 (N_8374,N_7404,N_5179);
xnor U8375 (N_8375,N_6442,N_5390);
nand U8376 (N_8376,N_5458,N_6558);
xnor U8377 (N_8377,N_5437,N_5810);
nor U8378 (N_8378,N_6362,N_6697);
and U8379 (N_8379,N_6454,N_5900);
and U8380 (N_8380,N_5322,N_5693);
or U8381 (N_8381,N_7007,N_7282);
xor U8382 (N_8382,N_5877,N_7368);
or U8383 (N_8383,N_6737,N_6472);
xnor U8384 (N_8384,N_6571,N_7133);
nand U8385 (N_8385,N_5874,N_5350);
or U8386 (N_8386,N_5418,N_6053);
nand U8387 (N_8387,N_6991,N_6077);
xnor U8388 (N_8388,N_5115,N_5894);
xnor U8389 (N_8389,N_6184,N_6274);
or U8390 (N_8390,N_5674,N_6987);
nor U8391 (N_8391,N_7481,N_6909);
nand U8392 (N_8392,N_5173,N_6120);
and U8393 (N_8393,N_6009,N_5610);
and U8394 (N_8394,N_6842,N_6404);
and U8395 (N_8395,N_5271,N_6067);
nor U8396 (N_8396,N_5950,N_5896);
nor U8397 (N_8397,N_7329,N_7252);
nor U8398 (N_8398,N_6238,N_5903);
or U8399 (N_8399,N_5504,N_7289);
nand U8400 (N_8400,N_5009,N_6349);
or U8401 (N_8401,N_6425,N_7095);
nand U8402 (N_8402,N_6916,N_7358);
xor U8403 (N_8403,N_7340,N_5866);
nand U8404 (N_8404,N_6693,N_5640);
and U8405 (N_8405,N_5295,N_5365);
xnor U8406 (N_8406,N_6878,N_5533);
xor U8407 (N_8407,N_6955,N_6420);
and U8408 (N_8408,N_5233,N_6551);
xor U8409 (N_8409,N_6005,N_7308);
or U8410 (N_8410,N_6156,N_6877);
xor U8411 (N_8411,N_6890,N_6029);
nand U8412 (N_8412,N_5720,N_5811);
xor U8413 (N_8413,N_5748,N_6374);
xnor U8414 (N_8414,N_7129,N_5534);
nor U8415 (N_8415,N_5442,N_5551);
nor U8416 (N_8416,N_7237,N_5187);
xnor U8417 (N_8417,N_6547,N_6615);
nand U8418 (N_8418,N_7243,N_5561);
xor U8419 (N_8419,N_5030,N_5389);
nor U8420 (N_8420,N_6014,N_5116);
nand U8421 (N_8421,N_6794,N_6310);
nor U8422 (N_8422,N_7043,N_5619);
nor U8423 (N_8423,N_7355,N_7386);
xnor U8424 (N_8424,N_7077,N_6012);
nand U8425 (N_8425,N_6921,N_5967);
or U8426 (N_8426,N_5251,N_6240);
xor U8427 (N_8427,N_7399,N_6200);
nand U8428 (N_8428,N_6715,N_6568);
nor U8429 (N_8429,N_5274,N_6879);
nand U8430 (N_8430,N_6512,N_7438);
nor U8431 (N_8431,N_5199,N_6704);
xor U8432 (N_8432,N_6859,N_5183);
or U8433 (N_8433,N_6584,N_6626);
and U8434 (N_8434,N_6753,N_5064);
and U8435 (N_8435,N_5249,N_5101);
and U8436 (N_8436,N_7366,N_5452);
and U8437 (N_8437,N_6510,N_6007);
xnor U8438 (N_8438,N_5232,N_5746);
xnor U8439 (N_8439,N_6629,N_6359);
nand U8440 (N_8440,N_6639,N_7472);
nand U8441 (N_8441,N_6261,N_6101);
xnor U8442 (N_8442,N_6413,N_6245);
nor U8443 (N_8443,N_6667,N_6375);
nand U8444 (N_8444,N_5541,N_6515);
nor U8445 (N_8445,N_7189,N_5684);
and U8446 (N_8446,N_7092,N_5686);
nor U8447 (N_8447,N_5512,N_5190);
or U8448 (N_8448,N_7270,N_5825);
nand U8449 (N_8449,N_6969,N_5555);
or U8450 (N_8450,N_6489,N_5787);
nand U8451 (N_8451,N_6303,N_7317);
and U8452 (N_8452,N_6893,N_5882);
nor U8453 (N_8453,N_5164,N_6266);
and U8454 (N_8454,N_7101,N_7441);
and U8455 (N_8455,N_6342,N_5771);
nor U8456 (N_8456,N_6797,N_7046);
and U8457 (N_8457,N_5067,N_6617);
and U8458 (N_8458,N_7014,N_5137);
xor U8459 (N_8459,N_7096,N_6260);
or U8460 (N_8460,N_5329,N_5887);
xor U8461 (N_8461,N_5034,N_5891);
xor U8462 (N_8462,N_6844,N_7363);
and U8463 (N_8463,N_6022,N_5338);
nor U8464 (N_8464,N_5602,N_6287);
or U8465 (N_8465,N_5244,N_5280);
nor U8466 (N_8466,N_5517,N_5767);
nand U8467 (N_8467,N_7187,N_5743);
or U8468 (N_8468,N_6696,N_5733);
and U8469 (N_8469,N_5934,N_7268);
nand U8470 (N_8470,N_6630,N_7343);
xor U8471 (N_8471,N_5984,N_7287);
or U8472 (N_8472,N_6656,N_5339);
and U8473 (N_8473,N_5460,N_5058);
xor U8474 (N_8474,N_5650,N_7088);
nand U8475 (N_8475,N_5609,N_5820);
xor U8476 (N_8476,N_6838,N_6385);
xor U8477 (N_8477,N_6883,N_6654);
or U8478 (N_8478,N_5848,N_5400);
nor U8479 (N_8479,N_5311,N_5677);
nand U8480 (N_8480,N_5996,N_5528);
nand U8481 (N_8481,N_5655,N_5577);
nand U8482 (N_8482,N_6599,N_5639);
xnor U8483 (N_8483,N_6531,N_5240);
or U8484 (N_8484,N_5607,N_6218);
nor U8485 (N_8485,N_5246,N_5074);
nor U8486 (N_8486,N_5468,N_6085);
and U8487 (N_8487,N_5549,N_7499);
nor U8488 (N_8488,N_6324,N_6269);
nor U8489 (N_8489,N_7110,N_7136);
xnor U8490 (N_8490,N_6776,N_6908);
nand U8491 (N_8491,N_6352,N_6003);
nand U8492 (N_8492,N_7422,N_5723);
nor U8493 (N_8493,N_6762,N_6444);
nor U8494 (N_8494,N_6075,N_6695);
or U8495 (N_8495,N_5595,N_5341);
or U8496 (N_8496,N_5989,N_7466);
or U8497 (N_8497,N_7286,N_6846);
xor U8498 (N_8498,N_7206,N_6354);
nand U8499 (N_8499,N_7130,N_5263);
nor U8500 (N_8500,N_6407,N_6507);
nand U8501 (N_8501,N_7125,N_6632);
or U8502 (N_8502,N_6338,N_5831);
xnor U8503 (N_8503,N_7371,N_6216);
or U8504 (N_8504,N_6236,N_5564);
nor U8505 (N_8505,N_5815,N_6785);
nor U8506 (N_8506,N_6984,N_6631);
xor U8507 (N_8507,N_6683,N_6415);
nand U8508 (N_8508,N_6983,N_5548);
or U8509 (N_8509,N_5926,N_6462);
nand U8510 (N_8510,N_5471,N_6768);
or U8511 (N_8511,N_6112,N_5860);
or U8512 (N_8512,N_6459,N_7487);
nand U8513 (N_8513,N_7062,N_6225);
nand U8514 (N_8514,N_6540,N_6370);
and U8515 (N_8515,N_5971,N_6922);
xnor U8516 (N_8516,N_6270,N_6296);
or U8517 (N_8517,N_6826,N_6450);
xor U8518 (N_8518,N_6092,N_7018);
nand U8519 (N_8519,N_7126,N_6443);
nor U8520 (N_8520,N_6641,N_6187);
or U8521 (N_8521,N_6179,N_6302);
xor U8522 (N_8522,N_7041,N_5912);
and U8523 (N_8523,N_6933,N_5858);
and U8524 (N_8524,N_7462,N_5479);
nand U8525 (N_8525,N_5051,N_6856);
nor U8526 (N_8526,N_6501,N_6919);
nor U8527 (N_8527,N_5111,N_7160);
or U8528 (N_8528,N_5425,N_6322);
nor U8529 (N_8529,N_6464,N_5142);
nand U8530 (N_8530,N_5473,N_7033);
and U8531 (N_8531,N_6514,N_7107);
and U8532 (N_8532,N_5371,N_6281);
xnor U8533 (N_8533,N_5669,N_6690);
and U8534 (N_8534,N_5732,N_5543);
xor U8535 (N_8535,N_5475,N_5824);
and U8536 (N_8536,N_5885,N_5444);
xnor U8537 (N_8537,N_6789,N_5108);
nor U8538 (N_8538,N_6841,N_5256);
and U8539 (N_8539,N_7356,N_5238);
xor U8540 (N_8540,N_6843,N_5914);
or U8541 (N_8541,N_6486,N_6380);
and U8542 (N_8542,N_5261,N_6196);
xor U8543 (N_8543,N_6016,N_5878);
or U8544 (N_8544,N_6665,N_6836);
and U8545 (N_8545,N_5443,N_5875);
nand U8546 (N_8546,N_6148,N_6226);
or U8547 (N_8547,N_5499,N_5178);
nor U8548 (N_8548,N_7178,N_5635);
nand U8549 (N_8549,N_6366,N_6435);
nand U8550 (N_8550,N_5215,N_6884);
nor U8551 (N_8551,N_5298,N_6971);
nor U8552 (N_8552,N_6465,N_5416);
and U8553 (N_8553,N_7066,N_6282);
or U8554 (N_8554,N_6252,N_5231);
nand U8555 (N_8555,N_7370,N_6664);
or U8556 (N_8556,N_6911,N_6628);
and U8557 (N_8557,N_7076,N_7194);
xor U8558 (N_8558,N_5236,N_5463);
or U8559 (N_8559,N_6701,N_6781);
nor U8560 (N_8560,N_7277,N_6351);
or U8561 (N_8561,N_7048,N_5087);
xor U8562 (N_8562,N_6256,N_6320);
or U8563 (N_8563,N_5809,N_5916);
nor U8564 (N_8564,N_7390,N_5880);
nor U8565 (N_8565,N_7205,N_5893);
or U8566 (N_8566,N_5117,N_5181);
and U8567 (N_8567,N_6692,N_6972);
nor U8568 (N_8568,N_7159,N_7465);
or U8569 (N_8569,N_6195,N_6853);
nand U8570 (N_8570,N_5260,N_5867);
nand U8571 (N_8571,N_6943,N_6833);
nor U8572 (N_8572,N_5358,N_6111);
nor U8573 (N_8573,N_7480,N_6847);
and U8574 (N_8574,N_6774,N_5219);
xnor U8575 (N_8575,N_6675,N_6244);
nor U8576 (N_8576,N_7104,N_5398);
or U8577 (N_8577,N_6163,N_6786);
and U8578 (N_8578,N_5630,N_6610);
or U8579 (N_8579,N_5203,N_6593);
nor U8580 (N_8580,N_5889,N_5268);
nor U8581 (N_8581,N_5019,N_6677);
xnor U8582 (N_8582,N_6199,N_5633);
nor U8583 (N_8583,N_5539,N_5378);
and U8584 (N_8584,N_6368,N_6084);
and U8585 (N_8585,N_6186,N_5537);
nor U8586 (N_8586,N_6076,N_6809);
and U8587 (N_8587,N_5214,N_6152);
or U8588 (N_8588,N_6416,N_5581);
nor U8589 (N_8589,N_6447,N_6397);
and U8590 (N_8590,N_5403,N_5780);
nor U8591 (N_8591,N_6441,N_5039);
and U8592 (N_8592,N_7320,N_6748);
nand U8593 (N_8593,N_5392,N_6072);
and U8594 (N_8594,N_5957,N_7174);
nand U8595 (N_8595,N_6212,N_5208);
nor U8596 (N_8596,N_5457,N_6666);
and U8597 (N_8597,N_6232,N_5136);
xor U8598 (N_8598,N_7253,N_6358);
and U8599 (N_8599,N_6223,N_5415);
nor U8600 (N_8600,N_5151,N_6364);
nor U8601 (N_8601,N_6021,N_5827);
or U8602 (N_8602,N_7473,N_6166);
or U8603 (N_8603,N_6295,N_7169);
and U8604 (N_8604,N_6498,N_7220);
and U8605 (N_8605,N_7378,N_7384);
nor U8606 (N_8606,N_5296,N_6323);
or U8607 (N_8607,N_5132,N_7297);
nor U8608 (N_8608,N_5532,N_5196);
or U8609 (N_8609,N_6140,N_6894);
or U8610 (N_8610,N_5775,N_6627);
xnor U8611 (N_8611,N_7245,N_5218);
or U8612 (N_8612,N_6304,N_5756);
nor U8613 (N_8613,N_6947,N_5688);
xor U8614 (N_8614,N_7251,N_5929);
nand U8615 (N_8615,N_5845,N_5166);
or U8616 (N_8616,N_5257,N_7065);
nor U8617 (N_8617,N_5570,N_7209);
and U8618 (N_8618,N_5973,N_6585);
xor U8619 (N_8619,N_6145,N_5773);
xor U8620 (N_8620,N_5854,N_5072);
nand U8621 (N_8621,N_5366,N_5315);
nor U8622 (N_8622,N_5227,N_7415);
and U8623 (N_8623,N_7467,N_6710);
or U8624 (N_8624,N_7166,N_7151);
and U8625 (N_8625,N_7455,N_7458);
nor U8626 (N_8626,N_6777,N_5558);
nand U8627 (N_8627,N_6329,N_5690);
xor U8628 (N_8628,N_7373,N_5149);
xnor U8629 (N_8629,N_5049,N_5265);
and U8630 (N_8630,N_5726,N_6574);
nand U8631 (N_8631,N_7468,N_7372);
xor U8632 (N_8632,N_5057,N_7167);
xor U8633 (N_8633,N_5562,N_5760);
xor U8634 (N_8634,N_5521,N_6161);
xnor U8635 (N_8635,N_6513,N_5500);
or U8636 (N_8636,N_6190,N_7491);
xor U8637 (N_8637,N_6142,N_5638);
and U8638 (N_8638,N_5487,N_5445);
or U8639 (N_8639,N_5494,N_6192);
nor U8640 (N_8640,N_6849,N_5740);
xnor U8641 (N_8641,N_5470,N_5920);
or U8642 (N_8642,N_6941,N_6755);
and U8643 (N_8643,N_5516,N_6267);
or U8644 (N_8644,N_7090,N_5917);
nand U8645 (N_8645,N_5188,N_5752);
nor U8646 (N_8646,N_6487,N_5857);
and U8647 (N_8647,N_6265,N_6592);
xor U8648 (N_8648,N_7012,N_5384);
xor U8649 (N_8649,N_5413,N_7079);
nor U8650 (N_8650,N_6070,N_6560);
nor U8651 (N_8651,N_5404,N_6220);
and U8652 (N_8652,N_6345,N_5182);
nor U8653 (N_8653,N_7074,N_5719);
xnor U8654 (N_8654,N_6063,N_5304);
nor U8655 (N_8655,N_7139,N_6530);
and U8656 (N_8656,N_7247,N_6308);
nand U8657 (N_8657,N_7279,N_6068);
xnor U8658 (N_8658,N_7457,N_5616);
nor U8659 (N_8659,N_6418,N_5198);
nand U8660 (N_8660,N_6573,N_5545);
nor U8661 (N_8661,N_6865,N_5424);
nand U8662 (N_8662,N_6170,N_6567);
and U8663 (N_8663,N_6928,N_5594);
nand U8664 (N_8664,N_7004,N_6104);
and U8665 (N_8665,N_7442,N_7053);
xnor U8666 (N_8666,N_5229,N_5205);
or U8667 (N_8667,N_6722,N_6348);
nand U8668 (N_8668,N_6839,N_7246);
and U8669 (N_8669,N_5071,N_6041);
xnor U8670 (N_8670,N_5269,N_5486);
and U8671 (N_8671,N_6333,N_5436);
or U8672 (N_8672,N_5972,N_7177);
xor U8673 (N_8673,N_7453,N_6453);
or U8674 (N_8674,N_5156,N_5987);
nor U8675 (N_8675,N_6106,N_6978);
nor U8676 (N_8676,N_6468,N_5519);
and U8677 (N_8677,N_5193,N_7081);
xor U8678 (N_8678,N_5580,N_5696);
or U8679 (N_8679,N_5816,N_5197);
nand U8680 (N_8680,N_6124,N_5118);
nor U8681 (N_8681,N_6906,N_6107);
nor U8682 (N_8682,N_6343,N_5351);
nand U8683 (N_8683,N_7086,N_5430);
nor U8684 (N_8684,N_5135,N_5645);
nand U8685 (N_8685,N_5368,N_6657);
nor U8686 (N_8686,N_7190,N_6914);
and U8687 (N_8687,N_7072,N_5946);
nand U8688 (N_8688,N_7248,N_5408);
nor U8689 (N_8689,N_5093,N_5092);
or U8690 (N_8690,N_6820,N_7424);
nand U8691 (N_8691,N_6905,N_6071);
nor U8692 (N_8692,N_6669,N_6806);
and U8693 (N_8693,N_5759,N_6648);
nor U8694 (N_8694,N_7440,N_6399);
or U8695 (N_8695,N_7315,N_7108);
nand U8696 (N_8696,N_7284,N_5123);
nand U8697 (N_8697,N_5711,N_6229);
or U8698 (N_8698,N_7228,N_5847);
and U8699 (N_8699,N_6155,N_6115);
and U8700 (N_8700,N_6765,N_6612);
nor U8701 (N_8701,N_6258,N_6467);
and U8702 (N_8702,N_6979,N_6159);
or U8703 (N_8703,N_6054,N_6391);
nand U8704 (N_8704,N_5103,N_5540);
xor U8705 (N_8705,N_5228,N_5426);
and U8706 (N_8706,N_5127,N_6533);
and U8707 (N_8707,N_6389,N_5059);
nor U8708 (N_8708,N_5439,N_5861);
or U8709 (N_8709,N_5666,N_7084);
xnor U8710 (N_8710,N_5778,N_6455);
xor U8711 (N_8711,N_5245,N_5849);
and U8712 (N_8712,N_6424,N_6131);
nor U8713 (N_8713,N_6892,N_5864);
xnor U8714 (N_8714,N_5382,N_5826);
nand U8715 (N_8715,N_5597,N_7215);
nor U8716 (N_8716,N_5285,N_6619);
nor U8717 (N_8717,N_5774,N_5995);
nand U8718 (N_8718,N_6023,N_5045);
or U8719 (N_8719,N_5601,N_7128);
or U8720 (N_8720,N_6171,N_5738);
nand U8721 (N_8721,N_5654,N_5239);
or U8722 (N_8722,N_7301,N_5966);
and U8723 (N_8723,N_7484,N_6563);
or U8724 (N_8724,N_6025,N_5491);
or U8725 (N_8725,N_6008,N_5804);
xnor U8726 (N_8726,N_6506,N_6052);
and U8727 (N_8727,N_5201,N_5331);
xor U8728 (N_8728,N_5333,N_6268);
nand U8729 (N_8729,N_5209,N_7038);
and U8730 (N_8730,N_7323,N_5952);
and U8731 (N_8731,N_7224,N_6782);
nor U8732 (N_8732,N_6508,N_5559);
nand U8733 (N_8733,N_6975,N_5818);
xnor U8734 (N_8734,N_6885,N_5081);
xnor U8735 (N_8735,N_5892,N_7233);
nand U8736 (N_8736,N_5637,N_6083);
and U8737 (N_8737,N_5708,N_6466);
nand U8738 (N_8738,N_6411,N_6799);
nand U8739 (N_8739,N_6254,N_6747);
nand U8740 (N_8740,N_6297,N_5872);
xnor U8741 (N_8741,N_6938,N_5507);
and U8742 (N_8742,N_6788,N_5974);
nor U8743 (N_8743,N_7336,N_5474);
nor U8744 (N_8744,N_6713,N_6827);
nor U8745 (N_8745,N_6253,N_5337);
and U8746 (N_8746,N_7179,N_5002);
nand U8747 (N_8747,N_5884,N_5224);
and U8748 (N_8748,N_6871,N_6102);
or U8749 (N_8749,N_5907,N_7002);
or U8750 (N_8750,N_7343,N_6268);
xnor U8751 (N_8751,N_7041,N_7359);
or U8752 (N_8752,N_6849,N_6571);
nand U8753 (N_8753,N_5538,N_6325);
xnor U8754 (N_8754,N_6998,N_5219);
nand U8755 (N_8755,N_6797,N_6644);
or U8756 (N_8756,N_7190,N_5349);
and U8757 (N_8757,N_5569,N_7251);
and U8758 (N_8758,N_5810,N_7220);
nand U8759 (N_8759,N_5687,N_5226);
nor U8760 (N_8760,N_6539,N_5937);
and U8761 (N_8761,N_7007,N_7389);
and U8762 (N_8762,N_6322,N_6804);
nand U8763 (N_8763,N_5741,N_7144);
nor U8764 (N_8764,N_6286,N_6865);
and U8765 (N_8765,N_7009,N_5843);
and U8766 (N_8766,N_7273,N_7297);
nand U8767 (N_8767,N_5477,N_6808);
xnor U8768 (N_8768,N_6693,N_7257);
or U8769 (N_8769,N_5738,N_6423);
nor U8770 (N_8770,N_5191,N_6790);
or U8771 (N_8771,N_6507,N_6506);
and U8772 (N_8772,N_5591,N_5864);
nand U8773 (N_8773,N_6075,N_5284);
and U8774 (N_8774,N_5389,N_6304);
and U8775 (N_8775,N_5021,N_5802);
xnor U8776 (N_8776,N_5302,N_5128);
xor U8777 (N_8777,N_5803,N_7052);
and U8778 (N_8778,N_6197,N_6867);
and U8779 (N_8779,N_6431,N_7095);
nand U8780 (N_8780,N_6459,N_5116);
or U8781 (N_8781,N_5362,N_7471);
nor U8782 (N_8782,N_5834,N_5012);
nand U8783 (N_8783,N_6667,N_7441);
xnor U8784 (N_8784,N_7119,N_5927);
or U8785 (N_8785,N_7268,N_6875);
and U8786 (N_8786,N_6358,N_6593);
or U8787 (N_8787,N_7170,N_5869);
or U8788 (N_8788,N_5527,N_7012);
and U8789 (N_8789,N_5281,N_5118);
nand U8790 (N_8790,N_5076,N_6893);
and U8791 (N_8791,N_5161,N_5306);
or U8792 (N_8792,N_5620,N_6456);
nor U8793 (N_8793,N_5594,N_6901);
xnor U8794 (N_8794,N_5828,N_5586);
xnor U8795 (N_8795,N_7259,N_5113);
xor U8796 (N_8796,N_5843,N_6164);
nor U8797 (N_8797,N_6634,N_5354);
nand U8798 (N_8798,N_5528,N_5755);
xnor U8799 (N_8799,N_7101,N_6977);
xnor U8800 (N_8800,N_5196,N_5584);
or U8801 (N_8801,N_6695,N_6321);
xnor U8802 (N_8802,N_7386,N_6518);
or U8803 (N_8803,N_5646,N_5996);
nand U8804 (N_8804,N_6929,N_7114);
xor U8805 (N_8805,N_7347,N_5494);
xor U8806 (N_8806,N_6336,N_5741);
nor U8807 (N_8807,N_6002,N_5202);
xor U8808 (N_8808,N_6260,N_5645);
nor U8809 (N_8809,N_6695,N_6178);
and U8810 (N_8810,N_6976,N_5353);
and U8811 (N_8811,N_6131,N_6948);
and U8812 (N_8812,N_5000,N_6880);
nand U8813 (N_8813,N_5441,N_6599);
xnor U8814 (N_8814,N_5938,N_5491);
xor U8815 (N_8815,N_6648,N_5689);
or U8816 (N_8816,N_6910,N_6881);
nand U8817 (N_8817,N_6315,N_6697);
nor U8818 (N_8818,N_5088,N_7156);
nor U8819 (N_8819,N_7142,N_5930);
xnor U8820 (N_8820,N_5935,N_5107);
and U8821 (N_8821,N_6336,N_5013);
nor U8822 (N_8822,N_5581,N_5824);
or U8823 (N_8823,N_5770,N_6395);
nand U8824 (N_8824,N_7449,N_6608);
and U8825 (N_8825,N_6155,N_5170);
nor U8826 (N_8826,N_6834,N_6116);
nor U8827 (N_8827,N_5291,N_5373);
xor U8828 (N_8828,N_7026,N_6775);
nand U8829 (N_8829,N_5990,N_5408);
and U8830 (N_8830,N_6589,N_5686);
or U8831 (N_8831,N_6109,N_6058);
nand U8832 (N_8832,N_5992,N_6126);
nor U8833 (N_8833,N_5152,N_6973);
xnor U8834 (N_8834,N_6821,N_5230);
or U8835 (N_8835,N_7376,N_5852);
or U8836 (N_8836,N_7472,N_7035);
and U8837 (N_8837,N_6688,N_5562);
and U8838 (N_8838,N_6315,N_6492);
and U8839 (N_8839,N_5294,N_5522);
nor U8840 (N_8840,N_5606,N_6563);
and U8841 (N_8841,N_7137,N_7160);
xnor U8842 (N_8842,N_5800,N_5397);
nor U8843 (N_8843,N_7372,N_6016);
xnor U8844 (N_8844,N_5287,N_5449);
and U8845 (N_8845,N_6662,N_6521);
nand U8846 (N_8846,N_7260,N_6078);
or U8847 (N_8847,N_6549,N_7203);
nand U8848 (N_8848,N_6180,N_6280);
and U8849 (N_8849,N_7187,N_7325);
xor U8850 (N_8850,N_5284,N_6538);
or U8851 (N_8851,N_7387,N_6599);
and U8852 (N_8852,N_6136,N_6104);
xor U8853 (N_8853,N_5438,N_5909);
or U8854 (N_8854,N_5993,N_7458);
xnor U8855 (N_8855,N_6021,N_7087);
and U8856 (N_8856,N_5318,N_6631);
xor U8857 (N_8857,N_7227,N_6847);
or U8858 (N_8858,N_5003,N_6216);
or U8859 (N_8859,N_5763,N_5332);
or U8860 (N_8860,N_5213,N_5425);
nor U8861 (N_8861,N_5533,N_5127);
or U8862 (N_8862,N_5880,N_7335);
xor U8863 (N_8863,N_7173,N_5889);
nor U8864 (N_8864,N_6470,N_7450);
xnor U8865 (N_8865,N_5627,N_5700);
or U8866 (N_8866,N_5285,N_6667);
or U8867 (N_8867,N_7088,N_6424);
nand U8868 (N_8868,N_6455,N_6698);
nor U8869 (N_8869,N_5647,N_7079);
or U8870 (N_8870,N_6458,N_6493);
and U8871 (N_8871,N_7343,N_5702);
or U8872 (N_8872,N_6192,N_6852);
or U8873 (N_8873,N_5208,N_5379);
nor U8874 (N_8874,N_5983,N_6490);
nand U8875 (N_8875,N_5454,N_5785);
and U8876 (N_8876,N_6991,N_7066);
nand U8877 (N_8877,N_5963,N_5780);
nand U8878 (N_8878,N_6362,N_6647);
or U8879 (N_8879,N_6134,N_5524);
and U8880 (N_8880,N_7011,N_5761);
and U8881 (N_8881,N_7158,N_5834);
xor U8882 (N_8882,N_6449,N_7304);
nand U8883 (N_8883,N_6578,N_7457);
and U8884 (N_8884,N_5050,N_7024);
nand U8885 (N_8885,N_5567,N_5202);
xnor U8886 (N_8886,N_6799,N_5161);
and U8887 (N_8887,N_5770,N_6499);
or U8888 (N_8888,N_5805,N_5667);
nand U8889 (N_8889,N_5161,N_5440);
nand U8890 (N_8890,N_6827,N_5038);
nand U8891 (N_8891,N_7111,N_7020);
nand U8892 (N_8892,N_6742,N_5710);
or U8893 (N_8893,N_6966,N_5582);
xor U8894 (N_8894,N_6037,N_6576);
or U8895 (N_8895,N_5525,N_5710);
or U8896 (N_8896,N_5370,N_5756);
nor U8897 (N_8897,N_6861,N_5473);
xor U8898 (N_8898,N_5394,N_6859);
and U8899 (N_8899,N_6913,N_5016);
or U8900 (N_8900,N_5527,N_6648);
or U8901 (N_8901,N_6820,N_5977);
nor U8902 (N_8902,N_7330,N_7365);
nor U8903 (N_8903,N_6812,N_7403);
and U8904 (N_8904,N_6228,N_7406);
xor U8905 (N_8905,N_6235,N_5439);
or U8906 (N_8906,N_7043,N_7168);
and U8907 (N_8907,N_6154,N_6885);
nand U8908 (N_8908,N_5125,N_5026);
and U8909 (N_8909,N_6543,N_6602);
nand U8910 (N_8910,N_5112,N_6752);
nor U8911 (N_8911,N_5105,N_7148);
or U8912 (N_8912,N_5869,N_7181);
xor U8913 (N_8913,N_5735,N_5268);
or U8914 (N_8914,N_5745,N_6887);
nand U8915 (N_8915,N_5349,N_7116);
nand U8916 (N_8916,N_5809,N_6972);
or U8917 (N_8917,N_6184,N_6728);
nor U8918 (N_8918,N_6013,N_5416);
nand U8919 (N_8919,N_7285,N_6141);
xor U8920 (N_8920,N_5605,N_5563);
xnor U8921 (N_8921,N_6094,N_5653);
xnor U8922 (N_8922,N_6849,N_6839);
nand U8923 (N_8923,N_7157,N_6087);
xor U8924 (N_8924,N_6961,N_5317);
nor U8925 (N_8925,N_6483,N_7108);
nor U8926 (N_8926,N_7079,N_6544);
nor U8927 (N_8927,N_5290,N_5549);
xnor U8928 (N_8928,N_6756,N_5963);
nand U8929 (N_8929,N_6281,N_5714);
or U8930 (N_8930,N_6745,N_6360);
or U8931 (N_8931,N_5773,N_6721);
and U8932 (N_8932,N_6497,N_5725);
or U8933 (N_8933,N_5963,N_6099);
and U8934 (N_8934,N_5515,N_5671);
xor U8935 (N_8935,N_7448,N_5125);
xor U8936 (N_8936,N_5037,N_6235);
or U8937 (N_8937,N_6205,N_6059);
xnor U8938 (N_8938,N_6296,N_6364);
and U8939 (N_8939,N_7366,N_7224);
nor U8940 (N_8940,N_5411,N_5657);
xnor U8941 (N_8941,N_7365,N_5405);
and U8942 (N_8942,N_7491,N_7346);
nand U8943 (N_8943,N_5587,N_5795);
or U8944 (N_8944,N_6992,N_5612);
xnor U8945 (N_8945,N_5689,N_5929);
xor U8946 (N_8946,N_6142,N_5420);
and U8947 (N_8947,N_5021,N_7047);
nand U8948 (N_8948,N_6410,N_6018);
and U8949 (N_8949,N_6173,N_7482);
xnor U8950 (N_8950,N_6194,N_5587);
and U8951 (N_8951,N_5778,N_6628);
xor U8952 (N_8952,N_6541,N_6387);
and U8953 (N_8953,N_6543,N_6851);
nor U8954 (N_8954,N_7226,N_7166);
and U8955 (N_8955,N_6203,N_7081);
nor U8956 (N_8956,N_6381,N_5366);
xnor U8957 (N_8957,N_7034,N_5768);
nor U8958 (N_8958,N_5775,N_7312);
or U8959 (N_8959,N_5335,N_6468);
xnor U8960 (N_8960,N_5095,N_6769);
and U8961 (N_8961,N_5269,N_5373);
xnor U8962 (N_8962,N_5357,N_5264);
xor U8963 (N_8963,N_6693,N_5897);
nand U8964 (N_8964,N_5071,N_6394);
xnor U8965 (N_8965,N_6698,N_5383);
nand U8966 (N_8966,N_5139,N_5121);
or U8967 (N_8967,N_7007,N_7293);
nand U8968 (N_8968,N_5502,N_5172);
nand U8969 (N_8969,N_5413,N_5644);
or U8970 (N_8970,N_5465,N_7265);
and U8971 (N_8971,N_7249,N_6001);
nand U8972 (N_8972,N_6211,N_6495);
or U8973 (N_8973,N_5233,N_5925);
nor U8974 (N_8974,N_6355,N_6683);
nand U8975 (N_8975,N_6766,N_5941);
xor U8976 (N_8976,N_7364,N_5940);
nor U8977 (N_8977,N_7130,N_5665);
nand U8978 (N_8978,N_5782,N_7030);
xnor U8979 (N_8979,N_6230,N_7018);
nand U8980 (N_8980,N_6964,N_6835);
nand U8981 (N_8981,N_5990,N_5421);
nand U8982 (N_8982,N_5577,N_7010);
and U8983 (N_8983,N_6079,N_6364);
xor U8984 (N_8984,N_7246,N_7229);
nand U8985 (N_8985,N_6780,N_5538);
and U8986 (N_8986,N_5103,N_6027);
or U8987 (N_8987,N_6528,N_6750);
and U8988 (N_8988,N_5741,N_5769);
and U8989 (N_8989,N_7332,N_6690);
xor U8990 (N_8990,N_6193,N_7303);
xor U8991 (N_8991,N_7296,N_5881);
nand U8992 (N_8992,N_5860,N_5757);
or U8993 (N_8993,N_7339,N_5778);
nand U8994 (N_8994,N_5418,N_6088);
nor U8995 (N_8995,N_5772,N_7428);
or U8996 (N_8996,N_7294,N_5847);
xnor U8997 (N_8997,N_6160,N_5532);
nand U8998 (N_8998,N_5748,N_7379);
or U8999 (N_8999,N_5293,N_7389);
xor U9000 (N_9000,N_6822,N_5871);
xor U9001 (N_9001,N_6698,N_6219);
or U9002 (N_9002,N_6189,N_7330);
or U9003 (N_9003,N_5373,N_5799);
nor U9004 (N_9004,N_7406,N_7405);
or U9005 (N_9005,N_5362,N_6615);
and U9006 (N_9006,N_7361,N_5393);
nand U9007 (N_9007,N_7378,N_7320);
nand U9008 (N_9008,N_5702,N_5180);
nor U9009 (N_9009,N_6794,N_5663);
and U9010 (N_9010,N_5198,N_7345);
xor U9011 (N_9011,N_5311,N_5093);
and U9012 (N_9012,N_5508,N_5634);
xnor U9013 (N_9013,N_5882,N_7211);
xnor U9014 (N_9014,N_5831,N_6361);
and U9015 (N_9015,N_6541,N_6143);
nor U9016 (N_9016,N_6940,N_5327);
nand U9017 (N_9017,N_6821,N_5389);
and U9018 (N_9018,N_5707,N_6769);
and U9019 (N_9019,N_6361,N_5655);
nor U9020 (N_9020,N_6401,N_6966);
nor U9021 (N_9021,N_6254,N_6936);
and U9022 (N_9022,N_5822,N_6664);
nand U9023 (N_9023,N_7003,N_5273);
xor U9024 (N_9024,N_6157,N_6067);
and U9025 (N_9025,N_6777,N_6546);
or U9026 (N_9026,N_6095,N_5885);
and U9027 (N_9027,N_5816,N_5162);
xor U9028 (N_9028,N_7101,N_5914);
xor U9029 (N_9029,N_6189,N_5431);
nor U9030 (N_9030,N_7305,N_6019);
xnor U9031 (N_9031,N_6040,N_5056);
or U9032 (N_9032,N_6080,N_5796);
and U9033 (N_9033,N_7308,N_6446);
and U9034 (N_9034,N_6595,N_5030);
or U9035 (N_9035,N_6740,N_7405);
or U9036 (N_9036,N_7422,N_6164);
nand U9037 (N_9037,N_6115,N_6453);
and U9038 (N_9038,N_5891,N_7427);
or U9039 (N_9039,N_6967,N_5252);
nand U9040 (N_9040,N_5755,N_7088);
and U9041 (N_9041,N_7374,N_6315);
or U9042 (N_9042,N_7131,N_7075);
nor U9043 (N_9043,N_7397,N_7052);
xnor U9044 (N_9044,N_6905,N_6259);
xnor U9045 (N_9045,N_5649,N_6805);
nand U9046 (N_9046,N_5517,N_5637);
nor U9047 (N_9047,N_6050,N_6454);
or U9048 (N_9048,N_7084,N_5543);
nor U9049 (N_9049,N_6070,N_5526);
or U9050 (N_9050,N_5017,N_6907);
nand U9051 (N_9051,N_5299,N_7059);
or U9052 (N_9052,N_5388,N_5149);
and U9053 (N_9053,N_5164,N_6261);
and U9054 (N_9054,N_6026,N_6574);
xnor U9055 (N_9055,N_6433,N_5061);
and U9056 (N_9056,N_6577,N_6914);
nor U9057 (N_9057,N_5993,N_6882);
nor U9058 (N_9058,N_6151,N_5922);
and U9059 (N_9059,N_5349,N_6534);
or U9060 (N_9060,N_5302,N_6967);
and U9061 (N_9061,N_5803,N_5897);
and U9062 (N_9062,N_6882,N_6331);
xnor U9063 (N_9063,N_6821,N_5610);
xnor U9064 (N_9064,N_6207,N_5819);
and U9065 (N_9065,N_5617,N_5021);
nand U9066 (N_9066,N_5210,N_6621);
or U9067 (N_9067,N_6727,N_6197);
or U9068 (N_9068,N_5605,N_7000);
or U9069 (N_9069,N_5497,N_6723);
xor U9070 (N_9070,N_6896,N_5300);
and U9071 (N_9071,N_5774,N_5453);
and U9072 (N_9072,N_6403,N_6535);
xnor U9073 (N_9073,N_7257,N_5467);
nor U9074 (N_9074,N_5847,N_5543);
xnor U9075 (N_9075,N_6791,N_5739);
nand U9076 (N_9076,N_6047,N_5189);
or U9077 (N_9077,N_6186,N_6554);
or U9078 (N_9078,N_7114,N_5240);
nor U9079 (N_9079,N_5428,N_5250);
or U9080 (N_9080,N_6069,N_5843);
nor U9081 (N_9081,N_5748,N_5250);
xor U9082 (N_9082,N_6778,N_6793);
nor U9083 (N_9083,N_6753,N_6550);
nor U9084 (N_9084,N_5323,N_5681);
nor U9085 (N_9085,N_5680,N_6608);
and U9086 (N_9086,N_6242,N_5753);
or U9087 (N_9087,N_5923,N_7150);
nor U9088 (N_9088,N_5374,N_7020);
xnor U9089 (N_9089,N_7337,N_7498);
xor U9090 (N_9090,N_6764,N_5173);
xor U9091 (N_9091,N_6302,N_6717);
or U9092 (N_9092,N_7144,N_6047);
xnor U9093 (N_9093,N_7151,N_5231);
xor U9094 (N_9094,N_5608,N_5673);
and U9095 (N_9095,N_6083,N_6115);
nand U9096 (N_9096,N_6511,N_7409);
and U9097 (N_9097,N_5723,N_5614);
xor U9098 (N_9098,N_5502,N_5976);
and U9099 (N_9099,N_6224,N_6460);
and U9100 (N_9100,N_7121,N_6969);
and U9101 (N_9101,N_6722,N_5408);
or U9102 (N_9102,N_6003,N_6951);
xnor U9103 (N_9103,N_5344,N_5491);
and U9104 (N_9104,N_7248,N_5771);
and U9105 (N_9105,N_6475,N_7148);
nand U9106 (N_9106,N_5429,N_5141);
xnor U9107 (N_9107,N_5023,N_5055);
and U9108 (N_9108,N_7490,N_5471);
or U9109 (N_9109,N_6004,N_6691);
xnor U9110 (N_9110,N_5241,N_5705);
nand U9111 (N_9111,N_6470,N_6466);
and U9112 (N_9112,N_5228,N_5169);
nand U9113 (N_9113,N_5676,N_6599);
xor U9114 (N_9114,N_7157,N_6082);
nor U9115 (N_9115,N_5986,N_6324);
and U9116 (N_9116,N_5217,N_5742);
xor U9117 (N_9117,N_6566,N_5634);
and U9118 (N_9118,N_7108,N_6973);
xnor U9119 (N_9119,N_5520,N_5404);
nand U9120 (N_9120,N_6480,N_5815);
nor U9121 (N_9121,N_6376,N_5311);
nand U9122 (N_9122,N_7133,N_7416);
and U9123 (N_9123,N_6516,N_6886);
and U9124 (N_9124,N_7262,N_6772);
nand U9125 (N_9125,N_7243,N_6525);
and U9126 (N_9126,N_5205,N_5628);
xor U9127 (N_9127,N_5640,N_6225);
and U9128 (N_9128,N_5831,N_5661);
nor U9129 (N_9129,N_7368,N_6722);
and U9130 (N_9130,N_5240,N_6802);
and U9131 (N_9131,N_7132,N_5324);
or U9132 (N_9132,N_5367,N_5195);
nand U9133 (N_9133,N_6507,N_6939);
and U9134 (N_9134,N_6202,N_5080);
nand U9135 (N_9135,N_6455,N_5033);
or U9136 (N_9136,N_6855,N_6723);
xor U9137 (N_9137,N_7438,N_6152);
nand U9138 (N_9138,N_5708,N_6501);
and U9139 (N_9139,N_7135,N_7342);
nand U9140 (N_9140,N_6080,N_6649);
or U9141 (N_9141,N_7472,N_6987);
nor U9142 (N_9142,N_5686,N_5662);
xnor U9143 (N_9143,N_5574,N_7449);
or U9144 (N_9144,N_5267,N_6402);
nor U9145 (N_9145,N_6555,N_7387);
xor U9146 (N_9146,N_7145,N_5522);
or U9147 (N_9147,N_6422,N_7447);
nand U9148 (N_9148,N_5804,N_5540);
nand U9149 (N_9149,N_5928,N_5688);
xnor U9150 (N_9150,N_7370,N_5152);
and U9151 (N_9151,N_5899,N_6987);
xnor U9152 (N_9152,N_6126,N_5824);
nand U9153 (N_9153,N_6807,N_5784);
nand U9154 (N_9154,N_7441,N_5525);
nand U9155 (N_9155,N_6879,N_7204);
nand U9156 (N_9156,N_7121,N_5100);
nor U9157 (N_9157,N_5368,N_6142);
xnor U9158 (N_9158,N_6135,N_5034);
xor U9159 (N_9159,N_6636,N_6702);
nor U9160 (N_9160,N_5396,N_6562);
nand U9161 (N_9161,N_6032,N_7014);
or U9162 (N_9162,N_5994,N_5777);
nand U9163 (N_9163,N_5960,N_5117);
or U9164 (N_9164,N_6485,N_5528);
or U9165 (N_9165,N_5325,N_5837);
and U9166 (N_9166,N_6326,N_7107);
or U9167 (N_9167,N_6805,N_6273);
and U9168 (N_9168,N_5837,N_6810);
or U9169 (N_9169,N_6403,N_7074);
nand U9170 (N_9170,N_5325,N_5025);
xor U9171 (N_9171,N_6107,N_5542);
or U9172 (N_9172,N_5109,N_5105);
xor U9173 (N_9173,N_5954,N_7129);
and U9174 (N_9174,N_5937,N_7111);
nor U9175 (N_9175,N_7103,N_5066);
and U9176 (N_9176,N_6598,N_6067);
nor U9177 (N_9177,N_5809,N_5548);
xnor U9178 (N_9178,N_5575,N_6208);
nand U9179 (N_9179,N_6011,N_5110);
or U9180 (N_9180,N_6028,N_6315);
and U9181 (N_9181,N_7239,N_6624);
or U9182 (N_9182,N_5788,N_5312);
or U9183 (N_9183,N_7451,N_6944);
nand U9184 (N_9184,N_5091,N_7428);
xor U9185 (N_9185,N_6796,N_7223);
nand U9186 (N_9186,N_7427,N_5653);
nor U9187 (N_9187,N_7067,N_6845);
and U9188 (N_9188,N_6623,N_7194);
nand U9189 (N_9189,N_5971,N_5342);
xor U9190 (N_9190,N_5662,N_6277);
nor U9191 (N_9191,N_6398,N_5491);
nor U9192 (N_9192,N_5894,N_5920);
nor U9193 (N_9193,N_6143,N_5615);
xor U9194 (N_9194,N_5474,N_5351);
nand U9195 (N_9195,N_5614,N_6257);
and U9196 (N_9196,N_5179,N_5316);
nor U9197 (N_9197,N_6102,N_6321);
nand U9198 (N_9198,N_6575,N_5282);
nand U9199 (N_9199,N_7291,N_6199);
or U9200 (N_9200,N_7490,N_6937);
and U9201 (N_9201,N_5067,N_6885);
or U9202 (N_9202,N_6216,N_5767);
nand U9203 (N_9203,N_5739,N_6267);
and U9204 (N_9204,N_5681,N_5882);
nor U9205 (N_9205,N_5589,N_7490);
or U9206 (N_9206,N_5911,N_7308);
or U9207 (N_9207,N_5527,N_5828);
or U9208 (N_9208,N_7485,N_5513);
and U9209 (N_9209,N_6661,N_6326);
nor U9210 (N_9210,N_7255,N_5647);
nor U9211 (N_9211,N_6833,N_6825);
or U9212 (N_9212,N_7156,N_6113);
or U9213 (N_9213,N_6103,N_5003);
xor U9214 (N_9214,N_5167,N_6426);
nand U9215 (N_9215,N_7312,N_7398);
xor U9216 (N_9216,N_5689,N_6880);
xnor U9217 (N_9217,N_7234,N_7306);
xor U9218 (N_9218,N_7215,N_6065);
and U9219 (N_9219,N_6115,N_6450);
and U9220 (N_9220,N_6510,N_5373);
xor U9221 (N_9221,N_5733,N_5723);
nand U9222 (N_9222,N_6612,N_6250);
xor U9223 (N_9223,N_7218,N_6042);
xnor U9224 (N_9224,N_5676,N_6433);
nor U9225 (N_9225,N_6571,N_5241);
nor U9226 (N_9226,N_6520,N_5989);
and U9227 (N_9227,N_6915,N_6541);
nor U9228 (N_9228,N_7117,N_5108);
or U9229 (N_9229,N_7257,N_5417);
nand U9230 (N_9230,N_6401,N_7399);
nand U9231 (N_9231,N_6668,N_6852);
nand U9232 (N_9232,N_6996,N_6630);
nor U9233 (N_9233,N_6150,N_6525);
or U9234 (N_9234,N_6516,N_5483);
and U9235 (N_9235,N_6252,N_7277);
and U9236 (N_9236,N_6848,N_5646);
xnor U9237 (N_9237,N_5958,N_5558);
and U9238 (N_9238,N_5326,N_7418);
and U9239 (N_9239,N_7072,N_5841);
nor U9240 (N_9240,N_6260,N_6076);
nor U9241 (N_9241,N_5965,N_6800);
xnor U9242 (N_9242,N_7066,N_7498);
nor U9243 (N_9243,N_6284,N_7326);
and U9244 (N_9244,N_7306,N_7440);
nand U9245 (N_9245,N_6709,N_6610);
xor U9246 (N_9246,N_5661,N_5161);
xor U9247 (N_9247,N_7391,N_5226);
nand U9248 (N_9248,N_7385,N_7450);
or U9249 (N_9249,N_7129,N_6136);
xor U9250 (N_9250,N_6602,N_6215);
nand U9251 (N_9251,N_5773,N_6355);
nor U9252 (N_9252,N_6276,N_5510);
nor U9253 (N_9253,N_5409,N_6158);
nor U9254 (N_9254,N_6990,N_6998);
nand U9255 (N_9255,N_5074,N_5207);
nand U9256 (N_9256,N_5904,N_7393);
or U9257 (N_9257,N_7321,N_5029);
nand U9258 (N_9258,N_6012,N_5297);
and U9259 (N_9259,N_5190,N_5964);
or U9260 (N_9260,N_6228,N_6046);
nand U9261 (N_9261,N_6939,N_5373);
and U9262 (N_9262,N_5467,N_7248);
or U9263 (N_9263,N_5834,N_5470);
nor U9264 (N_9264,N_5663,N_6366);
and U9265 (N_9265,N_7315,N_6825);
nor U9266 (N_9266,N_5550,N_6830);
nor U9267 (N_9267,N_7467,N_5701);
xnor U9268 (N_9268,N_5708,N_5946);
nand U9269 (N_9269,N_7399,N_5071);
xor U9270 (N_9270,N_7336,N_6049);
or U9271 (N_9271,N_6680,N_5878);
nor U9272 (N_9272,N_7219,N_7115);
or U9273 (N_9273,N_5033,N_5153);
nor U9274 (N_9274,N_6453,N_5348);
nand U9275 (N_9275,N_5021,N_7301);
nor U9276 (N_9276,N_5255,N_5998);
and U9277 (N_9277,N_6688,N_6795);
and U9278 (N_9278,N_6944,N_6816);
or U9279 (N_9279,N_7040,N_6472);
nor U9280 (N_9280,N_7238,N_5912);
xnor U9281 (N_9281,N_5128,N_7161);
nand U9282 (N_9282,N_5596,N_6383);
xor U9283 (N_9283,N_5516,N_7303);
xnor U9284 (N_9284,N_6228,N_7389);
nor U9285 (N_9285,N_6452,N_5605);
nor U9286 (N_9286,N_6877,N_7170);
nand U9287 (N_9287,N_7339,N_6320);
nand U9288 (N_9288,N_6963,N_6406);
nor U9289 (N_9289,N_5760,N_6761);
or U9290 (N_9290,N_5379,N_5556);
or U9291 (N_9291,N_7113,N_7439);
and U9292 (N_9292,N_6299,N_6633);
xor U9293 (N_9293,N_6011,N_5340);
nor U9294 (N_9294,N_7465,N_6225);
or U9295 (N_9295,N_7456,N_7356);
or U9296 (N_9296,N_6309,N_5948);
nor U9297 (N_9297,N_5775,N_6378);
nor U9298 (N_9298,N_7108,N_5501);
or U9299 (N_9299,N_6185,N_7180);
xnor U9300 (N_9300,N_7005,N_6782);
and U9301 (N_9301,N_6215,N_6941);
or U9302 (N_9302,N_6124,N_5889);
xor U9303 (N_9303,N_7324,N_6649);
xnor U9304 (N_9304,N_6121,N_5262);
nor U9305 (N_9305,N_5664,N_6147);
and U9306 (N_9306,N_5473,N_6116);
xnor U9307 (N_9307,N_5984,N_5840);
xor U9308 (N_9308,N_6635,N_6765);
xor U9309 (N_9309,N_6813,N_6994);
or U9310 (N_9310,N_6563,N_6177);
or U9311 (N_9311,N_5542,N_7315);
xnor U9312 (N_9312,N_6056,N_6272);
or U9313 (N_9313,N_7336,N_6110);
and U9314 (N_9314,N_5105,N_7071);
nor U9315 (N_9315,N_5548,N_6252);
and U9316 (N_9316,N_6003,N_5825);
or U9317 (N_9317,N_5963,N_6428);
or U9318 (N_9318,N_7313,N_5822);
xnor U9319 (N_9319,N_5834,N_6623);
and U9320 (N_9320,N_6206,N_6582);
xnor U9321 (N_9321,N_5918,N_6446);
and U9322 (N_9322,N_7311,N_7105);
or U9323 (N_9323,N_7053,N_5825);
nand U9324 (N_9324,N_7299,N_6472);
xnor U9325 (N_9325,N_6618,N_7091);
or U9326 (N_9326,N_6794,N_7165);
nor U9327 (N_9327,N_5334,N_5933);
or U9328 (N_9328,N_5247,N_7014);
or U9329 (N_9329,N_6550,N_6417);
and U9330 (N_9330,N_6271,N_5023);
and U9331 (N_9331,N_6429,N_6816);
nor U9332 (N_9332,N_6791,N_5411);
nor U9333 (N_9333,N_6107,N_6533);
xor U9334 (N_9334,N_7176,N_6608);
nand U9335 (N_9335,N_7442,N_6120);
nor U9336 (N_9336,N_7041,N_5620);
and U9337 (N_9337,N_6509,N_7273);
xor U9338 (N_9338,N_6127,N_5428);
and U9339 (N_9339,N_5683,N_6405);
or U9340 (N_9340,N_7151,N_6745);
nor U9341 (N_9341,N_7046,N_7275);
and U9342 (N_9342,N_5038,N_6322);
xnor U9343 (N_9343,N_5888,N_6743);
and U9344 (N_9344,N_5471,N_5504);
nor U9345 (N_9345,N_6133,N_6021);
nand U9346 (N_9346,N_5133,N_6527);
nor U9347 (N_9347,N_7443,N_6586);
nor U9348 (N_9348,N_6920,N_5874);
and U9349 (N_9349,N_6296,N_7339);
xnor U9350 (N_9350,N_6585,N_7243);
and U9351 (N_9351,N_7230,N_6832);
xor U9352 (N_9352,N_6472,N_6477);
xnor U9353 (N_9353,N_5067,N_7469);
nand U9354 (N_9354,N_5518,N_5112);
nand U9355 (N_9355,N_5400,N_5195);
nand U9356 (N_9356,N_5549,N_7321);
and U9357 (N_9357,N_5545,N_5702);
or U9358 (N_9358,N_5785,N_5970);
or U9359 (N_9359,N_7200,N_6421);
nor U9360 (N_9360,N_6905,N_5622);
nand U9361 (N_9361,N_6110,N_7391);
xor U9362 (N_9362,N_6358,N_6988);
nor U9363 (N_9363,N_5853,N_5287);
nand U9364 (N_9364,N_5775,N_6481);
xnor U9365 (N_9365,N_5998,N_7464);
nand U9366 (N_9366,N_7355,N_6317);
and U9367 (N_9367,N_6753,N_5634);
nor U9368 (N_9368,N_7248,N_5033);
xnor U9369 (N_9369,N_6918,N_5936);
and U9370 (N_9370,N_5341,N_5843);
xnor U9371 (N_9371,N_6815,N_5578);
xnor U9372 (N_9372,N_6693,N_6997);
nand U9373 (N_9373,N_5821,N_5958);
nand U9374 (N_9374,N_5944,N_6673);
or U9375 (N_9375,N_7293,N_6075);
or U9376 (N_9376,N_7244,N_5919);
and U9377 (N_9377,N_5342,N_6578);
and U9378 (N_9378,N_6666,N_7140);
nor U9379 (N_9379,N_6131,N_5801);
or U9380 (N_9380,N_6320,N_6354);
and U9381 (N_9381,N_5044,N_6693);
or U9382 (N_9382,N_6742,N_6037);
and U9383 (N_9383,N_6213,N_6864);
nor U9384 (N_9384,N_5440,N_5475);
and U9385 (N_9385,N_6860,N_5974);
nor U9386 (N_9386,N_6271,N_6042);
nor U9387 (N_9387,N_5918,N_5649);
and U9388 (N_9388,N_6285,N_5618);
xor U9389 (N_9389,N_6795,N_5432);
nor U9390 (N_9390,N_7329,N_6867);
nor U9391 (N_9391,N_7102,N_5582);
nor U9392 (N_9392,N_5721,N_6649);
xnor U9393 (N_9393,N_7462,N_7416);
nand U9394 (N_9394,N_6497,N_5312);
nor U9395 (N_9395,N_7198,N_5381);
nor U9396 (N_9396,N_6599,N_7181);
nor U9397 (N_9397,N_5706,N_6423);
and U9398 (N_9398,N_6968,N_5661);
nand U9399 (N_9399,N_6017,N_6562);
and U9400 (N_9400,N_6801,N_7389);
nor U9401 (N_9401,N_5299,N_5080);
nor U9402 (N_9402,N_5338,N_5016);
nor U9403 (N_9403,N_5065,N_5419);
xnor U9404 (N_9404,N_7212,N_6476);
xor U9405 (N_9405,N_5057,N_7090);
nor U9406 (N_9406,N_6053,N_5230);
xor U9407 (N_9407,N_6437,N_5134);
or U9408 (N_9408,N_5466,N_5856);
xnor U9409 (N_9409,N_5457,N_5191);
or U9410 (N_9410,N_5230,N_5248);
or U9411 (N_9411,N_7393,N_5324);
nand U9412 (N_9412,N_7138,N_6172);
and U9413 (N_9413,N_7493,N_6389);
xnor U9414 (N_9414,N_5164,N_7200);
or U9415 (N_9415,N_7270,N_6382);
nand U9416 (N_9416,N_7135,N_6548);
or U9417 (N_9417,N_7415,N_6020);
and U9418 (N_9418,N_6387,N_6009);
nand U9419 (N_9419,N_6506,N_7469);
nand U9420 (N_9420,N_7221,N_7471);
nand U9421 (N_9421,N_5272,N_6631);
xor U9422 (N_9422,N_5422,N_7069);
xnor U9423 (N_9423,N_6789,N_5372);
nor U9424 (N_9424,N_5003,N_5323);
and U9425 (N_9425,N_5549,N_6454);
nand U9426 (N_9426,N_6046,N_5151);
nor U9427 (N_9427,N_5616,N_7186);
xor U9428 (N_9428,N_7186,N_5544);
or U9429 (N_9429,N_7089,N_7447);
and U9430 (N_9430,N_7440,N_6655);
or U9431 (N_9431,N_6351,N_7328);
xor U9432 (N_9432,N_6991,N_5485);
or U9433 (N_9433,N_5284,N_5812);
and U9434 (N_9434,N_7121,N_7179);
nor U9435 (N_9435,N_6935,N_6553);
and U9436 (N_9436,N_5309,N_6480);
nand U9437 (N_9437,N_5888,N_6375);
and U9438 (N_9438,N_6457,N_6813);
nor U9439 (N_9439,N_6807,N_6477);
nand U9440 (N_9440,N_7415,N_5381);
or U9441 (N_9441,N_7178,N_6589);
or U9442 (N_9442,N_5060,N_5113);
nand U9443 (N_9443,N_6949,N_7189);
and U9444 (N_9444,N_5211,N_5360);
or U9445 (N_9445,N_5342,N_6600);
and U9446 (N_9446,N_7290,N_6892);
or U9447 (N_9447,N_5517,N_5436);
nor U9448 (N_9448,N_5973,N_6259);
nand U9449 (N_9449,N_5931,N_5484);
xor U9450 (N_9450,N_7217,N_7310);
and U9451 (N_9451,N_7213,N_7065);
or U9452 (N_9452,N_5689,N_7000);
nand U9453 (N_9453,N_6161,N_6010);
and U9454 (N_9454,N_5342,N_5060);
nand U9455 (N_9455,N_6605,N_6832);
xor U9456 (N_9456,N_5201,N_5873);
and U9457 (N_9457,N_7498,N_6296);
nor U9458 (N_9458,N_5164,N_6653);
and U9459 (N_9459,N_7431,N_6933);
nand U9460 (N_9460,N_6073,N_5270);
nor U9461 (N_9461,N_5789,N_5285);
or U9462 (N_9462,N_7344,N_5043);
or U9463 (N_9463,N_7105,N_6132);
xnor U9464 (N_9464,N_7371,N_6091);
xnor U9465 (N_9465,N_7136,N_7003);
and U9466 (N_9466,N_5681,N_7131);
nand U9467 (N_9467,N_6645,N_7493);
nor U9468 (N_9468,N_6684,N_6607);
and U9469 (N_9469,N_5621,N_7429);
xor U9470 (N_9470,N_5630,N_6898);
and U9471 (N_9471,N_5463,N_5967);
xor U9472 (N_9472,N_5769,N_5086);
xnor U9473 (N_9473,N_7196,N_6074);
and U9474 (N_9474,N_6207,N_6853);
nor U9475 (N_9475,N_7320,N_5873);
and U9476 (N_9476,N_6979,N_5364);
nor U9477 (N_9477,N_7282,N_6997);
xnor U9478 (N_9478,N_6828,N_7035);
nor U9479 (N_9479,N_6956,N_6835);
xnor U9480 (N_9480,N_5397,N_5985);
nor U9481 (N_9481,N_5776,N_6452);
nand U9482 (N_9482,N_5461,N_6855);
xor U9483 (N_9483,N_5578,N_5951);
nand U9484 (N_9484,N_6088,N_6008);
or U9485 (N_9485,N_6242,N_7388);
or U9486 (N_9486,N_6012,N_5542);
or U9487 (N_9487,N_5208,N_5051);
and U9488 (N_9488,N_6125,N_5223);
xnor U9489 (N_9489,N_7179,N_7186);
or U9490 (N_9490,N_5088,N_6631);
nand U9491 (N_9491,N_5520,N_6046);
xnor U9492 (N_9492,N_6713,N_5169);
nor U9493 (N_9493,N_7041,N_5028);
nor U9494 (N_9494,N_5684,N_7250);
xnor U9495 (N_9495,N_7344,N_6654);
xnor U9496 (N_9496,N_6397,N_7031);
nor U9497 (N_9497,N_6576,N_5948);
xor U9498 (N_9498,N_6073,N_5218);
or U9499 (N_9499,N_6159,N_5579);
nor U9500 (N_9500,N_6768,N_5923);
nand U9501 (N_9501,N_6257,N_6018);
nor U9502 (N_9502,N_5654,N_7368);
and U9503 (N_9503,N_7450,N_5648);
xor U9504 (N_9504,N_6219,N_6409);
nand U9505 (N_9505,N_5781,N_7494);
nor U9506 (N_9506,N_6466,N_6444);
xnor U9507 (N_9507,N_5271,N_5410);
nand U9508 (N_9508,N_6378,N_5236);
nand U9509 (N_9509,N_6700,N_7189);
xor U9510 (N_9510,N_5970,N_6498);
xnor U9511 (N_9511,N_5069,N_7416);
nand U9512 (N_9512,N_5088,N_5040);
nor U9513 (N_9513,N_5980,N_6914);
and U9514 (N_9514,N_7409,N_6270);
xnor U9515 (N_9515,N_6806,N_6606);
and U9516 (N_9516,N_7260,N_6768);
nor U9517 (N_9517,N_6969,N_5148);
nand U9518 (N_9518,N_7262,N_6728);
xor U9519 (N_9519,N_6362,N_6543);
nand U9520 (N_9520,N_6337,N_7029);
nand U9521 (N_9521,N_5013,N_6950);
or U9522 (N_9522,N_7348,N_5603);
nor U9523 (N_9523,N_6330,N_5022);
and U9524 (N_9524,N_5260,N_6192);
and U9525 (N_9525,N_7157,N_6380);
nor U9526 (N_9526,N_5340,N_5503);
and U9527 (N_9527,N_6545,N_6846);
nor U9528 (N_9528,N_6370,N_5464);
and U9529 (N_9529,N_5740,N_7113);
nand U9530 (N_9530,N_5267,N_5425);
nand U9531 (N_9531,N_5919,N_6176);
xnor U9532 (N_9532,N_5837,N_7359);
and U9533 (N_9533,N_5226,N_5844);
nand U9534 (N_9534,N_6392,N_5486);
nand U9535 (N_9535,N_6250,N_6943);
and U9536 (N_9536,N_5434,N_5491);
or U9537 (N_9537,N_5259,N_6436);
and U9538 (N_9538,N_6368,N_5075);
and U9539 (N_9539,N_5983,N_5560);
nand U9540 (N_9540,N_7094,N_6433);
or U9541 (N_9541,N_6497,N_7460);
and U9542 (N_9542,N_6029,N_5737);
xor U9543 (N_9543,N_5603,N_6873);
nand U9544 (N_9544,N_6579,N_6609);
nand U9545 (N_9545,N_7199,N_6534);
xor U9546 (N_9546,N_6348,N_5535);
and U9547 (N_9547,N_5439,N_6014);
nand U9548 (N_9548,N_7468,N_6756);
and U9549 (N_9549,N_6089,N_5186);
nor U9550 (N_9550,N_6739,N_6160);
and U9551 (N_9551,N_7357,N_5628);
nor U9552 (N_9552,N_6166,N_5359);
and U9553 (N_9553,N_7148,N_5621);
and U9554 (N_9554,N_7271,N_5226);
nand U9555 (N_9555,N_6045,N_7043);
nand U9556 (N_9556,N_7240,N_6313);
xor U9557 (N_9557,N_7020,N_5652);
or U9558 (N_9558,N_6718,N_5446);
nor U9559 (N_9559,N_7247,N_7307);
nor U9560 (N_9560,N_7109,N_6246);
and U9561 (N_9561,N_7243,N_6468);
or U9562 (N_9562,N_7193,N_6749);
xnor U9563 (N_9563,N_5613,N_6372);
and U9564 (N_9564,N_6683,N_6632);
and U9565 (N_9565,N_6312,N_7046);
nand U9566 (N_9566,N_6879,N_7065);
nor U9567 (N_9567,N_5514,N_5032);
nor U9568 (N_9568,N_6666,N_5956);
or U9569 (N_9569,N_6381,N_7083);
and U9570 (N_9570,N_6163,N_5770);
xnor U9571 (N_9571,N_5104,N_5621);
nand U9572 (N_9572,N_5479,N_6415);
and U9573 (N_9573,N_5456,N_6991);
and U9574 (N_9574,N_6180,N_5216);
nor U9575 (N_9575,N_6828,N_6390);
and U9576 (N_9576,N_5783,N_6558);
and U9577 (N_9577,N_7104,N_6801);
and U9578 (N_9578,N_7176,N_6052);
and U9579 (N_9579,N_7169,N_6360);
nand U9580 (N_9580,N_6277,N_6356);
xor U9581 (N_9581,N_6317,N_6027);
nor U9582 (N_9582,N_5921,N_5980);
nand U9583 (N_9583,N_5993,N_5745);
xor U9584 (N_9584,N_5579,N_6331);
or U9585 (N_9585,N_6242,N_5501);
xor U9586 (N_9586,N_7404,N_7176);
nor U9587 (N_9587,N_5572,N_6526);
or U9588 (N_9588,N_7249,N_6021);
nand U9589 (N_9589,N_6814,N_5911);
nor U9590 (N_9590,N_7434,N_5008);
nor U9591 (N_9591,N_5928,N_5862);
nor U9592 (N_9592,N_6797,N_5344);
nor U9593 (N_9593,N_5234,N_5208);
or U9594 (N_9594,N_6109,N_5743);
xnor U9595 (N_9595,N_6176,N_6844);
nand U9596 (N_9596,N_6544,N_5034);
nand U9597 (N_9597,N_6382,N_5164);
nor U9598 (N_9598,N_7113,N_6423);
and U9599 (N_9599,N_7417,N_6465);
and U9600 (N_9600,N_6447,N_6554);
and U9601 (N_9601,N_7071,N_5158);
or U9602 (N_9602,N_6903,N_5371);
xnor U9603 (N_9603,N_6663,N_5031);
nand U9604 (N_9604,N_6057,N_6985);
or U9605 (N_9605,N_6561,N_7288);
nor U9606 (N_9606,N_7001,N_7006);
and U9607 (N_9607,N_6307,N_5780);
or U9608 (N_9608,N_6888,N_5197);
xor U9609 (N_9609,N_6279,N_7009);
or U9610 (N_9610,N_6420,N_5831);
xor U9611 (N_9611,N_6306,N_5238);
xnor U9612 (N_9612,N_6154,N_7488);
and U9613 (N_9613,N_5069,N_5551);
nand U9614 (N_9614,N_5915,N_7069);
nand U9615 (N_9615,N_5631,N_5451);
nand U9616 (N_9616,N_6570,N_6629);
nor U9617 (N_9617,N_5551,N_5228);
nor U9618 (N_9618,N_5088,N_6872);
xnor U9619 (N_9619,N_5462,N_7290);
xnor U9620 (N_9620,N_5821,N_6728);
or U9621 (N_9621,N_6571,N_7098);
and U9622 (N_9622,N_6470,N_5648);
nor U9623 (N_9623,N_7404,N_6256);
nand U9624 (N_9624,N_7413,N_5627);
nor U9625 (N_9625,N_5143,N_6276);
nor U9626 (N_9626,N_5560,N_7384);
and U9627 (N_9627,N_5631,N_5841);
or U9628 (N_9628,N_5283,N_7241);
nand U9629 (N_9629,N_7259,N_6137);
nor U9630 (N_9630,N_6143,N_5216);
and U9631 (N_9631,N_6009,N_6584);
nand U9632 (N_9632,N_6621,N_6189);
nor U9633 (N_9633,N_5867,N_6483);
and U9634 (N_9634,N_6739,N_6481);
and U9635 (N_9635,N_6288,N_5614);
nor U9636 (N_9636,N_5161,N_6973);
and U9637 (N_9637,N_5544,N_5667);
nand U9638 (N_9638,N_6016,N_6388);
nand U9639 (N_9639,N_6968,N_6162);
nor U9640 (N_9640,N_6108,N_5260);
and U9641 (N_9641,N_7164,N_6969);
nor U9642 (N_9642,N_7035,N_6103);
xnor U9643 (N_9643,N_5044,N_6454);
and U9644 (N_9644,N_7327,N_6855);
nor U9645 (N_9645,N_7184,N_5350);
xnor U9646 (N_9646,N_5184,N_6008);
xor U9647 (N_9647,N_5838,N_7128);
and U9648 (N_9648,N_7372,N_6528);
xnor U9649 (N_9649,N_6630,N_6598);
nor U9650 (N_9650,N_5503,N_6580);
and U9651 (N_9651,N_5212,N_7226);
and U9652 (N_9652,N_7316,N_7231);
and U9653 (N_9653,N_6596,N_5350);
and U9654 (N_9654,N_6019,N_5993);
or U9655 (N_9655,N_5706,N_6088);
or U9656 (N_9656,N_7403,N_7404);
and U9657 (N_9657,N_5079,N_6790);
and U9658 (N_9658,N_6541,N_5211);
nand U9659 (N_9659,N_6794,N_7154);
nand U9660 (N_9660,N_5570,N_7123);
nor U9661 (N_9661,N_6103,N_7486);
or U9662 (N_9662,N_7166,N_5126);
and U9663 (N_9663,N_6553,N_5369);
nor U9664 (N_9664,N_6743,N_5692);
nand U9665 (N_9665,N_6355,N_5822);
or U9666 (N_9666,N_5790,N_5350);
xnor U9667 (N_9667,N_6285,N_6099);
nor U9668 (N_9668,N_6719,N_5342);
xnor U9669 (N_9669,N_5317,N_5795);
xnor U9670 (N_9670,N_5920,N_5281);
nor U9671 (N_9671,N_7149,N_5712);
nand U9672 (N_9672,N_7399,N_6655);
nor U9673 (N_9673,N_5234,N_6569);
xnor U9674 (N_9674,N_6470,N_5759);
or U9675 (N_9675,N_6601,N_5972);
and U9676 (N_9676,N_6985,N_5732);
xor U9677 (N_9677,N_7079,N_6904);
and U9678 (N_9678,N_7215,N_5422);
nor U9679 (N_9679,N_7234,N_5051);
nand U9680 (N_9680,N_6243,N_6198);
nor U9681 (N_9681,N_5338,N_7238);
nand U9682 (N_9682,N_7385,N_5869);
or U9683 (N_9683,N_7092,N_6098);
or U9684 (N_9684,N_6298,N_6871);
nand U9685 (N_9685,N_5555,N_5482);
nand U9686 (N_9686,N_6042,N_6590);
xor U9687 (N_9687,N_5062,N_6012);
nor U9688 (N_9688,N_5746,N_5342);
or U9689 (N_9689,N_7403,N_5070);
nand U9690 (N_9690,N_5864,N_7440);
and U9691 (N_9691,N_5413,N_7096);
xor U9692 (N_9692,N_6477,N_6926);
xnor U9693 (N_9693,N_6688,N_5265);
or U9694 (N_9694,N_5132,N_5692);
and U9695 (N_9695,N_6183,N_7050);
or U9696 (N_9696,N_5352,N_5324);
and U9697 (N_9697,N_6453,N_5034);
nand U9698 (N_9698,N_6935,N_6323);
xor U9699 (N_9699,N_6767,N_7287);
or U9700 (N_9700,N_7320,N_7097);
or U9701 (N_9701,N_5146,N_6665);
or U9702 (N_9702,N_5299,N_6781);
xnor U9703 (N_9703,N_5942,N_5160);
nor U9704 (N_9704,N_7393,N_5257);
and U9705 (N_9705,N_6729,N_6258);
xnor U9706 (N_9706,N_7077,N_6600);
xor U9707 (N_9707,N_7314,N_6197);
xor U9708 (N_9708,N_7230,N_7173);
or U9709 (N_9709,N_5955,N_7183);
xor U9710 (N_9710,N_6350,N_7381);
nor U9711 (N_9711,N_5364,N_6937);
nor U9712 (N_9712,N_5600,N_6855);
and U9713 (N_9713,N_5582,N_5112);
nor U9714 (N_9714,N_6989,N_7079);
nand U9715 (N_9715,N_6144,N_7042);
and U9716 (N_9716,N_5173,N_6311);
or U9717 (N_9717,N_5528,N_6462);
nand U9718 (N_9718,N_5447,N_5455);
xnor U9719 (N_9719,N_6180,N_5636);
or U9720 (N_9720,N_7202,N_7379);
nand U9721 (N_9721,N_6054,N_6189);
or U9722 (N_9722,N_5163,N_7491);
or U9723 (N_9723,N_5706,N_5134);
and U9724 (N_9724,N_5879,N_6575);
xnor U9725 (N_9725,N_5979,N_6590);
nand U9726 (N_9726,N_6988,N_6671);
or U9727 (N_9727,N_5449,N_5779);
and U9728 (N_9728,N_5895,N_5647);
nor U9729 (N_9729,N_7133,N_5592);
nand U9730 (N_9730,N_5458,N_7081);
and U9731 (N_9731,N_5652,N_6404);
and U9732 (N_9732,N_5012,N_5110);
or U9733 (N_9733,N_6287,N_5877);
nor U9734 (N_9734,N_6312,N_6369);
nor U9735 (N_9735,N_5245,N_6961);
xor U9736 (N_9736,N_5283,N_5946);
nor U9737 (N_9737,N_5674,N_6095);
or U9738 (N_9738,N_5423,N_5652);
nor U9739 (N_9739,N_7135,N_7431);
xnor U9740 (N_9740,N_5451,N_5056);
or U9741 (N_9741,N_5407,N_5977);
xor U9742 (N_9742,N_5506,N_6949);
or U9743 (N_9743,N_7335,N_7172);
nor U9744 (N_9744,N_5491,N_6621);
or U9745 (N_9745,N_7292,N_5786);
or U9746 (N_9746,N_5245,N_6558);
nand U9747 (N_9747,N_6752,N_7462);
nor U9748 (N_9748,N_5448,N_7089);
nand U9749 (N_9749,N_6623,N_6833);
nand U9750 (N_9750,N_5806,N_7317);
xnor U9751 (N_9751,N_5055,N_5128);
or U9752 (N_9752,N_5190,N_7045);
nand U9753 (N_9753,N_5803,N_7224);
nor U9754 (N_9754,N_5125,N_7280);
or U9755 (N_9755,N_5775,N_7160);
nor U9756 (N_9756,N_6283,N_5870);
nand U9757 (N_9757,N_6408,N_6296);
xor U9758 (N_9758,N_7356,N_6988);
xor U9759 (N_9759,N_6525,N_6480);
nand U9760 (N_9760,N_5794,N_5952);
or U9761 (N_9761,N_6009,N_6361);
or U9762 (N_9762,N_5084,N_6123);
xnor U9763 (N_9763,N_5831,N_5427);
xnor U9764 (N_9764,N_5849,N_5605);
and U9765 (N_9765,N_6669,N_6655);
xor U9766 (N_9766,N_7346,N_6849);
nand U9767 (N_9767,N_5753,N_6709);
or U9768 (N_9768,N_6722,N_7132);
nand U9769 (N_9769,N_7338,N_5693);
xor U9770 (N_9770,N_7047,N_6270);
and U9771 (N_9771,N_7161,N_5215);
nand U9772 (N_9772,N_5303,N_7254);
or U9773 (N_9773,N_5852,N_6078);
or U9774 (N_9774,N_5152,N_6382);
nor U9775 (N_9775,N_6691,N_5084);
nor U9776 (N_9776,N_6836,N_5383);
xnor U9777 (N_9777,N_5959,N_7359);
nor U9778 (N_9778,N_6705,N_5859);
and U9779 (N_9779,N_5155,N_6460);
xor U9780 (N_9780,N_6534,N_5973);
nor U9781 (N_9781,N_5618,N_5182);
nand U9782 (N_9782,N_5591,N_5605);
nor U9783 (N_9783,N_6102,N_7434);
nand U9784 (N_9784,N_6073,N_5351);
nand U9785 (N_9785,N_6976,N_5296);
or U9786 (N_9786,N_6507,N_6886);
or U9787 (N_9787,N_6148,N_6863);
nand U9788 (N_9788,N_5701,N_6975);
and U9789 (N_9789,N_5932,N_7356);
and U9790 (N_9790,N_6697,N_7402);
xnor U9791 (N_9791,N_5825,N_6875);
or U9792 (N_9792,N_7431,N_7028);
or U9793 (N_9793,N_7260,N_5861);
or U9794 (N_9794,N_6958,N_6844);
and U9795 (N_9795,N_6630,N_6799);
xnor U9796 (N_9796,N_7017,N_5827);
xnor U9797 (N_9797,N_6296,N_5049);
and U9798 (N_9798,N_7175,N_6053);
xnor U9799 (N_9799,N_5050,N_6589);
xor U9800 (N_9800,N_6488,N_5014);
nor U9801 (N_9801,N_7393,N_6782);
nor U9802 (N_9802,N_5868,N_5250);
or U9803 (N_9803,N_5653,N_6421);
and U9804 (N_9804,N_5358,N_5603);
and U9805 (N_9805,N_7408,N_6567);
nor U9806 (N_9806,N_7176,N_5876);
nor U9807 (N_9807,N_6564,N_6643);
xnor U9808 (N_9808,N_6964,N_5149);
nand U9809 (N_9809,N_5606,N_5705);
nor U9810 (N_9810,N_7295,N_7499);
nand U9811 (N_9811,N_5634,N_6292);
xor U9812 (N_9812,N_6754,N_5994);
nor U9813 (N_9813,N_7317,N_6649);
nor U9814 (N_9814,N_5279,N_6530);
or U9815 (N_9815,N_6439,N_6661);
nor U9816 (N_9816,N_6223,N_5562);
or U9817 (N_9817,N_5677,N_6506);
nand U9818 (N_9818,N_5578,N_6677);
nor U9819 (N_9819,N_6057,N_5792);
nor U9820 (N_9820,N_6631,N_6909);
nor U9821 (N_9821,N_7075,N_5265);
nor U9822 (N_9822,N_5430,N_5508);
nor U9823 (N_9823,N_6820,N_5698);
nor U9824 (N_9824,N_5493,N_6321);
nor U9825 (N_9825,N_5590,N_6545);
or U9826 (N_9826,N_6326,N_7265);
nand U9827 (N_9827,N_6119,N_6555);
nand U9828 (N_9828,N_6511,N_7136);
and U9829 (N_9829,N_6097,N_5668);
nor U9830 (N_9830,N_6136,N_5913);
nand U9831 (N_9831,N_6146,N_5256);
and U9832 (N_9832,N_5477,N_5957);
nor U9833 (N_9833,N_6294,N_6094);
xor U9834 (N_9834,N_6118,N_5486);
and U9835 (N_9835,N_6979,N_6351);
nor U9836 (N_9836,N_6201,N_6906);
xnor U9837 (N_9837,N_5932,N_5596);
xor U9838 (N_9838,N_6844,N_6351);
and U9839 (N_9839,N_5717,N_6983);
and U9840 (N_9840,N_6544,N_7475);
and U9841 (N_9841,N_5160,N_6818);
xnor U9842 (N_9842,N_7017,N_5495);
nor U9843 (N_9843,N_5675,N_6396);
nor U9844 (N_9844,N_5927,N_6198);
xor U9845 (N_9845,N_7157,N_6372);
or U9846 (N_9846,N_5059,N_6014);
xor U9847 (N_9847,N_6318,N_6350);
and U9848 (N_9848,N_6018,N_5459);
and U9849 (N_9849,N_6756,N_5374);
and U9850 (N_9850,N_7216,N_5076);
nor U9851 (N_9851,N_5595,N_5774);
nand U9852 (N_9852,N_5340,N_5381);
or U9853 (N_9853,N_6842,N_7179);
nand U9854 (N_9854,N_5161,N_6970);
xor U9855 (N_9855,N_6136,N_6717);
nand U9856 (N_9856,N_7330,N_5300);
or U9857 (N_9857,N_6656,N_5392);
nand U9858 (N_9858,N_6211,N_5862);
or U9859 (N_9859,N_5142,N_5562);
nand U9860 (N_9860,N_6419,N_5048);
xnor U9861 (N_9861,N_7189,N_5816);
or U9862 (N_9862,N_6300,N_5985);
nor U9863 (N_9863,N_6854,N_5045);
xnor U9864 (N_9864,N_5637,N_5282);
or U9865 (N_9865,N_5558,N_7056);
and U9866 (N_9866,N_6152,N_5358);
nand U9867 (N_9867,N_5519,N_7474);
and U9868 (N_9868,N_6693,N_6799);
xor U9869 (N_9869,N_5316,N_7379);
nand U9870 (N_9870,N_6731,N_7124);
or U9871 (N_9871,N_6826,N_6381);
or U9872 (N_9872,N_5141,N_5607);
and U9873 (N_9873,N_6653,N_6137);
xnor U9874 (N_9874,N_6070,N_7402);
nor U9875 (N_9875,N_5899,N_5253);
and U9876 (N_9876,N_6158,N_6547);
nor U9877 (N_9877,N_5152,N_6249);
xnor U9878 (N_9878,N_6995,N_7206);
nor U9879 (N_9879,N_6387,N_6858);
xor U9880 (N_9880,N_6978,N_6256);
nand U9881 (N_9881,N_6989,N_6384);
and U9882 (N_9882,N_6376,N_5538);
nand U9883 (N_9883,N_6484,N_6929);
nand U9884 (N_9884,N_6940,N_5847);
and U9885 (N_9885,N_6342,N_6651);
nor U9886 (N_9886,N_7016,N_6502);
or U9887 (N_9887,N_5710,N_6713);
or U9888 (N_9888,N_6680,N_5104);
nand U9889 (N_9889,N_7041,N_5248);
nor U9890 (N_9890,N_7049,N_6694);
or U9891 (N_9891,N_5447,N_6946);
or U9892 (N_9892,N_5314,N_6394);
xnor U9893 (N_9893,N_5131,N_5809);
nand U9894 (N_9894,N_5217,N_6658);
and U9895 (N_9895,N_6691,N_6305);
xnor U9896 (N_9896,N_6730,N_7314);
and U9897 (N_9897,N_6776,N_6607);
xnor U9898 (N_9898,N_6025,N_5496);
xnor U9899 (N_9899,N_6062,N_7004);
or U9900 (N_9900,N_6090,N_5561);
xor U9901 (N_9901,N_7189,N_7154);
and U9902 (N_9902,N_6039,N_5583);
nand U9903 (N_9903,N_6827,N_7396);
xnor U9904 (N_9904,N_6645,N_6692);
and U9905 (N_9905,N_5556,N_6068);
nand U9906 (N_9906,N_5791,N_6394);
nor U9907 (N_9907,N_6200,N_6378);
and U9908 (N_9908,N_7085,N_7142);
nand U9909 (N_9909,N_7325,N_6895);
nand U9910 (N_9910,N_5163,N_5821);
nor U9911 (N_9911,N_6376,N_5639);
nor U9912 (N_9912,N_5302,N_5178);
nor U9913 (N_9913,N_6877,N_5370);
nor U9914 (N_9914,N_6558,N_7244);
and U9915 (N_9915,N_7384,N_6868);
or U9916 (N_9916,N_5130,N_5437);
and U9917 (N_9917,N_6527,N_6116);
or U9918 (N_9918,N_7138,N_6022);
nor U9919 (N_9919,N_5822,N_6897);
nand U9920 (N_9920,N_7360,N_7404);
nand U9921 (N_9921,N_6856,N_5573);
nand U9922 (N_9922,N_6343,N_5532);
or U9923 (N_9923,N_6042,N_5301);
and U9924 (N_9924,N_7151,N_5186);
or U9925 (N_9925,N_7030,N_5239);
nand U9926 (N_9926,N_6265,N_7223);
nor U9927 (N_9927,N_6067,N_6109);
xor U9928 (N_9928,N_7209,N_7132);
xor U9929 (N_9929,N_7333,N_6801);
nand U9930 (N_9930,N_7449,N_6465);
nor U9931 (N_9931,N_5359,N_5653);
nand U9932 (N_9932,N_6673,N_6637);
xor U9933 (N_9933,N_7048,N_5190);
nor U9934 (N_9934,N_5283,N_5247);
or U9935 (N_9935,N_5739,N_7302);
or U9936 (N_9936,N_6096,N_6561);
xor U9937 (N_9937,N_6535,N_5472);
xnor U9938 (N_9938,N_5832,N_6414);
nor U9939 (N_9939,N_5787,N_5518);
nand U9940 (N_9940,N_6798,N_5868);
nor U9941 (N_9941,N_5931,N_5262);
nor U9942 (N_9942,N_5667,N_7211);
xor U9943 (N_9943,N_5644,N_5202);
xnor U9944 (N_9944,N_6486,N_6394);
and U9945 (N_9945,N_6613,N_6476);
or U9946 (N_9946,N_7488,N_5501);
or U9947 (N_9947,N_6916,N_6319);
nor U9948 (N_9948,N_7139,N_5725);
nor U9949 (N_9949,N_5562,N_6773);
and U9950 (N_9950,N_6396,N_6987);
nor U9951 (N_9951,N_7426,N_5003);
and U9952 (N_9952,N_6777,N_6315);
xor U9953 (N_9953,N_5915,N_6540);
or U9954 (N_9954,N_7416,N_7170);
xor U9955 (N_9955,N_5863,N_6917);
and U9956 (N_9956,N_7145,N_5487);
or U9957 (N_9957,N_7204,N_7102);
or U9958 (N_9958,N_7309,N_5422);
xnor U9959 (N_9959,N_5483,N_6512);
nor U9960 (N_9960,N_6128,N_6370);
or U9961 (N_9961,N_6819,N_6882);
or U9962 (N_9962,N_6997,N_7039);
and U9963 (N_9963,N_5944,N_5047);
xor U9964 (N_9964,N_6002,N_5479);
xor U9965 (N_9965,N_6275,N_7121);
nor U9966 (N_9966,N_6243,N_6241);
nand U9967 (N_9967,N_5010,N_5385);
xnor U9968 (N_9968,N_5607,N_6228);
and U9969 (N_9969,N_6740,N_6389);
nand U9970 (N_9970,N_6170,N_6503);
nor U9971 (N_9971,N_5429,N_5964);
or U9972 (N_9972,N_7367,N_7216);
nand U9973 (N_9973,N_6854,N_6763);
and U9974 (N_9974,N_6591,N_5358);
and U9975 (N_9975,N_5656,N_6279);
nand U9976 (N_9976,N_6437,N_5769);
and U9977 (N_9977,N_7058,N_6253);
xnor U9978 (N_9978,N_5612,N_5836);
and U9979 (N_9979,N_6330,N_5030);
nor U9980 (N_9980,N_5896,N_5359);
xor U9981 (N_9981,N_7403,N_7033);
or U9982 (N_9982,N_6381,N_5749);
xor U9983 (N_9983,N_7091,N_6817);
and U9984 (N_9984,N_7349,N_7277);
and U9985 (N_9985,N_5272,N_5740);
or U9986 (N_9986,N_6112,N_7289);
xor U9987 (N_9987,N_6573,N_5000);
or U9988 (N_9988,N_5548,N_5406);
or U9989 (N_9989,N_7383,N_5583);
and U9990 (N_9990,N_5221,N_5754);
or U9991 (N_9991,N_7456,N_6364);
nand U9992 (N_9992,N_5716,N_5105);
nor U9993 (N_9993,N_5786,N_6764);
nor U9994 (N_9994,N_6453,N_7460);
nor U9995 (N_9995,N_6559,N_7102);
and U9996 (N_9996,N_6842,N_7125);
and U9997 (N_9997,N_6310,N_5133);
or U9998 (N_9998,N_7264,N_5307);
nor U9999 (N_9999,N_6028,N_6837);
or UO_0 (O_0,N_9091,N_9138);
nor UO_1 (O_1,N_8000,N_8419);
or UO_2 (O_2,N_8022,N_9576);
xor UO_3 (O_3,N_7630,N_7831);
xor UO_4 (O_4,N_9467,N_8748);
and UO_5 (O_5,N_9646,N_7930);
nand UO_6 (O_6,N_9602,N_9167);
or UO_7 (O_7,N_8595,N_7523);
or UO_8 (O_8,N_9842,N_9964);
or UO_9 (O_9,N_9392,N_8439);
xor UO_10 (O_10,N_8798,N_9781);
nand UO_11 (O_11,N_9269,N_9724);
or UO_12 (O_12,N_7669,N_9375);
and UO_13 (O_13,N_8460,N_9861);
or UO_14 (O_14,N_9722,N_9175);
or UO_15 (O_15,N_8017,N_9839);
xor UO_16 (O_16,N_9761,N_8373);
or UO_17 (O_17,N_9624,N_7927);
xor UO_18 (O_18,N_9548,N_7609);
xnor UO_19 (O_19,N_8675,N_8942);
and UO_20 (O_20,N_8971,N_7598);
nand UO_21 (O_21,N_8176,N_9235);
xnor UO_22 (O_22,N_8926,N_9323);
and UO_23 (O_23,N_8768,N_8403);
xnor UO_24 (O_24,N_8384,N_8078);
xor UO_25 (O_25,N_9706,N_9018);
xnor UO_26 (O_26,N_7740,N_9391);
xor UO_27 (O_27,N_8536,N_7791);
nand UO_28 (O_28,N_8506,N_8507);
and UO_29 (O_29,N_8808,N_9741);
nor UO_30 (O_30,N_8092,N_8538);
and UO_31 (O_31,N_8446,N_9593);
and UO_32 (O_32,N_9912,N_9633);
and UO_33 (O_33,N_7522,N_9401);
or UO_34 (O_34,N_9952,N_7922);
nand UO_35 (O_35,N_9896,N_8090);
or UO_36 (O_36,N_8686,N_9219);
nor UO_37 (O_37,N_9238,N_8004);
xor UO_38 (O_38,N_8716,N_9798);
and UO_39 (O_39,N_9419,N_9082);
nor UO_40 (O_40,N_9844,N_9209);
and UO_41 (O_41,N_8993,N_9677);
and UO_42 (O_42,N_8572,N_8640);
or UO_43 (O_43,N_7730,N_8714);
or UO_44 (O_44,N_7769,N_7583);
and UO_45 (O_45,N_7586,N_8668);
or UO_46 (O_46,N_9133,N_9674);
or UO_47 (O_47,N_8645,N_8327);
xor UO_48 (O_48,N_8038,N_8979);
nand UO_49 (O_49,N_9108,N_9926);
nor UO_50 (O_50,N_9951,N_7815);
nor UO_51 (O_51,N_9411,N_8249);
nor UO_52 (O_52,N_7987,N_9754);
and UO_53 (O_53,N_9123,N_9112);
nor UO_54 (O_54,N_7883,N_9752);
and UO_55 (O_55,N_7649,N_9849);
and UO_56 (O_56,N_9594,N_8328);
nor UO_57 (O_57,N_8331,N_8435);
nor UO_58 (O_58,N_8309,N_8360);
nand UO_59 (O_59,N_9639,N_9815);
nor UO_60 (O_60,N_7868,N_8649);
or UO_61 (O_61,N_8034,N_9814);
xnor UO_62 (O_62,N_9196,N_7718);
nand UO_63 (O_63,N_9749,N_9380);
xnor UO_64 (O_64,N_7876,N_9879);
and UO_65 (O_65,N_9887,N_8262);
or UO_66 (O_66,N_9784,N_8486);
nand UO_67 (O_67,N_9239,N_8470);
and UO_68 (O_68,N_9397,N_9592);
xnor UO_69 (O_69,N_8573,N_9363);
xnor UO_70 (O_70,N_7549,N_8286);
or UO_71 (O_71,N_9284,N_7925);
nand UO_72 (O_72,N_8531,N_8459);
nor UO_73 (O_73,N_9880,N_9991);
nor UO_74 (O_74,N_9644,N_8651);
xnor UO_75 (O_75,N_8201,N_7741);
nor UO_76 (O_76,N_7541,N_8671);
nand UO_77 (O_77,N_9647,N_8024);
and UO_78 (O_78,N_8634,N_8530);
nor UO_79 (O_79,N_8518,N_8962);
nand UO_80 (O_80,N_9285,N_9210);
or UO_81 (O_81,N_8529,N_8233);
and UO_82 (O_82,N_9379,N_9514);
and UO_83 (O_83,N_9151,N_9162);
or UO_84 (O_84,N_9486,N_7879);
and UO_85 (O_85,N_8280,N_8468);
nor UO_86 (O_86,N_8397,N_7921);
or UO_87 (O_87,N_9746,N_8582);
nor UO_88 (O_88,N_9377,N_9782);
or UO_89 (O_89,N_9867,N_8293);
xnor UO_90 (O_90,N_7793,N_8289);
and UO_91 (O_91,N_8484,N_9110);
and UO_92 (O_92,N_9766,N_7811);
nand UO_93 (O_93,N_8626,N_9417);
xnor UO_94 (O_94,N_9308,N_7813);
nor UO_95 (O_95,N_9945,N_7555);
xnor UO_96 (O_96,N_8145,N_9111);
xnor UO_97 (O_97,N_9290,N_8516);
xnor UO_98 (O_98,N_7908,N_9141);
xnor UO_99 (O_99,N_8801,N_9885);
nand UO_100 (O_100,N_8298,N_9231);
or UO_101 (O_101,N_9818,N_7909);
nand UO_102 (O_102,N_8777,N_8455);
or UO_103 (O_103,N_9017,N_7988);
xnor UO_104 (O_104,N_8086,N_9805);
or UO_105 (O_105,N_8246,N_9172);
nor UO_106 (O_106,N_8786,N_7819);
or UO_107 (O_107,N_8259,N_8705);
and UO_108 (O_108,N_7881,N_9549);
nor UO_109 (O_109,N_9052,N_9266);
or UO_110 (O_110,N_8830,N_9399);
and UO_111 (O_111,N_9464,N_8909);
xor UO_112 (O_112,N_8782,N_8731);
or UO_113 (O_113,N_8810,N_9989);
xor UO_114 (O_114,N_9581,N_9526);
nor UO_115 (O_115,N_8179,N_9618);
and UO_116 (O_116,N_8108,N_9902);
and UO_117 (O_117,N_7980,N_7842);
or UO_118 (O_118,N_9140,N_9037);
and UO_119 (O_119,N_8365,N_8407);
xnor UO_120 (O_120,N_9946,N_8134);
nand UO_121 (O_121,N_9097,N_9718);
and UO_122 (O_122,N_9029,N_9640);
nor UO_123 (O_123,N_7857,N_8995);
nand UO_124 (O_124,N_8733,N_8010);
xor UO_125 (O_125,N_7771,N_8127);
xnor UO_126 (O_126,N_9543,N_9685);
and UO_127 (O_127,N_8140,N_9364);
nor UO_128 (O_128,N_9918,N_8305);
nor UO_129 (O_129,N_8522,N_7898);
nand UO_130 (O_130,N_9919,N_7888);
xnor UO_131 (O_131,N_9039,N_9160);
and UO_132 (O_132,N_9744,N_8014);
nor UO_133 (O_133,N_7914,N_7851);
xor UO_134 (O_134,N_7652,N_9700);
nor UO_135 (O_135,N_9811,N_8823);
or UO_136 (O_136,N_9872,N_9499);
xnor UO_137 (O_137,N_7850,N_8137);
and UO_138 (O_138,N_8725,N_8167);
xnor UO_139 (O_139,N_9109,N_9770);
nand UO_140 (O_140,N_9928,N_9400);
nor UO_141 (O_141,N_8214,N_8866);
nand UO_142 (O_142,N_8272,N_7854);
and UO_143 (O_143,N_7701,N_8363);
xor UO_144 (O_144,N_9121,N_7786);
and UO_145 (O_145,N_7915,N_9947);
or UO_146 (O_146,N_8553,N_8292);
xnor UO_147 (O_147,N_8059,N_8586);
and UO_148 (O_148,N_7845,N_8661);
and UO_149 (O_149,N_7720,N_9985);
and UO_150 (O_150,N_8527,N_8098);
nand UO_151 (O_151,N_8647,N_9404);
nor UO_152 (O_152,N_9041,N_9775);
and UO_153 (O_153,N_8805,N_9698);
nor UO_154 (O_154,N_7633,N_9652);
or UO_155 (O_155,N_9228,N_7818);
or UO_156 (O_156,N_8421,N_8213);
nand UO_157 (O_157,N_9451,N_9779);
and UO_158 (O_158,N_9636,N_7911);
and UO_159 (O_159,N_9575,N_8975);
nand UO_160 (O_160,N_9130,N_7852);
nor UO_161 (O_161,N_8018,N_9398);
xor UO_162 (O_162,N_7521,N_9243);
nand UO_163 (O_163,N_8597,N_9932);
nor UO_164 (O_164,N_9855,N_7995);
nand UO_165 (O_165,N_7654,N_9957);
or UO_166 (O_166,N_9200,N_8961);
and UO_167 (O_167,N_9475,N_8390);
nor UO_168 (O_168,N_8035,N_9071);
xnor UO_169 (O_169,N_8245,N_9673);
and UO_170 (O_170,N_9521,N_8237);
xor UO_171 (O_171,N_8229,N_8225);
and UO_172 (O_172,N_8555,N_9054);
and UO_173 (O_173,N_8771,N_9281);
and UO_174 (O_174,N_7723,N_8515);
nor UO_175 (O_175,N_7961,N_8741);
xnor UO_176 (O_176,N_9739,N_8875);
nor UO_177 (O_177,N_7899,N_8936);
nor UO_178 (O_178,N_9743,N_8520);
nand UO_179 (O_179,N_8410,N_7903);
nor UO_180 (O_180,N_9664,N_8291);
xor UO_181 (O_181,N_8182,N_8713);
nand UO_182 (O_182,N_9653,N_9613);
nand UO_183 (O_183,N_9783,N_7639);
xnor UO_184 (O_184,N_9019,N_8477);
xor UO_185 (O_185,N_8006,N_8711);
xnor UO_186 (O_186,N_9073,N_7958);
xor UO_187 (O_187,N_8665,N_8130);
xnor UO_188 (O_188,N_9596,N_8575);
nand UO_189 (O_189,N_8488,N_8211);
or UO_190 (O_190,N_7690,N_9878);
nand UO_191 (O_191,N_7802,N_9667);
nor UO_192 (O_192,N_8697,N_7862);
nor UO_193 (O_193,N_9709,N_7974);
and UO_194 (O_194,N_9503,N_7564);
xnor UO_195 (O_195,N_8541,N_8223);
and UO_196 (O_196,N_8769,N_9390);
nor UO_197 (O_197,N_7890,N_9552);
nor UO_198 (O_198,N_9634,N_8613);
nor UO_199 (O_199,N_9505,N_7918);
or UO_200 (O_200,N_7686,N_9291);
or UO_201 (O_201,N_7936,N_8738);
nor UO_202 (O_202,N_8903,N_9627);
nand UO_203 (O_203,N_8348,N_9736);
and UO_204 (O_204,N_9453,N_8336);
or UO_205 (O_205,N_9977,N_8157);
nand UO_206 (O_206,N_9448,N_8907);
nand UO_207 (O_207,N_9190,N_8386);
xnor UO_208 (O_208,N_8894,N_8030);
and UO_209 (O_209,N_9871,N_8948);
or UO_210 (O_210,N_7810,N_8217);
nor UO_211 (O_211,N_9745,N_7948);
nand UO_212 (O_212,N_7924,N_9980);
nand UO_213 (O_213,N_8955,N_8324);
or UO_214 (O_214,N_7542,N_8248);
nor UO_215 (O_215,N_9892,N_9309);
and UO_216 (O_216,N_8800,N_8196);
and UO_217 (O_217,N_8587,N_9742);
nand UO_218 (O_218,N_8204,N_9333);
nor UO_219 (O_219,N_9599,N_7685);
xnor UO_220 (O_220,N_8062,N_9642);
xor UO_221 (O_221,N_8822,N_9445);
and UO_222 (O_222,N_7975,N_7833);
or UO_223 (O_223,N_8193,N_8126);
and UO_224 (O_224,N_9043,N_8170);
nor UO_225 (O_225,N_9758,N_8474);
nand UO_226 (O_226,N_7806,N_9950);
xnor UO_227 (O_227,N_8036,N_8791);
nor UO_228 (O_228,N_9960,N_8736);
or UO_229 (O_229,N_8231,N_8749);
nor UO_230 (O_230,N_8897,N_9354);
xor UO_231 (O_231,N_8700,N_7792);
or UO_232 (O_232,N_8760,N_7646);
xor UO_233 (O_233,N_9296,N_8911);
and UO_234 (O_234,N_8774,N_7999);
nor UO_235 (O_235,N_7984,N_8026);
nor UO_236 (O_236,N_8954,N_8815);
or UO_237 (O_237,N_9697,N_8547);
and UO_238 (O_238,N_9971,N_8499);
and UO_239 (O_239,N_7976,N_9788);
nor UO_240 (O_240,N_9315,N_8556);
nor UO_241 (O_241,N_9293,N_9619);
or UO_242 (O_242,N_7543,N_9355);
or UO_243 (O_243,N_9776,N_8202);
or UO_244 (O_244,N_9579,N_8118);
nand UO_245 (O_245,N_8462,N_8133);
or UO_246 (O_246,N_9649,N_9428);
and UO_247 (O_247,N_7869,N_9298);
nand UO_248 (O_248,N_9403,N_7629);
and UO_249 (O_249,N_8187,N_8471);
or UO_250 (O_250,N_8780,N_8652);
xor UO_251 (O_251,N_7981,N_9626);
and UO_252 (O_252,N_9997,N_7785);
and UO_253 (O_253,N_9164,N_9310);
and UO_254 (O_254,N_8779,N_7788);
nand UO_255 (O_255,N_9488,N_8047);
xnor UO_256 (O_256,N_9894,N_8696);
or UO_257 (O_257,N_8161,N_9873);
xnor UO_258 (O_258,N_7547,N_7755);
xor UO_259 (O_259,N_8189,N_8584);
or UO_260 (O_260,N_7680,N_9895);
nand UO_261 (O_261,N_8021,N_9276);
or UO_262 (O_262,N_9192,N_8230);
nand UO_263 (O_263,N_8091,N_9180);
xor UO_264 (O_264,N_8242,N_7559);
or UO_265 (O_265,N_8638,N_8637);
nand UO_266 (O_266,N_7506,N_9802);
xnor UO_267 (O_267,N_9711,N_7526);
or UO_268 (O_268,N_7977,N_7711);
nand UO_269 (O_269,N_9103,N_8497);
nor UO_270 (O_270,N_8226,N_9611);
nor UO_271 (O_271,N_8087,N_8743);
nor UO_272 (O_272,N_8253,N_9324);
nor UO_273 (O_273,N_8496,N_8073);
xor UO_274 (O_274,N_8267,N_9936);
nor UO_275 (O_275,N_8860,N_7913);
or UO_276 (O_276,N_7971,N_9676);
xor UO_277 (O_277,N_8260,N_8889);
or UO_278 (O_278,N_9049,N_8591);
nand UO_279 (O_279,N_8312,N_7839);
nand UO_280 (O_280,N_8630,N_8349);
or UO_281 (O_281,N_8687,N_8337);
xor UO_282 (O_282,N_8500,N_8831);
nand UO_283 (O_283,N_8680,N_7929);
nand UO_284 (O_284,N_9513,N_7619);
and UO_285 (O_285,N_9424,N_7699);
nor UO_286 (O_286,N_9906,N_9455);
nor UO_287 (O_287,N_9412,N_9929);
or UO_288 (O_288,N_7878,N_8052);
and UO_289 (O_289,N_8055,N_8632);
nor UO_290 (O_290,N_8041,N_8306);
or UO_291 (O_291,N_8027,N_9641);
xnor UO_292 (O_292,N_9565,N_8834);
nor UO_293 (O_293,N_9074,N_9778);
and UO_294 (O_294,N_9125,N_9440);
or UO_295 (O_295,N_8788,N_9129);
or UO_296 (O_296,N_9940,N_8071);
and UO_297 (O_297,N_9365,N_7837);
xnor UO_298 (O_298,N_9139,N_9657);
or UO_299 (O_299,N_9574,N_9114);
and UO_300 (O_300,N_9004,N_9833);
or UO_301 (O_301,N_7614,N_8915);
or UO_302 (O_302,N_9427,N_8552);
or UO_303 (O_303,N_7779,N_7530);
nand UO_304 (O_304,N_8356,N_9289);
nand UO_305 (O_305,N_9396,N_9635);
or UO_306 (O_306,N_8431,N_8031);
or UO_307 (O_307,N_9679,N_7902);
xor UO_308 (O_308,N_8729,N_8846);
nor UO_309 (O_309,N_8882,N_8315);
or UO_310 (O_310,N_8409,N_8984);
nand UO_311 (O_311,N_8667,N_9036);
and UO_312 (O_312,N_9590,N_9601);
or UO_313 (O_313,N_9368,N_8358);
xor UO_314 (O_314,N_9346,N_8722);
and UO_315 (O_315,N_8674,N_9208);
xor UO_316 (O_316,N_7638,N_9322);
and UO_317 (O_317,N_8762,N_9142);
nor UO_318 (O_318,N_9482,N_7570);
nor UO_319 (O_319,N_8561,N_9406);
xor UO_320 (O_320,N_9913,N_9925);
or UO_321 (O_321,N_8141,N_8482);
nor UO_322 (O_322,N_8678,N_8119);
nor UO_323 (O_323,N_7518,N_8143);
xnor UO_324 (O_324,N_9714,N_8601);
and UO_325 (O_325,N_9267,N_9155);
xnor UO_326 (O_326,N_9517,N_8585);
nor UO_327 (O_327,N_9810,N_7861);
or UO_328 (O_328,N_7863,N_7765);
and UO_329 (O_329,N_9215,N_7693);
and UO_330 (O_330,N_8156,N_8311);
and UO_331 (O_331,N_9948,N_8967);
xnor UO_332 (O_332,N_9113,N_7551);
nor UO_333 (O_333,N_8072,N_7858);
xor UO_334 (O_334,N_9645,N_7799);
or UO_335 (O_335,N_8812,N_8296);
nand UO_336 (O_336,N_7737,N_9185);
and UO_337 (O_337,N_8717,N_9003);
xnor UO_338 (O_338,N_8162,N_9351);
and UO_339 (O_339,N_8827,N_8691);
xor UO_340 (O_340,N_9825,N_9812);
nor UO_341 (O_341,N_9477,N_8599);
xor UO_342 (O_342,N_9566,N_7529);
nand UO_343 (O_343,N_9546,N_7886);
and UO_344 (O_344,N_8326,N_9528);
nor UO_345 (O_345,N_7893,N_9212);
xor UO_346 (O_346,N_9569,N_8746);
nor UO_347 (O_347,N_7956,N_7885);
nor UO_348 (O_348,N_9863,N_9450);
or UO_349 (O_349,N_8060,N_8183);
or UO_350 (O_350,N_9921,N_8930);
xnor UO_351 (O_351,N_7590,N_8533);
nor UO_352 (O_352,N_8617,N_9661);
and UO_353 (O_353,N_8347,N_9369);
or UO_354 (O_354,N_8151,N_9437);
nor UO_355 (O_355,N_7954,N_7783);
xor UO_356 (O_356,N_9485,N_9413);
xnor UO_357 (O_357,N_8646,N_9699);
and UO_358 (O_358,N_9001,N_7678);
or UO_359 (O_359,N_7795,N_8111);
nand UO_360 (O_360,N_9502,N_8783);
and UO_361 (O_361,N_8608,N_8982);
nand UO_362 (O_362,N_7662,N_9944);
xor UO_363 (O_363,N_9556,N_8512);
nand UO_364 (O_364,N_7772,N_7834);
and UO_365 (O_365,N_8235,N_8672);
or UO_366 (O_366,N_8745,N_9146);
or UO_367 (O_367,N_8913,N_9067);
nand UO_368 (O_368,N_8372,N_8841);
nor UO_369 (O_369,N_8952,N_8195);
xnor UO_370 (O_370,N_7955,N_8949);
or UO_371 (O_371,N_7683,N_7964);
and UO_372 (O_372,N_7606,N_7968);
or UO_373 (O_373,N_9834,N_9553);
and UO_374 (O_374,N_8432,N_8519);
and UO_375 (O_375,N_7658,N_8469);
xnor UO_376 (O_376,N_8557,N_8723);
xnor UO_377 (O_377,N_7928,N_8602);
nor UO_378 (O_378,N_9735,N_9609);
nor UO_379 (O_379,N_8220,N_8040);
nand UO_380 (O_380,N_9804,N_9727);
and UO_381 (O_381,N_7768,N_7571);
xor UO_382 (O_382,N_8106,N_7962);
and UO_383 (O_383,N_8956,N_9102);
or UO_384 (O_384,N_9432,N_9253);
xor UO_385 (O_385,N_7528,N_8169);
xnor UO_386 (O_386,N_9005,N_9442);
nor UO_387 (O_387,N_9223,N_8346);
xnor UO_388 (O_388,N_9311,N_8428);
or UO_389 (O_389,N_9621,N_8394);
nor UO_390 (O_390,N_9530,N_9524);
and UO_391 (O_391,N_9149,N_9096);
and UO_392 (O_392,N_9076,N_8404);
nor UO_393 (O_393,N_8863,N_8898);
or UO_394 (O_394,N_7937,N_7660);
and UO_395 (O_395,N_7731,N_9459);
or UO_396 (O_396,N_8284,N_9717);
nor UO_397 (O_397,N_7998,N_8423);
nor UO_398 (O_398,N_8013,N_8063);
nor UO_399 (O_399,N_8611,N_8593);
xnor UO_400 (O_400,N_8932,N_9669);
nand UO_401 (O_401,N_9246,N_8906);
nor UO_402 (O_402,N_9836,N_9360);
xnor UO_403 (O_403,N_9047,N_8139);
xnor UO_404 (O_404,N_8657,N_8510);
nand UO_405 (O_405,N_8124,N_8789);
xor UO_406 (O_406,N_9462,N_9319);
xor UO_407 (O_407,N_9327,N_9170);
nor UO_408 (O_408,N_9961,N_9764);
nor UO_409 (O_409,N_8692,N_7777);
nand UO_410 (O_410,N_9725,N_9682);
or UO_411 (O_411,N_8895,N_8174);
and UO_412 (O_412,N_9194,N_9118);
and UO_413 (O_413,N_8603,N_9509);
nand UO_414 (O_414,N_7826,N_8828);
nor UO_415 (O_415,N_9429,N_7982);
nand UO_416 (O_416,N_7610,N_9979);
nand UO_417 (O_417,N_8994,N_8250);
xnor UO_418 (O_418,N_8159,N_7517);
xor UO_419 (O_419,N_9010,N_8401);
or UO_420 (O_420,N_9738,N_8379);
nand UO_421 (O_421,N_8802,N_8116);
nor UO_422 (O_422,N_7666,N_8444);
xor UO_423 (O_423,N_8391,N_9072);
and UO_424 (O_424,N_9542,N_8131);
xnor UO_425 (O_425,N_9765,N_8149);
xnor UO_426 (O_426,N_8929,N_8304);
or UO_427 (O_427,N_9325,N_8258);
and UO_428 (O_428,N_9807,N_8732);
or UO_429 (O_429,N_9507,N_8198);
and UO_430 (O_430,N_9760,N_9808);
and UO_431 (O_431,N_9430,N_9981);
xnor UO_432 (O_432,N_9608,N_8685);
or UO_433 (O_433,N_9382,N_9183);
and UO_434 (O_434,N_7965,N_8343);
or UO_435 (O_435,N_9173,N_8544);
xor UO_436 (O_436,N_8325,N_9152);
xnor UO_437 (O_437,N_9658,N_9470);
nor UO_438 (O_438,N_8473,N_7847);
and UO_439 (O_439,N_9115,N_7556);
or UO_440 (O_440,N_8726,N_8387);
xor UO_441 (O_441,N_9583,N_9614);
nor UO_442 (O_442,N_8412,N_9539);
and UO_443 (O_443,N_8252,N_9344);
or UO_444 (O_444,N_8307,N_8891);
xor UO_445 (O_445,N_7940,N_8988);
xnor UO_446 (O_446,N_7695,N_8043);
and UO_447 (O_447,N_9550,N_7794);
xnor UO_448 (O_448,N_9572,N_8065);
nor UO_449 (O_449,N_8438,N_8709);
and UO_450 (O_450,N_9837,N_9903);
or UO_451 (O_451,N_9777,N_8345);
or UO_452 (O_452,N_8208,N_8933);
or UO_453 (O_453,N_9119,N_9137);
or UO_454 (O_454,N_9234,N_9708);
or UO_455 (O_455,N_7626,N_9350);
nor UO_456 (O_456,N_9233,N_8592);
or UO_457 (O_457,N_9793,N_9817);
and UO_458 (O_458,N_9342,N_9933);
or UO_459 (O_459,N_7673,N_9527);
nor UO_460 (O_460,N_7891,N_8163);
or UO_461 (O_461,N_9300,N_8795);
or UO_462 (O_462,N_9630,N_9230);
and UO_463 (O_463,N_8752,N_8445);
and UO_464 (O_464,N_8992,N_7679);
and UO_465 (O_465,N_7882,N_9931);
nor UO_466 (O_466,N_7803,N_9156);
nor UO_467 (O_467,N_8974,N_8644);
or UO_468 (O_468,N_9637,N_9066);
and UO_469 (O_469,N_9862,N_8178);
nor UO_470 (O_470,N_9358,N_8494);
nor UO_471 (O_471,N_8580,N_8148);
or UO_472 (O_472,N_9573,N_9381);
nand UO_473 (O_473,N_8845,N_7565);
xor UO_474 (O_474,N_8867,N_8596);
nand UO_475 (O_475,N_8276,N_8851);
xor UO_476 (O_476,N_7822,N_8767);
and UO_477 (O_477,N_7643,N_8766);
nor UO_478 (O_478,N_8684,N_9943);
nor UO_479 (O_479,N_9265,N_8388);
xor UO_480 (O_480,N_9910,N_9127);
or UO_481 (O_481,N_8045,N_8425);
or UO_482 (O_482,N_9225,N_8138);
or UO_483 (O_483,N_8747,N_9923);
nand UO_484 (O_484,N_7504,N_7616);
and UO_485 (O_485,N_8919,N_9288);
xor UO_486 (O_486,N_9438,N_8941);
nand UO_487 (O_487,N_9726,N_9461);
and UO_488 (O_488,N_8793,N_7817);
xor UO_489 (O_489,N_8775,N_9983);
nand UO_490 (O_490,N_7624,N_8662);
nand UO_491 (O_491,N_9881,N_8648);
nand UO_492 (O_492,N_8853,N_7696);
xor UO_493 (O_493,N_7966,N_9302);
xor UO_494 (O_494,N_7738,N_8429);
xnor UO_495 (O_495,N_8335,N_9386);
or UO_496 (O_496,N_8465,N_9260);
nand UO_497 (O_497,N_9089,N_9100);
nor UO_498 (O_498,N_7709,N_7726);
and UO_499 (O_499,N_8980,N_8938);
xor UO_500 (O_500,N_8890,N_9249);
and UO_501 (O_501,N_8283,N_8466);
or UO_502 (O_502,N_9532,N_9084);
or UO_503 (O_503,N_8670,N_7887);
xnor UO_504 (O_504,N_8069,N_8479);
and UO_505 (O_505,N_9914,N_8666);
xnor UO_506 (O_506,N_9870,N_9965);
nand UO_507 (O_507,N_8492,N_9651);
nand UO_508 (O_508,N_8383,N_9975);
or UO_509 (O_509,N_9480,N_7787);
xnor UO_510 (O_510,N_9853,N_7935);
nor UO_511 (O_511,N_8682,N_7951);
xnor UO_512 (O_512,N_9740,N_9261);
and UO_513 (O_513,N_8160,N_8058);
and UO_514 (O_514,N_8101,N_9934);
and UO_515 (O_515,N_7724,N_7744);
or UO_516 (O_516,N_9996,N_9510);
xor UO_517 (O_517,N_8570,N_8228);
xnor UO_518 (O_518,N_8150,N_9730);
nand UO_519 (O_519,N_7939,N_7515);
xor UO_520 (O_520,N_9680,N_8718);
xnor UO_521 (O_521,N_9719,N_9889);
and UO_522 (O_522,N_9320,N_9191);
nand UO_523 (O_523,N_9193,N_8877);
nor UO_524 (O_524,N_9489,N_9168);
xnor UO_525 (O_525,N_9062,N_8344);
nor UO_526 (O_526,N_9080,N_9723);
or UO_527 (O_527,N_9122,N_9105);
and UO_528 (O_528,N_8338,N_8212);
and UO_529 (O_529,N_8374,N_8781);
xor UO_530 (O_530,N_7748,N_7760);
nand UO_531 (O_531,N_7872,N_8856);
nand UO_532 (O_532,N_7641,N_8790);
or UO_533 (O_533,N_8415,N_9686);
nand UO_534 (O_534,N_8825,N_9508);
nor UO_535 (O_535,N_7809,N_8643);
nor UO_536 (O_536,N_8303,N_7501);
nand UO_537 (O_537,N_9900,N_8254);
nand UO_538 (O_538,N_9395,N_7767);
xor UO_539 (O_539,N_7747,N_7659);
xor UO_540 (O_540,N_9762,N_8614);
nand UO_541 (O_541,N_9328,N_9515);
xnor UO_542 (O_542,N_9620,N_9226);
xnor UO_543 (O_543,N_8676,N_9240);
nand UO_544 (O_544,N_9966,N_8535);
nor UO_545 (O_545,N_7705,N_9188);
and UO_546 (O_546,N_9984,N_7603);
xor UO_547 (O_547,N_7855,N_9562);
nor UO_548 (O_548,N_7519,N_8064);
or UO_549 (O_549,N_9728,N_8194);
nor UO_550 (O_550,N_7527,N_9035);
nor UO_551 (O_551,N_7566,N_8112);
nor UO_552 (O_552,N_8203,N_8330);
nand UO_553 (O_553,N_8414,N_9707);
xnor UO_554 (O_554,N_7920,N_9441);
xnor UO_555 (O_555,N_8442,N_8977);
nor UO_556 (O_556,N_8615,N_9568);
xor UO_557 (O_557,N_8107,N_9854);
and UO_558 (O_558,N_9969,N_8009);
and UO_559 (O_559,N_8664,N_8753);
and UO_560 (O_560,N_9538,N_8096);
nor UO_561 (O_561,N_9660,N_9245);
and UO_562 (O_562,N_9959,N_7969);
nand UO_563 (O_563,N_9163,N_7625);
or UO_564 (O_564,N_8785,N_9241);
nor UO_565 (O_565,N_7990,N_8317);
nor UO_566 (O_566,N_8965,N_9081);
and UO_567 (O_567,N_9962,N_8837);
nand UO_568 (O_568,N_7944,N_9454);
and UO_569 (O_569,N_9790,N_9312);
nand UO_570 (O_570,N_8489,N_9835);
nor UO_571 (O_571,N_8461,N_7715);
nor UO_572 (O_572,N_7880,N_8872);
nand UO_573 (O_573,N_8144,N_9898);
or UO_574 (O_574,N_7587,N_9688);
and UO_575 (O_575,N_8256,N_9988);
xnor UO_576 (O_576,N_8257,N_8540);
xnor UO_577 (O_577,N_8180,N_7665);
and UO_578 (O_578,N_7617,N_8703);
nor UO_579 (O_579,N_9478,N_8490);
nor UO_580 (O_580,N_8263,N_9877);
and UO_581 (O_581,N_8011,N_9446);
xnor UO_582 (O_582,N_8023,N_8986);
xor UO_583 (O_583,N_8609,N_7864);
nor UO_584 (O_584,N_9169,N_8168);
or UO_585 (O_585,N_8215,N_8776);
and UO_586 (O_586,N_8270,N_9032);
and UO_587 (O_587,N_8854,N_8454);
nor UO_588 (O_588,N_8318,N_9787);
or UO_589 (O_589,N_8865,N_7681);
xor UO_590 (O_590,N_7591,N_8184);
or UO_591 (O_591,N_8068,N_7963);
nand UO_592 (O_592,N_8624,N_8185);
xnor UO_593 (O_593,N_8219,N_7808);
or UO_594 (O_594,N_8839,N_8997);
or UO_595 (O_595,N_8007,N_9306);
xor UO_596 (O_596,N_9058,N_9045);
nor UO_597 (O_597,N_9415,N_9751);
or UO_598 (O_598,N_8945,N_9471);
or UO_599 (O_599,N_8173,N_9055);
xnor UO_600 (O_600,N_9824,N_9525);
nand UO_601 (O_601,N_8991,N_9287);
or UO_602 (O_602,N_9493,N_9610);
and UO_603 (O_603,N_9580,N_7996);
nand UO_604 (O_604,N_8612,N_8061);
and UO_605 (O_605,N_8067,N_8079);
and UO_606 (O_606,N_8051,N_9484);
xor UO_607 (O_607,N_9710,N_9343);
nor UO_608 (O_608,N_8528,N_7502);
and UO_609 (O_609,N_9083,N_8050);
xnor UO_610 (O_610,N_7620,N_9332);
nor UO_611 (O_611,N_9632,N_9859);
and UO_612 (O_612,N_9147,N_8048);
nand UO_613 (O_613,N_9326,N_9638);
nor UO_614 (O_614,N_9813,N_8105);
or UO_615 (O_615,N_8158,N_7923);
or UO_616 (O_616,N_7781,N_9274);
nor UO_617 (O_617,N_9023,N_9547);
nand UO_618 (O_618,N_8339,N_9909);
or UO_619 (O_619,N_9251,N_9314);
nand UO_620 (O_620,N_9520,N_9244);
nor UO_621 (O_621,N_8757,N_8281);
nand UO_622 (O_622,N_9042,N_9882);
nor UO_623 (O_623,N_8803,N_8128);
and UO_624 (O_624,N_8146,N_9447);
and UO_625 (O_625,N_9978,N_9838);
and UO_626 (O_626,N_7994,N_8835);
and UO_627 (O_627,N_8015,N_8963);
nand UO_628 (O_628,N_7823,N_8693);
and UO_629 (O_629,N_8770,N_9031);
xnor UO_630 (O_630,N_7943,N_8702);
nand UO_631 (O_631,N_9270,N_9207);
xor UO_632 (O_632,N_9967,N_7581);
nor UO_633 (O_633,N_8524,N_8402);
xor UO_634 (O_634,N_8655,N_9494);
nand UO_635 (O_635,N_8842,N_9048);
nor UO_636 (O_636,N_9886,N_8829);
or UO_637 (O_637,N_9356,N_9993);
and UO_638 (O_638,N_9819,N_7554);
nor UO_639 (O_639,N_9874,N_9656);
and UO_640 (O_640,N_7601,N_8422);
or UO_641 (O_641,N_8285,N_9654);
xnor UO_642 (O_642,N_7644,N_8294);
nor UO_643 (O_643,N_8452,N_8310);
nand UO_644 (O_644,N_9692,N_9000);
xor UO_645 (O_645,N_8457,N_8434);
xnor UO_646 (O_646,N_8396,N_9540);
nand UO_647 (O_647,N_8698,N_8029);
nand UO_648 (O_648,N_8885,N_8165);
or UO_649 (O_649,N_9025,N_7722);
xnor UO_650 (O_650,N_9942,N_8641);
nand UO_651 (O_651,N_8209,N_9571);
nand UO_652 (O_652,N_8663,N_7736);
or UO_653 (O_653,N_9065,N_7784);
and UO_654 (O_654,N_9015,N_8550);
xor UO_655 (O_655,N_8417,N_8721);
nand UO_656 (O_656,N_8920,N_9629);
xnor UO_657 (O_657,N_9307,N_9598);
nand UO_658 (O_658,N_7766,N_7829);
or UO_659 (O_659,N_7578,N_9750);
or UO_660 (O_660,N_7916,N_7797);
or UO_661 (O_661,N_7894,N_8689);
xnor UO_662 (O_662,N_7828,N_9237);
and UO_663 (O_663,N_7545,N_8940);
nand UO_664 (O_664,N_8175,N_7946);
nor UO_665 (O_665,N_8103,N_9026);
nor UO_666 (O_666,N_8241,N_8493);
nand UO_667 (O_667,N_8924,N_8334);
nor UO_668 (O_668,N_7933,N_8861);
or UO_669 (O_669,N_9721,N_8082);
nand UO_670 (O_670,N_9953,N_9387);
or UO_671 (O_671,N_8804,N_9075);
xor UO_672 (O_672,N_8826,N_7687);
or UO_673 (O_673,N_9182,N_8917);
or UO_674 (O_674,N_7582,N_7682);
nand UO_675 (O_675,N_9545,N_8074);
xnor UO_676 (O_676,N_7592,N_9278);
or UO_677 (O_677,N_9154,N_8393);
xnor UO_678 (O_678,N_7796,N_9715);
nand UO_679 (O_679,N_9483,N_7513);
nand UO_680 (O_680,N_7550,N_8392);
xnor UO_681 (O_681,N_9968,N_8588);
and UO_682 (O_682,N_7952,N_8764);
nor UO_683 (O_683,N_9876,N_7628);
or UO_684 (O_684,N_7867,N_9949);
and UO_685 (O_685,N_8951,N_9737);
nor UO_686 (O_686,N_9904,N_8809);
nor UO_687 (O_687,N_8110,N_8759);
and UO_688 (O_688,N_7580,N_9301);
nand UO_689 (O_689,N_8135,N_9786);
nor UO_690 (O_690,N_9405,N_8049);
nand UO_691 (O_691,N_7732,N_7503);
nor UO_692 (O_692,N_8970,N_9008);
nor UO_693 (O_693,N_7650,N_9797);
nand UO_694 (O_694,N_9832,N_7983);
or UO_695 (O_695,N_8261,N_8218);
nand UO_696 (O_696,N_9143,N_8778);
nand UO_697 (O_697,N_9518,N_9186);
or UO_698 (O_698,N_7763,N_7553);
or UO_699 (O_699,N_8405,N_9443);
nor UO_700 (O_700,N_9299,N_7538);
and UO_701 (O_701,N_8990,N_7653);
nor UO_702 (O_702,N_7840,N_9329);
and UO_703 (O_703,N_8308,N_7849);
or UO_704 (O_704,N_8234,N_7531);
nor UO_705 (O_705,N_7563,N_8987);
and UO_706 (O_706,N_8534,N_9028);
nand UO_707 (O_707,N_8847,N_9659);
and UO_708 (O_708,N_8673,N_8511);
and UO_709 (O_709,N_8715,N_9623);
xor UO_710 (O_710,N_9535,N_9203);
nand UO_711 (O_711,N_8205,N_8548);
nor UO_712 (O_712,N_9145,N_9816);
or UO_713 (O_713,N_7941,N_9822);
or UO_714 (O_714,N_8152,N_8563);
nand UO_715 (O_715,N_7656,N_8734);
and UO_716 (O_716,N_9131,N_7919);
or UO_717 (O_717,N_8453,N_9930);
xor UO_718 (O_718,N_7827,N_7733);
nand UO_719 (O_719,N_9334,N_8005);
or UO_720 (O_720,N_9040,N_9171);
nand UO_721 (O_721,N_8627,N_7634);
nand UO_722 (O_722,N_7572,N_8577);
and UO_723 (O_723,N_8427,N_8355);
or UO_724 (O_724,N_8288,N_8707);
nand UO_725 (O_725,N_9794,N_7611);
xnor UO_726 (O_726,N_8724,N_9009);
and UO_727 (O_727,N_9436,N_7596);
or UO_728 (O_728,N_9491,N_8567);
or UO_729 (O_729,N_7700,N_8199);
xor UO_730 (O_730,N_9731,N_9057);
nand UO_731 (O_731,N_9449,N_9850);
and UO_732 (O_732,N_7753,N_9201);
and UO_733 (O_733,N_9668,N_9220);
or UO_734 (O_734,N_9789,N_8513);
nand UO_735 (O_735,N_8947,N_8660);
and UO_736 (O_736,N_8758,N_8622);
nor UO_737 (O_737,N_7904,N_9560);
or UO_738 (O_738,N_7514,N_7841);
nand UO_739 (O_739,N_9214,N_8735);
nand UO_740 (O_740,N_8342,N_7759);
xor UO_741 (O_741,N_8695,N_9561);
or UO_742 (O_742,N_9273,N_7622);
and UO_743 (O_743,N_9687,N_9374);
or UO_744 (O_744,N_8416,N_9211);
xor UO_745 (O_745,N_9098,N_8546);
or UO_746 (O_746,N_9435,N_8843);
or UO_747 (O_747,N_7674,N_9829);
xor UO_748 (O_748,N_8081,N_7717);
nor UO_749 (O_749,N_8605,N_7993);
or UO_750 (O_750,N_8569,N_7636);
xnor UO_751 (O_751,N_8265,N_9555);
and UO_752 (O_752,N_8299,N_9456);
xnor UO_753 (O_753,N_9033,N_9189);
or UO_754 (O_754,N_8683,N_9079);
nor UO_755 (O_755,N_8273,N_7585);
or UO_756 (O_756,N_8554,N_7897);
nor UO_757 (O_757,N_9282,N_9695);
nand UO_758 (O_758,N_8020,N_8032);
and UO_759 (O_759,N_8850,N_9013);
xor UO_760 (O_760,N_7821,N_9372);
nand UO_761 (O_761,N_9117,N_8287);
or UO_762 (O_762,N_9227,N_9402);
nand UO_763 (O_763,N_9992,N_8447);
or UO_764 (O_764,N_9606,N_9178);
and UO_765 (O_765,N_7967,N_8192);
xor UO_766 (O_766,N_9252,N_8656);
xor UO_767 (O_767,N_7860,N_7900);
xnor UO_768 (O_768,N_7607,N_8750);
or UO_769 (O_769,N_8240,N_9753);
xnor UO_770 (O_770,N_9516,N_9107);
and UO_771 (O_771,N_9523,N_7938);
xor UO_772 (O_772,N_9589,N_9148);
xor UO_773 (O_773,N_9297,N_9481);
and UO_774 (O_774,N_8862,N_7684);
xor UO_775 (O_775,N_9254,N_8154);
and UO_776 (O_776,N_9099,N_7569);
nand UO_777 (O_777,N_9922,N_9085);
or UO_778 (O_778,N_8606,N_9529);
and UO_779 (O_779,N_9166,N_9277);
nor UO_780 (O_780,N_8236,N_9452);
nand UO_781 (O_781,N_7510,N_8451);
nor UO_782 (O_782,N_7838,N_8361);
or UO_783 (O_783,N_9875,N_9317);
nor UO_784 (O_784,N_9020,N_8398);
or UO_785 (O_785,N_8996,N_7579);
or UO_786 (O_786,N_9232,N_7568);
xor UO_787 (O_787,N_7907,N_9321);
nand UO_788 (O_788,N_8080,N_9337);
xor UO_789 (O_789,N_9986,N_9116);
or UO_790 (O_790,N_7874,N_8277);
xnor UO_791 (O_791,N_9670,N_8893);
and UO_792 (O_792,N_7835,N_8620);
nand UO_793 (O_793,N_7728,N_7615);
and UO_794 (O_794,N_8902,N_7832);
and UO_795 (O_795,N_8799,N_7746);
xnor UO_796 (O_796,N_8450,N_8905);
nor UO_797 (O_797,N_9883,N_8811);
nor UO_798 (O_798,N_8565,N_8794);
nor UO_799 (O_799,N_7500,N_7642);
or UO_800 (O_800,N_9841,N_9612);
nor UO_801 (O_801,N_9955,N_9248);
nor UO_802 (O_802,N_7655,N_7595);
or UO_803 (O_803,N_9376,N_9426);
and UO_804 (O_804,N_7697,N_7754);
and UO_805 (O_805,N_8636,N_7561);
xnor UO_806 (O_806,N_8706,N_9027);
or UO_807 (O_807,N_8366,N_9558);
nor UO_808 (O_808,N_8362,N_9704);
xor UO_809 (O_809,N_9897,N_7631);
nor UO_810 (O_810,N_8164,N_9869);
and UO_811 (O_811,N_8818,N_8937);
or UO_812 (O_812,N_8132,N_8629);
and UO_813 (O_813,N_8899,N_8268);
xor UO_814 (O_814,N_9763,N_9002);
xnor UO_815 (O_815,N_9177,N_8579);
nor UO_816 (O_816,N_8282,N_9463);
or UO_817 (O_817,N_7668,N_8456);
and UO_818 (O_818,N_8302,N_9803);
or UO_819 (O_819,N_7704,N_9671);
or UO_820 (O_820,N_8819,N_9418);
nand UO_821 (O_821,N_8480,N_9643);
xor UO_822 (O_822,N_8012,N_8376);
xor UO_823 (O_823,N_9973,N_8498);
nand UO_824 (O_824,N_8378,N_9512);
nand UO_825 (O_825,N_7713,N_9756);
nand UO_826 (O_826,N_9022,N_7775);
xor UO_827 (O_827,N_8681,N_9187);
and UO_828 (O_828,N_7895,N_8558);
or UO_829 (O_829,N_7664,N_7756);
and UO_830 (O_830,N_7645,N_8892);
and UO_831 (O_831,N_9472,N_9422);
nand UO_832 (O_832,N_9990,N_8395);
or UO_833 (O_833,N_8737,N_8232);
nand UO_834 (O_834,N_9174,N_8003);
and UO_835 (O_835,N_7991,N_9567);
nor UO_836 (O_836,N_9283,N_8568);
or UO_837 (O_837,N_8476,N_7950);
and UO_838 (O_838,N_9600,N_9531);
nand UO_839 (O_839,N_8881,N_9262);
or UO_840 (O_840,N_9068,N_8491);
and UO_841 (O_841,N_9856,N_8832);
nand UO_842 (O_842,N_7804,N_7780);
or UO_843 (O_843,N_8244,N_9421);
nor UO_844 (O_844,N_9487,N_8197);
nand UO_845 (O_845,N_9622,N_7870);
and UO_846 (O_846,N_8247,N_8316);
nor UO_847 (O_847,N_8744,N_9534);
or UO_848 (O_848,N_8981,N_9857);
xor UO_849 (O_849,N_7676,N_8094);
or UO_850 (O_850,N_7960,N_8985);
nor UO_851 (O_851,N_9204,N_7716);
nor UO_852 (O_852,N_7507,N_9690);
xnor UO_853 (O_853,N_7770,N_9134);
nand UO_854 (O_854,N_9264,N_9420);
nand UO_855 (O_855,N_8102,N_7725);
nor UO_856 (O_856,N_8857,N_9941);
and UO_857 (O_857,N_9963,N_9349);
nor UO_858 (O_858,N_7670,N_8056);
and UO_859 (O_859,N_7805,N_8549);
and UO_860 (O_860,N_8046,N_9585);
nor UO_861 (O_861,N_8042,N_9551);
xor UO_862 (O_862,N_7535,N_8545);
or UO_863 (O_863,N_7536,N_9858);
and UO_864 (O_864,N_9927,N_7520);
or UO_865 (O_865,N_9492,N_9069);
xor UO_866 (O_866,N_8436,N_9864);
and UO_867 (O_867,N_8517,N_8319);
or UO_868 (O_868,N_8177,N_8968);
xnor UO_869 (O_869,N_8594,N_7912);
and UO_870 (O_870,N_9559,N_9034);
and UO_871 (O_871,N_9335,N_9662);
nand UO_872 (O_872,N_9759,N_9665);
and UO_873 (O_873,N_8844,N_8275);
and UO_874 (O_874,N_8943,N_9729);
or UO_875 (O_875,N_7774,N_9361);
nand UO_876 (O_876,N_8274,N_8619);
nand UO_877 (O_877,N_7706,N_9801);
xor UO_878 (O_878,N_8514,N_7820);
and UO_879 (O_879,N_8840,N_9460);
and UO_880 (O_880,N_7751,N_7698);
and UO_881 (O_881,N_7997,N_9087);
and UO_882 (O_882,N_8380,N_8123);
or UO_883 (O_883,N_9383,N_8125);
xnor UO_884 (O_884,N_9791,N_9747);
nor UO_885 (O_885,N_7884,N_8551);
nor UO_886 (O_886,N_9769,N_8772);
and UO_887 (O_887,N_9366,N_9255);
xnor UO_888 (O_888,N_8278,N_8973);
and UO_889 (O_889,N_9533,N_8271);
xnor UO_890 (O_890,N_9995,N_7573);
xnor UO_891 (O_891,N_8578,N_8998);
and UO_892 (O_892,N_9416,N_8960);
and UO_893 (O_893,N_7589,N_7548);
xnor UO_894 (O_894,N_9347,N_7932);
xor UO_895 (O_895,N_9106,N_9823);
and UO_896 (O_896,N_9827,N_8600);
or UO_897 (O_897,N_8904,N_8884);
or UO_898 (O_898,N_7558,N_8719);
nand UO_899 (O_899,N_8406,N_9648);
and UO_900 (O_900,N_8756,N_7970);
and UO_901 (O_901,N_7745,N_7534);
and UO_902 (O_902,N_9357,N_7734);
nand UO_903 (O_903,N_8057,N_9384);
and UO_904 (O_904,N_8095,N_7557);
nand UO_905 (O_905,N_8382,N_9586);
and UO_906 (O_906,N_8437,N_9313);
nand UO_907 (O_907,N_7972,N_9908);
nor UO_908 (O_908,N_9316,N_7877);
or UO_909 (O_909,N_8701,N_8503);
nand UO_910 (O_910,N_8564,N_8147);
and UO_911 (O_911,N_8426,N_8495);
nor UO_912 (O_912,N_8269,N_8109);
nor UO_913 (O_913,N_8371,N_7575);
nor UO_914 (O_914,N_7648,N_8922);
nor UO_915 (O_915,N_7599,N_9410);
nand UO_916 (O_916,N_8353,N_7593);
xnor UO_917 (O_917,N_9378,N_8654);
or UO_918 (O_918,N_8370,N_7798);
nor UO_919 (O_919,N_8690,N_8566);
nand UO_920 (O_920,N_8039,N_7905);
or UO_921 (O_921,N_7871,N_9628);
nand UO_922 (O_922,N_8054,N_8999);
or UO_923 (O_923,N_8859,N_9393);
xnor UO_924 (O_924,N_9901,N_8816);
or UO_925 (O_925,N_8509,N_9304);
xnor UO_926 (O_926,N_9733,N_9597);
or UO_927 (O_927,N_8677,N_9359);
nand UO_928 (O_928,N_8297,N_8730);
xnor UO_929 (O_929,N_8181,N_7816);
nand UO_930 (O_930,N_8953,N_8631);
or UO_931 (O_931,N_9217,N_7776);
nand UO_932 (O_932,N_8066,N_8508);
and UO_933 (O_933,N_9060,N_7576);
xor UO_934 (O_934,N_9425,N_7712);
nor UO_935 (O_935,N_8122,N_7604);
or UO_936 (O_936,N_9468,N_9124);
and UO_937 (O_937,N_9748,N_9757);
xor UO_938 (O_938,N_8449,N_7647);
or UO_939 (O_939,N_9584,N_9271);
and UO_940 (O_940,N_9891,N_7584);
nand UO_941 (O_941,N_8016,N_7623);
nor UO_942 (O_942,N_9070,N_8313);
or UO_943 (O_943,N_7901,N_9479);
nand UO_944 (O_944,N_8879,N_9077);
xnor UO_945 (O_945,N_9338,N_8222);
xor UO_946 (O_946,N_9498,N_9974);
xnor UO_947 (O_947,N_8033,N_8848);
and UO_948 (O_948,N_9884,N_7675);
nand UO_949 (O_949,N_9570,N_9434);
xnor UO_950 (O_950,N_8037,N_9195);
nor UO_951 (O_951,N_9678,N_7608);
nand UO_952 (O_952,N_7953,N_9496);
or UO_953 (O_953,N_8523,N_9497);
or UO_954 (O_954,N_8525,N_8478);
and UO_955 (O_955,N_8076,N_8251);
nor UO_956 (O_956,N_9681,N_9433);
nor UO_957 (O_957,N_7508,N_9078);
xor UO_958 (O_958,N_9213,N_9617);
or UO_959 (O_959,N_9615,N_8399);
xor UO_960 (O_960,N_8085,N_8443);
nand UO_961 (O_961,N_7661,N_8755);
nand UO_962 (O_962,N_8836,N_9161);
and UO_963 (O_963,N_9198,N_9286);
nand UO_964 (O_964,N_9092,N_7663);
and UO_965 (O_965,N_9905,N_7688);
xnor UO_966 (O_966,N_9495,N_8623);
xnor UO_967 (O_967,N_9331,N_9890);
nand UO_968 (O_968,N_9158,N_9275);
xor UO_969 (O_969,N_9457,N_9294);
nor UO_970 (O_970,N_8359,N_9536);
nor UO_971 (O_971,N_9132,N_9280);
and UO_972 (O_972,N_9772,N_7525);
nand UO_973 (O_973,N_8969,N_9336);
or UO_974 (O_974,N_7719,N_7979);
nand UO_975 (O_975,N_8191,N_9848);
nor UO_976 (O_976,N_9165,N_7945);
or UO_977 (O_977,N_7812,N_9616);
nand UO_978 (O_978,N_8728,N_9353);
nor UO_979 (O_979,N_9053,N_7613);
nand UO_980 (O_980,N_9755,N_8712);
xor UO_981 (O_981,N_9809,N_8332);
or UO_982 (O_982,N_9705,N_8820);
or UO_983 (O_983,N_9093,N_8001);
nand UO_984 (O_984,N_8852,N_9352);
and UO_985 (O_985,N_9050,N_8186);
nand UO_986 (O_986,N_9295,N_7708);
and UO_987 (O_987,N_8784,N_7830);
and UO_988 (O_988,N_7567,N_8876);
nor UO_989 (O_989,N_8077,N_7942);
and UO_990 (O_990,N_9683,N_8243);
xor UO_991 (O_991,N_7764,N_8910);
nand UO_992 (O_992,N_7926,N_9159);
or UO_993 (O_993,N_9920,N_7807);
nand UO_994 (O_994,N_9394,N_8928);
nor UO_995 (O_995,N_8333,N_9522);
nand UO_996 (O_996,N_9511,N_7721);
nor UO_997 (O_997,N_9830,N_8255);
nor UO_998 (O_998,N_7577,N_7692);
or UO_999 (O_999,N_9094,N_8166);
or UO_1000 (O_1000,N_7773,N_8321);
nand UO_1001 (O_1001,N_8008,N_9655);
xor UO_1002 (O_1002,N_7866,N_9631);
nor UO_1003 (O_1003,N_8481,N_7727);
nand UO_1004 (O_1004,N_7758,N_8504);
or UO_1005 (O_1005,N_8773,N_9935);
nor UO_1006 (O_1006,N_9197,N_8053);
and UO_1007 (O_1007,N_8505,N_8916);
or UO_1008 (O_1008,N_9150,N_9954);
nand UO_1009 (O_1009,N_7800,N_8413);
nand UO_1010 (O_1010,N_8389,N_9063);
nand UO_1011 (O_1011,N_7632,N_9976);
and UO_1012 (O_1012,N_7594,N_8400);
xnor UO_1013 (O_1013,N_8351,N_8487);
and UO_1014 (O_1014,N_7959,N_9557);
or UO_1015 (O_1015,N_8870,N_9916);
xor UO_1016 (O_1016,N_8957,N_9519);
nor UO_1017 (O_1017,N_7560,N_7836);
xnor UO_1018 (O_1018,N_9970,N_8295);
xnor UO_1019 (O_1019,N_9490,N_9153);
nand UO_1020 (O_1020,N_7848,N_9466);
xnor UO_1021 (O_1021,N_7505,N_8925);
or UO_1022 (O_1022,N_7637,N_8598);
nor UO_1023 (O_1023,N_8868,N_8279);
and UO_1024 (O_1024,N_9917,N_8618);
xor UO_1025 (O_1025,N_8833,N_8607);
xnor UO_1026 (O_1026,N_8966,N_8463);
and UO_1027 (O_1027,N_9915,N_8560);
and UO_1028 (O_1028,N_8921,N_8239);
and UO_1029 (O_1029,N_8787,N_8120);
nand UO_1030 (O_1030,N_9272,N_9625);
or UO_1031 (O_1031,N_8129,N_9544);
xnor UO_1032 (O_1032,N_9828,N_9907);
and UO_1033 (O_1033,N_8742,N_7691);
and UO_1034 (O_1034,N_8002,N_8464);
xor UO_1035 (O_1035,N_9474,N_9501);
and UO_1036 (O_1036,N_8659,N_9059);
nand UO_1037 (O_1037,N_9771,N_9184);
nand UO_1038 (O_1038,N_8385,N_8238);
and UO_1039 (O_1039,N_8369,N_7978);
nor UO_1040 (O_1040,N_9684,N_8950);
nor UO_1041 (O_1041,N_8807,N_9767);
or UO_1042 (O_1042,N_8441,N_8976);
and UO_1043 (O_1043,N_7544,N_8089);
xor UO_1044 (O_1044,N_9090,N_8935);
nor UO_1045 (O_1045,N_8440,N_8543);
nor UO_1046 (O_1046,N_9292,N_8610);
nor UO_1047 (O_1047,N_9373,N_9408);
and UO_1048 (O_1048,N_8377,N_9469);
xor UO_1049 (O_1049,N_8117,N_9016);
nor UO_1050 (O_1050,N_8458,N_9982);
and UO_1051 (O_1051,N_7588,N_7761);
nor UO_1052 (O_1052,N_8100,N_9157);
nand UO_1053 (O_1053,N_8761,N_7778);
xnor UO_1054 (O_1054,N_9554,N_8084);
nand UO_1055 (O_1055,N_9720,N_8710);
xnor UO_1056 (O_1056,N_7762,N_7562);
or UO_1057 (O_1057,N_7789,N_7516);
xnor UO_1058 (O_1058,N_8633,N_7749);
and UO_1059 (O_1059,N_7873,N_8989);
nand UO_1060 (O_1060,N_8207,N_7533);
nor UO_1061 (O_1061,N_9821,N_9582);
xnor UO_1062 (O_1062,N_9795,N_8502);
nor UO_1063 (O_1063,N_7889,N_9362);
nor UO_1064 (O_1064,N_9120,N_9537);
xor UO_1065 (O_1065,N_8542,N_9956);
and UO_1066 (O_1066,N_9126,N_8886);
xnor UO_1067 (O_1067,N_8589,N_8028);
nand UO_1068 (O_1068,N_8153,N_9840);
xnor UO_1069 (O_1069,N_8341,N_8694);
nand UO_1070 (O_1070,N_7844,N_7790);
or UO_1071 (O_1071,N_7511,N_8821);
nand UO_1072 (O_1072,N_8314,N_8367);
xnor UO_1073 (O_1073,N_7702,N_7856);
and UO_1074 (O_1074,N_8475,N_8838);
xor UO_1075 (O_1075,N_9044,N_8571);
nor UO_1076 (O_1076,N_7689,N_9506);
nor UO_1077 (O_1077,N_8699,N_8368);
nand UO_1078 (O_1078,N_9423,N_8765);
nor UO_1079 (O_1079,N_8375,N_9414);
nor UO_1080 (O_1080,N_7710,N_8172);
nand UO_1081 (O_1081,N_7986,N_8357);
xnor UO_1082 (O_1082,N_9303,N_8322);
and UO_1083 (O_1083,N_8574,N_8972);
or UO_1084 (O_1084,N_9998,N_9409);
xnor UO_1085 (O_1085,N_9101,N_9095);
and UO_1086 (O_1086,N_8628,N_8763);
or UO_1087 (O_1087,N_9006,N_9202);
nand UO_1088 (O_1088,N_8206,N_8526);
or UO_1089 (O_1089,N_9843,N_8044);
or UO_1090 (O_1090,N_8190,N_8025);
nor UO_1091 (O_1091,N_9367,N_7537);
nor UO_1092 (O_1092,N_7931,N_7989);
or UO_1093 (O_1093,N_9716,N_7875);
xnor UO_1094 (O_1094,N_8467,N_7750);
nor UO_1095 (O_1095,N_8958,N_9999);
nor UO_1096 (O_1096,N_9064,N_8727);
nand UO_1097 (O_1097,N_7651,N_8320);
or UO_1098 (O_1098,N_9229,N_8688);
nor UO_1099 (O_1099,N_9831,N_9256);
xor UO_1100 (O_1100,N_8323,N_8888);
or UO_1101 (O_1101,N_7612,N_9144);
xnor UO_1102 (O_1102,N_8381,N_9389);
and UO_1103 (O_1103,N_8869,N_9768);
xnor UO_1104 (O_1104,N_9056,N_8720);
nand UO_1105 (O_1105,N_9800,N_8864);
nor UO_1106 (O_1106,N_8070,N_7509);
and UO_1107 (O_1107,N_9222,N_9563);
and UO_1108 (O_1108,N_9860,N_7910);
nor UO_1109 (O_1109,N_8874,N_8959);
xor UO_1110 (O_1110,N_7742,N_9504);
or UO_1111 (O_1111,N_7973,N_8604);
nand UO_1112 (O_1112,N_8408,N_9994);
and UO_1113 (O_1113,N_8751,N_9218);
and UO_1114 (O_1114,N_8939,N_9780);
and UO_1115 (O_1115,N_8104,N_9038);
and UO_1116 (O_1116,N_9666,N_9205);
or UO_1117 (O_1117,N_8944,N_9136);
and UO_1118 (O_1118,N_8639,N_7602);
xnor UO_1119 (O_1119,N_9911,N_9541);
and UO_1120 (O_1120,N_9046,N_8880);
nand UO_1121 (O_1121,N_8300,N_8581);
or UO_1122 (O_1122,N_9242,N_8934);
xnor UO_1123 (O_1123,N_9216,N_9444);
nor UO_1124 (O_1124,N_7532,N_9663);
nand UO_1125 (O_1125,N_8740,N_9024);
xor UO_1126 (O_1126,N_8227,N_8113);
xor UO_1127 (O_1127,N_9702,N_9785);
and UO_1128 (O_1128,N_9799,N_9458);
and UO_1129 (O_1129,N_8411,N_9135);
nand UO_1130 (O_1130,N_9713,N_8813);
nor UO_1131 (O_1131,N_8931,N_7627);
and UO_1132 (O_1132,N_9701,N_8485);
nor UO_1133 (O_1133,N_8099,N_9866);
nand UO_1134 (O_1134,N_8171,N_8093);
nor UO_1135 (O_1135,N_7621,N_8908);
nor UO_1136 (O_1136,N_8559,N_7671);
nand UO_1137 (O_1137,N_9030,N_9206);
or UO_1138 (O_1138,N_9250,N_8883);
or UO_1139 (O_1139,N_8472,N_8887);
and UO_1140 (O_1140,N_7703,N_8155);
xor UO_1141 (O_1141,N_8521,N_7694);
and UO_1142 (O_1142,N_7949,N_8797);
nor UO_1143 (O_1143,N_9578,N_9577);
nor UO_1144 (O_1144,N_9605,N_7957);
nor UO_1145 (O_1145,N_9696,N_9987);
or UO_1146 (O_1146,N_8625,N_8329);
nand UO_1147 (O_1147,N_9088,N_9007);
xnor UO_1148 (O_1148,N_9341,N_7757);
and UO_1149 (O_1149,N_8088,N_9603);
nor UO_1150 (O_1150,N_8539,N_7906);
and UO_1151 (O_1151,N_9128,N_9330);
or UO_1152 (O_1152,N_9845,N_7814);
or UO_1153 (O_1153,N_9591,N_9851);
nor UO_1154 (O_1154,N_9257,N_7824);
or UO_1155 (O_1155,N_9937,N_7657);
or UO_1156 (O_1156,N_8824,N_7635);
xor UO_1157 (O_1157,N_7934,N_8266);
and UO_1158 (O_1158,N_8704,N_9061);
xnor UO_1159 (O_1159,N_8340,N_7896);
nand UO_1160 (O_1160,N_8420,N_8653);
nand UO_1161 (O_1161,N_8858,N_9385);
nand UO_1162 (O_1162,N_9820,N_7853);
xnor UO_1163 (O_1163,N_9689,N_8635);
or UO_1164 (O_1164,N_8621,N_9500);
nand UO_1165 (O_1165,N_9263,N_8983);
nand UO_1166 (O_1166,N_8901,N_9588);
nand UO_1167 (O_1167,N_9407,N_9958);
nor UO_1168 (O_1168,N_8900,N_8210);
nor UO_1169 (O_1169,N_9473,N_8354);
or UO_1170 (O_1170,N_8978,N_7739);
and UO_1171 (O_1171,N_8264,N_9476);
and UO_1172 (O_1172,N_8224,N_8878);
xnor UO_1173 (O_1173,N_9011,N_9650);
nor UO_1174 (O_1174,N_9691,N_9852);
or UO_1175 (O_1175,N_8817,N_9236);
nand UO_1176 (O_1176,N_8583,N_8424);
nor UO_1177 (O_1177,N_8075,N_9339);
nor UO_1178 (O_1178,N_9939,N_7597);
xnor UO_1179 (O_1179,N_8115,N_7540);
or UO_1180 (O_1180,N_8221,N_9258);
nor UO_1181 (O_1181,N_7574,N_8142);
nor UO_1182 (O_1182,N_8562,N_9268);
and UO_1183 (O_1183,N_9021,N_9847);
nor UO_1184 (O_1184,N_7512,N_8796);
and UO_1185 (O_1185,N_8912,N_8448);
or UO_1186 (O_1186,N_8136,N_7667);
nor UO_1187 (O_1187,N_9259,N_9318);
or UO_1188 (O_1188,N_8708,N_9224);
nor UO_1189 (O_1189,N_9199,N_9348);
nor UO_1190 (O_1190,N_7714,N_7865);
and UO_1191 (O_1191,N_7605,N_8352);
nand UO_1192 (O_1192,N_9247,N_8739);
nand UO_1193 (O_1193,N_9899,N_9924);
xor UO_1194 (O_1194,N_7546,N_7947);
nand UO_1195 (O_1195,N_9607,N_9712);
nand UO_1196 (O_1196,N_7524,N_8532);
xor UO_1197 (O_1197,N_7729,N_9051);
or UO_1198 (O_1198,N_8097,N_9865);
nor UO_1199 (O_1199,N_8918,N_8364);
xor UO_1200 (O_1200,N_9888,N_9345);
nand UO_1201 (O_1201,N_8301,N_9694);
xnor UO_1202 (O_1202,N_7707,N_7801);
nor UO_1203 (O_1203,N_7552,N_7640);
nor UO_1204 (O_1204,N_8188,N_9305);
xnor UO_1205 (O_1205,N_8873,N_9734);
and UO_1206 (O_1206,N_9340,N_7917);
nand UO_1207 (O_1207,N_7743,N_9587);
nand UO_1208 (O_1208,N_9893,N_7735);
or UO_1209 (O_1209,N_9868,N_8114);
xor UO_1210 (O_1210,N_9370,N_9176);
or UO_1211 (O_1211,N_8537,N_8806);
and UO_1212 (O_1212,N_9972,N_7892);
nand UO_1213 (O_1213,N_8350,N_9806);
nand UO_1214 (O_1214,N_9774,N_8914);
or UO_1215 (O_1215,N_9221,N_8658);
or UO_1216 (O_1216,N_8642,N_8483);
nor UO_1217 (O_1217,N_8669,N_9086);
nor UO_1218 (O_1218,N_7859,N_7846);
and UO_1219 (O_1219,N_8679,N_9773);
nand UO_1220 (O_1220,N_8946,N_7677);
or UO_1221 (O_1221,N_9846,N_9675);
nor UO_1222 (O_1222,N_9014,N_9604);
or UO_1223 (O_1223,N_8433,N_9792);
xnor UO_1224 (O_1224,N_9465,N_9388);
nand UO_1225 (O_1225,N_9279,N_8576);
nor UO_1226 (O_1226,N_8083,N_9595);
or UO_1227 (O_1227,N_9693,N_8650);
and UO_1228 (O_1228,N_8896,N_8418);
nor UO_1229 (O_1229,N_9439,N_8927);
xnor UO_1230 (O_1230,N_9179,N_8121);
or UO_1231 (O_1231,N_7985,N_9796);
nor UO_1232 (O_1232,N_8754,N_9431);
and UO_1233 (O_1233,N_8590,N_7825);
nand UO_1234 (O_1234,N_8871,N_8216);
xor UO_1235 (O_1235,N_7843,N_8200);
or UO_1236 (O_1236,N_9826,N_9564);
nand UO_1237 (O_1237,N_7752,N_9104);
or UO_1238 (O_1238,N_7782,N_8430);
and UO_1239 (O_1239,N_8501,N_8792);
xor UO_1240 (O_1240,N_8290,N_7539);
nand UO_1241 (O_1241,N_9732,N_8814);
nor UO_1242 (O_1242,N_9012,N_7672);
and UO_1243 (O_1243,N_8616,N_7618);
nor UO_1244 (O_1244,N_9672,N_9938);
xnor UO_1245 (O_1245,N_7600,N_9371);
and UO_1246 (O_1246,N_7992,N_9181);
nor UO_1247 (O_1247,N_8855,N_8849);
xor UO_1248 (O_1248,N_8019,N_8964);
nand UO_1249 (O_1249,N_8923,N_9703);
and UO_1250 (O_1250,N_8217,N_8866);
and UO_1251 (O_1251,N_9349,N_9653);
or UO_1252 (O_1252,N_8872,N_7839);
and UO_1253 (O_1253,N_7814,N_9631);
xnor UO_1254 (O_1254,N_9539,N_8700);
and UO_1255 (O_1255,N_7956,N_9264);
nor UO_1256 (O_1256,N_8823,N_8555);
or UO_1257 (O_1257,N_9432,N_8348);
or UO_1258 (O_1258,N_9791,N_8795);
xor UO_1259 (O_1259,N_8675,N_8032);
or UO_1260 (O_1260,N_9473,N_8514);
nand UO_1261 (O_1261,N_9299,N_9424);
or UO_1262 (O_1262,N_9159,N_9273);
xnor UO_1263 (O_1263,N_7641,N_8442);
or UO_1264 (O_1264,N_9382,N_8636);
xnor UO_1265 (O_1265,N_9077,N_9067);
and UO_1266 (O_1266,N_9597,N_9924);
nand UO_1267 (O_1267,N_9346,N_7586);
nand UO_1268 (O_1268,N_9894,N_7642);
or UO_1269 (O_1269,N_8799,N_9986);
and UO_1270 (O_1270,N_8093,N_8849);
and UO_1271 (O_1271,N_8789,N_7720);
nand UO_1272 (O_1272,N_7537,N_9315);
nor UO_1273 (O_1273,N_8800,N_8648);
nand UO_1274 (O_1274,N_7798,N_7616);
or UO_1275 (O_1275,N_9901,N_9464);
nor UO_1276 (O_1276,N_8709,N_8453);
nor UO_1277 (O_1277,N_8177,N_9596);
and UO_1278 (O_1278,N_8583,N_8749);
nor UO_1279 (O_1279,N_8956,N_7710);
xor UO_1280 (O_1280,N_7769,N_9101);
or UO_1281 (O_1281,N_9351,N_7682);
nand UO_1282 (O_1282,N_7845,N_9614);
nand UO_1283 (O_1283,N_8217,N_8945);
xnor UO_1284 (O_1284,N_9901,N_7601);
or UO_1285 (O_1285,N_9710,N_9859);
nor UO_1286 (O_1286,N_9169,N_9726);
or UO_1287 (O_1287,N_8212,N_9154);
nor UO_1288 (O_1288,N_8209,N_8954);
xor UO_1289 (O_1289,N_8992,N_9160);
nor UO_1290 (O_1290,N_9050,N_9765);
xnor UO_1291 (O_1291,N_8971,N_9648);
nor UO_1292 (O_1292,N_9441,N_9324);
xnor UO_1293 (O_1293,N_7669,N_7865);
and UO_1294 (O_1294,N_7582,N_8677);
nor UO_1295 (O_1295,N_9137,N_7929);
or UO_1296 (O_1296,N_8329,N_9585);
xnor UO_1297 (O_1297,N_8323,N_7719);
nor UO_1298 (O_1298,N_8702,N_9772);
and UO_1299 (O_1299,N_9110,N_9787);
nor UO_1300 (O_1300,N_9553,N_9980);
and UO_1301 (O_1301,N_7564,N_9347);
or UO_1302 (O_1302,N_9846,N_8140);
xor UO_1303 (O_1303,N_7954,N_8980);
nand UO_1304 (O_1304,N_8505,N_9569);
and UO_1305 (O_1305,N_9054,N_9158);
or UO_1306 (O_1306,N_7720,N_8538);
xnor UO_1307 (O_1307,N_9185,N_9551);
nor UO_1308 (O_1308,N_7913,N_7982);
nand UO_1309 (O_1309,N_9946,N_8757);
and UO_1310 (O_1310,N_7991,N_9978);
or UO_1311 (O_1311,N_9012,N_9949);
xnor UO_1312 (O_1312,N_8368,N_7715);
or UO_1313 (O_1313,N_9611,N_8636);
nand UO_1314 (O_1314,N_8968,N_9214);
or UO_1315 (O_1315,N_8058,N_9518);
xnor UO_1316 (O_1316,N_8052,N_9459);
xnor UO_1317 (O_1317,N_9817,N_9092);
nand UO_1318 (O_1318,N_7616,N_9854);
xnor UO_1319 (O_1319,N_9976,N_8576);
nor UO_1320 (O_1320,N_8463,N_9713);
nand UO_1321 (O_1321,N_9874,N_7980);
nor UO_1322 (O_1322,N_9982,N_8041);
nand UO_1323 (O_1323,N_9257,N_8328);
nor UO_1324 (O_1324,N_7666,N_8421);
or UO_1325 (O_1325,N_9432,N_9552);
nor UO_1326 (O_1326,N_7705,N_8824);
and UO_1327 (O_1327,N_8486,N_9951);
nand UO_1328 (O_1328,N_9751,N_8767);
and UO_1329 (O_1329,N_8889,N_8902);
nor UO_1330 (O_1330,N_9816,N_8229);
nand UO_1331 (O_1331,N_8796,N_9639);
nor UO_1332 (O_1332,N_8072,N_9098);
and UO_1333 (O_1333,N_7973,N_8993);
or UO_1334 (O_1334,N_7867,N_9561);
xor UO_1335 (O_1335,N_8919,N_9935);
nand UO_1336 (O_1336,N_7815,N_8476);
nor UO_1337 (O_1337,N_9605,N_9206);
and UO_1338 (O_1338,N_9144,N_8235);
and UO_1339 (O_1339,N_9401,N_9610);
and UO_1340 (O_1340,N_8548,N_7568);
and UO_1341 (O_1341,N_8285,N_7625);
xnor UO_1342 (O_1342,N_9887,N_8887);
and UO_1343 (O_1343,N_9440,N_9584);
or UO_1344 (O_1344,N_7525,N_9856);
xnor UO_1345 (O_1345,N_9741,N_9312);
nor UO_1346 (O_1346,N_8756,N_9645);
nand UO_1347 (O_1347,N_9577,N_8911);
and UO_1348 (O_1348,N_8435,N_8223);
nor UO_1349 (O_1349,N_8162,N_9743);
xnor UO_1350 (O_1350,N_9177,N_9173);
nor UO_1351 (O_1351,N_8141,N_9034);
and UO_1352 (O_1352,N_9908,N_8224);
xnor UO_1353 (O_1353,N_9923,N_8085);
and UO_1354 (O_1354,N_9228,N_8018);
nor UO_1355 (O_1355,N_8110,N_8431);
and UO_1356 (O_1356,N_7747,N_9120);
nor UO_1357 (O_1357,N_9277,N_7770);
and UO_1358 (O_1358,N_8433,N_9778);
nand UO_1359 (O_1359,N_7513,N_8248);
nand UO_1360 (O_1360,N_7982,N_8041);
and UO_1361 (O_1361,N_8742,N_8855);
and UO_1362 (O_1362,N_9764,N_9647);
xor UO_1363 (O_1363,N_9160,N_9313);
nand UO_1364 (O_1364,N_8806,N_8695);
and UO_1365 (O_1365,N_7702,N_8585);
nor UO_1366 (O_1366,N_7832,N_8467);
and UO_1367 (O_1367,N_8257,N_8818);
xor UO_1368 (O_1368,N_8267,N_9220);
or UO_1369 (O_1369,N_8987,N_9007);
nand UO_1370 (O_1370,N_9709,N_8082);
or UO_1371 (O_1371,N_8979,N_7840);
nand UO_1372 (O_1372,N_8581,N_9492);
xnor UO_1373 (O_1373,N_8830,N_9835);
and UO_1374 (O_1374,N_9876,N_9825);
xnor UO_1375 (O_1375,N_8998,N_8029);
xor UO_1376 (O_1376,N_7754,N_8930);
and UO_1377 (O_1377,N_9427,N_7797);
xor UO_1378 (O_1378,N_7941,N_8843);
nor UO_1379 (O_1379,N_7932,N_7532);
nand UO_1380 (O_1380,N_9532,N_7762);
or UO_1381 (O_1381,N_9635,N_9416);
or UO_1382 (O_1382,N_8726,N_7668);
and UO_1383 (O_1383,N_8857,N_8110);
xor UO_1384 (O_1384,N_9701,N_9992);
and UO_1385 (O_1385,N_9979,N_7633);
nand UO_1386 (O_1386,N_9183,N_7609);
nand UO_1387 (O_1387,N_9944,N_8262);
and UO_1388 (O_1388,N_9133,N_9591);
or UO_1389 (O_1389,N_9863,N_9100);
xor UO_1390 (O_1390,N_8923,N_9269);
xnor UO_1391 (O_1391,N_9714,N_8569);
or UO_1392 (O_1392,N_9250,N_9963);
xor UO_1393 (O_1393,N_8709,N_8021);
or UO_1394 (O_1394,N_9128,N_9065);
xnor UO_1395 (O_1395,N_9237,N_7986);
nor UO_1396 (O_1396,N_9463,N_9018);
xor UO_1397 (O_1397,N_7550,N_7564);
xnor UO_1398 (O_1398,N_9326,N_7579);
xor UO_1399 (O_1399,N_7857,N_8962);
xor UO_1400 (O_1400,N_8987,N_9411);
nand UO_1401 (O_1401,N_9698,N_8135);
or UO_1402 (O_1402,N_9172,N_8360);
nor UO_1403 (O_1403,N_9846,N_8061);
nor UO_1404 (O_1404,N_9949,N_8332);
or UO_1405 (O_1405,N_9431,N_9893);
xnor UO_1406 (O_1406,N_9123,N_9508);
or UO_1407 (O_1407,N_7593,N_8126);
nor UO_1408 (O_1408,N_9301,N_9646);
or UO_1409 (O_1409,N_7886,N_9057);
nand UO_1410 (O_1410,N_8035,N_8822);
nand UO_1411 (O_1411,N_9707,N_8598);
nor UO_1412 (O_1412,N_8441,N_7633);
or UO_1413 (O_1413,N_8204,N_7543);
nor UO_1414 (O_1414,N_9163,N_7588);
nand UO_1415 (O_1415,N_9830,N_8401);
nand UO_1416 (O_1416,N_8644,N_8910);
and UO_1417 (O_1417,N_7785,N_8228);
nor UO_1418 (O_1418,N_9179,N_9210);
and UO_1419 (O_1419,N_9400,N_7921);
and UO_1420 (O_1420,N_9698,N_8031);
or UO_1421 (O_1421,N_8765,N_9465);
and UO_1422 (O_1422,N_8798,N_9389);
xnor UO_1423 (O_1423,N_9254,N_7865);
or UO_1424 (O_1424,N_8899,N_9876);
and UO_1425 (O_1425,N_7856,N_9059);
and UO_1426 (O_1426,N_9780,N_8790);
or UO_1427 (O_1427,N_8333,N_8198);
xor UO_1428 (O_1428,N_8828,N_8178);
xnor UO_1429 (O_1429,N_7785,N_9329);
nor UO_1430 (O_1430,N_8041,N_7930);
xor UO_1431 (O_1431,N_9000,N_8749);
nand UO_1432 (O_1432,N_8015,N_9208);
and UO_1433 (O_1433,N_8610,N_9554);
nor UO_1434 (O_1434,N_9850,N_8833);
nand UO_1435 (O_1435,N_8632,N_7840);
nand UO_1436 (O_1436,N_9306,N_8843);
and UO_1437 (O_1437,N_8835,N_9340);
or UO_1438 (O_1438,N_8060,N_9363);
nand UO_1439 (O_1439,N_8097,N_7513);
nor UO_1440 (O_1440,N_7701,N_9845);
and UO_1441 (O_1441,N_8116,N_9770);
nand UO_1442 (O_1442,N_9981,N_8338);
or UO_1443 (O_1443,N_9679,N_9033);
or UO_1444 (O_1444,N_8356,N_9022);
nor UO_1445 (O_1445,N_9574,N_9910);
and UO_1446 (O_1446,N_7779,N_9919);
or UO_1447 (O_1447,N_8587,N_7818);
nand UO_1448 (O_1448,N_9009,N_9422);
and UO_1449 (O_1449,N_8688,N_8073);
xor UO_1450 (O_1450,N_9562,N_8889);
xnor UO_1451 (O_1451,N_8955,N_9127);
nor UO_1452 (O_1452,N_9021,N_9491);
or UO_1453 (O_1453,N_9387,N_8848);
xnor UO_1454 (O_1454,N_8950,N_7642);
nor UO_1455 (O_1455,N_8902,N_9824);
or UO_1456 (O_1456,N_9250,N_9379);
xnor UO_1457 (O_1457,N_7545,N_7943);
and UO_1458 (O_1458,N_9147,N_9329);
or UO_1459 (O_1459,N_8133,N_9115);
and UO_1460 (O_1460,N_9069,N_9273);
and UO_1461 (O_1461,N_7652,N_9651);
and UO_1462 (O_1462,N_8555,N_9257);
and UO_1463 (O_1463,N_8058,N_8608);
nor UO_1464 (O_1464,N_9220,N_8886);
nor UO_1465 (O_1465,N_8157,N_8900);
or UO_1466 (O_1466,N_7653,N_8191);
nor UO_1467 (O_1467,N_9017,N_8529);
or UO_1468 (O_1468,N_8421,N_8588);
or UO_1469 (O_1469,N_9518,N_7574);
nor UO_1470 (O_1470,N_9757,N_9557);
nor UO_1471 (O_1471,N_7833,N_9119);
xor UO_1472 (O_1472,N_9056,N_9371);
and UO_1473 (O_1473,N_9103,N_9511);
nor UO_1474 (O_1474,N_7652,N_9363);
and UO_1475 (O_1475,N_9713,N_9425);
nor UO_1476 (O_1476,N_7973,N_7995);
xor UO_1477 (O_1477,N_8890,N_9631);
nand UO_1478 (O_1478,N_9164,N_8620);
nor UO_1479 (O_1479,N_9783,N_9623);
nand UO_1480 (O_1480,N_8139,N_9612);
and UO_1481 (O_1481,N_9512,N_8173);
or UO_1482 (O_1482,N_9908,N_9438);
nor UO_1483 (O_1483,N_9713,N_8930);
and UO_1484 (O_1484,N_7861,N_7953);
or UO_1485 (O_1485,N_8195,N_9761);
and UO_1486 (O_1486,N_9549,N_8203);
or UO_1487 (O_1487,N_8632,N_8841);
and UO_1488 (O_1488,N_9906,N_7720);
or UO_1489 (O_1489,N_9059,N_9873);
nand UO_1490 (O_1490,N_9501,N_8470);
xnor UO_1491 (O_1491,N_8037,N_8806);
xnor UO_1492 (O_1492,N_7743,N_8415);
xor UO_1493 (O_1493,N_8098,N_8712);
or UO_1494 (O_1494,N_8402,N_8052);
nand UO_1495 (O_1495,N_8199,N_7859);
nor UO_1496 (O_1496,N_7748,N_8826);
nand UO_1497 (O_1497,N_8184,N_7570);
and UO_1498 (O_1498,N_7719,N_7661);
nor UO_1499 (O_1499,N_9436,N_8024);
endmodule