module basic_1000_10000_1500_100_levels_5xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
xnor U0 (N_0,In_736,In_785);
nand U1 (N_1,In_871,In_241);
or U2 (N_2,In_727,In_971);
nor U3 (N_3,In_208,In_349);
nand U4 (N_4,In_520,In_395);
and U5 (N_5,In_403,In_632);
nand U6 (N_6,In_321,In_501);
and U7 (N_7,In_825,In_153);
nor U8 (N_8,In_938,In_546);
or U9 (N_9,In_570,In_442);
nor U10 (N_10,In_393,In_148);
or U11 (N_11,In_571,In_246);
or U12 (N_12,In_866,In_230);
or U13 (N_13,In_596,In_214);
xnor U14 (N_14,In_455,In_243);
and U15 (N_15,In_933,In_821);
nand U16 (N_16,In_942,In_118);
xor U17 (N_17,In_444,In_575);
and U18 (N_18,In_223,In_239);
nor U19 (N_19,In_616,In_647);
nand U20 (N_20,In_244,In_702);
nor U21 (N_21,In_591,In_334);
or U22 (N_22,In_629,In_946);
and U23 (N_23,In_749,In_965);
and U24 (N_24,In_401,In_906);
and U25 (N_25,In_672,In_402);
and U26 (N_26,In_220,In_495);
nand U27 (N_27,In_276,In_492);
nor U28 (N_28,In_792,In_469);
or U29 (N_29,In_253,In_994);
or U30 (N_30,In_394,In_878);
or U31 (N_31,In_294,In_648);
and U32 (N_32,In_592,In_304);
nor U33 (N_33,In_112,In_113);
or U34 (N_34,In_751,In_265);
and U35 (N_35,In_865,In_614);
xnor U36 (N_36,In_756,In_860);
and U37 (N_37,In_200,In_108);
or U38 (N_38,In_360,In_932);
nor U39 (N_39,In_264,In_149);
nor U40 (N_40,In_445,In_977);
nand U41 (N_41,In_679,In_436);
nor U42 (N_42,In_896,In_982);
nor U43 (N_43,In_630,In_165);
nand U44 (N_44,In_519,In_275);
nand U45 (N_45,In_964,In_453);
or U46 (N_46,In_920,In_595);
or U47 (N_47,In_370,In_375);
and U48 (N_48,In_891,In_615);
nand U49 (N_49,In_27,In_178);
or U50 (N_50,In_653,In_837);
or U51 (N_51,In_64,In_85);
nand U52 (N_52,In_30,In_398);
nor U53 (N_53,In_717,In_24);
and U54 (N_54,In_659,In_564);
and U55 (N_55,In_651,In_735);
xor U56 (N_56,In_236,In_586);
nand U57 (N_57,In_611,In_386);
nand U58 (N_58,In_836,In_274);
and U59 (N_59,In_449,In_28);
xnor U60 (N_60,In_251,In_119);
and U61 (N_61,In_888,In_911);
nand U62 (N_62,In_950,In_376);
or U63 (N_63,In_867,In_598);
xnor U64 (N_64,In_104,In_768);
or U65 (N_65,In_904,In_432);
nor U66 (N_66,In_279,In_183);
nor U67 (N_67,In_284,In_995);
and U68 (N_68,In_103,In_325);
nor U69 (N_69,In_195,In_56);
nor U70 (N_70,In_844,In_714);
nand U71 (N_71,In_905,In_340);
or U72 (N_72,In_159,In_59);
nand U73 (N_73,In_677,In_926);
or U74 (N_74,In_743,In_824);
or U75 (N_75,In_74,In_799);
nand U76 (N_76,In_823,In_635);
nor U77 (N_77,In_790,In_468);
nand U78 (N_78,In_310,In_431);
nor U79 (N_79,In_706,In_428);
nor U80 (N_80,In_527,In_408);
and U81 (N_81,In_34,In_228);
nand U82 (N_82,In_288,In_175);
and U83 (N_83,In_271,In_357);
and U84 (N_84,In_345,In_471);
nor U85 (N_85,In_801,In_76);
or U86 (N_86,In_126,In_140);
nand U87 (N_87,In_914,In_36);
nor U88 (N_88,In_259,In_86);
and U89 (N_89,In_561,In_354);
nor U90 (N_90,In_503,In_480);
nor U91 (N_91,In_681,In_332);
and U92 (N_92,In_212,In_855);
or U93 (N_93,In_700,In_634);
and U94 (N_94,In_948,In_999);
nand U95 (N_95,In_122,In_723);
nand U96 (N_96,In_897,In_68);
nand U97 (N_97,In_473,In_405);
nand U98 (N_98,In_231,In_806);
or U99 (N_99,In_956,In_922);
nand U100 (N_100,In_441,In_998);
nand U101 (N_101,In_524,In_72);
nand U102 (N_102,In_568,In_752);
nand U103 (N_103,In_516,In_606);
nor U104 (N_104,In_397,In_880);
nor U105 (N_105,In_990,In_757);
xnor U106 (N_106,In_141,In_923);
and U107 (N_107,In_205,In_301);
xnor U108 (N_108,N_43,In_822);
or U109 (N_109,In_767,In_350);
and U110 (N_110,In_188,In_708);
nor U111 (N_111,In_868,In_795);
nor U112 (N_112,N_26,In_777);
nand U113 (N_113,In_830,In_551);
or U114 (N_114,N_51,In_302);
and U115 (N_115,In_879,In_580);
or U116 (N_116,In_160,In_158);
and U117 (N_117,In_798,N_58);
nor U118 (N_118,In_222,In_784);
and U119 (N_119,In_423,In_486);
or U120 (N_120,N_92,In_960);
nor U121 (N_121,In_710,In_45);
nor U122 (N_122,In_996,In_381);
and U123 (N_123,In_762,In_989);
nand U124 (N_124,In_957,In_523);
nor U125 (N_125,In_23,In_831);
xnor U126 (N_126,In_399,N_64);
nand U127 (N_127,In_931,In_556);
nor U128 (N_128,N_67,In_721);
nor U129 (N_129,N_65,N_1);
nand U130 (N_130,N_25,N_46);
nor U131 (N_131,In_627,In_162);
nor U132 (N_132,In_364,In_840);
and U133 (N_133,N_59,In_48);
or U134 (N_134,In_98,In_882);
and U135 (N_135,In_992,In_881);
nor U136 (N_136,In_384,N_90);
and U137 (N_137,In_430,In_796);
and U138 (N_138,In_300,In_37);
nor U139 (N_139,In_572,In_216);
nor U140 (N_140,In_587,In_440);
xor U141 (N_141,In_322,In_377);
xor U142 (N_142,In_176,In_603);
nor U143 (N_143,In_715,N_72);
nor U144 (N_144,In_125,In_578);
and U145 (N_145,In_505,N_99);
nor U146 (N_146,In_248,In_704);
nand U147 (N_147,In_850,In_202);
nor U148 (N_148,In_373,In_323);
or U149 (N_149,N_61,In_552);
and U150 (N_150,In_111,In_820);
xor U151 (N_151,In_686,In_335);
nor U152 (N_152,In_641,N_37);
and U153 (N_153,In_380,In_565);
nand U154 (N_154,In_15,In_963);
nor U155 (N_155,In_429,In_389);
xnor U156 (N_156,In_167,In_314);
or U157 (N_157,In_229,In_387);
and U158 (N_158,In_936,In_156);
or U159 (N_159,In_260,In_233);
nand U160 (N_160,In_538,In_585);
nor U161 (N_161,In_512,N_9);
or U162 (N_162,In_50,In_161);
nor U163 (N_163,In_414,In_984);
nand U164 (N_164,N_48,In_297);
nor U165 (N_165,N_60,In_548);
or U166 (N_166,In_739,N_4);
or U167 (N_167,N_70,In_780);
or U168 (N_168,In_579,N_3);
nand U169 (N_169,In_741,In_907);
or U170 (N_170,In_346,In_975);
or U171 (N_171,In_351,In_312);
nor U172 (N_172,In_899,In_813);
nor U173 (N_173,N_98,In_978);
and U174 (N_174,In_848,In_811);
or U175 (N_175,In_818,In_128);
or U176 (N_176,In_734,In_789);
nand U177 (N_177,In_769,In_65);
or U178 (N_178,In_529,In_192);
or U179 (N_179,In_262,In_307);
nand U180 (N_180,In_885,In_604);
nor U181 (N_181,In_191,In_225);
or U182 (N_182,N_45,In_863);
nand U183 (N_183,In_759,In_462);
or U184 (N_184,In_53,N_34);
nor U185 (N_185,In_418,In_477);
nor U186 (N_186,In_249,In_410);
nand U187 (N_187,In_326,In_282);
xor U188 (N_188,In_658,In_182);
nand U189 (N_189,In_290,In_664);
xor U190 (N_190,In_26,In_481);
xor U191 (N_191,In_569,In_698);
xor U192 (N_192,In_170,In_391);
xnor U193 (N_193,In_18,In_99);
nor U194 (N_194,In_943,In_81);
xor U195 (N_195,In_110,In_55);
nor U196 (N_196,In_594,In_466);
nand U197 (N_197,In_242,In_525);
and U198 (N_198,In_77,N_38);
nor U199 (N_199,N_66,In_600);
xor U200 (N_200,In_333,N_18);
or U201 (N_201,N_160,In_925);
and U202 (N_202,N_137,In_227);
nor U203 (N_203,In_839,In_625);
nor U204 (N_204,In_261,In_232);
nand U205 (N_205,In_371,In_201);
and U206 (N_206,N_123,In_20);
and U207 (N_207,N_178,N_186);
nand U208 (N_208,In_774,In_940);
and U209 (N_209,N_68,N_85);
xnor U210 (N_210,N_96,In_452);
and U211 (N_211,In_947,In_497);
and U212 (N_212,In_668,In_67);
and U213 (N_213,In_138,N_69);
xnor U214 (N_214,In_786,N_112);
nand U215 (N_215,In_2,In_915);
xor U216 (N_216,In_114,N_195);
or U217 (N_217,In_152,In_47);
or U218 (N_218,In_857,In_890);
and U219 (N_219,N_194,In_46);
or U220 (N_220,In_203,N_102);
nor U221 (N_221,N_78,In_691);
nand U222 (N_222,In_235,In_134);
nor U223 (N_223,In_478,In_16);
or U224 (N_224,In_667,In_808);
nand U225 (N_225,N_42,N_0);
and U226 (N_226,In_535,N_88);
and U227 (N_227,In_210,In_489);
xor U228 (N_228,In_256,In_355);
nor U229 (N_229,In_139,In_819);
nor U230 (N_230,In_547,In_910);
and U231 (N_231,In_221,In_130);
nand U232 (N_232,In_908,In_102);
nor U233 (N_233,In_21,In_12);
and U234 (N_234,In_463,N_179);
xnor U235 (N_235,In_859,In_645);
nand U236 (N_236,N_164,In_883);
nand U237 (N_237,In_804,In_35);
nand U238 (N_238,In_456,N_93);
and U239 (N_239,In_198,In_448);
xnor U240 (N_240,In_690,N_55);
and U241 (N_241,In_928,In_218);
and U242 (N_242,In_439,N_97);
and U243 (N_243,In_107,N_13);
and U244 (N_244,N_24,In_1);
or U245 (N_245,In_601,In_404);
xor U246 (N_246,In_487,N_124);
nor U247 (N_247,N_20,In_268);
nor U248 (N_248,In_316,N_152);
xnor U249 (N_249,In_422,N_63);
or U250 (N_250,In_577,N_30);
or U251 (N_251,In_317,In_245);
and U252 (N_252,In_842,In_919);
and U253 (N_253,N_82,In_509);
nand U254 (N_254,N_157,N_148);
and U255 (N_255,In_726,In_562);
or U256 (N_256,In_873,In_419);
and U257 (N_257,N_135,N_126);
nand U258 (N_258,N_163,In_609);
and U259 (N_259,In_83,In_461);
nand U260 (N_260,In_266,In_522);
or U261 (N_261,In_378,In_411);
and U262 (N_262,In_286,In_973);
and U263 (N_263,In_802,In_754);
nand U264 (N_264,In_135,In_967);
and U265 (N_265,In_318,In_460);
and U266 (N_266,In_713,In_238);
and U267 (N_267,N_151,N_106);
nand U268 (N_268,N_73,In_44);
xnor U269 (N_269,In_699,In_961);
and U270 (N_270,In_952,In_289);
nand U271 (N_271,In_631,In_909);
nor U272 (N_272,In_412,In_764);
or U273 (N_273,In_530,In_589);
nand U274 (N_274,In_738,N_27);
nor U275 (N_275,In_898,In_293);
nor U276 (N_276,N_153,In_413);
nor U277 (N_277,In_966,In_90);
or U278 (N_278,In_320,In_545);
or U279 (N_279,In_674,N_108);
nor U280 (N_280,N_138,In_13);
nor U281 (N_281,N_169,In_215);
or U282 (N_282,In_646,In_750);
or U283 (N_283,In_793,In_61);
or U284 (N_284,In_313,In_788);
nor U285 (N_285,In_273,In_84);
nor U286 (N_286,In_147,N_122);
or U287 (N_287,In_272,N_174);
nand U288 (N_288,In_935,In_356);
or U289 (N_289,In_117,In_582);
nand U290 (N_290,In_532,N_117);
or U291 (N_291,N_136,N_105);
nand U292 (N_292,In_144,In_748);
xnor U293 (N_293,N_7,In_540);
or U294 (N_294,In_6,N_29);
nand U295 (N_295,In_969,In_979);
nand U296 (N_296,In_237,In_94);
or U297 (N_297,In_91,In_917);
xnor U298 (N_298,N_191,In_278);
and U299 (N_299,N_104,In_347);
or U300 (N_300,In_337,N_272);
xnor U301 (N_301,In_42,N_183);
nor U302 (N_302,In_683,In_490);
nand U303 (N_303,In_918,N_259);
nor U304 (N_304,In_800,In_19);
nand U305 (N_305,In_675,N_285);
or U306 (N_306,In_164,In_981);
nand U307 (N_307,In_157,N_12);
or U308 (N_308,In_746,N_41);
xor U309 (N_309,In_892,In_760);
and U310 (N_310,In_772,In_513);
nand U311 (N_311,N_262,N_220);
xor U312 (N_312,N_75,In_776);
nand U313 (N_313,In_531,N_16);
xor U314 (N_314,In_396,N_172);
and U315 (N_315,In_88,In_833);
and U316 (N_316,N_265,In_687);
xor U317 (N_317,In_281,In_362);
nand U318 (N_318,N_227,In_678);
xnor U319 (N_319,N_103,In_0);
and U320 (N_320,In_199,In_435);
xnor U321 (N_321,In_299,N_280);
or U322 (N_322,In_464,In_78);
nand U323 (N_323,In_816,N_166);
nand U324 (N_324,In_184,N_260);
nand U325 (N_325,N_213,In_287);
or U326 (N_326,In_382,In_311);
or U327 (N_327,In_189,In_916);
nand U328 (N_328,In_851,In_719);
nor U329 (N_329,In_331,In_602);
or U330 (N_330,In_96,In_425);
or U331 (N_331,N_94,In_902);
nor U332 (N_332,In_330,In_987);
nand U333 (N_333,In_877,N_297);
nor U334 (N_334,In_458,In_959);
or U335 (N_335,In_493,N_33);
or U336 (N_336,N_222,N_197);
xnor U337 (N_337,In_541,N_147);
nor U338 (N_338,N_199,In_163);
and U339 (N_339,N_32,In_845);
and U340 (N_340,In_204,In_385);
and U341 (N_341,N_168,N_76);
and U342 (N_342,In_180,In_177);
or U343 (N_343,In_955,N_276);
nor U344 (N_344,N_253,N_238);
xnor U345 (N_345,In_951,N_39);
or U346 (N_346,In_433,In_753);
and U347 (N_347,In_115,In_500);
and U348 (N_348,In_544,In_549);
nor U349 (N_349,N_236,In_705);
xor U350 (N_350,In_367,N_266);
nand U351 (N_351,In_31,In_129);
and U352 (N_352,In_876,In_559);
and U353 (N_353,In_617,In_958);
or U354 (N_354,N_2,N_167);
and U355 (N_355,In_567,In_680);
nor U356 (N_356,N_275,N_44);
or U357 (N_357,In_665,N_80);
nor U358 (N_358,In_41,In_426);
nand U359 (N_359,In_470,N_6);
nand U360 (N_360,In_32,In_841);
nor U361 (N_361,In_709,In_584);
nor U362 (N_362,N_14,In_224);
and U363 (N_363,In_11,N_294);
and U364 (N_364,N_291,In_49);
and U365 (N_365,In_344,In_894);
nor U366 (N_366,N_133,In_359);
and U367 (N_367,In_689,In_63);
nor U368 (N_368,N_216,In_269);
nor U369 (N_369,In_974,N_279);
or U370 (N_370,In_69,N_22);
and U371 (N_371,N_118,N_212);
and U372 (N_372,In_869,N_228);
nand U373 (N_373,In_427,In_146);
nand U374 (N_374,N_114,In_716);
and U375 (N_375,N_261,N_221);
or U376 (N_376,N_209,In_744);
nor U377 (N_377,In_517,In_137);
nor U378 (N_378,In_849,In_619);
or U379 (N_379,N_182,In_54);
nor U380 (N_380,N_237,N_91);
or U381 (N_381,In_962,In_25);
nor U382 (N_382,N_15,In_758);
nand U383 (N_383,In_70,In_476);
and U384 (N_384,N_143,N_35);
nand U385 (N_385,In_339,N_284);
xor U386 (N_386,In_610,In_729);
nor U387 (N_387,N_251,In_720);
xor U388 (N_388,In_725,In_573);
or U389 (N_389,In_874,In_624);
and U390 (N_390,N_217,N_290);
and U391 (N_391,In_660,In_930);
or U392 (N_392,In_60,N_175);
and U393 (N_393,N_154,In_475);
and U394 (N_394,In_639,In_57);
nand U395 (N_395,In_652,In_847);
and U396 (N_396,N_264,In_4);
nor U397 (N_397,In_353,In_543);
or U398 (N_398,N_77,N_125);
or U399 (N_399,In_252,N_159);
or U400 (N_400,N_358,N_231);
nand U401 (N_401,In_366,In_379);
nor U402 (N_402,In_219,N_301);
and U403 (N_403,N_326,N_319);
and U404 (N_404,In_763,N_232);
and U405 (N_405,In_765,N_52);
nor U406 (N_406,N_158,In_447);
nand U407 (N_407,In_406,In_654);
nor U408 (N_408,In_887,N_339);
and U409 (N_409,N_11,N_374);
and U410 (N_410,N_161,In_858);
nand U411 (N_411,In_781,In_508);
and U412 (N_412,In_638,N_363);
or U413 (N_413,In_132,In_695);
and U414 (N_414,In_608,In_187);
xor U415 (N_415,N_17,N_371);
xnor U416 (N_416,In_515,In_181);
nor U417 (N_417,N_344,N_81);
and U418 (N_418,In_536,In_526);
nor U419 (N_419,N_360,In_701);
nor U420 (N_420,In_79,N_338);
nand U421 (N_421,In_770,In_217);
and U422 (N_422,In_737,N_170);
nor U423 (N_423,In_852,In_75);
or U424 (N_424,In_451,In_901);
and U425 (N_425,In_82,In_438);
or U426 (N_426,N_377,N_203);
or U427 (N_427,In_291,In_250);
nor U428 (N_428,N_367,N_254);
nor U429 (N_429,N_187,N_269);
xor U430 (N_430,In_296,In_136);
xnor U431 (N_431,In_179,In_929);
nand U432 (N_432,In_870,N_248);
nand U433 (N_433,In_518,In_563);
or U434 (N_434,N_388,In_688);
or U435 (N_435,N_113,N_373);
nor U436 (N_436,N_79,N_270);
nor U437 (N_437,In_694,In_853);
or U438 (N_438,N_318,In_213);
or U439 (N_439,In_711,In_174);
nand U440 (N_440,N_111,In_383);
nand U441 (N_441,In_986,In_937);
or U442 (N_442,In_742,N_36);
xor U443 (N_443,In_829,In_446);
and U444 (N_444,N_115,N_246);
nand U445 (N_445,In_479,In_434);
and U446 (N_446,In_194,In_968);
or U447 (N_447,In_502,N_299);
or U448 (N_448,In_566,N_395);
nand U449 (N_449,In_854,N_389);
nand U450 (N_450,In_605,In_663);
xor U451 (N_451,In_109,In_150);
and U452 (N_452,N_323,In_612);
or U453 (N_453,N_349,In_87);
nor U454 (N_454,N_206,In_173);
or U455 (N_455,In_766,N_139);
or U456 (N_456,In_172,In_620);
nor U457 (N_457,In_787,N_140);
and U458 (N_458,In_498,N_193);
or U459 (N_459,In_484,In_496);
nand U460 (N_460,In_557,In_327);
or U461 (N_461,In_812,N_235);
xor U462 (N_462,In_558,N_256);
nand U463 (N_463,In_731,In_483);
or U464 (N_464,In_73,N_119);
xor U465 (N_465,In_169,N_271);
nand U466 (N_466,N_352,In_537);
nand U467 (N_467,In_782,In_722);
nand U468 (N_468,In_953,N_19);
and U469 (N_469,In_732,In_247);
or U470 (N_470,N_354,In_666);
and U471 (N_471,In_832,In_843);
nor U472 (N_472,In_778,N_165);
and U473 (N_473,N_333,N_83);
nand U474 (N_474,N_226,In_939);
nor U475 (N_475,In_661,N_53);
nand U476 (N_476,In_671,In_636);
and U477 (N_477,In_123,N_234);
nor U478 (N_478,N_295,N_258);
and U479 (N_479,In_196,In_171);
or U480 (N_480,In_454,In_991);
and U481 (N_481,In_542,N_386);
and U482 (N_482,In_306,In_640);
or U483 (N_483,N_132,In_416);
nand U484 (N_484,In_309,In_685);
or U485 (N_485,In_618,In_151);
or U486 (N_486,In_338,In_93);
xor U487 (N_487,N_257,N_336);
xnor U488 (N_488,N_343,In_924);
nand U489 (N_489,In_539,In_485);
and U490 (N_490,N_177,N_28);
nor U491 (N_491,N_288,N_121);
nand U492 (N_492,N_289,N_243);
nand U493 (N_493,In_343,In_437);
nor U494 (N_494,In_305,In_89);
nor U495 (N_495,In_593,In_794);
and U496 (N_496,In_388,In_555);
nand U497 (N_497,N_365,In_491);
and U498 (N_498,In_17,In_814);
and U499 (N_499,N_278,In_903);
nand U500 (N_500,N_313,N_120);
and U501 (N_501,In_482,N_460);
nand U502 (N_502,N_431,N_414);
nand U503 (N_503,N_325,N_381);
or U504 (N_504,N_317,In_106);
and U505 (N_505,In_682,N_230);
nand U506 (N_506,N_71,In_997);
nor U507 (N_507,N_376,In_193);
nand U508 (N_508,In_417,N_345);
nand U509 (N_509,In_40,N_412);
and U510 (N_510,In_358,In_263);
nor U511 (N_511,In_315,In_211);
nor U512 (N_512,N_202,N_327);
nor U513 (N_513,In_409,N_463);
nand U514 (N_514,In_155,In_550);
and U515 (N_515,In_197,In_257);
nor U516 (N_516,In_657,N_54);
nor U517 (N_517,In_828,In_590);
nor U518 (N_518,In_101,N_171);
nor U519 (N_519,In_697,N_293);
or U520 (N_520,In_33,In_809);
nand U521 (N_521,In_872,N_413);
nor U522 (N_522,N_127,N_454);
nand U523 (N_523,N_334,N_347);
nand U524 (N_524,In_670,N_335);
nor U525 (N_525,N_449,In_3);
and U526 (N_526,In_921,N_477);
nor U527 (N_527,N_445,N_283);
and U528 (N_528,In_361,N_341);
xnor U529 (N_529,N_404,N_459);
and U530 (N_530,In_127,In_644);
nor U531 (N_531,N_240,In_712);
nor U532 (N_532,N_21,N_87);
or U533 (N_533,N_210,N_31);
nand U534 (N_534,N_428,In_886);
and U535 (N_535,In_420,In_39);
or U536 (N_536,In_457,N_252);
or U537 (N_537,N_205,N_415);
nand U538 (N_538,In_807,N_348);
and U539 (N_539,In_95,In_29);
or U540 (N_540,In_14,In_267);
nand U541 (N_541,In_43,In_143);
and U542 (N_542,N_130,N_478);
nand U543 (N_543,N_383,In_528);
xor U544 (N_544,In_8,N_473);
nand U545 (N_545,N_405,N_201);
xnor U546 (N_546,N_305,In_893);
and U547 (N_547,N_263,N_485);
or U548 (N_548,N_350,In_207);
nand U549 (N_549,N_368,N_218);
nand U550 (N_550,In_5,In_941);
or U551 (N_551,In_669,In_38);
nand U552 (N_552,In_142,In_728);
or U553 (N_553,N_292,N_397);
or U554 (N_554,N_464,In_993);
and U555 (N_555,In_145,N_211);
nand U556 (N_556,N_493,In_254);
or U557 (N_557,N_155,N_380);
nand U558 (N_558,N_393,In_10);
nand U559 (N_559,In_655,In_190);
and U560 (N_560,N_200,N_467);
or U561 (N_561,In_168,N_145);
and U562 (N_562,In_988,In_718);
nor U563 (N_563,In_861,In_588);
and U564 (N_564,N_223,In_58);
or U565 (N_565,N_56,In_875);
nand U566 (N_566,In_693,In_912);
nor U567 (N_567,N_402,In_583);
nand U568 (N_568,N_483,N_322);
or U569 (N_569,In_206,N_382);
and U570 (N_570,In_499,N_375);
and U571 (N_571,N_312,In_465);
xnor U572 (N_572,In_467,N_469);
nor U573 (N_573,N_10,In_703);
and U574 (N_574,N_439,In_415);
nand U575 (N_575,In_328,In_424);
xnor U576 (N_576,N_173,In_944);
or U577 (N_577,N_311,In_707);
xnor U578 (N_578,In_954,N_109);
or U579 (N_579,N_324,N_489);
xor U580 (N_580,N_392,N_487);
nand U581 (N_581,In_154,In_626);
nand U582 (N_582,In_116,N_315);
or U583 (N_583,N_364,In_673);
and U584 (N_584,In_348,N_314);
nand U585 (N_585,In_443,N_129);
and U586 (N_586,In_797,N_255);
and U587 (N_587,N_426,N_224);
nor U588 (N_588,N_23,N_62);
nor U589 (N_589,N_398,N_408);
and U590 (N_590,N_357,N_427);
nand U591 (N_591,N_50,In_186);
nand U592 (N_592,In_185,N_451);
nor U593 (N_593,In_649,In_650);
xor U594 (N_594,In_319,In_884);
nor U595 (N_595,N_273,N_146);
and U596 (N_596,N_162,In_623);
or U597 (N_597,N_250,N_47);
nor U598 (N_598,N_369,N_452);
xnor U599 (N_599,In_372,N_387);
or U600 (N_600,N_528,In_510);
nor U601 (N_601,N_543,In_363);
and U602 (N_602,In_120,In_637);
or U603 (N_603,In_970,In_934);
xnor U604 (N_604,N_497,N_517);
or U605 (N_605,N_541,N_575);
nor U606 (N_606,N_462,N_274);
or U607 (N_607,In_656,In_324);
and U608 (N_608,In_277,N_286);
nand U609 (N_609,N_446,In_392);
and U610 (N_610,In_972,In_7);
or U611 (N_611,N_551,N_438);
nand U612 (N_612,In_696,In_166);
nand U613 (N_613,In_643,N_321);
and U614 (N_614,In_369,In_506);
or U615 (N_615,N_593,N_556);
or U616 (N_616,N_337,In_511);
and U617 (N_617,N_569,In_226);
nand U618 (N_618,N_8,N_384);
xor U619 (N_619,In_298,N_482);
nor U620 (N_620,N_188,N_141);
and U621 (N_621,N_577,N_508);
nor U622 (N_622,In_308,In_773);
and U623 (N_623,N_474,In_783);
and U624 (N_624,In_66,N_421);
or U625 (N_625,N_245,In_105);
nand U626 (N_626,In_827,N_189);
nand U627 (N_627,N_116,N_442);
or U628 (N_628,N_547,In_270);
xor U629 (N_629,N_559,In_864);
nor U630 (N_630,In_805,N_535);
nor U631 (N_631,N_244,In_581);
xnor U632 (N_632,In_62,In_80);
and U633 (N_633,N_531,N_180);
or U634 (N_634,In_642,N_553);
or U635 (N_635,N_391,N_530);
nand U636 (N_636,N_550,N_310);
nand U637 (N_637,In_949,N_308);
nor U638 (N_638,In_507,In_234);
or U639 (N_639,N_307,N_198);
and U640 (N_640,N_479,In_815);
nand U641 (N_641,N_142,N_342);
and U642 (N_642,N_409,N_331);
nand U643 (N_643,N_595,N_481);
nor U644 (N_644,N_434,In_121);
and U645 (N_645,N_444,In_775);
and U646 (N_646,In_52,N_501);
nand U647 (N_647,N_586,N_330);
and U648 (N_648,N_521,N_510);
xor U649 (N_649,In_494,N_468);
nand U650 (N_650,N_500,N_407);
or U651 (N_651,N_353,In_862);
and U652 (N_652,N_490,In_791);
nor U653 (N_653,N_494,N_557);
nor U654 (N_654,N_239,N_588);
or U655 (N_655,In_745,N_503);
or U656 (N_656,N_562,In_779);
nor U657 (N_657,N_576,N_568);
nand U658 (N_658,N_400,N_359);
or U659 (N_659,In_597,In_817);
nand U660 (N_660,In_889,N_456);
nor U661 (N_661,N_536,N_150);
nor U662 (N_662,N_356,N_511);
and U663 (N_663,N_399,N_249);
nand U664 (N_664,N_519,In_628);
or U665 (N_665,N_522,N_329);
and U666 (N_666,N_196,N_340);
nor U667 (N_667,N_385,In_534);
or U668 (N_668,N_100,N_300);
or U669 (N_669,N_268,N_525);
xor U670 (N_670,N_563,N_567);
xor U671 (N_671,N_471,N_598);
and U672 (N_672,N_440,In_621);
and U673 (N_673,N_424,N_580);
or U674 (N_674,N_570,In_662);
or U675 (N_675,N_491,N_394);
nand U676 (N_676,In_342,In_368);
or U677 (N_677,N_296,N_472);
nor U678 (N_678,N_507,In_560);
and U679 (N_679,In_554,In_533);
or U680 (N_680,N_514,N_554);
xor U681 (N_681,N_589,N_309);
or U682 (N_682,N_131,N_74);
and U683 (N_683,N_509,In_913);
nor U684 (N_684,N_219,In_724);
nor U685 (N_685,N_476,N_190);
nor U686 (N_686,N_351,N_578);
xor U687 (N_687,N_443,In_622);
and U688 (N_688,N_492,N_144);
and U689 (N_689,N_355,N_320);
nand U690 (N_690,In_352,N_585);
and U691 (N_691,N_523,In_283);
or U692 (N_692,N_527,N_524);
or U693 (N_693,In_421,In_553);
xor U694 (N_694,N_488,In_895);
and U695 (N_695,N_95,N_480);
or U696 (N_696,N_539,N_579);
nor U697 (N_697,In_740,N_184);
nand U698 (N_698,N_215,N_429);
or U699 (N_699,N_450,In_574);
xor U700 (N_700,In_927,N_448);
or U701 (N_701,In_131,In_985);
and U702 (N_702,N_518,N_558);
or U703 (N_703,N_526,N_520);
nand U704 (N_704,N_5,N_484);
or U705 (N_705,In_747,N_626);
or U706 (N_706,N_649,N_57);
nand U707 (N_707,N_411,N_470);
and U708 (N_708,N_540,N_625);
nor U709 (N_709,N_502,N_181);
nand U710 (N_710,In_295,N_622);
and U711 (N_711,N_689,N_691);
nand U712 (N_712,N_538,N_692);
nand U713 (N_713,In_390,In_576);
nor U714 (N_714,N_214,In_733);
or U715 (N_715,In_51,N_583);
and U716 (N_716,N_654,N_549);
nor U717 (N_717,N_619,N_677);
or U718 (N_718,N_561,In_285);
nor U719 (N_719,N_546,N_242);
nor U720 (N_720,In_450,N_657);
and U721 (N_721,N_86,In_684);
or U722 (N_722,N_378,N_698);
nand U723 (N_723,In_838,N_645);
nor U724 (N_724,N_466,N_552);
and U725 (N_725,N_634,N_613);
xor U726 (N_726,In_124,N_495);
nand U727 (N_727,N_612,N_611);
nand U728 (N_728,N_686,N_632);
xnor U729 (N_729,N_134,N_298);
nor U730 (N_730,N_422,In_945);
or U731 (N_731,In_133,N_581);
nand U732 (N_732,N_461,N_542);
nand U733 (N_733,N_417,In_9);
xnor U734 (N_734,In_976,N_332);
or U735 (N_735,In_692,N_648);
or U736 (N_736,N_208,In_292);
and U737 (N_737,N_419,N_697);
nand U738 (N_738,N_603,N_669);
nor U739 (N_739,N_627,N_587);
nand U740 (N_740,In_303,N_682);
nor U741 (N_741,N_638,In_488);
nand U742 (N_742,N_633,N_694);
or U743 (N_743,N_596,N_652);
nor U744 (N_744,In_761,N_513);
xor U745 (N_745,N_566,In_676);
or U746 (N_746,In_755,In_240);
and U747 (N_747,N_403,N_433);
nand U748 (N_748,N_396,In_846);
or U749 (N_749,N_600,In_771);
and U750 (N_750,N_653,N_465);
nand U751 (N_751,N_673,N_571);
nor U752 (N_752,In_459,N_496);
nand U753 (N_753,N_663,In_599);
nor U754 (N_754,N_545,N_533);
or U755 (N_755,N_233,In_336);
or U756 (N_756,N_447,N_688);
nand U757 (N_757,N_229,In_329);
and U758 (N_758,N_149,In_209);
xnor U759 (N_759,N_277,N_537);
and U760 (N_760,N_685,N_668);
nand U761 (N_761,N_670,N_89);
or U762 (N_762,N_420,In_856);
and U763 (N_763,N_695,N_379);
nor U764 (N_764,N_624,N_287);
or U765 (N_765,In_280,N_660);
nand U766 (N_766,N_582,N_656);
xnor U767 (N_767,In_514,In_983);
or U768 (N_768,In_365,N_534);
nand U769 (N_769,N_591,N_630);
and U770 (N_770,N_597,N_441);
nor U771 (N_771,N_302,N_486);
xor U772 (N_772,N_281,In_900);
xor U773 (N_773,N_498,N_516);
nand U774 (N_774,N_675,N_564);
nand U775 (N_775,N_156,N_436);
xor U776 (N_776,N_101,N_693);
nor U777 (N_777,N_604,N_650);
or U778 (N_778,N_453,N_610);
nor U779 (N_779,N_505,N_573);
xor U780 (N_780,In_810,N_555);
or U781 (N_781,In_400,N_207);
xnor U782 (N_782,N_641,N_608);
nand U783 (N_783,N_609,N_681);
or U784 (N_784,N_687,In_835);
or U785 (N_785,In_92,N_667);
and U786 (N_786,In_607,N_225);
nand U787 (N_787,In_374,N_606);
or U788 (N_788,N_457,N_672);
nor U789 (N_789,N_599,N_362);
nor U790 (N_790,N_602,N_416);
and U791 (N_791,N_615,N_410);
nor U792 (N_792,N_437,N_590);
and U793 (N_793,N_328,N_644);
and U794 (N_794,N_594,N_176);
nand U795 (N_795,N_40,In_521);
nor U796 (N_796,N_548,N_661);
or U797 (N_797,In_474,N_241);
or U798 (N_798,N_601,N_631);
nor U799 (N_799,N_674,In_980);
xor U800 (N_800,In_633,N_713);
nand U801 (N_801,N_623,N_737);
nor U802 (N_802,N_748,N_797);
or U803 (N_803,N_794,N_430);
nor U804 (N_804,In_22,N_758);
nand U805 (N_805,N_757,N_775);
or U806 (N_806,N_679,N_702);
or U807 (N_807,N_607,N_761);
or U808 (N_808,N_684,In_97);
nand U809 (N_809,N_709,N_346);
nand U810 (N_810,N_370,N_734);
nand U811 (N_811,N_706,N_790);
xnor U812 (N_812,N_512,N_719);
nand U813 (N_813,N_584,N_185);
and U814 (N_814,N_728,N_662);
and U815 (N_815,N_791,N_777);
nor U816 (N_816,N_544,N_458);
nand U817 (N_817,In_255,N_741);
and U818 (N_818,N_640,N_744);
nor U819 (N_819,N_730,N_764);
nor U820 (N_820,In_71,N_204);
and U821 (N_821,N_680,N_192);
and U822 (N_822,N_707,N_592);
nor U823 (N_823,N_708,N_701);
or U824 (N_824,N_788,N_770);
nor U825 (N_825,N_755,N_747);
nor U826 (N_826,N_372,N_637);
nor U827 (N_827,N_718,N_781);
nor U828 (N_828,N_795,N_784);
or U829 (N_829,N_799,N_406);
xor U830 (N_830,N_798,N_671);
and U831 (N_831,N_678,N_390);
and U832 (N_832,N_723,N_642);
xnor U833 (N_833,N_789,N_636);
or U834 (N_834,N_729,In_826);
nand U835 (N_835,N_756,N_751);
nor U836 (N_836,N_714,N_727);
xor U837 (N_837,N_664,N_617);
and U838 (N_838,In_504,N_665);
nand U839 (N_839,N_773,N_304);
and U840 (N_840,N_731,N_418);
or U841 (N_841,N_704,In_100);
and U842 (N_842,N_743,N_504);
nand U843 (N_843,N_763,N_720);
nand U844 (N_844,N_532,N_766);
nand U845 (N_845,N_303,N_774);
nand U846 (N_846,N_455,N_110);
nor U847 (N_847,N_724,N_683);
nand U848 (N_848,N_772,N_716);
nand U849 (N_849,N_722,N_696);
nor U850 (N_850,N_786,N_621);
or U851 (N_851,N_776,N_749);
and U852 (N_852,N_628,N_506);
and U853 (N_853,N_401,N_760);
xor U854 (N_854,N_738,N_759);
or U855 (N_855,N_425,N_658);
or U856 (N_856,N_616,In_834);
and U857 (N_857,N_676,N_752);
and U858 (N_858,N_635,N_762);
or U859 (N_859,N_316,N_742);
xnor U860 (N_860,N_629,N_745);
nand U861 (N_861,N_618,N_750);
and U862 (N_862,In_258,N_792);
nor U863 (N_863,N_643,N_574);
nand U864 (N_864,N_515,N_782);
nand U865 (N_865,N_560,N_647);
and U866 (N_866,N_646,N_361);
or U867 (N_867,N_666,N_740);
nand U868 (N_868,N_499,N_785);
nor U869 (N_869,N_778,N_710);
nand U870 (N_870,N_49,N_780);
or U871 (N_871,In_613,In_803);
or U872 (N_872,N_726,N_736);
nor U873 (N_873,N_771,N_793);
nand U874 (N_874,N_717,N_739);
nand U875 (N_875,N_475,N_435);
nor U876 (N_876,N_620,N_699);
nand U877 (N_877,N_768,N_267);
nor U878 (N_878,N_306,N_715);
or U879 (N_879,N_614,N_423);
nand U880 (N_880,N_690,In_472);
or U881 (N_881,N_721,N_529);
and U882 (N_882,In_730,N_765);
nor U883 (N_883,N_572,N_705);
and U884 (N_884,N_753,N_107);
nand U885 (N_885,N_767,N_247);
nor U886 (N_886,N_712,N_796);
and U887 (N_887,N_651,N_779);
or U888 (N_888,N_703,N_659);
and U889 (N_889,N_639,N_700);
nand U890 (N_890,N_128,N_605);
and U891 (N_891,N_783,N_565);
nor U892 (N_892,N_746,N_732);
nor U893 (N_893,N_711,N_787);
nor U894 (N_894,N_366,N_733);
or U895 (N_895,N_84,In_341);
nand U896 (N_896,N_725,N_769);
or U897 (N_897,N_282,N_432);
nor U898 (N_898,N_754,N_735);
or U899 (N_899,N_655,In_407);
or U900 (N_900,N_821,N_884);
xor U901 (N_901,N_852,N_871);
nand U902 (N_902,N_811,N_835);
nor U903 (N_903,N_843,N_814);
or U904 (N_904,N_897,N_822);
and U905 (N_905,N_893,N_807);
nor U906 (N_906,N_818,N_803);
nand U907 (N_907,N_868,N_834);
nor U908 (N_908,N_869,N_805);
xnor U909 (N_909,N_828,N_889);
or U910 (N_910,N_827,N_820);
or U911 (N_911,N_846,N_860);
nand U912 (N_912,N_881,N_882);
nand U913 (N_913,N_837,N_844);
nor U914 (N_914,N_865,N_812);
and U915 (N_915,N_898,N_873);
and U916 (N_916,N_887,N_806);
and U917 (N_917,N_875,N_853);
and U918 (N_918,N_857,N_892);
or U919 (N_919,N_878,N_872);
or U920 (N_920,N_817,N_883);
or U921 (N_921,N_855,N_801);
nor U922 (N_922,N_819,N_867);
and U923 (N_923,N_841,N_829);
and U924 (N_924,N_886,N_816);
nand U925 (N_925,N_856,N_832);
nand U926 (N_926,N_809,N_880);
nand U927 (N_927,N_863,N_833);
nor U928 (N_928,N_862,N_858);
nand U929 (N_929,N_839,N_845);
nand U930 (N_930,N_808,N_890);
nand U931 (N_931,N_888,N_879);
xnor U932 (N_932,N_815,N_877);
and U933 (N_933,N_831,N_836);
nand U934 (N_934,N_825,N_864);
or U935 (N_935,N_851,N_894);
xnor U936 (N_936,N_802,N_859);
or U937 (N_937,N_840,N_899);
or U938 (N_938,N_874,N_838);
and U939 (N_939,N_800,N_830);
xor U940 (N_940,N_826,N_876);
nor U941 (N_941,N_849,N_891);
nand U942 (N_942,N_804,N_810);
nand U943 (N_943,N_870,N_861);
nor U944 (N_944,N_885,N_896);
nand U945 (N_945,N_854,N_866);
nand U946 (N_946,N_895,N_842);
nor U947 (N_947,N_823,N_848);
and U948 (N_948,N_824,N_847);
nor U949 (N_949,N_850,N_813);
and U950 (N_950,N_894,N_872);
nor U951 (N_951,N_879,N_862);
nand U952 (N_952,N_893,N_839);
nand U953 (N_953,N_848,N_878);
and U954 (N_954,N_848,N_816);
and U955 (N_955,N_880,N_866);
nor U956 (N_956,N_803,N_838);
and U957 (N_957,N_898,N_847);
nor U958 (N_958,N_852,N_875);
nand U959 (N_959,N_859,N_813);
or U960 (N_960,N_812,N_803);
nand U961 (N_961,N_800,N_850);
or U962 (N_962,N_895,N_819);
nand U963 (N_963,N_895,N_808);
and U964 (N_964,N_810,N_887);
and U965 (N_965,N_826,N_849);
or U966 (N_966,N_884,N_842);
nand U967 (N_967,N_899,N_872);
and U968 (N_968,N_873,N_827);
nand U969 (N_969,N_895,N_886);
xnor U970 (N_970,N_822,N_885);
and U971 (N_971,N_884,N_815);
nor U972 (N_972,N_811,N_802);
nor U973 (N_973,N_813,N_862);
and U974 (N_974,N_889,N_851);
and U975 (N_975,N_804,N_839);
nand U976 (N_976,N_827,N_818);
and U977 (N_977,N_897,N_828);
and U978 (N_978,N_861,N_809);
and U979 (N_979,N_843,N_895);
and U980 (N_980,N_829,N_849);
nand U981 (N_981,N_818,N_811);
nor U982 (N_982,N_861,N_852);
and U983 (N_983,N_862,N_868);
nand U984 (N_984,N_880,N_842);
xnor U985 (N_985,N_888,N_845);
or U986 (N_986,N_855,N_809);
or U987 (N_987,N_846,N_842);
and U988 (N_988,N_824,N_827);
nand U989 (N_989,N_801,N_816);
nand U990 (N_990,N_865,N_892);
or U991 (N_991,N_878,N_866);
nand U992 (N_992,N_840,N_837);
and U993 (N_993,N_867,N_897);
nor U994 (N_994,N_817,N_891);
or U995 (N_995,N_808,N_882);
nand U996 (N_996,N_866,N_805);
or U997 (N_997,N_824,N_801);
nand U998 (N_998,N_859,N_892);
and U999 (N_999,N_897,N_847);
or U1000 (N_1000,N_919,N_935);
and U1001 (N_1001,N_948,N_941);
nor U1002 (N_1002,N_960,N_977);
and U1003 (N_1003,N_959,N_925);
nor U1004 (N_1004,N_921,N_934);
and U1005 (N_1005,N_988,N_901);
xor U1006 (N_1006,N_932,N_980);
nand U1007 (N_1007,N_916,N_947);
and U1008 (N_1008,N_965,N_931);
or U1009 (N_1009,N_990,N_969);
or U1010 (N_1010,N_930,N_974);
or U1011 (N_1011,N_979,N_910);
and U1012 (N_1012,N_995,N_942);
xor U1013 (N_1013,N_984,N_961);
nor U1014 (N_1014,N_968,N_900);
and U1015 (N_1015,N_983,N_992);
xor U1016 (N_1016,N_972,N_994);
xnor U1017 (N_1017,N_964,N_907);
or U1018 (N_1018,N_993,N_998);
or U1019 (N_1019,N_970,N_943);
nand U1020 (N_1020,N_962,N_952);
nor U1021 (N_1021,N_966,N_963);
nand U1022 (N_1022,N_996,N_967);
nor U1023 (N_1023,N_957,N_986);
nand U1024 (N_1024,N_905,N_955);
nor U1025 (N_1025,N_973,N_913);
and U1026 (N_1026,N_956,N_949);
or U1027 (N_1027,N_953,N_923);
nor U1028 (N_1028,N_971,N_909);
xnor U1029 (N_1029,N_918,N_939);
or U1030 (N_1030,N_999,N_914);
xor U1031 (N_1031,N_920,N_912);
or U1032 (N_1032,N_926,N_904);
nand U1033 (N_1033,N_987,N_997);
and U1034 (N_1034,N_981,N_906);
nand U1035 (N_1035,N_991,N_917);
nand U1036 (N_1036,N_911,N_958);
nor U1037 (N_1037,N_915,N_938);
xor U1038 (N_1038,N_936,N_902);
or U1039 (N_1039,N_922,N_950);
xnor U1040 (N_1040,N_978,N_945);
nand U1041 (N_1041,N_940,N_989);
xor U1042 (N_1042,N_903,N_929);
nor U1043 (N_1043,N_946,N_937);
and U1044 (N_1044,N_954,N_985);
nor U1045 (N_1045,N_975,N_927);
nand U1046 (N_1046,N_976,N_951);
or U1047 (N_1047,N_982,N_924);
and U1048 (N_1048,N_908,N_944);
nor U1049 (N_1049,N_933,N_928);
and U1050 (N_1050,N_905,N_936);
and U1051 (N_1051,N_936,N_993);
nor U1052 (N_1052,N_949,N_997);
nand U1053 (N_1053,N_928,N_916);
xnor U1054 (N_1054,N_980,N_922);
nor U1055 (N_1055,N_992,N_905);
xor U1056 (N_1056,N_938,N_968);
nand U1057 (N_1057,N_965,N_936);
or U1058 (N_1058,N_912,N_944);
or U1059 (N_1059,N_989,N_974);
nor U1060 (N_1060,N_918,N_931);
and U1061 (N_1061,N_974,N_926);
or U1062 (N_1062,N_937,N_976);
or U1063 (N_1063,N_977,N_938);
nor U1064 (N_1064,N_939,N_940);
xor U1065 (N_1065,N_989,N_997);
and U1066 (N_1066,N_959,N_969);
nor U1067 (N_1067,N_930,N_945);
nor U1068 (N_1068,N_906,N_910);
nand U1069 (N_1069,N_939,N_924);
nor U1070 (N_1070,N_966,N_929);
nor U1071 (N_1071,N_960,N_922);
nor U1072 (N_1072,N_916,N_905);
nand U1073 (N_1073,N_962,N_905);
or U1074 (N_1074,N_908,N_905);
and U1075 (N_1075,N_985,N_952);
nand U1076 (N_1076,N_998,N_966);
and U1077 (N_1077,N_982,N_949);
or U1078 (N_1078,N_984,N_978);
nand U1079 (N_1079,N_979,N_976);
or U1080 (N_1080,N_907,N_962);
or U1081 (N_1081,N_934,N_978);
or U1082 (N_1082,N_989,N_921);
or U1083 (N_1083,N_941,N_914);
nor U1084 (N_1084,N_944,N_925);
or U1085 (N_1085,N_908,N_936);
nand U1086 (N_1086,N_969,N_939);
or U1087 (N_1087,N_948,N_939);
or U1088 (N_1088,N_956,N_984);
and U1089 (N_1089,N_906,N_912);
or U1090 (N_1090,N_906,N_937);
or U1091 (N_1091,N_969,N_979);
nor U1092 (N_1092,N_912,N_947);
nor U1093 (N_1093,N_942,N_985);
nand U1094 (N_1094,N_958,N_939);
or U1095 (N_1095,N_994,N_977);
xor U1096 (N_1096,N_910,N_935);
or U1097 (N_1097,N_931,N_954);
and U1098 (N_1098,N_974,N_986);
nor U1099 (N_1099,N_948,N_915);
nand U1100 (N_1100,N_1030,N_1008);
xor U1101 (N_1101,N_1065,N_1076);
or U1102 (N_1102,N_1086,N_1035);
nor U1103 (N_1103,N_1027,N_1012);
and U1104 (N_1104,N_1098,N_1038);
nor U1105 (N_1105,N_1017,N_1049);
or U1106 (N_1106,N_1009,N_1059);
xor U1107 (N_1107,N_1089,N_1062);
nor U1108 (N_1108,N_1056,N_1084);
and U1109 (N_1109,N_1051,N_1010);
nand U1110 (N_1110,N_1071,N_1001);
nand U1111 (N_1111,N_1079,N_1082);
and U1112 (N_1112,N_1075,N_1078);
nand U1113 (N_1113,N_1094,N_1093);
nor U1114 (N_1114,N_1053,N_1020);
and U1115 (N_1115,N_1042,N_1007);
and U1116 (N_1116,N_1097,N_1057);
xnor U1117 (N_1117,N_1045,N_1021);
nand U1118 (N_1118,N_1074,N_1024);
and U1119 (N_1119,N_1083,N_1028);
and U1120 (N_1120,N_1044,N_1011);
nor U1121 (N_1121,N_1014,N_1032);
nor U1122 (N_1122,N_1013,N_1060);
nand U1123 (N_1123,N_1002,N_1066);
or U1124 (N_1124,N_1088,N_1099);
nand U1125 (N_1125,N_1054,N_1064);
nand U1126 (N_1126,N_1046,N_1073);
or U1127 (N_1127,N_1077,N_1063);
nand U1128 (N_1128,N_1095,N_1067);
nor U1129 (N_1129,N_1003,N_1061);
nor U1130 (N_1130,N_1096,N_1031);
xnor U1131 (N_1131,N_1033,N_1040);
nand U1132 (N_1132,N_1068,N_1091);
and U1133 (N_1133,N_1005,N_1050);
xnor U1134 (N_1134,N_1058,N_1090);
nor U1135 (N_1135,N_1023,N_1055);
or U1136 (N_1136,N_1004,N_1052);
nand U1137 (N_1137,N_1087,N_1070);
nand U1138 (N_1138,N_1048,N_1022);
and U1139 (N_1139,N_1043,N_1081);
and U1140 (N_1140,N_1018,N_1025);
and U1141 (N_1141,N_1006,N_1019);
nor U1142 (N_1142,N_1039,N_1085);
or U1143 (N_1143,N_1047,N_1037);
xor U1144 (N_1144,N_1069,N_1080);
or U1145 (N_1145,N_1015,N_1041);
or U1146 (N_1146,N_1029,N_1000);
and U1147 (N_1147,N_1092,N_1034);
xnor U1148 (N_1148,N_1016,N_1072);
nor U1149 (N_1149,N_1026,N_1036);
and U1150 (N_1150,N_1039,N_1021);
nor U1151 (N_1151,N_1002,N_1028);
nand U1152 (N_1152,N_1063,N_1039);
or U1153 (N_1153,N_1071,N_1045);
nor U1154 (N_1154,N_1052,N_1033);
nand U1155 (N_1155,N_1045,N_1092);
or U1156 (N_1156,N_1025,N_1079);
nor U1157 (N_1157,N_1056,N_1082);
and U1158 (N_1158,N_1008,N_1095);
nand U1159 (N_1159,N_1015,N_1092);
and U1160 (N_1160,N_1062,N_1055);
nand U1161 (N_1161,N_1005,N_1000);
or U1162 (N_1162,N_1006,N_1032);
nand U1163 (N_1163,N_1024,N_1053);
nor U1164 (N_1164,N_1011,N_1031);
or U1165 (N_1165,N_1038,N_1022);
or U1166 (N_1166,N_1091,N_1049);
xnor U1167 (N_1167,N_1014,N_1089);
nor U1168 (N_1168,N_1017,N_1062);
nand U1169 (N_1169,N_1016,N_1076);
or U1170 (N_1170,N_1055,N_1059);
or U1171 (N_1171,N_1034,N_1027);
or U1172 (N_1172,N_1010,N_1086);
or U1173 (N_1173,N_1039,N_1081);
or U1174 (N_1174,N_1064,N_1069);
nor U1175 (N_1175,N_1021,N_1097);
nand U1176 (N_1176,N_1087,N_1001);
xnor U1177 (N_1177,N_1066,N_1029);
nor U1178 (N_1178,N_1086,N_1041);
xnor U1179 (N_1179,N_1014,N_1042);
xnor U1180 (N_1180,N_1050,N_1004);
nand U1181 (N_1181,N_1060,N_1087);
nor U1182 (N_1182,N_1007,N_1056);
and U1183 (N_1183,N_1005,N_1059);
nand U1184 (N_1184,N_1044,N_1072);
nor U1185 (N_1185,N_1020,N_1084);
nand U1186 (N_1186,N_1001,N_1053);
nor U1187 (N_1187,N_1003,N_1092);
nand U1188 (N_1188,N_1062,N_1007);
nand U1189 (N_1189,N_1000,N_1017);
nand U1190 (N_1190,N_1014,N_1097);
or U1191 (N_1191,N_1087,N_1019);
nor U1192 (N_1192,N_1039,N_1080);
and U1193 (N_1193,N_1074,N_1055);
or U1194 (N_1194,N_1061,N_1035);
xor U1195 (N_1195,N_1062,N_1015);
xnor U1196 (N_1196,N_1005,N_1061);
xnor U1197 (N_1197,N_1026,N_1033);
nand U1198 (N_1198,N_1015,N_1073);
xnor U1199 (N_1199,N_1041,N_1052);
nor U1200 (N_1200,N_1137,N_1131);
and U1201 (N_1201,N_1162,N_1144);
nand U1202 (N_1202,N_1102,N_1157);
xor U1203 (N_1203,N_1192,N_1114);
nand U1204 (N_1204,N_1152,N_1161);
or U1205 (N_1205,N_1110,N_1125);
nor U1206 (N_1206,N_1181,N_1141);
nor U1207 (N_1207,N_1138,N_1163);
nor U1208 (N_1208,N_1169,N_1197);
nor U1209 (N_1209,N_1118,N_1107);
nor U1210 (N_1210,N_1104,N_1146);
and U1211 (N_1211,N_1120,N_1122);
and U1212 (N_1212,N_1160,N_1196);
or U1213 (N_1213,N_1158,N_1178);
xor U1214 (N_1214,N_1101,N_1124);
nor U1215 (N_1215,N_1147,N_1130);
and U1216 (N_1216,N_1139,N_1119);
or U1217 (N_1217,N_1182,N_1113);
or U1218 (N_1218,N_1167,N_1186);
nand U1219 (N_1219,N_1155,N_1176);
or U1220 (N_1220,N_1126,N_1142);
nor U1221 (N_1221,N_1194,N_1188);
nand U1222 (N_1222,N_1135,N_1154);
nand U1223 (N_1223,N_1173,N_1136);
xnor U1224 (N_1224,N_1150,N_1195);
nand U1225 (N_1225,N_1121,N_1183);
xor U1226 (N_1226,N_1189,N_1184);
nand U1227 (N_1227,N_1174,N_1140);
nand U1228 (N_1228,N_1132,N_1123);
nor U1229 (N_1229,N_1159,N_1199);
nor U1230 (N_1230,N_1166,N_1111);
nor U1231 (N_1231,N_1148,N_1100);
or U1232 (N_1232,N_1145,N_1193);
nor U1233 (N_1233,N_1180,N_1187);
nor U1234 (N_1234,N_1156,N_1117);
nand U1235 (N_1235,N_1143,N_1168);
and U1236 (N_1236,N_1103,N_1175);
or U1237 (N_1237,N_1116,N_1149);
or U1238 (N_1238,N_1106,N_1177);
or U1239 (N_1239,N_1109,N_1134);
xor U1240 (N_1240,N_1127,N_1179);
and U1241 (N_1241,N_1191,N_1185);
nand U1242 (N_1242,N_1128,N_1170);
and U1243 (N_1243,N_1171,N_1164);
and U1244 (N_1244,N_1105,N_1190);
and U1245 (N_1245,N_1115,N_1153);
nand U1246 (N_1246,N_1172,N_1165);
or U1247 (N_1247,N_1151,N_1129);
or U1248 (N_1248,N_1112,N_1198);
nor U1249 (N_1249,N_1108,N_1133);
and U1250 (N_1250,N_1132,N_1106);
nand U1251 (N_1251,N_1196,N_1186);
nand U1252 (N_1252,N_1141,N_1156);
xor U1253 (N_1253,N_1131,N_1178);
or U1254 (N_1254,N_1140,N_1163);
nor U1255 (N_1255,N_1156,N_1149);
nor U1256 (N_1256,N_1197,N_1134);
or U1257 (N_1257,N_1146,N_1181);
or U1258 (N_1258,N_1174,N_1171);
nand U1259 (N_1259,N_1138,N_1179);
and U1260 (N_1260,N_1159,N_1125);
or U1261 (N_1261,N_1131,N_1190);
or U1262 (N_1262,N_1117,N_1115);
nand U1263 (N_1263,N_1102,N_1165);
nor U1264 (N_1264,N_1143,N_1195);
or U1265 (N_1265,N_1125,N_1151);
or U1266 (N_1266,N_1154,N_1127);
or U1267 (N_1267,N_1134,N_1151);
or U1268 (N_1268,N_1133,N_1110);
or U1269 (N_1269,N_1168,N_1174);
nor U1270 (N_1270,N_1155,N_1108);
and U1271 (N_1271,N_1162,N_1113);
nand U1272 (N_1272,N_1170,N_1176);
xnor U1273 (N_1273,N_1156,N_1194);
and U1274 (N_1274,N_1134,N_1112);
nor U1275 (N_1275,N_1109,N_1187);
nor U1276 (N_1276,N_1173,N_1125);
nor U1277 (N_1277,N_1132,N_1133);
nand U1278 (N_1278,N_1188,N_1162);
or U1279 (N_1279,N_1145,N_1142);
nand U1280 (N_1280,N_1147,N_1104);
nand U1281 (N_1281,N_1178,N_1155);
or U1282 (N_1282,N_1170,N_1173);
nand U1283 (N_1283,N_1167,N_1118);
nor U1284 (N_1284,N_1146,N_1165);
or U1285 (N_1285,N_1187,N_1106);
xor U1286 (N_1286,N_1149,N_1150);
and U1287 (N_1287,N_1160,N_1191);
or U1288 (N_1288,N_1183,N_1139);
nand U1289 (N_1289,N_1107,N_1165);
or U1290 (N_1290,N_1178,N_1146);
or U1291 (N_1291,N_1139,N_1174);
nor U1292 (N_1292,N_1105,N_1173);
or U1293 (N_1293,N_1187,N_1181);
or U1294 (N_1294,N_1171,N_1135);
nor U1295 (N_1295,N_1124,N_1126);
or U1296 (N_1296,N_1108,N_1104);
nand U1297 (N_1297,N_1190,N_1128);
nand U1298 (N_1298,N_1146,N_1186);
or U1299 (N_1299,N_1105,N_1103);
and U1300 (N_1300,N_1232,N_1297);
nand U1301 (N_1301,N_1224,N_1216);
and U1302 (N_1302,N_1288,N_1272);
and U1303 (N_1303,N_1226,N_1299);
and U1304 (N_1304,N_1236,N_1286);
nor U1305 (N_1305,N_1238,N_1265);
and U1306 (N_1306,N_1260,N_1240);
and U1307 (N_1307,N_1208,N_1212);
nor U1308 (N_1308,N_1231,N_1263);
nand U1309 (N_1309,N_1283,N_1270);
and U1310 (N_1310,N_1243,N_1278);
nand U1311 (N_1311,N_1284,N_1215);
nand U1312 (N_1312,N_1275,N_1280);
or U1313 (N_1313,N_1201,N_1266);
xor U1314 (N_1314,N_1252,N_1293);
or U1315 (N_1315,N_1214,N_1273);
or U1316 (N_1316,N_1298,N_1217);
and U1317 (N_1317,N_1279,N_1237);
or U1318 (N_1318,N_1250,N_1295);
and U1319 (N_1319,N_1230,N_1229);
nor U1320 (N_1320,N_1251,N_1213);
nand U1321 (N_1321,N_1239,N_1207);
nor U1322 (N_1322,N_1267,N_1228);
and U1323 (N_1323,N_1245,N_1223);
or U1324 (N_1324,N_1248,N_1285);
nor U1325 (N_1325,N_1294,N_1247);
and U1326 (N_1326,N_1204,N_1206);
or U1327 (N_1327,N_1222,N_1233);
and U1328 (N_1328,N_1209,N_1292);
nand U1329 (N_1329,N_1220,N_1210);
or U1330 (N_1330,N_1287,N_1211);
and U1331 (N_1331,N_1244,N_1289);
nand U1332 (N_1332,N_1202,N_1246);
nor U1333 (N_1333,N_1218,N_1254);
xor U1334 (N_1334,N_1281,N_1221);
and U1335 (N_1335,N_1271,N_1277);
nor U1336 (N_1336,N_1268,N_1249);
or U1337 (N_1337,N_1269,N_1225);
xor U1338 (N_1338,N_1296,N_1291);
and U1339 (N_1339,N_1264,N_1242);
or U1340 (N_1340,N_1258,N_1200);
and U1341 (N_1341,N_1235,N_1241);
nand U1342 (N_1342,N_1262,N_1259);
nor U1343 (N_1343,N_1257,N_1255);
and U1344 (N_1344,N_1253,N_1282);
and U1345 (N_1345,N_1276,N_1274);
nor U1346 (N_1346,N_1219,N_1234);
nand U1347 (N_1347,N_1256,N_1205);
nor U1348 (N_1348,N_1203,N_1261);
or U1349 (N_1349,N_1290,N_1227);
nor U1350 (N_1350,N_1273,N_1271);
or U1351 (N_1351,N_1211,N_1291);
xor U1352 (N_1352,N_1201,N_1289);
or U1353 (N_1353,N_1207,N_1274);
xnor U1354 (N_1354,N_1256,N_1276);
nor U1355 (N_1355,N_1227,N_1263);
or U1356 (N_1356,N_1273,N_1208);
nor U1357 (N_1357,N_1285,N_1220);
nor U1358 (N_1358,N_1256,N_1200);
nand U1359 (N_1359,N_1211,N_1255);
or U1360 (N_1360,N_1220,N_1211);
nor U1361 (N_1361,N_1200,N_1231);
nor U1362 (N_1362,N_1292,N_1298);
and U1363 (N_1363,N_1241,N_1207);
and U1364 (N_1364,N_1269,N_1204);
xnor U1365 (N_1365,N_1202,N_1227);
or U1366 (N_1366,N_1253,N_1208);
nor U1367 (N_1367,N_1285,N_1269);
nand U1368 (N_1368,N_1209,N_1241);
or U1369 (N_1369,N_1226,N_1244);
or U1370 (N_1370,N_1221,N_1202);
and U1371 (N_1371,N_1263,N_1235);
nand U1372 (N_1372,N_1279,N_1208);
xnor U1373 (N_1373,N_1224,N_1227);
or U1374 (N_1374,N_1231,N_1258);
nand U1375 (N_1375,N_1218,N_1246);
and U1376 (N_1376,N_1291,N_1247);
nor U1377 (N_1377,N_1275,N_1281);
xnor U1378 (N_1378,N_1248,N_1260);
nor U1379 (N_1379,N_1264,N_1260);
and U1380 (N_1380,N_1265,N_1212);
or U1381 (N_1381,N_1269,N_1233);
nand U1382 (N_1382,N_1270,N_1297);
nor U1383 (N_1383,N_1222,N_1227);
nor U1384 (N_1384,N_1264,N_1224);
nand U1385 (N_1385,N_1272,N_1281);
nor U1386 (N_1386,N_1277,N_1212);
nand U1387 (N_1387,N_1242,N_1229);
nor U1388 (N_1388,N_1251,N_1228);
and U1389 (N_1389,N_1234,N_1283);
xnor U1390 (N_1390,N_1209,N_1277);
nand U1391 (N_1391,N_1237,N_1218);
nor U1392 (N_1392,N_1220,N_1295);
or U1393 (N_1393,N_1251,N_1247);
xor U1394 (N_1394,N_1219,N_1278);
xnor U1395 (N_1395,N_1274,N_1239);
nor U1396 (N_1396,N_1237,N_1204);
nor U1397 (N_1397,N_1252,N_1256);
nor U1398 (N_1398,N_1201,N_1244);
nor U1399 (N_1399,N_1291,N_1288);
or U1400 (N_1400,N_1316,N_1390);
or U1401 (N_1401,N_1342,N_1318);
nand U1402 (N_1402,N_1393,N_1338);
xor U1403 (N_1403,N_1310,N_1352);
nand U1404 (N_1404,N_1351,N_1382);
nor U1405 (N_1405,N_1337,N_1364);
or U1406 (N_1406,N_1388,N_1372);
or U1407 (N_1407,N_1325,N_1391);
nor U1408 (N_1408,N_1341,N_1367);
nand U1409 (N_1409,N_1339,N_1327);
nor U1410 (N_1410,N_1326,N_1347);
and U1411 (N_1411,N_1362,N_1378);
nor U1412 (N_1412,N_1392,N_1356);
and U1413 (N_1413,N_1389,N_1321);
and U1414 (N_1414,N_1331,N_1376);
nand U1415 (N_1415,N_1303,N_1317);
or U1416 (N_1416,N_1377,N_1346);
or U1417 (N_1417,N_1343,N_1366);
and U1418 (N_1418,N_1361,N_1323);
nor U1419 (N_1419,N_1320,N_1330);
or U1420 (N_1420,N_1396,N_1328);
and U1421 (N_1421,N_1334,N_1309);
or U1422 (N_1422,N_1313,N_1332);
nor U1423 (N_1423,N_1302,N_1319);
nand U1424 (N_1424,N_1394,N_1363);
xor U1425 (N_1425,N_1311,N_1322);
and U1426 (N_1426,N_1345,N_1359);
xnor U1427 (N_1427,N_1355,N_1373);
nand U1428 (N_1428,N_1387,N_1375);
nand U1429 (N_1429,N_1384,N_1354);
nor U1430 (N_1430,N_1348,N_1357);
xor U1431 (N_1431,N_1386,N_1370);
xnor U1432 (N_1432,N_1301,N_1314);
nand U1433 (N_1433,N_1312,N_1300);
nor U1434 (N_1434,N_1381,N_1333);
and U1435 (N_1435,N_1383,N_1335);
nand U1436 (N_1436,N_1374,N_1308);
or U1437 (N_1437,N_1350,N_1397);
nor U1438 (N_1438,N_1371,N_1306);
and U1439 (N_1439,N_1380,N_1385);
nor U1440 (N_1440,N_1336,N_1395);
nor U1441 (N_1441,N_1368,N_1353);
and U1442 (N_1442,N_1379,N_1305);
or U1443 (N_1443,N_1307,N_1365);
or U1444 (N_1444,N_1398,N_1329);
nor U1445 (N_1445,N_1315,N_1324);
nor U1446 (N_1446,N_1369,N_1360);
or U1447 (N_1447,N_1349,N_1340);
nand U1448 (N_1448,N_1304,N_1399);
and U1449 (N_1449,N_1344,N_1358);
nor U1450 (N_1450,N_1304,N_1366);
nor U1451 (N_1451,N_1303,N_1391);
nor U1452 (N_1452,N_1395,N_1323);
nor U1453 (N_1453,N_1316,N_1310);
nand U1454 (N_1454,N_1399,N_1366);
xor U1455 (N_1455,N_1399,N_1349);
nand U1456 (N_1456,N_1380,N_1376);
nor U1457 (N_1457,N_1304,N_1335);
nand U1458 (N_1458,N_1339,N_1392);
and U1459 (N_1459,N_1364,N_1389);
and U1460 (N_1460,N_1307,N_1352);
nor U1461 (N_1461,N_1386,N_1319);
nor U1462 (N_1462,N_1343,N_1311);
and U1463 (N_1463,N_1338,N_1387);
and U1464 (N_1464,N_1337,N_1396);
nor U1465 (N_1465,N_1352,N_1328);
or U1466 (N_1466,N_1338,N_1395);
or U1467 (N_1467,N_1359,N_1382);
xnor U1468 (N_1468,N_1336,N_1319);
and U1469 (N_1469,N_1334,N_1364);
nor U1470 (N_1470,N_1331,N_1371);
xnor U1471 (N_1471,N_1350,N_1304);
and U1472 (N_1472,N_1396,N_1342);
nand U1473 (N_1473,N_1332,N_1354);
xnor U1474 (N_1474,N_1369,N_1301);
nand U1475 (N_1475,N_1344,N_1324);
and U1476 (N_1476,N_1313,N_1339);
or U1477 (N_1477,N_1301,N_1367);
or U1478 (N_1478,N_1343,N_1395);
nand U1479 (N_1479,N_1356,N_1326);
nand U1480 (N_1480,N_1355,N_1347);
xnor U1481 (N_1481,N_1371,N_1368);
nand U1482 (N_1482,N_1354,N_1320);
nor U1483 (N_1483,N_1328,N_1315);
or U1484 (N_1484,N_1335,N_1362);
and U1485 (N_1485,N_1302,N_1381);
and U1486 (N_1486,N_1396,N_1364);
or U1487 (N_1487,N_1377,N_1392);
nor U1488 (N_1488,N_1316,N_1377);
nand U1489 (N_1489,N_1321,N_1393);
nor U1490 (N_1490,N_1340,N_1392);
xnor U1491 (N_1491,N_1312,N_1362);
nor U1492 (N_1492,N_1369,N_1377);
nand U1493 (N_1493,N_1319,N_1358);
nor U1494 (N_1494,N_1368,N_1389);
and U1495 (N_1495,N_1326,N_1308);
and U1496 (N_1496,N_1346,N_1345);
nand U1497 (N_1497,N_1343,N_1383);
nand U1498 (N_1498,N_1365,N_1327);
nor U1499 (N_1499,N_1378,N_1305);
and U1500 (N_1500,N_1413,N_1485);
or U1501 (N_1501,N_1416,N_1407);
nand U1502 (N_1502,N_1450,N_1451);
and U1503 (N_1503,N_1441,N_1477);
and U1504 (N_1504,N_1467,N_1435);
or U1505 (N_1505,N_1418,N_1432);
or U1506 (N_1506,N_1404,N_1405);
nand U1507 (N_1507,N_1480,N_1482);
and U1508 (N_1508,N_1411,N_1447);
or U1509 (N_1509,N_1481,N_1440);
nor U1510 (N_1510,N_1491,N_1421);
or U1511 (N_1511,N_1490,N_1452);
and U1512 (N_1512,N_1408,N_1483);
and U1513 (N_1513,N_1436,N_1409);
and U1514 (N_1514,N_1433,N_1493);
and U1515 (N_1515,N_1479,N_1438);
nand U1516 (N_1516,N_1494,N_1406);
nand U1517 (N_1517,N_1496,N_1424);
xor U1518 (N_1518,N_1458,N_1499);
nand U1519 (N_1519,N_1446,N_1464);
nand U1520 (N_1520,N_1484,N_1442);
and U1521 (N_1521,N_1455,N_1417);
xor U1522 (N_1522,N_1437,N_1469);
nor U1523 (N_1523,N_1456,N_1466);
and U1524 (N_1524,N_1401,N_1462);
or U1525 (N_1525,N_1448,N_1453);
nand U1526 (N_1526,N_1486,N_1412);
or U1527 (N_1527,N_1423,N_1495);
nand U1528 (N_1528,N_1402,N_1431);
xor U1529 (N_1529,N_1430,N_1470);
and U1530 (N_1530,N_1465,N_1434);
and U1531 (N_1531,N_1475,N_1410);
nand U1532 (N_1532,N_1445,N_1474);
or U1533 (N_1533,N_1415,N_1403);
and U1534 (N_1534,N_1463,N_1422);
nand U1535 (N_1535,N_1443,N_1428);
and U1536 (N_1536,N_1487,N_1449);
nand U1537 (N_1537,N_1444,N_1439);
nor U1538 (N_1538,N_1457,N_1492);
nand U1539 (N_1539,N_1497,N_1489);
xor U1540 (N_1540,N_1472,N_1429);
or U1541 (N_1541,N_1425,N_1468);
nor U1542 (N_1542,N_1426,N_1488);
xnor U1543 (N_1543,N_1476,N_1454);
xnor U1544 (N_1544,N_1419,N_1420);
nor U1545 (N_1545,N_1414,N_1471);
nor U1546 (N_1546,N_1473,N_1400);
nor U1547 (N_1547,N_1460,N_1427);
or U1548 (N_1548,N_1498,N_1461);
xor U1549 (N_1549,N_1459,N_1478);
or U1550 (N_1550,N_1408,N_1405);
and U1551 (N_1551,N_1452,N_1406);
and U1552 (N_1552,N_1459,N_1468);
nor U1553 (N_1553,N_1413,N_1482);
nand U1554 (N_1554,N_1456,N_1465);
nor U1555 (N_1555,N_1414,N_1450);
and U1556 (N_1556,N_1456,N_1464);
nor U1557 (N_1557,N_1492,N_1493);
nand U1558 (N_1558,N_1404,N_1482);
nor U1559 (N_1559,N_1478,N_1466);
and U1560 (N_1560,N_1499,N_1429);
or U1561 (N_1561,N_1454,N_1401);
and U1562 (N_1562,N_1491,N_1452);
or U1563 (N_1563,N_1435,N_1443);
nor U1564 (N_1564,N_1435,N_1497);
or U1565 (N_1565,N_1488,N_1429);
and U1566 (N_1566,N_1463,N_1472);
and U1567 (N_1567,N_1436,N_1487);
and U1568 (N_1568,N_1492,N_1461);
or U1569 (N_1569,N_1495,N_1478);
and U1570 (N_1570,N_1406,N_1488);
or U1571 (N_1571,N_1456,N_1452);
nor U1572 (N_1572,N_1427,N_1493);
xnor U1573 (N_1573,N_1413,N_1417);
or U1574 (N_1574,N_1424,N_1407);
nor U1575 (N_1575,N_1408,N_1415);
and U1576 (N_1576,N_1423,N_1402);
nor U1577 (N_1577,N_1415,N_1440);
and U1578 (N_1578,N_1441,N_1455);
and U1579 (N_1579,N_1497,N_1436);
or U1580 (N_1580,N_1454,N_1492);
nand U1581 (N_1581,N_1484,N_1463);
nand U1582 (N_1582,N_1416,N_1475);
nor U1583 (N_1583,N_1444,N_1443);
nand U1584 (N_1584,N_1489,N_1438);
nor U1585 (N_1585,N_1490,N_1496);
or U1586 (N_1586,N_1437,N_1420);
or U1587 (N_1587,N_1483,N_1429);
nand U1588 (N_1588,N_1477,N_1423);
or U1589 (N_1589,N_1473,N_1433);
nor U1590 (N_1590,N_1438,N_1493);
or U1591 (N_1591,N_1456,N_1458);
nor U1592 (N_1592,N_1481,N_1430);
nor U1593 (N_1593,N_1409,N_1459);
nand U1594 (N_1594,N_1480,N_1424);
nor U1595 (N_1595,N_1442,N_1473);
nor U1596 (N_1596,N_1411,N_1468);
nand U1597 (N_1597,N_1437,N_1409);
and U1598 (N_1598,N_1425,N_1418);
and U1599 (N_1599,N_1487,N_1413);
nand U1600 (N_1600,N_1591,N_1554);
nor U1601 (N_1601,N_1576,N_1571);
nand U1602 (N_1602,N_1569,N_1579);
nand U1603 (N_1603,N_1529,N_1505);
or U1604 (N_1604,N_1553,N_1548);
nand U1605 (N_1605,N_1557,N_1504);
or U1606 (N_1606,N_1561,N_1560);
nor U1607 (N_1607,N_1530,N_1573);
nand U1608 (N_1608,N_1552,N_1516);
and U1609 (N_1609,N_1590,N_1500);
nor U1610 (N_1610,N_1501,N_1531);
nor U1611 (N_1611,N_1563,N_1517);
or U1612 (N_1612,N_1580,N_1595);
xnor U1613 (N_1613,N_1518,N_1506);
or U1614 (N_1614,N_1533,N_1585);
or U1615 (N_1615,N_1551,N_1593);
nor U1616 (N_1616,N_1578,N_1509);
nand U1617 (N_1617,N_1583,N_1503);
or U1618 (N_1618,N_1574,N_1538);
nor U1619 (N_1619,N_1592,N_1514);
or U1620 (N_1620,N_1555,N_1586);
nor U1621 (N_1621,N_1542,N_1547);
nand U1622 (N_1622,N_1568,N_1577);
nor U1623 (N_1623,N_1526,N_1537);
nand U1624 (N_1624,N_1508,N_1599);
or U1625 (N_1625,N_1594,N_1582);
nor U1626 (N_1626,N_1549,N_1556);
nor U1627 (N_1627,N_1546,N_1507);
or U1628 (N_1628,N_1545,N_1543);
and U1629 (N_1629,N_1598,N_1550);
and U1630 (N_1630,N_1572,N_1567);
or U1631 (N_1631,N_1513,N_1511);
nand U1632 (N_1632,N_1559,N_1521);
xnor U1633 (N_1633,N_1558,N_1589);
and U1634 (N_1634,N_1564,N_1512);
and U1635 (N_1635,N_1566,N_1541);
nand U1636 (N_1636,N_1525,N_1536);
nand U1637 (N_1637,N_1523,N_1539);
nand U1638 (N_1638,N_1588,N_1532);
or U1639 (N_1639,N_1562,N_1534);
nor U1640 (N_1640,N_1584,N_1527);
or U1641 (N_1641,N_1522,N_1519);
nand U1642 (N_1642,N_1520,N_1524);
nor U1643 (N_1643,N_1587,N_1535);
nand U1644 (N_1644,N_1565,N_1510);
nor U1645 (N_1645,N_1596,N_1544);
nand U1646 (N_1646,N_1502,N_1528);
or U1647 (N_1647,N_1575,N_1515);
nor U1648 (N_1648,N_1540,N_1581);
and U1649 (N_1649,N_1597,N_1570);
nand U1650 (N_1650,N_1560,N_1502);
and U1651 (N_1651,N_1597,N_1549);
xor U1652 (N_1652,N_1581,N_1592);
nor U1653 (N_1653,N_1541,N_1546);
nand U1654 (N_1654,N_1530,N_1588);
and U1655 (N_1655,N_1589,N_1534);
xor U1656 (N_1656,N_1594,N_1536);
nor U1657 (N_1657,N_1519,N_1597);
nor U1658 (N_1658,N_1586,N_1544);
and U1659 (N_1659,N_1592,N_1557);
nand U1660 (N_1660,N_1576,N_1593);
or U1661 (N_1661,N_1521,N_1583);
and U1662 (N_1662,N_1547,N_1523);
nand U1663 (N_1663,N_1542,N_1555);
nand U1664 (N_1664,N_1511,N_1510);
nor U1665 (N_1665,N_1543,N_1512);
nor U1666 (N_1666,N_1566,N_1544);
and U1667 (N_1667,N_1570,N_1571);
nand U1668 (N_1668,N_1549,N_1566);
xor U1669 (N_1669,N_1531,N_1537);
or U1670 (N_1670,N_1523,N_1592);
nand U1671 (N_1671,N_1536,N_1592);
or U1672 (N_1672,N_1512,N_1579);
nand U1673 (N_1673,N_1571,N_1573);
or U1674 (N_1674,N_1538,N_1592);
nand U1675 (N_1675,N_1528,N_1521);
nor U1676 (N_1676,N_1597,N_1561);
or U1677 (N_1677,N_1515,N_1538);
or U1678 (N_1678,N_1509,N_1501);
or U1679 (N_1679,N_1590,N_1527);
nand U1680 (N_1680,N_1572,N_1568);
xnor U1681 (N_1681,N_1598,N_1577);
xnor U1682 (N_1682,N_1532,N_1534);
and U1683 (N_1683,N_1514,N_1521);
or U1684 (N_1684,N_1525,N_1557);
nand U1685 (N_1685,N_1516,N_1525);
and U1686 (N_1686,N_1510,N_1591);
and U1687 (N_1687,N_1583,N_1581);
or U1688 (N_1688,N_1526,N_1540);
nand U1689 (N_1689,N_1559,N_1578);
nor U1690 (N_1690,N_1517,N_1599);
and U1691 (N_1691,N_1562,N_1512);
and U1692 (N_1692,N_1521,N_1571);
nand U1693 (N_1693,N_1570,N_1516);
nor U1694 (N_1694,N_1572,N_1578);
or U1695 (N_1695,N_1560,N_1584);
nand U1696 (N_1696,N_1582,N_1513);
nor U1697 (N_1697,N_1500,N_1505);
nand U1698 (N_1698,N_1569,N_1597);
nand U1699 (N_1699,N_1564,N_1525);
or U1700 (N_1700,N_1687,N_1619);
nand U1701 (N_1701,N_1603,N_1672);
nand U1702 (N_1702,N_1606,N_1639);
nand U1703 (N_1703,N_1651,N_1636);
nand U1704 (N_1704,N_1654,N_1690);
or U1705 (N_1705,N_1679,N_1677);
nand U1706 (N_1706,N_1683,N_1634);
or U1707 (N_1707,N_1646,N_1617);
nand U1708 (N_1708,N_1668,N_1608);
and U1709 (N_1709,N_1645,N_1631);
or U1710 (N_1710,N_1680,N_1694);
nand U1711 (N_1711,N_1650,N_1689);
and U1712 (N_1712,N_1691,N_1620);
or U1713 (N_1713,N_1655,N_1616);
nor U1714 (N_1714,N_1660,N_1670);
nand U1715 (N_1715,N_1686,N_1649);
and U1716 (N_1716,N_1662,N_1632);
nor U1717 (N_1717,N_1607,N_1625);
or U1718 (N_1718,N_1613,N_1614);
nor U1719 (N_1719,N_1652,N_1610);
or U1720 (N_1720,N_1669,N_1673);
or U1721 (N_1721,N_1629,N_1653);
nand U1722 (N_1722,N_1656,N_1692);
and U1723 (N_1723,N_1615,N_1600);
nand U1724 (N_1724,N_1644,N_1648);
nand U1725 (N_1725,N_1633,N_1621);
nor U1726 (N_1726,N_1685,N_1623);
and U1727 (N_1727,N_1643,N_1671);
nor U1728 (N_1728,N_1693,N_1627);
or U1729 (N_1729,N_1618,N_1661);
or U1730 (N_1730,N_1602,N_1684);
or U1731 (N_1731,N_1674,N_1605);
nor U1732 (N_1732,N_1647,N_1681);
nand U1733 (N_1733,N_1667,N_1638);
or U1734 (N_1734,N_1698,N_1628);
and U1735 (N_1735,N_1640,N_1696);
or U1736 (N_1736,N_1630,N_1637);
nor U1737 (N_1737,N_1676,N_1675);
nor U1738 (N_1738,N_1678,N_1604);
and U1739 (N_1739,N_1609,N_1665);
or U1740 (N_1740,N_1664,N_1666);
and U1741 (N_1741,N_1699,N_1624);
or U1742 (N_1742,N_1697,N_1601);
nor U1743 (N_1743,N_1641,N_1635);
or U1744 (N_1744,N_1688,N_1642);
or U1745 (N_1745,N_1657,N_1659);
or U1746 (N_1746,N_1611,N_1612);
and U1747 (N_1747,N_1658,N_1695);
nor U1748 (N_1748,N_1682,N_1622);
or U1749 (N_1749,N_1626,N_1663);
and U1750 (N_1750,N_1677,N_1615);
or U1751 (N_1751,N_1612,N_1639);
xor U1752 (N_1752,N_1672,N_1651);
or U1753 (N_1753,N_1666,N_1607);
nor U1754 (N_1754,N_1648,N_1642);
or U1755 (N_1755,N_1627,N_1697);
nand U1756 (N_1756,N_1649,N_1695);
or U1757 (N_1757,N_1695,N_1651);
nand U1758 (N_1758,N_1656,N_1688);
or U1759 (N_1759,N_1660,N_1612);
nor U1760 (N_1760,N_1608,N_1656);
or U1761 (N_1761,N_1663,N_1658);
nor U1762 (N_1762,N_1615,N_1668);
or U1763 (N_1763,N_1672,N_1666);
or U1764 (N_1764,N_1656,N_1617);
or U1765 (N_1765,N_1641,N_1638);
nand U1766 (N_1766,N_1644,N_1693);
or U1767 (N_1767,N_1617,N_1608);
nand U1768 (N_1768,N_1683,N_1695);
nor U1769 (N_1769,N_1651,N_1619);
nand U1770 (N_1770,N_1637,N_1605);
and U1771 (N_1771,N_1622,N_1684);
and U1772 (N_1772,N_1671,N_1621);
or U1773 (N_1773,N_1695,N_1621);
or U1774 (N_1774,N_1608,N_1643);
or U1775 (N_1775,N_1636,N_1641);
nand U1776 (N_1776,N_1680,N_1635);
nand U1777 (N_1777,N_1628,N_1645);
nor U1778 (N_1778,N_1614,N_1638);
nor U1779 (N_1779,N_1653,N_1609);
nor U1780 (N_1780,N_1612,N_1678);
nand U1781 (N_1781,N_1625,N_1693);
or U1782 (N_1782,N_1643,N_1656);
xor U1783 (N_1783,N_1602,N_1625);
and U1784 (N_1784,N_1650,N_1627);
xnor U1785 (N_1785,N_1632,N_1646);
and U1786 (N_1786,N_1621,N_1662);
nand U1787 (N_1787,N_1691,N_1607);
nor U1788 (N_1788,N_1639,N_1647);
nor U1789 (N_1789,N_1662,N_1670);
nand U1790 (N_1790,N_1631,N_1628);
and U1791 (N_1791,N_1666,N_1605);
nand U1792 (N_1792,N_1658,N_1604);
or U1793 (N_1793,N_1692,N_1619);
nand U1794 (N_1794,N_1687,N_1636);
and U1795 (N_1795,N_1675,N_1660);
and U1796 (N_1796,N_1636,N_1613);
and U1797 (N_1797,N_1629,N_1647);
nand U1798 (N_1798,N_1650,N_1659);
nand U1799 (N_1799,N_1619,N_1603);
nor U1800 (N_1800,N_1754,N_1743);
nor U1801 (N_1801,N_1762,N_1747);
or U1802 (N_1802,N_1791,N_1710);
or U1803 (N_1803,N_1775,N_1740);
nand U1804 (N_1804,N_1795,N_1719);
nor U1805 (N_1805,N_1750,N_1727);
or U1806 (N_1806,N_1730,N_1772);
and U1807 (N_1807,N_1767,N_1738);
or U1808 (N_1808,N_1702,N_1739);
nor U1809 (N_1809,N_1703,N_1737);
nor U1810 (N_1810,N_1777,N_1779);
nand U1811 (N_1811,N_1715,N_1735);
nand U1812 (N_1812,N_1780,N_1761);
nor U1813 (N_1813,N_1786,N_1749);
or U1814 (N_1814,N_1793,N_1717);
nand U1815 (N_1815,N_1760,N_1785);
nand U1816 (N_1816,N_1701,N_1764);
nor U1817 (N_1817,N_1763,N_1755);
and U1818 (N_1818,N_1714,N_1778);
and U1819 (N_1819,N_1757,N_1783);
nand U1820 (N_1820,N_1751,N_1742);
or U1821 (N_1821,N_1797,N_1729);
nand U1822 (N_1822,N_1724,N_1713);
or U1823 (N_1823,N_1799,N_1728);
nand U1824 (N_1824,N_1711,N_1771);
nor U1825 (N_1825,N_1752,N_1723);
nand U1826 (N_1826,N_1741,N_1790);
and U1827 (N_1827,N_1781,N_1700);
or U1828 (N_1828,N_1758,N_1712);
and U1829 (N_1829,N_1722,N_1734);
xor U1830 (N_1830,N_1746,N_1748);
and U1831 (N_1831,N_1716,N_1753);
nand U1832 (N_1832,N_1756,N_1725);
nor U1833 (N_1833,N_1705,N_1707);
xor U1834 (N_1834,N_1773,N_1792);
nand U1835 (N_1835,N_1759,N_1789);
or U1836 (N_1836,N_1709,N_1788);
nor U1837 (N_1837,N_1798,N_1721);
and U1838 (N_1838,N_1784,N_1796);
nand U1839 (N_1839,N_1787,N_1706);
and U1840 (N_1840,N_1745,N_1708);
nand U1841 (N_1841,N_1769,N_1765);
and U1842 (N_1842,N_1726,N_1720);
or U1843 (N_1843,N_1733,N_1704);
xnor U1844 (N_1844,N_1770,N_1731);
nor U1845 (N_1845,N_1794,N_1766);
and U1846 (N_1846,N_1768,N_1776);
and U1847 (N_1847,N_1744,N_1718);
nor U1848 (N_1848,N_1736,N_1782);
xnor U1849 (N_1849,N_1732,N_1774);
or U1850 (N_1850,N_1778,N_1728);
or U1851 (N_1851,N_1775,N_1754);
nand U1852 (N_1852,N_1753,N_1766);
xor U1853 (N_1853,N_1763,N_1746);
nor U1854 (N_1854,N_1788,N_1722);
and U1855 (N_1855,N_1764,N_1777);
or U1856 (N_1856,N_1796,N_1706);
nor U1857 (N_1857,N_1782,N_1740);
nor U1858 (N_1858,N_1787,N_1774);
or U1859 (N_1859,N_1727,N_1752);
nand U1860 (N_1860,N_1786,N_1723);
nand U1861 (N_1861,N_1797,N_1763);
and U1862 (N_1862,N_1712,N_1736);
nand U1863 (N_1863,N_1779,N_1712);
or U1864 (N_1864,N_1751,N_1795);
and U1865 (N_1865,N_1769,N_1700);
nor U1866 (N_1866,N_1774,N_1758);
or U1867 (N_1867,N_1732,N_1714);
nor U1868 (N_1868,N_1779,N_1776);
xnor U1869 (N_1869,N_1702,N_1774);
nor U1870 (N_1870,N_1708,N_1752);
nor U1871 (N_1871,N_1739,N_1794);
and U1872 (N_1872,N_1783,N_1730);
nand U1873 (N_1873,N_1767,N_1701);
nor U1874 (N_1874,N_1753,N_1740);
or U1875 (N_1875,N_1754,N_1739);
and U1876 (N_1876,N_1766,N_1723);
and U1877 (N_1877,N_1798,N_1770);
nand U1878 (N_1878,N_1716,N_1738);
xnor U1879 (N_1879,N_1746,N_1773);
or U1880 (N_1880,N_1703,N_1738);
nor U1881 (N_1881,N_1716,N_1780);
nor U1882 (N_1882,N_1795,N_1780);
and U1883 (N_1883,N_1792,N_1783);
and U1884 (N_1884,N_1713,N_1782);
nand U1885 (N_1885,N_1759,N_1724);
nor U1886 (N_1886,N_1740,N_1786);
or U1887 (N_1887,N_1728,N_1724);
xor U1888 (N_1888,N_1724,N_1762);
nor U1889 (N_1889,N_1714,N_1799);
or U1890 (N_1890,N_1758,N_1715);
nand U1891 (N_1891,N_1713,N_1784);
or U1892 (N_1892,N_1749,N_1738);
and U1893 (N_1893,N_1747,N_1717);
nor U1894 (N_1894,N_1714,N_1771);
or U1895 (N_1895,N_1729,N_1734);
nor U1896 (N_1896,N_1733,N_1712);
or U1897 (N_1897,N_1704,N_1753);
nor U1898 (N_1898,N_1796,N_1715);
nand U1899 (N_1899,N_1728,N_1732);
nand U1900 (N_1900,N_1846,N_1851);
or U1901 (N_1901,N_1807,N_1890);
and U1902 (N_1902,N_1873,N_1863);
and U1903 (N_1903,N_1877,N_1837);
and U1904 (N_1904,N_1875,N_1835);
and U1905 (N_1905,N_1819,N_1832);
and U1906 (N_1906,N_1874,N_1827);
nand U1907 (N_1907,N_1880,N_1852);
xor U1908 (N_1908,N_1810,N_1865);
xnor U1909 (N_1909,N_1850,N_1828);
nor U1910 (N_1910,N_1879,N_1858);
and U1911 (N_1911,N_1885,N_1844);
nand U1912 (N_1912,N_1887,N_1840);
nand U1913 (N_1913,N_1894,N_1817);
nor U1914 (N_1914,N_1889,N_1843);
and U1915 (N_1915,N_1859,N_1866);
or U1916 (N_1916,N_1861,N_1898);
nor U1917 (N_1917,N_1871,N_1860);
nand U1918 (N_1918,N_1842,N_1882);
or U1919 (N_1919,N_1811,N_1809);
nor U1920 (N_1920,N_1870,N_1803);
nor U1921 (N_1921,N_1823,N_1814);
and U1922 (N_1922,N_1896,N_1855);
xnor U1923 (N_1923,N_1822,N_1824);
xor U1924 (N_1924,N_1899,N_1820);
and U1925 (N_1925,N_1833,N_1825);
nand U1926 (N_1926,N_1848,N_1826);
and U1927 (N_1927,N_1853,N_1862);
nand U1928 (N_1928,N_1867,N_1872);
nor U1929 (N_1929,N_1805,N_1888);
nor U1930 (N_1930,N_1800,N_1864);
nand U1931 (N_1931,N_1801,N_1808);
nor U1932 (N_1932,N_1804,N_1815);
or U1933 (N_1933,N_1895,N_1836);
nor U1934 (N_1934,N_1816,N_1802);
xnor U1935 (N_1935,N_1829,N_1892);
xnor U1936 (N_1936,N_1838,N_1884);
and U1937 (N_1937,N_1821,N_1886);
nand U1938 (N_1938,N_1806,N_1891);
or U1939 (N_1939,N_1897,N_1868);
nor U1940 (N_1940,N_1878,N_1845);
nor U1941 (N_1941,N_1881,N_1857);
and U1942 (N_1942,N_1876,N_1847);
xor U1943 (N_1943,N_1856,N_1812);
nand U1944 (N_1944,N_1869,N_1839);
and U1945 (N_1945,N_1841,N_1849);
or U1946 (N_1946,N_1883,N_1893);
or U1947 (N_1947,N_1834,N_1813);
nand U1948 (N_1948,N_1830,N_1818);
nand U1949 (N_1949,N_1854,N_1831);
nand U1950 (N_1950,N_1809,N_1838);
nor U1951 (N_1951,N_1843,N_1875);
xnor U1952 (N_1952,N_1847,N_1813);
nor U1953 (N_1953,N_1877,N_1830);
nor U1954 (N_1954,N_1800,N_1849);
xor U1955 (N_1955,N_1846,N_1811);
xor U1956 (N_1956,N_1896,N_1891);
nand U1957 (N_1957,N_1866,N_1891);
nor U1958 (N_1958,N_1881,N_1845);
and U1959 (N_1959,N_1866,N_1868);
xnor U1960 (N_1960,N_1857,N_1808);
or U1961 (N_1961,N_1835,N_1806);
xnor U1962 (N_1962,N_1810,N_1878);
or U1963 (N_1963,N_1868,N_1832);
and U1964 (N_1964,N_1879,N_1836);
and U1965 (N_1965,N_1830,N_1808);
nand U1966 (N_1966,N_1863,N_1886);
nand U1967 (N_1967,N_1805,N_1871);
and U1968 (N_1968,N_1861,N_1850);
nor U1969 (N_1969,N_1893,N_1874);
nand U1970 (N_1970,N_1875,N_1842);
nand U1971 (N_1971,N_1888,N_1873);
nor U1972 (N_1972,N_1866,N_1855);
nand U1973 (N_1973,N_1843,N_1806);
or U1974 (N_1974,N_1834,N_1865);
xnor U1975 (N_1975,N_1882,N_1877);
nor U1976 (N_1976,N_1895,N_1870);
nor U1977 (N_1977,N_1863,N_1809);
nor U1978 (N_1978,N_1855,N_1881);
nand U1979 (N_1979,N_1838,N_1871);
nand U1980 (N_1980,N_1890,N_1832);
or U1981 (N_1981,N_1851,N_1819);
nand U1982 (N_1982,N_1839,N_1865);
and U1983 (N_1983,N_1866,N_1822);
and U1984 (N_1984,N_1826,N_1801);
nor U1985 (N_1985,N_1815,N_1809);
or U1986 (N_1986,N_1877,N_1887);
nor U1987 (N_1987,N_1881,N_1820);
nand U1988 (N_1988,N_1882,N_1853);
xnor U1989 (N_1989,N_1878,N_1818);
and U1990 (N_1990,N_1890,N_1822);
and U1991 (N_1991,N_1853,N_1884);
nand U1992 (N_1992,N_1851,N_1854);
or U1993 (N_1993,N_1824,N_1849);
nor U1994 (N_1994,N_1804,N_1832);
nand U1995 (N_1995,N_1856,N_1832);
or U1996 (N_1996,N_1871,N_1835);
and U1997 (N_1997,N_1804,N_1840);
nor U1998 (N_1998,N_1850,N_1871);
xnor U1999 (N_1999,N_1860,N_1869);
nor U2000 (N_2000,N_1959,N_1983);
or U2001 (N_2001,N_1939,N_1972);
or U2002 (N_2002,N_1994,N_1985);
or U2003 (N_2003,N_1936,N_1931);
nand U2004 (N_2004,N_1919,N_1927);
and U2005 (N_2005,N_1998,N_1904);
nand U2006 (N_2006,N_1925,N_1960);
xnor U2007 (N_2007,N_1981,N_1943);
nor U2008 (N_2008,N_1911,N_1977);
nand U2009 (N_2009,N_1963,N_1918);
nor U2010 (N_2010,N_1995,N_1949);
and U2011 (N_2011,N_1986,N_1988);
nor U2012 (N_2012,N_1954,N_1956);
xor U2013 (N_2013,N_1948,N_1934);
and U2014 (N_2014,N_1958,N_1913);
nand U2015 (N_2015,N_1915,N_1924);
or U2016 (N_2016,N_1908,N_1928);
nand U2017 (N_2017,N_1951,N_1987);
nor U2018 (N_2018,N_1999,N_1974);
nand U2019 (N_2019,N_1905,N_1990);
or U2020 (N_2020,N_1969,N_1976);
or U2021 (N_2021,N_1947,N_1957);
nor U2022 (N_2022,N_1970,N_1978);
or U2023 (N_2023,N_1980,N_1968);
xnor U2024 (N_2024,N_1993,N_1902);
nand U2025 (N_2025,N_1920,N_1965);
or U2026 (N_2026,N_1966,N_1942);
or U2027 (N_2027,N_1991,N_1944);
nand U2028 (N_2028,N_1982,N_1901);
nor U2029 (N_2029,N_1940,N_1929);
or U2030 (N_2030,N_1906,N_1945);
nor U2031 (N_2031,N_1933,N_1967);
nand U2032 (N_2032,N_1932,N_1909);
and U2033 (N_2033,N_1941,N_1910);
nand U2034 (N_2034,N_1926,N_1914);
nand U2035 (N_2035,N_1922,N_1907);
or U2036 (N_2036,N_1973,N_1971);
nor U2037 (N_2037,N_1996,N_1903);
xor U2038 (N_2038,N_1917,N_1950);
nand U2039 (N_2039,N_1979,N_1900);
or U2040 (N_2040,N_1953,N_1992);
and U2041 (N_2041,N_1912,N_1984);
nand U2042 (N_2042,N_1930,N_1997);
nand U2043 (N_2043,N_1975,N_1921);
xor U2044 (N_2044,N_1946,N_1961);
nand U2045 (N_2045,N_1923,N_1952);
nor U2046 (N_2046,N_1964,N_1938);
or U2047 (N_2047,N_1916,N_1989);
xnor U2048 (N_2048,N_1937,N_1962);
xor U2049 (N_2049,N_1955,N_1935);
nand U2050 (N_2050,N_1963,N_1914);
or U2051 (N_2051,N_1909,N_1905);
xor U2052 (N_2052,N_1905,N_1944);
and U2053 (N_2053,N_1930,N_1959);
nor U2054 (N_2054,N_1985,N_1936);
or U2055 (N_2055,N_1977,N_1948);
and U2056 (N_2056,N_1988,N_1910);
nor U2057 (N_2057,N_1946,N_1981);
nand U2058 (N_2058,N_1949,N_1986);
xor U2059 (N_2059,N_1930,N_1979);
and U2060 (N_2060,N_1935,N_1957);
nor U2061 (N_2061,N_1946,N_1901);
or U2062 (N_2062,N_1916,N_1920);
and U2063 (N_2063,N_1962,N_1991);
nor U2064 (N_2064,N_1944,N_1955);
nor U2065 (N_2065,N_1913,N_1928);
and U2066 (N_2066,N_1990,N_1935);
nor U2067 (N_2067,N_1995,N_1900);
or U2068 (N_2068,N_1998,N_1958);
nand U2069 (N_2069,N_1918,N_1924);
or U2070 (N_2070,N_1963,N_1967);
nor U2071 (N_2071,N_1995,N_1985);
nor U2072 (N_2072,N_1929,N_1971);
nor U2073 (N_2073,N_1937,N_1980);
or U2074 (N_2074,N_1988,N_1959);
or U2075 (N_2075,N_1973,N_1996);
nand U2076 (N_2076,N_1901,N_1921);
xnor U2077 (N_2077,N_1963,N_1950);
or U2078 (N_2078,N_1969,N_1989);
nor U2079 (N_2079,N_1947,N_1922);
or U2080 (N_2080,N_1948,N_1939);
nand U2081 (N_2081,N_1975,N_1960);
nor U2082 (N_2082,N_1918,N_1973);
or U2083 (N_2083,N_1980,N_1914);
nand U2084 (N_2084,N_1942,N_1989);
or U2085 (N_2085,N_1929,N_1910);
xnor U2086 (N_2086,N_1917,N_1965);
and U2087 (N_2087,N_1983,N_1966);
or U2088 (N_2088,N_1991,N_1946);
nor U2089 (N_2089,N_1986,N_1913);
nand U2090 (N_2090,N_1963,N_1958);
and U2091 (N_2091,N_1937,N_1955);
nand U2092 (N_2092,N_1939,N_1969);
nor U2093 (N_2093,N_1975,N_1907);
nand U2094 (N_2094,N_1980,N_1955);
and U2095 (N_2095,N_1943,N_1978);
nand U2096 (N_2096,N_1915,N_1912);
nor U2097 (N_2097,N_1919,N_1908);
xnor U2098 (N_2098,N_1908,N_1985);
and U2099 (N_2099,N_1971,N_1957);
xor U2100 (N_2100,N_2085,N_2045);
nor U2101 (N_2101,N_2074,N_2095);
and U2102 (N_2102,N_2010,N_2071);
xnor U2103 (N_2103,N_2082,N_2033);
or U2104 (N_2104,N_2043,N_2064);
nor U2105 (N_2105,N_2072,N_2056);
nor U2106 (N_2106,N_2097,N_2011);
and U2107 (N_2107,N_2069,N_2087);
and U2108 (N_2108,N_2009,N_2005);
nand U2109 (N_2109,N_2031,N_2070);
and U2110 (N_2110,N_2037,N_2057);
nand U2111 (N_2111,N_2025,N_2023);
and U2112 (N_2112,N_2013,N_2049);
and U2113 (N_2113,N_2054,N_2039);
and U2114 (N_2114,N_2008,N_2076);
or U2115 (N_2115,N_2066,N_2090);
and U2116 (N_2116,N_2035,N_2002);
nor U2117 (N_2117,N_2044,N_2040);
xor U2118 (N_2118,N_2047,N_2073);
nand U2119 (N_2119,N_2038,N_2019);
or U2120 (N_2120,N_2065,N_2021);
or U2121 (N_2121,N_2015,N_2012);
and U2122 (N_2122,N_2028,N_2081);
and U2123 (N_2123,N_2006,N_2093);
xor U2124 (N_2124,N_2022,N_2094);
xor U2125 (N_2125,N_2032,N_2079);
nor U2126 (N_2126,N_2061,N_2014);
or U2127 (N_2127,N_2001,N_2000);
nor U2128 (N_2128,N_2003,N_2041);
xor U2129 (N_2129,N_2083,N_2098);
nand U2130 (N_2130,N_2018,N_2067);
nor U2131 (N_2131,N_2016,N_2096);
nand U2132 (N_2132,N_2092,N_2060);
or U2133 (N_2133,N_2075,N_2029);
or U2134 (N_2134,N_2091,N_2046);
nor U2135 (N_2135,N_2080,N_2059);
and U2136 (N_2136,N_2050,N_2020);
and U2137 (N_2137,N_2017,N_2030);
and U2138 (N_2138,N_2099,N_2024);
nor U2139 (N_2139,N_2055,N_2034);
or U2140 (N_2140,N_2027,N_2004);
nand U2141 (N_2141,N_2063,N_2089);
xnor U2142 (N_2142,N_2088,N_2084);
or U2143 (N_2143,N_2042,N_2053);
and U2144 (N_2144,N_2052,N_2051);
nor U2145 (N_2145,N_2086,N_2078);
or U2146 (N_2146,N_2007,N_2058);
and U2147 (N_2147,N_2036,N_2048);
xor U2148 (N_2148,N_2068,N_2077);
nor U2149 (N_2149,N_2062,N_2026);
or U2150 (N_2150,N_2007,N_2073);
or U2151 (N_2151,N_2092,N_2039);
or U2152 (N_2152,N_2054,N_2061);
xor U2153 (N_2153,N_2018,N_2030);
nand U2154 (N_2154,N_2087,N_2054);
nand U2155 (N_2155,N_2037,N_2026);
nand U2156 (N_2156,N_2029,N_2066);
and U2157 (N_2157,N_2080,N_2044);
nor U2158 (N_2158,N_2053,N_2044);
or U2159 (N_2159,N_2081,N_2014);
or U2160 (N_2160,N_2063,N_2040);
nand U2161 (N_2161,N_2018,N_2011);
nand U2162 (N_2162,N_2029,N_2087);
xor U2163 (N_2163,N_2029,N_2051);
or U2164 (N_2164,N_2036,N_2002);
nand U2165 (N_2165,N_2094,N_2017);
nor U2166 (N_2166,N_2054,N_2080);
nand U2167 (N_2167,N_2060,N_2057);
or U2168 (N_2168,N_2077,N_2096);
nand U2169 (N_2169,N_2045,N_2060);
nand U2170 (N_2170,N_2064,N_2075);
and U2171 (N_2171,N_2029,N_2036);
or U2172 (N_2172,N_2001,N_2076);
nand U2173 (N_2173,N_2022,N_2061);
and U2174 (N_2174,N_2058,N_2033);
or U2175 (N_2175,N_2014,N_2021);
xnor U2176 (N_2176,N_2052,N_2059);
nand U2177 (N_2177,N_2003,N_2015);
and U2178 (N_2178,N_2072,N_2079);
or U2179 (N_2179,N_2068,N_2078);
nand U2180 (N_2180,N_2066,N_2053);
nor U2181 (N_2181,N_2012,N_2085);
nor U2182 (N_2182,N_2033,N_2004);
xor U2183 (N_2183,N_2098,N_2013);
nor U2184 (N_2184,N_2082,N_2042);
nand U2185 (N_2185,N_2004,N_2028);
or U2186 (N_2186,N_2020,N_2041);
nor U2187 (N_2187,N_2049,N_2024);
xor U2188 (N_2188,N_2039,N_2006);
nor U2189 (N_2189,N_2009,N_2052);
nand U2190 (N_2190,N_2034,N_2017);
nor U2191 (N_2191,N_2075,N_2069);
nor U2192 (N_2192,N_2040,N_2070);
nand U2193 (N_2193,N_2028,N_2090);
and U2194 (N_2194,N_2080,N_2023);
or U2195 (N_2195,N_2089,N_2037);
and U2196 (N_2196,N_2043,N_2031);
or U2197 (N_2197,N_2036,N_2066);
nand U2198 (N_2198,N_2093,N_2088);
and U2199 (N_2199,N_2014,N_2065);
nor U2200 (N_2200,N_2156,N_2113);
nor U2201 (N_2201,N_2116,N_2131);
or U2202 (N_2202,N_2138,N_2137);
nor U2203 (N_2203,N_2129,N_2177);
nand U2204 (N_2204,N_2141,N_2183);
nand U2205 (N_2205,N_2162,N_2161);
and U2206 (N_2206,N_2186,N_2102);
or U2207 (N_2207,N_2193,N_2174);
nand U2208 (N_2208,N_2139,N_2195);
xnor U2209 (N_2209,N_2172,N_2115);
nor U2210 (N_2210,N_2119,N_2112);
nor U2211 (N_2211,N_2160,N_2198);
or U2212 (N_2212,N_2110,N_2180);
or U2213 (N_2213,N_2151,N_2150);
nor U2214 (N_2214,N_2144,N_2120);
nor U2215 (N_2215,N_2104,N_2179);
or U2216 (N_2216,N_2101,N_2142);
nor U2217 (N_2217,N_2126,N_2192);
nor U2218 (N_2218,N_2128,N_2197);
and U2219 (N_2219,N_2136,N_2103);
nor U2220 (N_2220,N_2149,N_2178);
and U2221 (N_2221,N_2145,N_2134);
nand U2222 (N_2222,N_2148,N_2168);
and U2223 (N_2223,N_2164,N_2130);
and U2224 (N_2224,N_2171,N_2127);
nand U2225 (N_2225,N_2196,N_2158);
nor U2226 (N_2226,N_2143,N_2199);
nand U2227 (N_2227,N_2167,N_2191);
xor U2228 (N_2228,N_2169,N_2163);
or U2229 (N_2229,N_2118,N_2117);
nor U2230 (N_2230,N_2122,N_2182);
and U2231 (N_2231,N_2140,N_2100);
and U2232 (N_2232,N_2157,N_2106);
nand U2233 (N_2233,N_2133,N_2107);
nand U2234 (N_2234,N_2154,N_2108);
or U2235 (N_2235,N_2185,N_2189);
and U2236 (N_2236,N_2155,N_2173);
or U2237 (N_2237,N_2147,N_2109);
xor U2238 (N_2238,N_2146,N_2132);
xor U2239 (N_2239,N_2123,N_2124);
and U2240 (N_2240,N_2114,N_2176);
or U2241 (N_2241,N_2111,N_2105);
or U2242 (N_2242,N_2187,N_2170);
or U2243 (N_2243,N_2184,N_2121);
nor U2244 (N_2244,N_2190,N_2153);
xnor U2245 (N_2245,N_2152,N_2135);
or U2246 (N_2246,N_2166,N_2165);
or U2247 (N_2247,N_2181,N_2194);
nor U2248 (N_2248,N_2188,N_2175);
nor U2249 (N_2249,N_2125,N_2159);
nand U2250 (N_2250,N_2158,N_2135);
nor U2251 (N_2251,N_2136,N_2185);
or U2252 (N_2252,N_2104,N_2162);
nand U2253 (N_2253,N_2123,N_2161);
nand U2254 (N_2254,N_2140,N_2165);
or U2255 (N_2255,N_2184,N_2116);
nor U2256 (N_2256,N_2129,N_2143);
xnor U2257 (N_2257,N_2188,N_2102);
xor U2258 (N_2258,N_2194,N_2151);
or U2259 (N_2259,N_2100,N_2146);
nand U2260 (N_2260,N_2147,N_2131);
nand U2261 (N_2261,N_2160,N_2156);
and U2262 (N_2262,N_2189,N_2180);
and U2263 (N_2263,N_2172,N_2189);
nor U2264 (N_2264,N_2109,N_2151);
and U2265 (N_2265,N_2154,N_2161);
and U2266 (N_2266,N_2153,N_2198);
nor U2267 (N_2267,N_2185,N_2143);
or U2268 (N_2268,N_2183,N_2185);
nor U2269 (N_2269,N_2175,N_2100);
nand U2270 (N_2270,N_2111,N_2110);
and U2271 (N_2271,N_2111,N_2156);
and U2272 (N_2272,N_2191,N_2184);
nor U2273 (N_2273,N_2198,N_2173);
nand U2274 (N_2274,N_2138,N_2147);
nor U2275 (N_2275,N_2149,N_2123);
xor U2276 (N_2276,N_2134,N_2183);
and U2277 (N_2277,N_2165,N_2112);
and U2278 (N_2278,N_2118,N_2114);
nand U2279 (N_2279,N_2171,N_2139);
or U2280 (N_2280,N_2112,N_2181);
and U2281 (N_2281,N_2163,N_2189);
and U2282 (N_2282,N_2103,N_2169);
or U2283 (N_2283,N_2138,N_2142);
and U2284 (N_2284,N_2172,N_2151);
nand U2285 (N_2285,N_2108,N_2125);
nor U2286 (N_2286,N_2196,N_2118);
nor U2287 (N_2287,N_2198,N_2122);
or U2288 (N_2288,N_2190,N_2142);
nor U2289 (N_2289,N_2175,N_2186);
or U2290 (N_2290,N_2129,N_2190);
and U2291 (N_2291,N_2180,N_2167);
and U2292 (N_2292,N_2105,N_2171);
and U2293 (N_2293,N_2138,N_2114);
nor U2294 (N_2294,N_2197,N_2136);
nand U2295 (N_2295,N_2153,N_2138);
nor U2296 (N_2296,N_2181,N_2136);
and U2297 (N_2297,N_2197,N_2102);
nor U2298 (N_2298,N_2128,N_2144);
or U2299 (N_2299,N_2162,N_2152);
nor U2300 (N_2300,N_2204,N_2209);
or U2301 (N_2301,N_2268,N_2235);
or U2302 (N_2302,N_2232,N_2221);
xor U2303 (N_2303,N_2286,N_2203);
and U2304 (N_2304,N_2295,N_2274);
nor U2305 (N_2305,N_2243,N_2256);
nor U2306 (N_2306,N_2292,N_2213);
xnor U2307 (N_2307,N_2251,N_2255);
nand U2308 (N_2308,N_2212,N_2237);
and U2309 (N_2309,N_2219,N_2290);
nand U2310 (N_2310,N_2228,N_2293);
and U2311 (N_2311,N_2201,N_2229);
and U2312 (N_2312,N_2246,N_2210);
nor U2313 (N_2313,N_2298,N_2214);
and U2314 (N_2314,N_2269,N_2260);
nor U2315 (N_2315,N_2283,N_2264);
and U2316 (N_2316,N_2225,N_2288);
nand U2317 (N_2317,N_2216,N_2267);
and U2318 (N_2318,N_2206,N_2249);
nor U2319 (N_2319,N_2270,N_2224);
or U2320 (N_2320,N_2257,N_2220);
nor U2321 (N_2321,N_2223,N_2244);
nand U2322 (N_2322,N_2297,N_2287);
or U2323 (N_2323,N_2245,N_2266);
nand U2324 (N_2324,N_2236,N_2252);
nand U2325 (N_2325,N_2200,N_2233);
xnor U2326 (N_2326,N_2215,N_2231);
and U2327 (N_2327,N_2280,N_2222);
nor U2328 (N_2328,N_2226,N_2272);
nor U2329 (N_2329,N_2211,N_2227);
and U2330 (N_2330,N_2294,N_2230);
nand U2331 (N_2331,N_2207,N_2202);
nor U2332 (N_2332,N_2265,N_2218);
nor U2333 (N_2333,N_2259,N_2234);
nand U2334 (N_2334,N_2238,N_2253);
or U2335 (N_2335,N_2277,N_2258);
nor U2336 (N_2336,N_2271,N_2279);
nand U2337 (N_2337,N_2278,N_2296);
nor U2338 (N_2338,N_2242,N_2273);
xnor U2339 (N_2339,N_2239,N_2240);
and U2340 (N_2340,N_2248,N_2208);
nand U2341 (N_2341,N_2250,N_2275);
or U2342 (N_2342,N_2217,N_2299);
nand U2343 (N_2343,N_2291,N_2261);
xor U2344 (N_2344,N_2276,N_2262);
and U2345 (N_2345,N_2205,N_2247);
or U2346 (N_2346,N_2281,N_2289);
nand U2347 (N_2347,N_2282,N_2241);
or U2348 (N_2348,N_2284,N_2254);
nor U2349 (N_2349,N_2263,N_2285);
nor U2350 (N_2350,N_2251,N_2282);
nor U2351 (N_2351,N_2265,N_2251);
nor U2352 (N_2352,N_2265,N_2230);
and U2353 (N_2353,N_2271,N_2292);
and U2354 (N_2354,N_2255,N_2264);
or U2355 (N_2355,N_2220,N_2214);
xor U2356 (N_2356,N_2227,N_2208);
nor U2357 (N_2357,N_2263,N_2264);
and U2358 (N_2358,N_2257,N_2281);
nand U2359 (N_2359,N_2269,N_2250);
or U2360 (N_2360,N_2235,N_2210);
and U2361 (N_2361,N_2225,N_2268);
nand U2362 (N_2362,N_2265,N_2231);
nand U2363 (N_2363,N_2260,N_2241);
nand U2364 (N_2364,N_2299,N_2249);
and U2365 (N_2365,N_2225,N_2224);
xor U2366 (N_2366,N_2288,N_2249);
nand U2367 (N_2367,N_2206,N_2267);
nor U2368 (N_2368,N_2242,N_2256);
nand U2369 (N_2369,N_2235,N_2248);
or U2370 (N_2370,N_2204,N_2284);
xnor U2371 (N_2371,N_2266,N_2298);
nand U2372 (N_2372,N_2267,N_2268);
and U2373 (N_2373,N_2216,N_2219);
and U2374 (N_2374,N_2271,N_2224);
nand U2375 (N_2375,N_2259,N_2202);
and U2376 (N_2376,N_2264,N_2275);
xnor U2377 (N_2377,N_2296,N_2204);
and U2378 (N_2378,N_2231,N_2288);
nand U2379 (N_2379,N_2264,N_2242);
nor U2380 (N_2380,N_2237,N_2242);
nand U2381 (N_2381,N_2274,N_2297);
and U2382 (N_2382,N_2266,N_2234);
nand U2383 (N_2383,N_2252,N_2270);
nor U2384 (N_2384,N_2259,N_2263);
or U2385 (N_2385,N_2250,N_2233);
and U2386 (N_2386,N_2243,N_2284);
and U2387 (N_2387,N_2258,N_2234);
and U2388 (N_2388,N_2231,N_2216);
and U2389 (N_2389,N_2298,N_2292);
nor U2390 (N_2390,N_2255,N_2202);
or U2391 (N_2391,N_2254,N_2216);
and U2392 (N_2392,N_2207,N_2237);
and U2393 (N_2393,N_2241,N_2221);
and U2394 (N_2394,N_2295,N_2277);
nor U2395 (N_2395,N_2209,N_2242);
or U2396 (N_2396,N_2262,N_2244);
nand U2397 (N_2397,N_2201,N_2239);
and U2398 (N_2398,N_2220,N_2275);
or U2399 (N_2399,N_2254,N_2239);
or U2400 (N_2400,N_2325,N_2310);
nor U2401 (N_2401,N_2324,N_2386);
nor U2402 (N_2402,N_2351,N_2391);
nand U2403 (N_2403,N_2347,N_2397);
nand U2404 (N_2404,N_2329,N_2312);
and U2405 (N_2405,N_2363,N_2335);
and U2406 (N_2406,N_2321,N_2350);
nor U2407 (N_2407,N_2346,N_2328);
nor U2408 (N_2408,N_2374,N_2365);
nand U2409 (N_2409,N_2364,N_2361);
nand U2410 (N_2410,N_2306,N_2339);
and U2411 (N_2411,N_2326,N_2368);
and U2412 (N_2412,N_2341,N_2392);
nor U2413 (N_2413,N_2385,N_2319);
and U2414 (N_2414,N_2332,N_2372);
and U2415 (N_2415,N_2349,N_2311);
nand U2416 (N_2416,N_2384,N_2331);
and U2417 (N_2417,N_2302,N_2333);
nor U2418 (N_2418,N_2334,N_2356);
and U2419 (N_2419,N_2398,N_2303);
nor U2420 (N_2420,N_2399,N_2301);
xnor U2421 (N_2421,N_2393,N_2353);
or U2422 (N_2422,N_2323,N_2344);
nand U2423 (N_2423,N_2387,N_2366);
nand U2424 (N_2424,N_2354,N_2313);
or U2425 (N_2425,N_2300,N_2367);
nand U2426 (N_2426,N_2369,N_2343);
nor U2427 (N_2427,N_2360,N_2394);
nor U2428 (N_2428,N_2304,N_2377);
xor U2429 (N_2429,N_2305,N_2395);
xor U2430 (N_2430,N_2373,N_2314);
and U2431 (N_2431,N_2309,N_2340);
and U2432 (N_2432,N_2342,N_2315);
and U2433 (N_2433,N_2308,N_2316);
nand U2434 (N_2434,N_2337,N_2338);
or U2435 (N_2435,N_2357,N_2388);
xor U2436 (N_2436,N_2322,N_2348);
xnor U2437 (N_2437,N_2376,N_2380);
and U2438 (N_2438,N_2330,N_2336);
xnor U2439 (N_2439,N_2358,N_2327);
nand U2440 (N_2440,N_2379,N_2307);
nor U2441 (N_2441,N_2375,N_2355);
nand U2442 (N_2442,N_2370,N_2318);
nor U2443 (N_2443,N_2382,N_2378);
or U2444 (N_2444,N_2371,N_2396);
nor U2445 (N_2445,N_2390,N_2352);
nor U2446 (N_2446,N_2383,N_2359);
xnor U2447 (N_2447,N_2389,N_2345);
nand U2448 (N_2448,N_2320,N_2381);
nor U2449 (N_2449,N_2317,N_2362);
and U2450 (N_2450,N_2353,N_2367);
or U2451 (N_2451,N_2378,N_2361);
nand U2452 (N_2452,N_2366,N_2357);
nand U2453 (N_2453,N_2392,N_2385);
or U2454 (N_2454,N_2364,N_2389);
nor U2455 (N_2455,N_2349,N_2366);
and U2456 (N_2456,N_2373,N_2308);
nand U2457 (N_2457,N_2373,N_2301);
or U2458 (N_2458,N_2372,N_2373);
nor U2459 (N_2459,N_2359,N_2354);
nor U2460 (N_2460,N_2390,N_2360);
or U2461 (N_2461,N_2376,N_2361);
nand U2462 (N_2462,N_2385,N_2362);
or U2463 (N_2463,N_2366,N_2325);
and U2464 (N_2464,N_2336,N_2327);
nand U2465 (N_2465,N_2354,N_2339);
xnor U2466 (N_2466,N_2312,N_2349);
and U2467 (N_2467,N_2365,N_2391);
and U2468 (N_2468,N_2369,N_2335);
nand U2469 (N_2469,N_2358,N_2387);
or U2470 (N_2470,N_2366,N_2324);
and U2471 (N_2471,N_2379,N_2327);
nand U2472 (N_2472,N_2369,N_2302);
nand U2473 (N_2473,N_2393,N_2344);
nand U2474 (N_2474,N_2386,N_2378);
and U2475 (N_2475,N_2388,N_2309);
nor U2476 (N_2476,N_2390,N_2363);
and U2477 (N_2477,N_2363,N_2365);
xnor U2478 (N_2478,N_2383,N_2363);
or U2479 (N_2479,N_2382,N_2392);
nor U2480 (N_2480,N_2354,N_2390);
nor U2481 (N_2481,N_2356,N_2350);
or U2482 (N_2482,N_2320,N_2394);
nor U2483 (N_2483,N_2391,N_2332);
nor U2484 (N_2484,N_2347,N_2369);
and U2485 (N_2485,N_2361,N_2325);
and U2486 (N_2486,N_2387,N_2354);
and U2487 (N_2487,N_2321,N_2349);
nor U2488 (N_2488,N_2304,N_2367);
xor U2489 (N_2489,N_2324,N_2391);
xor U2490 (N_2490,N_2387,N_2342);
nor U2491 (N_2491,N_2335,N_2394);
nand U2492 (N_2492,N_2379,N_2304);
nor U2493 (N_2493,N_2308,N_2359);
and U2494 (N_2494,N_2369,N_2336);
nand U2495 (N_2495,N_2329,N_2349);
nor U2496 (N_2496,N_2374,N_2325);
xor U2497 (N_2497,N_2388,N_2394);
or U2498 (N_2498,N_2345,N_2348);
xor U2499 (N_2499,N_2335,N_2338);
xnor U2500 (N_2500,N_2497,N_2441);
and U2501 (N_2501,N_2456,N_2427);
nand U2502 (N_2502,N_2410,N_2444);
nor U2503 (N_2503,N_2461,N_2473);
nand U2504 (N_2504,N_2486,N_2459);
and U2505 (N_2505,N_2475,N_2404);
or U2506 (N_2506,N_2478,N_2460);
nand U2507 (N_2507,N_2464,N_2426);
or U2508 (N_2508,N_2436,N_2429);
or U2509 (N_2509,N_2453,N_2403);
nand U2510 (N_2510,N_2412,N_2498);
or U2511 (N_2511,N_2407,N_2472);
nand U2512 (N_2512,N_2458,N_2471);
nor U2513 (N_2513,N_2493,N_2484);
or U2514 (N_2514,N_2420,N_2482);
nor U2515 (N_2515,N_2433,N_2443);
and U2516 (N_2516,N_2476,N_2416);
nand U2517 (N_2517,N_2431,N_2415);
nor U2518 (N_2518,N_2422,N_2445);
or U2519 (N_2519,N_2432,N_2489);
and U2520 (N_2520,N_2468,N_2450);
nand U2521 (N_2521,N_2409,N_2439);
and U2522 (N_2522,N_2469,N_2406);
or U2523 (N_2523,N_2435,N_2417);
and U2524 (N_2524,N_2400,N_2401);
or U2525 (N_2525,N_2425,N_2440);
xor U2526 (N_2526,N_2462,N_2448);
xor U2527 (N_2527,N_2423,N_2499);
or U2528 (N_2528,N_2479,N_2414);
or U2529 (N_2529,N_2496,N_2408);
and U2530 (N_2530,N_2424,N_2491);
and U2531 (N_2531,N_2494,N_2488);
and U2532 (N_2532,N_2428,N_2438);
nor U2533 (N_2533,N_2465,N_2480);
or U2534 (N_2534,N_2467,N_2419);
nand U2535 (N_2535,N_2455,N_2437);
and U2536 (N_2536,N_2446,N_2454);
nor U2537 (N_2537,N_2487,N_2466);
or U2538 (N_2538,N_2457,N_2405);
and U2539 (N_2539,N_2411,N_2495);
nand U2540 (N_2540,N_2483,N_2463);
and U2541 (N_2541,N_2477,N_2492);
and U2542 (N_2542,N_2430,N_2449);
nand U2543 (N_2543,N_2474,N_2481);
or U2544 (N_2544,N_2490,N_2452);
and U2545 (N_2545,N_2413,N_2421);
nor U2546 (N_2546,N_2485,N_2470);
nand U2547 (N_2547,N_2447,N_2402);
and U2548 (N_2548,N_2442,N_2451);
xnor U2549 (N_2549,N_2434,N_2418);
xor U2550 (N_2550,N_2473,N_2400);
xor U2551 (N_2551,N_2437,N_2435);
nand U2552 (N_2552,N_2474,N_2492);
nor U2553 (N_2553,N_2490,N_2436);
or U2554 (N_2554,N_2476,N_2498);
nand U2555 (N_2555,N_2437,N_2413);
nand U2556 (N_2556,N_2441,N_2472);
or U2557 (N_2557,N_2444,N_2405);
nor U2558 (N_2558,N_2446,N_2411);
nand U2559 (N_2559,N_2404,N_2413);
and U2560 (N_2560,N_2462,N_2473);
or U2561 (N_2561,N_2471,N_2413);
or U2562 (N_2562,N_2410,N_2435);
and U2563 (N_2563,N_2452,N_2499);
nand U2564 (N_2564,N_2458,N_2422);
or U2565 (N_2565,N_2475,N_2470);
or U2566 (N_2566,N_2474,N_2450);
nand U2567 (N_2567,N_2437,N_2490);
and U2568 (N_2568,N_2432,N_2487);
nand U2569 (N_2569,N_2455,N_2477);
and U2570 (N_2570,N_2401,N_2499);
and U2571 (N_2571,N_2441,N_2420);
and U2572 (N_2572,N_2477,N_2406);
nor U2573 (N_2573,N_2490,N_2428);
xor U2574 (N_2574,N_2400,N_2427);
xor U2575 (N_2575,N_2402,N_2404);
nor U2576 (N_2576,N_2448,N_2445);
or U2577 (N_2577,N_2476,N_2440);
or U2578 (N_2578,N_2433,N_2422);
xor U2579 (N_2579,N_2457,N_2441);
or U2580 (N_2580,N_2425,N_2406);
nor U2581 (N_2581,N_2475,N_2472);
nor U2582 (N_2582,N_2418,N_2401);
nand U2583 (N_2583,N_2466,N_2470);
nor U2584 (N_2584,N_2405,N_2453);
and U2585 (N_2585,N_2460,N_2458);
nand U2586 (N_2586,N_2485,N_2454);
nand U2587 (N_2587,N_2483,N_2496);
nand U2588 (N_2588,N_2429,N_2464);
or U2589 (N_2589,N_2404,N_2441);
or U2590 (N_2590,N_2400,N_2402);
nor U2591 (N_2591,N_2431,N_2419);
and U2592 (N_2592,N_2497,N_2487);
or U2593 (N_2593,N_2447,N_2469);
nor U2594 (N_2594,N_2453,N_2443);
and U2595 (N_2595,N_2407,N_2431);
nor U2596 (N_2596,N_2421,N_2425);
nand U2597 (N_2597,N_2406,N_2453);
nor U2598 (N_2598,N_2427,N_2495);
and U2599 (N_2599,N_2414,N_2495);
nand U2600 (N_2600,N_2549,N_2525);
or U2601 (N_2601,N_2580,N_2524);
or U2602 (N_2602,N_2581,N_2537);
nand U2603 (N_2603,N_2576,N_2555);
nor U2604 (N_2604,N_2558,N_2539);
nor U2605 (N_2605,N_2535,N_2544);
or U2606 (N_2606,N_2519,N_2565);
and U2607 (N_2607,N_2503,N_2598);
and U2608 (N_2608,N_2512,N_2507);
nor U2609 (N_2609,N_2574,N_2570);
or U2610 (N_2610,N_2522,N_2585);
nand U2611 (N_2611,N_2556,N_2527);
or U2612 (N_2612,N_2528,N_2548);
nor U2613 (N_2613,N_2587,N_2541);
or U2614 (N_2614,N_2530,N_2542);
nor U2615 (N_2615,N_2501,N_2554);
and U2616 (N_2616,N_2567,N_2508);
and U2617 (N_2617,N_2560,N_2563);
or U2618 (N_2618,N_2561,N_2591);
or U2619 (N_2619,N_2599,N_2550);
nor U2620 (N_2620,N_2594,N_2589);
and U2621 (N_2621,N_2551,N_2595);
nor U2622 (N_2622,N_2578,N_2583);
and U2623 (N_2623,N_2505,N_2575);
nand U2624 (N_2624,N_2564,N_2593);
nor U2625 (N_2625,N_2509,N_2513);
or U2626 (N_2626,N_2540,N_2526);
and U2627 (N_2627,N_2579,N_2547);
nor U2628 (N_2628,N_2504,N_2566);
nor U2629 (N_2629,N_2559,N_2586);
or U2630 (N_2630,N_2543,N_2534);
and U2631 (N_2631,N_2506,N_2546);
nor U2632 (N_2632,N_2500,N_2569);
or U2633 (N_2633,N_2518,N_2577);
and U2634 (N_2634,N_2582,N_2517);
nand U2635 (N_2635,N_2572,N_2516);
or U2636 (N_2636,N_2523,N_2562);
nor U2637 (N_2637,N_2515,N_2568);
and U2638 (N_2638,N_2592,N_2553);
nand U2639 (N_2639,N_2597,N_2590);
nand U2640 (N_2640,N_2584,N_2511);
nand U2641 (N_2641,N_2529,N_2510);
nand U2642 (N_2642,N_2588,N_2545);
and U2643 (N_2643,N_2531,N_2514);
or U2644 (N_2644,N_2521,N_2573);
nor U2645 (N_2645,N_2552,N_2520);
xnor U2646 (N_2646,N_2596,N_2538);
nand U2647 (N_2647,N_2532,N_2533);
or U2648 (N_2648,N_2571,N_2536);
nor U2649 (N_2649,N_2502,N_2557);
or U2650 (N_2650,N_2524,N_2552);
or U2651 (N_2651,N_2533,N_2542);
nand U2652 (N_2652,N_2521,N_2511);
nor U2653 (N_2653,N_2552,N_2584);
xor U2654 (N_2654,N_2560,N_2598);
or U2655 (N_2655,N_2583,N_2517);
or U2656 (N_2656,N_2516,N_2566);
nand U2657 (N_2657,N_2541,N_2593);
nor U2658 (N_2658,N_2561,N_2580);
or U2659 (N_2659,N_2506,N_2516);
and U2660 (N_2660,N_2576,N_2505);
nor U2661 (N_2661,N_2542,N_2527);
or U2662 (N_2662,N_2542,N_2508);
and U2663 (N_2663,N_2567,N_2547);
nand U2664 (N_2664,N_2514,N_2576);
or U2665 (N_2665,N_2552,N_2565);
nor U2666 (N_2666,N_2586,N_2539);
and U2667 (N_2667,N_2528,N_2536);
and U2668 (N_2668,N_2541,N_2501);
or U2669 (N_2669,N_2596,N_2543);
or U2670 (N_2670,N_2508,N_2550);
nand U2671 (N_2671,N_2584,N_2555);
and U2672 (N_2672,N_2520,N_2560);
xor U2673 (N_2673,N_2506,N_2567);
nor U2674 (N_2674,N_2592,N_2578);
or U2675 (N_2675,N_2588,N_2569);
xnor U2676 (N_2676,N_2583,N_2597);
nor U2677 (N_2677,N_2581,N_2593);
and U2678 (N_2678,N_2563,N_2514);
or U2679 (N_2679,N_2548,N_2566);
nor U2680 (N_2680,N_2542,N_2506);
nand U2681 (N_2681,N_2599,N_2541);
nor U2682 (N_2682,N_2564,N_2522);
and U2683 (N_2683,N_2504,N_2530);
or U2684 (N_2684,N_2575,N_2585);
and U2685 (N_2685,N_2525,N_2539);
nor U2686 (N_2686,N_2586,N_2587);
and U2687 (N_2687,N_2509,N_2502);
nand U2688 (N_2688,N_2596,N_2561);
nand U2689 (N_2689,N_2537,N_2522);
nand U2690 (N_2690,N_2528,N_2560);
nor U2691 (N_2691,N_2543,N_2573);
nor U2692 (N_2692,N_2504,N_2533);
or U2693 (N_2693,N_2530,N_2553);
nand U2694 (N_2694,N_2524,N_2592);
or U2695 (N_2695,N_2504,N_2568);
xor U2696 (N_2696,N_2500,N_2576);
xnor U2697 (N_2697,N_2590,N_2587);
xor U2698 (N_2698,N_2525,N_2561);
xor U2699 (N_2699,N_2502,N_2538);
and U2700 (N_2700,N_2649,N_2607);
and U2701 (N_2701,N_2686,N_2633);
nand U2702 (N_2702,N_2636,N_2632);
and U2703 (N_2703,N_2670,N_2660);
or U2704 (N_2704,N_2639,N_2616);
or U2705 (N_2705,N_2601,N_2621);
and U2706 (N_2706,N_2662,N_2638);
or U2707 (N_2707,N_2653,N_2658);
or U2708 (N_2708,N_2620,N_2609);
nor U2709 (N_2709,N_2651,N_2613);
nand U2710 (N_2710,N_2685,N_2696);
or U2711 (N_2711,N_2664,N_2684);
nand U2712 (N_2712,N_2640,N_2650);
nor U2713 (N_2713,N_2600,N_2682);
or U2714 (N_2714,N_2626,N_2668);
or U2715 (N_2715,N_2666,N_2643);
nor U2716 (N_2716,N_2665,N_2648);
and U2717 (N_2717,N_2610,N_2687);
or U2718 (N_2718,N_2622,N_2605);
nor U2719 (N_2719,N_2683,N_2669);
nand U2720 (N_2720,N_2630,N_2697);
nor U2721 (N_2721,N_2628,N_2608);
nor U2722 (N_2722,N_2641,N_2617);
and U2723 (N_2723,N_2606,N_2679);
or U2724 (N_2724,N_2681,N_2693);
nand U2725 (N_2725,N_2672,N_2635);
nand U2726 (N_2726,N_2677,N_2642);
nand U2727 (N_2727,N_2629,N_2602);
and U2728 (N_2728,N_2611,N_2623);
nor U2729 (N_2729,N_2699,N_2614);
nand U2730 (N_2730,N_2612,N_2688);
and U2731 (N_2731,N_2675,N_2655);
nand U2732 (N_2732,N_2698,N_2652);
nand U2733 (N_2733,N_2678,N_2618);
or U2734 (N_2734,N_2647,N_2692);
and U2735 (N_2735,N_2627,N_2657);
xnor U2736 (N_2736,N_2695,N_2644);
nand U2737 (N_2737,N_2661,N_2689);
nand U2738 (N_2738,N_2603,N_2680);
or U2739 (N_2739,N_2604,N_2667);
and U2740 (N_2740,N_2631,N_2637);
nor U2741 (N_2741,N_2690,N_2671);
nand U2742 (N_2742,N_2659,N_2615);
and U2743 (N_2743,N_2625,N_2646);
nor U2744 (N_2744,N_2676,N_2645);
and U2745 (N_2745,N_2654,N_2674);
or U2746 (N_2746,N_2656,N_2663);
and U2747 (N_2747,N_2673,N_2694);
or U2748 (N_2748,N_2691,N_2634);
or U2749 (N_2749,N_2624,N_2619);
nand U2750 (N_2750,N_2667,N_2666);
and U2751 (N_2751,N_2671,N_2695);
nor U2752 (N_2752,N_2697,N_2689);
nor U2753 (N_2753,N_2623,N_2674);
and U2754 (N_2754,N_2619,N_2615);
or U2755 (N_2755,N_2647,N_2630);
nor U2756 (N_2756,N_2621,N_2678);
and U2757 (N_2757,N_2695,N_2624);
nand U2758 (N_2758,N_2631,N_2605);
and U2759 (N_2759,N_2666,N_2629);
and U2760 (N_2760,N_2689,N_2654);
nand U2761 (N_2761,N_2620,N_2650);
xor U2762 (N_2762,N_2672,N_2608);
and U2763 (N_2763,N_2682,N_2687);
nor U2764 (N_2764,N_2653,N_2613);
and U2765 (N_2765,N_2674,N_2647);
nand U2766 (N_2766,N_2612,N_2665);
and U2767 (N_2767,N_2695,N_2638);
xnor U2768 (N_2768,N_2604,N_2633);
and U2769 (N_2769,N_2628,N_2605);
nand U2770 (N_2770,N_2646,N_2658);
nand U2771 (N_2771,N_2620,N_2699);
or U2772 (N_2772,N_2676,N_2690);
nand U2773 (N_2773,N_2662,N_2696);
nor U2774 (N_2774,N_2650,N_2657);
or U2775 (N_2775,N_2695,N_2664);
and U2776 (N_2776,N_2655,N_2652);
nand U2777 (N_2777,N_2619,N_2676);
nor U2778 (N_2778,N_2621,N_2631);
or U2779 (N_2779,N_2668,N_2673);
and U2780 (N_2780,N_2615,N_2614);
or U2781 (N_2781,N_2630,N_2623);
and U2782 (N_2782,N_2623,N_2663);
and U2783 (N_2783,N_2685,N_2610);
nor U2784 (N_2784,N_2640,N_2661);
or U2785 (N_2785,N_2658,N_2649);
nor U2786 (N_2786,N_2625,N_2679);
and U2787 (N_2787,N_2662,N_2654);
and U2788 (N_2788,N_2692,N_2674);
nor U2789 (N_2789,N_2661,N_2651);
or U2790 (N_2790,N_2639,N_2623);
nand U2791 (N_2791,N_2654,N_2624);
and U2792 (N_2792,N_2678,N_2622);
nor U2793 (N_2793,N_2688,N_2624);
and U2794 (N_2794,N_2654,N_2602);
nand U2795 (N_2795,N_2662,N_2653);
or U2796 (N_2796,N_2682,N_2697);
nor U2797 (N_2797,N_2636,N_2641);
nand U2798 (N_2798,N_2654,N_2613);
nand U2799 (N_2799,N_2659,N_2622);
or U2800 (N_2800,N_2793,N_2739);
nor U2801 (N_2801,N_2707,N_2760);
nor U2802 (N_2802,N_2790,N_2745);
xor U2803 (N_2803,N_2784,N_2743);
or U2804 (N_2804,N_2729,N_2721);
nand U2805 (N_2805,N_2751,N_2781);
and U2806 (N_2806,N_2747,N_2722);
nand U2807 (N_2807,N_2737,N_2772);
nor U2808 (N_2808,N_2779,N_2746);
and U2809 (N_2809,N_2771,N_2720);
or U2810 (N_2810,N_2715,N_2768);
nor U2811 (N_2811,N_2712,N_2706);
nand U2812 (N_2812,N_2782,N_2773);
nor U2813 (N_2813,N_2785,N_2718);
nand U2814 (N_2814,N_2769,N_2789);
nor U2815 (N_2815,N_2799,N_2774);
or U2816 (N_2816,N_2758,N_2762);
or U2817 (N_2817,N_2732,N_2792);
nand U2818 (N_2818,N_2701,N_2756);
and U2819 (N_2819,N_2749,N_2703);
or U2820 (N_2820,N_2757,N_2741);
nor U2821 (N_2821,N_2750,N_2778);
or U2822 (N_2822,N_2704,N_2726);
nor U2823 (N_2823,N_2702,N_2730);
nor U2824 (N_2824,N_2740,N_2766);
xnor U2825 (N_2825,N_2763,N_2736);
and U2826 (N_2826,N_2717,N_2744);
nand U2827 (N_2827,N_2752,N_2775);
xor U2828 (N_2828,N_2798,N_2786);
nor U2829 (N_2829,N_2755,N_2791);
and U2830 (N_2830,N_2765,N_2727);
nor U2831 (N_2831,N_2742,N_2770);
nand U2832 (N_2832,N_2795,N_2714);
or U2833 (N_2833,N_2794,N_2767);
nand U2834 (N_2834,N_2748,N_2764);
and U2835 (N_2835,N_2734,N_2724);
nand U2836 (N_2836,N_2733,N_2716);
nor U2837 (N_2837,N_2788,N_2708);
or U2838 (N_2838,N_2759,N_2797);
nor U2839 (N_2839,N_2761,N_2783);
or U2840 (N_2840,N_2753,N_2731);
and U2841 (N_2841,N_2777,N_2780);
and U2842 (N_2842,N_2738,N_2735);
xnor U2843 (N_2843,N_2796,N_2776);
nor U2844 (N_2844,N_2713,N_2709);
or U2845 (N_2845,N_2700,N_2710);
nor U2846 (N_2846,N_2723,N_2787);
or U2847 (N_2847,N_2719,N_2711);
nand U2848 (N_2848,N_2728,N_2754);
xnor U2849 (N_2849,N_2725,N_2705);
nor U2850 (N_2850,N_2710,N_2757);
nor U2851 (N_2851,N_2737,N_2703);
or U2852 (N_2852,N_2709,N_2719);
or U2853 (N_2853,N_2788,N_2794);
and U2854 (N_2854,N_2711,N_2782);
and U2855 (N_2855,N_2766,N_2711);
nand U2856 (N_2856,N_2715,N_2783);
nand U2857 (N_2857,N_2763,N_2705);
nand U2858 (N_2858,N_2729,N_2791);
or U2859 (N_2859,N_2728,N_2772);
nand U2860 (N_2860,N_2725,N_2735);
and U2861 (N_2861,N_2722,N_2748);
xor U2862 (N_2862,N_2701,N_2762);
and U2863 (N_2863,N_2711,N_2715);
or U2864 (N_2864,N_2703,N_2739);
or U2865 (N_2865,N_2717,N_2735);
nor U2866 (N_2866,N_2787,N_2740);
or U2867 (N_2867,N_2760,N_2718);
or U2868 (N_2868,N_2733,N_2732);
nor U2869 (N_2869,N_2772,N_2700);
or U2870 (N_2870,N_2798,N_2721);
nand U2871 (N_2871,N_2790,N_2798);
nor U2872 (N_2872,N_2762,N_2725);
nand U2873 (N_2873,N_2719,N_2743);
xor U2874 (N_2874,N_2757,N_2797);
and U2875 (N_2875,N_2786,N_2737);
or U2876 (N_2876,N_2780,N_2776);
or U2877 (N_2877,N_2745,N_2752);
nor U2878 (N_2878,N_2739,N_2758);
nand U2879 (N_2879,N_2750,N_2732);
or U2880 (N_2880,N_2796,N_2791);
xnor U2881 (N_2881,N_2770,N_2797);
and U2882 (N_2882,N_2754,N_2726);
and U2883 (N_2883,N_2772,N_2769);
and U2884 (N_2884,N_2732,N_2777);
and U2885 (N_2885,N_2706,N_2717);
nand U2886 (N_2886,N_2741,N_2733);
nand U2887 (N_2887,N_2781,N_2785);
or U2888 (N_2888,N_2701,N_2771);
and U2889 (N_2889,N_2743,N_2715);
xor U2890 (N_2890,N_2773,N_2784);
and U2891 (N_2891,N_2728,N_2799);
or U2892 (N_2892,N_2722,N_2765);
nand U2893 (N_2893,N_2781,N_2708);
xnor U2894 (N_2894,N_2796,N_2732);
or U2895 (N_2895,N_2737,N_2707);
and U2896 (N_2896,N_2709,N_2731);
nand U2897 (N_2897,N_2772,N_2761);
xor U2898 (N_2898,N_2735,N_2782);
and U2899 (N_2899,N_2778,N_2701);
xor U2900 (N_2900,N_2843,N_2832);
nor U2901 (N_2901,N_2873,N_2878);
nor U2902 (N_2902,N_2895,N_2812);
xor U2903 (N_2903,N_2893,N_2825);
or U2904 (N_2904,N_2824,N_2883);
and U2905 (N_2905,N_2861,N_2854);
and U2906 (N_2906,N_2882,N_2879);
or U2907 (N_2907,N_2867,N_2809);
xor U2908 (N_2908,N_2876,N_2885);
and U2909 (N_2909,N_2887,N_2816);
nand U2910 (N_2910,N_2833,N_2871);
nand U2911 (N_2911,N_2891,N_2890);
and U2912 (N_2912,N_2875,N_2815);
nand U2913 (N_2913,N_2850,N_2889);
or U2914 (N_2914,N_2822,N_2829);
nor U2915 (N_2915,N_2813,N_2845);
nor U2916 (N_2916,N_2865,N_2868);
nor U2917 (N_2917,N_2859,N_2872);
and U2918 (N_2918,N_2842,N_2874);
and U2919 (N_2919,N_2877,N_2803);
or U2920 (N_2920,N_2858,N_2852);
xnor U2921 (N_2921,N_2800,N_2827);
nand U2922 (N_2922,N_2804,N_2836);
xor U2923 (N_2923,N_2818,N_2834);
and U2924 (N_2924,N_2863,N_2888);
and U2925 (N_2925,N_2880,N_2892);
or U2926 (N_2926,N_2896,N_2884);
nor U2927 (N_2927,N_2830,N_2805);
nand U2928 (N_2928,N_2839,N_2886);
nor U2929 (N_2929,N_2819,N_2897);
nand U2930 (N_2930,N_2841,N_2828);
nor U2931 (N_2931,N_2862,N_2807);
or U2932 (N_2932,N_2801,N_2806);
and U2933 (N_2933,N_2853,N_2881);
nand U2934 (N_2934,N_2831,N_2821);
and U2935 (N_2935,N_2802,N_2847);
or U2936 (N_2936,N_2838,N_2810);
nand U2937 (N_2937,N_2894,N_2870);
xor U2938 (N_2938,N_2860,N_2866);
nor U2939 (N_2939,N_2849,N_2899);
nand U2940 (N_2940,N_2835,N_2846);
nor U2941 (N_2941,N_2817,N_2898);
nor U2942 (N_2942,N_2848,N_2820);
xnor U2943 (N_2943,N_2855,N_2826);
nor U2944 (N_2944,N_2840,N_2808);
or U2945 (N_2945,N_2864,N_2837);
and U2946 (N_2946,N_2857,N_2823);
and U2947 (N_2947,N_2844,N_2851);
nor U2948 (N_2948,N_2856,N_2811);
and U2949 (N_2949,N_2869,N_2814);
and U2950 (N_2950,N_2895,N_2807);
nand U2951 (N_2951,N_2886,N_2868);
nor U2952 (N_2952,N_2870,N_2813);
or U2953 (N_2953,N_2879,N_2848);
nor U2954 (N_2954,N_2882,N_2865);
and U2955 (N_2955,N_2837,N_2882);
nor U2956 (N_2956,N_2829,N_2834);
xor U2957 (N_2957,N_2839,N_2833);
and U2958 (N_2958,N_2827,N_2870);
and U2959 (N_2959,N_2834,N_2836);
and U2960 (N_2960,N_2877,N_2836);
and U2961 (N_2961,N_2846,N_2828);
nand U2962 (N_2962,N_2834,N_2854);
and U2963 (N_2963,N_2850,N_2855);
nand U2964 (N_2964,N_2885,N_2872);
nand U2965 (N_2965,N_2807,N_2802);
and U2966 (N_2966,N_2890,N_2804);
nand U2967 (N_2967,N_2831,N_2870);
or U2968 (N_2968,N_2850,N_2843);
xor U2969 (N_2969,N_2829,N_2887);
xnor U2970 (N_2970,N_2877,N_2810);
and U2971 (N_2971,N_2851,N_2893);
and U2972 (N_2972,N_2872,N_2840);
nor U2973 (N_2973,N_2887,N_2881);
and U2974 (N_2974,N_2837,N_2813);
nand U2975 (N_2975,N_2883,N_2819);
nor U2976 (N_2976,N_2825,N_2829);
xor U2977 (N_2977,N_2809,N_2860);
and U2978 (N_2978,N_2803,N_2847);
or U2979 (N_2979,N_2880,N_2830);
and U2980 (N_2980,N_2882,N_2822);
nand U2981 (N_2981,N_2830,N_2835);
nor U2982 (N_2982,N_2803,N_2802);
nor U2983 (N_2983,N_2801,N_2835);
and U2984 (N_2984,N_2892,N_2870);
and U2985 (N_2985,N_2881,N_2856);
nand U2986 (N_2986,N_2885,N_2865);
and U2987 (N_2987,N_2858,N_2810);
xor U2988 (N_2988,N_2868,N_2883);
xor U2989 (N_2989,N_2879,N_2824);
or U2990 (N_2990,N_2832,N_2801);
or U2991 (N_2991,N_2892,N_2808);
nor U2992 (N_2992,N_2885,N_2832);
nand U2993 (N_2993,N_2851,N_2898);
xnor U2994 (N_2994,N_2892,N_2874);
nand U2995 (N_2995,N_2813,N_2823);
and U2996 (N_2996,N_2873,N_2898);
nor U2997 (N_2997,N_2819,N_2804);
nor U2998 (N_2998,N_2867,N_2897);
or U2999 (N_2999,N_2846,N_2881);
nor U3000 (N_3000,N_2976,N_2907);
xor U3001 (N_3001,N_2951,N_2904);
nand U3002 (N_3002,N_2941,N_2975);
and U3003 (N_3003,N_2943,N_2930);
or U3004 (N_3004,N_2966,N_2995);
nand U3005 (N_3005,N_2998,N_2910);
nand U3006 (N_3006,N_2988,N_2921);
nand U3007 (N_3007,N_2900,N_2905);
nor U3008 (N_3008,N_2969,N_2947);
nor U3009 (N_3009,N_2902,N_2985);
and U3010 (N_3010,N_2963,N_2929);
and U3011 (N_3011,N_2979,N_2952);
or U3012 (N_3012,N_2953,N_2964);
or U3013 (N_3013,N_2962,N_2993);
and U3014 (N_3014,N_2997,N_2949);
and U3015 (N_3015,N_2956,N_2954);
nor U3016 (N_3016,N_2984,N_2970);
and U3017 (N_3017,N_2923,N_2914);
nor U3018 (N_3018,N_2926,N_2948);
and U3019 (N_3019,N_2944,N_2917);
or U3020 (N_3020,N_2990,N_2967);
or U3021 (N_3021,N_2940,N_2937);
xnor U3022 (N_3022,N_2942,N_2992);
xnor U3023 (N_3023,N_2903,N_2931);
nand U3024 (N_3024,N_2945,N_2974);
xor U3025 (N_3025,N_2996,N_2922);
nand U3026 (N_3026,N_2978,N_2928);
and U3027 (N_3027,N_2906,N_2957);
nand U3028 (N_3028,N_2918,N_2915);
nor U3029 (N_3029,N_2971,N_2920);
nor U3030 (N_3030,N_2908,N_2961);
nor U3031 (N_3031,N_2983,N_2939);
and U3032 (N_3032,N_2913,N_2912);
nand U3033 (N_3033,N_2933,N_2925);
and U3034 (N_3034,N_2959,N_2973);
nand U3035 (N_3035,N_2935,N_2936);
or U3036 (N_3036,N_2968,N_2965);
xor U3037 (N_3037,N_2989,N_2981);
nor U3038 (N_3038,N_2911,N_2916);
nor U3039 (N_3039,N_2924,N_2934);
nor U3040 (N_3040,N_2955,N_2994);
xor U3041 (N_3041,N_2972,N_2932);
nor U3042 (N_3042,N_2938,N_2982);
nand U3043 (N_3043,N_2960,N_2909);
and U3044 (N_3044,N_2901,N_2950);
or U3045 (N_3045,N_2977,N_2987);
nor U3046 (N_3046,N_2999,N_2986);
or U3047 (N_3047,N_2958,N_2980);
nand U3048 (N_3048,N_2946,N_2919);
xor U3049 (N_3049,N_2927,N_2991);
nand U3050 (N_3050,N_2976,N_2922);
and U3051 (N_3051,N_2976,N_2934);
and U3052 (N_3052,N_2922,N_2986);
nand U3053 (N_3053,N_2936,N_2905);
nand U3054 (N_3054,N_2955,N_2968);
xor U3055 (N_3055,N_2946,N_2954);
nand U3056 (N_3056,N_2955,N_2981);
or U3057 (N_3057,N_2906,N_2945);
and U3058 (N_3058,N_2926,N_2942);
and U3059 (N_3059,N_2902,N_2923);
or U3060 (N_3060,N_2999,N_2916);
nor U3061 (N_3061,N_2942,N_2974);
or U3062 (N_3062,N_2930,N_2970);
and U3063 (N_3063,N_2941,N_2942);
nor U3064 (N_3064,N_2970,N_2980);
and U3065 (N_3065,N_2987,N_2928);
or U3066 (N_3066,N_2967,N_2978);
and U3067 (N_3067,N_2991,N_2963);
xor U3068 (N_3068,N_2902,N_2964);
nor U3069 (N_3069,N_2913,N_2924);
or U3070 (N_3070,N_2929,N_2938);
nor U3071 (N_3071,N_2969,N_2953);
and U3072 (N_3072,N_2983,N_2967);
nor U3073 (N_3073,N_2999,N_2918);
or U3074 (N_3074,N_2985,N_2999);
nor U3075 (N_3075,N_2992,N_2999);
nor U3076 (N_3076,N_2994,N_2936);
nand U3077 (N_3077,N_2922,N_2921);
nand U3078 (N_3078,N_2909,N_2975);
or U3079 (N_3079,N_2970,N_2926);
and U3080 (N_3080,N_2958,N_2974);
nor U3081 (N_3081,N_2984,N_2915);
and U3082 (N_3082,N_2954,N_2914);
and U3083 (N_3083,N_2993,N_2991);
or U3084 (N_3084,N_2976,N_2931);
or U3085 (N_3085,N_2979,N_2944);
nor U3086 (N_3086,N_2935,N_2969);
or U3087 (N_3087,N_2905,N_2933);
or U3088 (N_3088,N_2929,N_2960);
or U3089 (N_3089,N_2986,N_2991);
xor U3090 (N_3090,N_2942,N_2903);
and U3091 (N_3091,N_2961,N_2976);
or U3092 (N_3092,N_2973,N_2948);
and U3093 (N_3093,N_2944,N_2905);
nand U3094 (N_3094,N_2938,N_2972);
nand U3095 (N_3095,N_2994,N_2902);
or U3096 (N_3096,N_2932,N_2994);
or U3097 (N_3097,N_2969,N_2971);
xnor U3098 (N_3098,N_2904,N_2942);
and U3099 (N_3099,N_2962,N_2921);
xor U3100 (N_3100,N_3037,N_3085);
nand U3101 (N_3101,N_3020,N_3048);
nand U3102 (N_3102,N_3052,N_3021);
or U3103 (N_3103,N_3007,N_3084);
nand U3104 (N_3104,N_3008,N_3029);
xnor U3105 (N_3105,N_3001,N_3047);
or U3106 (N_3106,N_3097,N_3009);
or U3107 (N_3107,N_3063,N_3003);
nor U3108 (N_3108,N_3077,N_3043);
xnor U3109 (N_3109,N_3050,N_3016);
nand U3110 (N_3110,N_3046,N_3098);
and U3111 (N_3111,N_3053,N_3059);
nor U3112 (N_3112,N_3074,N_3004);
or U3113 (N_3113,N_3011,N_3041);
or U3114 (N_3114,N_3078,N_3006);
and U3115 (N_3115,N_3000,N_3034);
and U3116 (N_3116,N_3094,N_3068);
nand U3117 (N_3117,N_3023,N_3018);
or U3118 (N_3118,N_3012,N_3089);
nand U3119 (N_3119,N_3076,N_3027);
or U3120 (N_3120,N_3035,N_3099);
nand U3121 (N_3121,N_3057,N_3080);
nand U3122 (N_3122,N_3049,N_3025);
nor U3123 (N_3123,N_3070,N_3026);
or U3124 (N_3124,N_3071,N_3036);
nor U3125 (N_3125,N_3073,N_3058);
nor U3126 (N_3126,N_3005,N_3030);
or U3127 (N_3127,N_3038,N_3010);
nor U3128 (N_3128,N_3022,N_3040);
nor U3129 (N_3129,N_3039,N_3013);
nand U3130 (N_3130,N_3095,N_3017);
xor U3131 (N_3131,N_3055,N_3019);
or U3132 (N_3132,N_3014,N_3054);
xnor U3133 (N_3133,N_3086,N_3044);
and U3134 (N_3134,N_3087,N_3091);
nor U3135 (N_3135,N_3079,N_3081);
xor U3136 (N_3136,N_3082,N_3067);
nor U3137 (N_3137,N_3066,N_3093);
or U3138 (N_3138,N_3051,N_3032);
or U3139 (N_3139,N_3065,N_3075);
nand U3140 (N_3140,N_3061,N_3064);
nand U3141 (N_3141,N_3088,N_3069);
xor U3142 (N_3142,N_3072,N_3092);
or U3143 (N_3143,N_3083,N_3033);
and U3144 (N_3144,N_3045,N_3002);
nor U3145 (N_3145,N_3028,N_3042);
and U3146 (N_3146,N_3031,N_3096);
nand U3147 (N_3147,N_3015,N_3090);
and U3148 (N_3148,N_3060,N_3024);
nor U3149 (N_3149,N_3062,N_3056);
nand U3150 (N_3150,N_3073,N_3031);
nor U3151 (N_3151,N_3045,N_3036);
xnor U3152 (N_3152,N_3074,N_3019);
nand U3153 (N_3153,N_3087,N_3096);
and U3154 (N_3154,N_3058,N_3069);
or U3155 (N_3155,N_3050,N_3030);
nor U3156 (N_3156,N_3044,N_3075);
or U3157 (N_3157,N_3049,N_3016);
nand U3158 (N_3158,N_3078,N_3032);
and U3159 (N_3159,N_3031,N_3097);
nand U3160 (N_3160,N_3015,N_3017);
and U3161 (N_3161,N_3097,N_3021);
xor U3162 (N_3162,N_3068,N_3087);
nor U3163 (N_3163,N_3059,N_3036);
nor U3164 (N_3164,N_3057,N_3086);
or U3165 (N_3165,N_3018,N_3084);
or U3166 (N_3166,N_3003,N_3065);
nand U3167 (N_3167,N_3089,N_3032);
or U3168 (N_3168,N_3081,N_3083);
nor U3169 (N_3169,N_3084,N_3063);
nor U3170 (N_3170,N_3032,N_3017);
and U3171 (N_3171,N_3016,N_3003);
xor U3172 (N_3172,N_3074,N_3045);
or U3173 (N_3173,N_3025,N_3040);
or U3174 (N_3174,N_3076,N_3095);
or U3175 (N_3175,N_3025,N_3031);
nor U3176 (N_3176,N_3076,N_3044);
or U3177 (N_3177,N_3045,N_3032);
nand U3178 (N_3178,N_3052,N_3037);
xor U3179 (N_3179,N_3007,N_3031);
or U3180 (N_3180,N_3088,N_3093);
and U3181 (N_3181,N_3041,N_3061);
nor U3182 (N_3182,N_3041,N_3015);
nor U3183 (N_3183,N_3044,N_3079);
nand U3184 (N_3184,N_3076,N_3051);
and U3185 (N_3185,N_3026,N_3095);
or U3186 (N_3186,N_3057,N_3022);
or U3187 (N_3187,N_3005,N_3018);
and U3188 (N_3188,N_3048,N_3085);
nand U3189 (N_3189,N_3078,N_3063);
xor U3190 (N_3190,N_3079,N_3039);
or U3191 (N_3191,N_3003,N_3038);
and U3192 (N_3192,N_3078,N_3070);
and U3193 (N_3193,N_3024,N_3071);
nor U3194 (N_3194,N_3072,N_3079);
nand U3195 (N_3195,N_3008,N_3066);
xor U3196 (N_3196,N_3012,N_3044);
or U3197 (N_3197,N_3015,N_3018);
or U3198 (N_3198,N_3069,N_3046);
or U3199 (N_3199,N_3089,N_3086);
and U3200 (N_3200,N_3146,N_3151);
and U3201 (N_3201,N_3170,N_3101);
and U3202 (N_3202,N_3193,N_3111);
nor U3203 (N_3203,N_3173,N_3153);
xnor U3204 (N_3204,N_3150,N_3115);
xnor U3205 (N_3205,N_3106,N_3103);
and U3206 (N_3206,N_3158,N_3136);
nor U3207 (N_3207,N_3166,N_3129);
and U3208 (N_3208,N_3122,N_3142);
xor U3209 (N_3209,N_3138,N_3184);
nand U3210 (N_3210,N_3143,N_3190);
nor U3211 (N_3211,N_3196,N_3160);
and U3212 (N_3212,N_3172,N_3167);
nand U3213 (N_3213,N_3118,N_3148);
and U3214 (N_3214,N_3189,N_3165);
xor U3215 (N_3215,N_3132,N_3185);
and U3216 (N_3216,N_3171,N_3168);
or U3217 (N_3217,N_3175,N_3145);
or U3218 (N_3218,N_3104,N_3178);
and U3219 (N_3219,N_3179,N_3113);
nor U3220 (N_3220,N_3131,N_3102);
nand U3221 (N_3221,N_3139,N_3187);
or U3222 (N_3222,N_3109,N_3162);
nand U3223 (N_3223,N_3155,N_3110);
or U3224 (N_3224,N_3112,N_3156);
xor U3225 (N_3225,N_3116,N_3174);
nand U3226 (N_3226,N_3117,N_3108);
nand U3227 (N_3227,N_3197,N_3192);
nor U3228 (N_3228,N_3191,N_3147);
and U3229 (N_3229,N_3128,N_3133);
xor U3230 (N_3230,N_3140,N_3164);
and U3231 (N_3231,N_3134,N_3149);
nand U3232 (N_3232,N_3141,N_3126);
nor U3233 (N_3233,N_3195,N_3157);
or U3234 (N_3234,N_3120,N_3198);
and U3235 (N_3235,N_3154,N_3127);
nor U3236 (N_3236,N_3124,N_3137);
nand U3237 (N_3237,N_3199,N_3176);
and U3238 (N_3238,N_3183,N_3188);
nor U3239 (N_3239,N_3177,N_3130);
and U3240 (N_3240,N_3144,N_3105);
nand U3241 (N_3241,N_3125,N_3182);
nor U3242 (N_3242,N_3121,N_3186);
or U3243 (N_3243,N_3100,N_3169);
nand U3244 (N_3244,N_3114,N_3159);
nand U3245 (N_3245,N_3181,N_3180);
nand U3246 (N_3246,N_3123,N_3161);
nor U3247 (N_3247,N_3135,N_3194);
nand U3248 (N_3248,N_3119,N_3152);
or U3249 (N_3249,N_3163,N_3107);
and U3250 (N_3250,N_3112,N_3165);
and U3251 (N_3251,N_3199,N_3105);
and U3252 (N_3252,N_3148,N_3135);
or U3253 (N_3253,N_3182,N_3109);
or U3254 (N_3254,N_3120,N_3121);
nor U3255 (N_3255,N_3172,N_3107);
and U3256 (N_3256,N_3175,N_3195);
nand U3257 (N_3257,N_3135,N_3197);
and U3258 (N_3258,N_3109,N_3194);
or U3259 (N_3259,N_3157,N_3114);
nor U3260 (N_3260,N_3177,N_3174);
and U3261 (N_3261,N_3133,N_3108);
or U3262 (N_3262,N_3135,N_3146);
or U3263 (N_3263,N_3189,N_3141);
nor U3264 (N_3264,N_3106,N_3165);
or U3265 (N_3265,N_3114,N_3149);
nand U3266 (N_3266,N_3123,N_3167);
or U3267 (N_3267,N_3136,N_3110);
or U3268 (N_3268,N_3184,N_3103);
and U3269 (N_3269,N_3100,N_3191);
xor U3270 (N_3270,N_3141,N_3148);
and U3271 (N_3271,N_3176,N_3168);
and U3272 (N_3272,N_3185,N_3169);
and U3273 (N_3273,N_3108,N_3178);
and U3274 (N_3274,N_3118,N_3107);
nand U3275 (N_3275,N_3112,N_3127);
nand U3276 (N_3276,N_3115,N_3162);
xnor U3277 (N_3277,N_3162,N_3148);
nor U3278 (N_3278,N_3101,N_3103);
xor U3279 (N_3279,N_3162,N_3164);
nand U3280 (N_3280,N_3177,N_3188);
nand U3281 (N_3281,N_3173,N_3110);
nand U3282 (N_3282,N_3183,N_3141);
or U3283 (N_3283,N_3160,N_3102);
xnor U3284 (N_3284,N_3153,N_3148);
and U3285 (N_3285,N_3109,N_3134);
and U3286 (N_3286,N_3113,N_3144);
or U3287 (N_3287,N_3189,N_3133);
nor U3288 (N_3288,N_3184,N_3175);
nand U3289 (N_3289,N_3135,N_3168);
nor U3290 (N_3290,N_3100,N_3113);
nor U3291 (N_3291,N_3195,N_3126);
or U3292 (N_3292,N_3107,N_3146);
nand U3293 (N_3293,N_3149,N_3146);
nand U3294 (N_3294,N_3109,N_3181);
nand U3295 (N_3295,N_3193,N_3150);
nand U3296 (N_3296,N_3134,N_3117);
xnor U3297 (N_3297,N_3172,N_3178);
and U3298 (N_3298,N_3113,N_3120);
nand U3299 (N_3299,N_3149,N_3172);
or U3300 (N_3300,N_3268,N_3258);
and U3301 (N_3301,N_3245,N_3271);
nand U3302 (N_3302,N_3216,N_3203);
nor U3303 (N_3303,N_3242,N_3202);
nand U3304 (N_3304,N_3296,N_3207);
nor U3305 (N_3305,N_3251,N_3252);
nand U3306 (N_3306,N_3243,N_3262);
nor U3307 (N_3307,N_3276,N_3297);
or U3308 (N_3308,N_3255,N_3248);
nand U3309 (N_3309,N_3233,N_3261);
or U3310 (N_3310,N_3299,N_3294);
or U3311 (N_3311,N_3201,N_3236);
or U3312 (N_3312,N_3291,N_3244);
or U3313 (N_3313,N_3227,N_3225);
nor U3314 (N_3314,N_3257,N_3238);
or U3315 (N_3315,N_3275,N_3278);
nor U3316 (N_3316,N_3283,N_3265);
nand U3317 (N_3317,N_3247,N_3217);
nand U3318 (N_3318,N_3237,N_3228);
and U3319 (N_3319,N_3208,N_3249);
nor U3320 (N_3320,N_3289,N_3230);
and U3321 (N_3321,N_3209,N_3266);
xor U3322 (N_3322,N_3260,N_3282);
and U3323 (N_3323,N_3293,N_3210);
nor U3324 (N_3324,N_3250,N_3288);
nand U3325 (N_3325,N_3298,N_3239);
nand U3326 (N_3326,N_3264,N_3222);
nand U3327 (N_3327,N_3240,N_3256);
or U3328 (N_3328,N_3223,N_3224);
nor U3329 (N_3329,N_3281,N_3211);
and U3330 (N_3330,N_3254,N_3221);
nor U3331 (N_3331,N_3279,N_3246);
or U3332 (N_3332,N_3290,N_3263);
and U3333 (N_3333,N_3274,N_3295);
and U3334 (N_3334,N_3214,N_3229);
and U3335 (N_3335,N_3213,N_3219);
nor U3336 (N_3336,N_3287,N_3292);
nor U3337 (N_3337,N_3253,N_3205);
and U3338 (N_3338,N_3204,N_3272);
xor U3339 (N_3339,N_3212,N_3269);
or U3340 (N_3340,N_3220,N_3285);
xnor U3341 (N_3341,N_3259,N_3215);
and U3342 (N_3342,N_3267,N_3241);
or U3343 (N_3343,N_3270,N_3232);
nor U3344 (N_3344,N_3273,N_3284);
xor U3345 (N_3345,N_3218,N_3280);
nor U3346 (N_3346,N_3277,N_3231);
nor U3347 (N_3347,N_3206,N_3234);
nand U3348 (N_3348,N_3286,N_3235);
nor U3349 (N_3349,N_3226,N_3200);
nor U3350 (N_3350,N_3215,N_3200);
or U3351 (N_3351,N_3285,N_3299);
nand U3352 (N_3352,N_3228,N_3270);
and U3353 (N_3353,N_3294,N_3214);
and U3354 (N_3354,N_3278,N_3286);
nand U3355 (N_3355,N_3226,N_3289);
nand U3356 (N_3356,N_3278,N_3269);
or U3357 (N_3357,N_3262,N_3297);
and U3358 (N_3358,N_3266,N_3235);
nor U3359 (N_3359,N_3235,N_3267);
or U3360 (N_3360,N_3255,N_3219);
nand U3361 (N_3361,N_3262,N_3229);
nand U3362 (N_3362,N_3261,N_3219);
nor U3363 (N_3363,N_3298,N_3263);
and U3364 (N_3364,N_3201,N_3241);
or U3365 (N_3365,N_3228,N_3251);
nor U3366 (N_3366,N_3286,N_3272);
and U3367 (N_3367,N_3272,N_3297);
and U3368 (N_3368,N_3270,N_3267);
nor U3369 (N_3369,N_3294,N_3202);
and U3370 (N_3370,N_3260,N_3243);
and U3371 (N_3371,N_3215,N_3212);
nor U3372 (N_3372,N_3277,N_3244);
nor U3373 (N_3373,N_3258,N_3272);
or U3374 (N_3374,N_3266,N_3257);
xor U3375 (N_3375,N_3288,N_3242);
nand U3376 (N_3376,N_3215,N_3248);
and U3377 (N_3377,N_3209,N_3277);
and U3378 (N_3378,N_3229,N_3295);
xnor U3379 (N_3379,N_3263,N_3239);
nand U3380 (N_3380,N_3276,N_3273);
nand U3381 (N_3381,N_3230,N_3285);
or U3382 (N_3382,N_3222,N_3290);
and U3383 (N_3383,N_3227,N_3296);
or U3384 (N_3384,N_3271,N_3226);
nand U3385 (N_3385,N_3235,N_3270);
and U3386 (N_3386,N_3256,N_3293);
or U3387 (N_3387,N_3230,N_3295);
nand U3388 (N_3388,N_3259,N_3249);
xor U3389 (N_3389,N_3288,N_3220);
or U3390 (N_3390,N_3235,N_3211);
and U3391 (N_3391,N_3263,N_3219);
and U3392 (N_3392,N_3263,N_3277);
or U3393 (N_3393,N_3206,N_3240);
nor U3394 (N_3394,N_3286,N_3209);
and U3395 (N_3395,N_3208,N_3239);
xor U3396 (N_3396,N_3221,N_3212);
xnor U3397 (N_3397,N_3237,N_3253);
nor U3398 (N_3398,N_3284,N_3212);
and U3399 (N_3399,N_3229,N_3284);
and U3400 (N_3400,N_3345,N_3339);
and U3401 (N_3401,N_3357,N_3330);
and U3402 (N_3402,N_3340,N_3394);
or U3403 (N_3403,N_3337,N_3335);
or U3404 (N_3404,N_3309,N_3397);
nor U3405 (N_3405,N_3388,N_3379);
xor U3406 (N_3406,N_3304,N_3361);
nor U3407 (N_3407,N_3331,N_3377);
and U3408 (N_3408,N_3329,N_3323);
or U3409 (N_3409,N_3327,N_3355);
and U3410 (N_3410,N_3368,N_3369);
or U3411 (N_3411,N_3343,N_3386);
nor U3412 (N_3412,N_3312,N_3350);
nor U3413 (N_3413,N_3389,N_3303);
or U3414 (N_3414,N_3367,N_3338);
xnor U3415 (N_3415,N_3378,N_3346);
nand U3416 (N_3416,N_3358,N_3370);
and U3417 (N_3417,N_3307,N_3362);
nand U3418 (N_3418,N_3310,N_3306);
nand U3419 (N_3419,N_3376,N_3311);
nor U3420 (N_3420,N_3399,N_3344);
nand U3421 (N_3421,N_3371,N_3320);
nand U3422 (N_3422,N_3349,N_3325);
or U3423 (N_3423,N_3351,N_3313);
and U3424 (N_3424,N_3342,N_3353);
nand U3425 (N_3425,N_3393,N_3347);
nor U3426 (N_3426,N_3324,N_3336);
and U3427 (N_3427,N_3374,N_3392);
nand U3428 (N_3428,N_3364,N_3305);
xor U3429 (N_3429,N_3301,N_3308);
or U3430 (N_3430,N_3385,N_3372);
nand U3431 (N_3431,N_3334,N_3373);
xor U3432 (N_3432,N_3366,N_3333);
or U3433 (N_3433,N_3314,N_3363);
nor U3434 (N_3434,N_3315,N_3387);
xor U3435 (N_3435,N_3322,N_3395);
xnor U3436 (N_3436,N_3300,N_3383);
nor U3437 (N_3437,N_3356,N_3321);
xnor U3438 (N_3438,N_3359,N_3326);
and U3439 (N_3439,N_3390,N_3384);
nand U3440 (N_3440,N_3341,N_3382);
nand U3441 (N_3441,N_3317,N_3381);
nor U3442 (N_3442,N_3398,N_3391);
nand U3443 (N_3443,N_3316,N_3354);
nor U3444 (N_3444,N_3302,N_3348);
or U3445 (N_3445,N_3380,N_3365);
nand U3446 (N_3446,N_3328,N_3352);
or U3447 (N_3447,N_3360,N_3319);
or U3448 (N_3448,N_3375,N_3396);
nand U3449 (N_3449,N_3332,N_3318);
nand U3450 (N_3450,N_3386,N_3333);
or U3451 (N_3451,N_3320,N_3347);
nand U3452 (N_3452,N_3337,N_3393);
nor U3453 (N_3453,N_3327,N_3305);
nor U3454 (N_3454,N_3355,N_3317);
nand U3455 (N_3455,N_3364,N_3300);
and U3456 (N_3456,N_3366,N_3328);
or U3457 (N_3457,N_3305,N_3317);
or U3458 (N_3458,N_3346,N_3330);
nor U3459 (N_3459,N_3333,N_3392);
and U3460 (N_3460,N_3337,N_3319);
and U3461 (N_3461,N_3318,N_3307);
nand U3462 (N_3462,N_3394,N_3307);
nor U3463 (N_3463,N_3334,N_3341);
nor U3464 (N_3464,N_3357,N_3345);
and U3465 (N_3465,N_3348,N_3372);
nor U3466 (N_3466,N_3318,N_3368);
xor U3467 (N_3467,N_3312,N_3322);
or U3468 (N_3468,N_3367,N_3309);
and U3469 (N_3469,N_3319,N_3358);
or U3470 (N_3470,N_3361,N_3339);
nand U3471 (N_3471,N_3318,N_3392);
nand U3472 (N_3472,N_3380,N_3391);
or U3473 (N_3473,N_3321,N_3339);
xor U3474 (N_3474,N_3343,N_3310);
nand U3475 (N_3475,N_3312,N_3345);
and U3476 (N_3476,N_3318,N_3348);
nor U3477 (N_3477,N_3399,N_3397);
or U3478 (N_3478,N_3314,N_3383);
or U3479 (N_3479,N_3393,N_3385);
nor U3480 (N_3480,N_3324,N_3398);
nor U3481 (N_3481,N_3320,N_3362);
nand U3482 (N_3482,N_3300,N_3327);
and U3483 (N_3483,N_3325,N_3384);
nor U3484 (N_3484,N_3397,N_3314);
and U3485 (N_3485,N_3368,N_3371);
nand U3486 (N_3486,N_3367,N_3348);
and U3487 (N_3487,N_3353,N_3374);
nand U3488 (N_3488,N_3351,N_3328);
nand U3489 (N_3489,N_3325,N_3395);
nand U3490 (N_3490,N_3385,N_3319);
nor U3491 (N_3491,N_3383,N_3303);
or U3492 (N_3492,N_3344,N_3325);
and U3493 (N_3493,N_3391,N_3378);
nand U3494 (N_3494,N_3381,N_3341);
and U3495 (N_3495,N_3399,N_3381);
nand U3496 (N_3496,N_3342,N_3346);
and U3497 (N_3497,N_3318,N_3319);
nand U3498 (N_3498,N_3366,N_3350);
xnor U3499 (N_3499,N_3369,N_3328);
and U3500 (N_3500,N_3428,N_3418);
nor U3501 (N_3501,N_3459,N_3437);
xnor U3502 (N_3502,N_3482,N_3414);
or U3503 (N_3503,N_3430,N_3486);
nand U3504 (N_3504,N_3450,N_3460);
nor U3505 (N_3505,N_3404,N_3484);
or U3506 (N_3506,N_3415,N_3444);
and U3507 (N_3507,N_3452,N_3467);
nor U3508 (N_3508,N_3488,N_3416);
xnor U3509 (N_3509,N_3462,N_3433);
xor U3510 (N_3510,N_3473,N_3498);
nand U3511 (N_3511,N_3439,N_3407);
nand U3512 (N_3512,N_3491,N_3455);
nor U3513 (N_3513,N_3499,N_3409);
and U3514 (N_3514,N_3410,N_3435);
xor U3515 (N_3515,N_3497,N_3489);
nor U3516 (N_3516,N_3417,N_3487);
nand U3517 (N_3517,N_3472,N_3412);
nand U3518 (N_3518,N_3432,N_3448);
nor U3519 (N_3519,N_3449,N_3478);
nor U3520 (N_3520,N_3421,N_3494);
or U3521 (N_3521,N_3481,N_3456);
xnor U3522 (N_3522,N_3445,N_3492);
nand U3523 (N_3523,N_3468,N_3447);
nand U3524 (N_3524,N_3464,N_3438);
or U3525 (N_3525,N_3475,N_3442);
nor U3526 (N_3526,N_3451,N_3441);
nand U3527 (N_3527,N_3479,N_3443);
xor U3528 (N_3528,N_3413,N_3496);
and U3529 (N_3529,N_3408,N_3495);
nand U3530 (N_3530,N_3476,N_3440);
xor U3531 (N_3531,N_3425,N_3411);
and U3532 (N_3532,N_3400,N_3461);
nor U3533 (N_3533,N_3426,N_3427);
nor U3534 (N_3534,N_3471,N_3454);
nand U3535 (N_3535,N_3405,N_3466);
or U3536 (N_3536,N_3401,N_3406);
or U3537 (N_3537,N_3424,N_3490);
nand U3538 (N_3538,N_3402,N_3458);
nand U3539 (N_3539,N_3434,N_3493);
xor U3540 (N_3540,N_3429,N_3463);
xor U3541 (N_3541,N_3446,N_3457);
xnor U3542 (N_3542,N_3423,N_3436);
or U3543 (N_3543,N_3419,N_3453);
nand U3544 (N_3544,N_3469,N_3431);
nand U3545 (N_3545,N_3477,N_3465);
nand U3546 (N_3546,N_3474,N_3422);
nor U3547 (N_3547,N_3480,N_3420);
nor U3548 (N_3548,N_3470,N_3483);
nand U3549 (N_3549,N_3485,N_3403);
and U3550 (N_3550,N_3485,N_3484);
nor U3551 (N_3551,N_3486,N_3491);
nand U3552 (N_3552,N_3444,N_3472);
nand U3553 (N_3553,N_3438,N_3404);
nor U3554 (N_3554,N_3408,N_3451);
nand U3555 (N_3555,N_3402,N_3474);
and U3556 (N_3556,N_3482,N_3402);
nand U3557 (N_3557,N_3423,N_3444);
and U3558 (N_3558,N_3437,N_3454);
nand U3559 (N_3559,N_3431,N_3498);
nor U3560 (N_3560,N_3411,N_3467);
nand U3561 (N_3561,N_3408,N_3437);
xnor U3562 (N_3562,N_3470,N_3411);
and U3563 (N_3563,N_3499,N_3403);
nand U3564 (N_3564,N_3448,N_3464);
or U3565 (N_3565,N_3494,N_3495);
nand U3566 (N_3566,N_3413,N_3477);
or U3567 (N_3567,N_3497,N_3451);
and U3568 (N_3568,N_3464,N_3433);
nand U3569 (N_3569,N_3423,N_3491);
nand U3570 (N_3570,N_3469,N_3484);
nor U3571 (N_3571,N_3464,N_3417);
nand U3572 (N_3572,N_3492,N_3402);
nand U3573 (N_3573,N_3423,N_3465);
nor U3574 (N_3574,N_3406,N_3410);
xor U3575 (N_3575,N_3485,N_3497);
or U3576 (N_3576,N_3407,N_3476);
or U3577 (N_3577,N_3443,N_3483);
nor U3578 (N_3578,N_3413,N_3402);
nand U3579 (N_3579,N_3453,N_3466);
and U3580 (N_3580,N_3431,N_3428);
or U3581 (N_3581,N_3418,N_3471);
nor U3582 (N_3582,N_3421,N_3437);
nor U3583 (N_3583,N_3433,N_3440);
and U3584 (N_3584,N_3403,N_3441);
or U3585 (N_3585,N_3494,N_3482);
nand U3586 (N_3586,N_3432,N_3415);
and U3587 (N_3587,N_3450,N_3459);
nor U3588 (N_3588,N_3470,N_3466);
xnor U3589 (N_3589,N_3417,N_3427);
nor U3590 (N_3590,N_3480,N_3445);
or U3591 (N_3591,N_3415,N_3410);
nor U3592 (N_3592,N_3412,N_3438);
nor U3593 (N_3593,N_3489,N_3440);
nand U3594 (N_3594,N_3439,N_3406);
xnor U3595 (N_3595,N_3459,N_3438);
xnor U3596 (N_3596,N_3405,N_3484);
nand U3597 (N_3597,N_3497,N_3419);
or U3598 (N_3598,N_3425,N_3440);
and U3599 (N_3599,N_3488,N_3417);
or U3600 (N_3600,N_3573,N_3560);
nand U3601 (N_3601,N_3537,N_3574);
xor U3602 (N_3602,N_3503,N_3589);
nor U3603 (N_3603,N_3533,N_3599);
or U3604 (N_3604,N_3523,N_3552);
and U3605 (N_3605,N_3506,N_3513);
nand U3606 (N_3606,N_3571,N_3567);
xnor U3607 (N_3607,N_3588,N_3595);
nor U3608 (N_3608,N_3505,N_3592);
nor U3609 (N_3609,N_3550,N_3556);
or U3610 (N_3610,N_3508,N_3545);
and U3611 (N_3611,N_3579,N_3565);
and U3612 (N_3612,N_3546,N_3570);
or U3613 (N_3613,N_3572,N_3568);
xnor U3614 (N_3614,N_3581,N_3511);
nor U3615 (N_3615,N_3519,N_3585);
and U3616 (N_3616,N_3516,N_3578);
xnor U3617 (N_3617,N_3544,N_3569);
or U3618 (N_3618,N_3526,N_3518);
nand U3619 (N_3619,N_3597,N_3535);
nand U3620 (N_3620,N_3514,N_3598);
and U3621 (N_3621,N_3559,N_3541);
xor U3622 (N_3622,N_3591,N_3540);
nand U3623 (N_3623,N_3557,N_3596);
nor U3624 (N_3624,N_3566,N_3582);
and U3625 (N_3625,N_3587,N_3530);
or U3626 (N_3626,N_3580,N_3586);
and U3627 (N_3627,N_3553,N_3562);
and U3628 (N_3628,N_3521,N_3510);
and U3629 (N_3629,N_3542,N_3534);
xor U3630 (N_3630,N_3575,N_3539);
or U3631 (N_3631,N_3551,N_3524);
nand U3632 (N_3632,N_3583,N_3512);
and U3633 (N_3633,N_3522,N_3501);
and U3634 (N_3634,N_3584,N_3576);
nand U3635 (N_3635,N_3561,N_3502);
nor U3636 (N_3636,N_3536,N_3563);
xor U3637 (N_3637,N_3515,N_3590);
or U3638 (N_3638,N_3558,N_3564);
nand U3639 (N_3639,N_3500,N_3509);
or U3640 (N_3640,N_3593,N_3549);
nand U3641 (N_3641,N_3529,N_3527);
and U3642 (N_3642,N_3543,N_3525);
nor U3643 (N_3643,N_3577,N_3520);
or U3644 (N_3644,N_3548,N_3547);
nor U3645 (N_3645,N_3538,N_3555);
or U3646 (N_3646,N_3504,N_3517);
nor U3647 (N_3647,N_3532,N_3528);
or U3648 (N_3648,N_3531,N_3507);
nand U3649 (N_3649,N_3594,N_3554);
or U3650 (N_3650,N_3552,N_3578);
nor U3651 (N_3651,N_3544,N_3598);
and U3652 (N_3652,N_3573,N_3564);
and U3653 (N_3653,N_3599,N_3588);
nand U3654 (N_3654,N_3595,N_3581);
and U3655 (N_3655,N_3544,N_3579);
or U3656 (N_3656,N_3539,N_3527);
nor U3657 (N_3657,N_3549,N_3512);
nor U3658 (N_3658,N_3530,N_3539);
nor U3659 (N_3659,N_3570,N_3568);
nand U3660 (N_3660,N_3580,N_3515);
or U3661 (N_3661,N_3501,N_3577);
nand U3662 (N_3662,N_3547,N_3553);
nand U3663 (N_3663,N_3523,N_3508);
xor U3664 (N_3664,N_3587,N_3567);
nand U3665 (N_3665,N_3544,N_3507);
nand U3666 (N_3666,N_3585,N_3539);
nand U3667 (N_3667,N_3546,N_3528);
nor U3668 (N_3668,N_3542,N_3517);
and U3669 (N_3669,N_3525,N_3580);
nand U3670 (N_3670,N_3572,N_3589);
or U3671 (N_3671,N_3541,N_3594);
and U3672 (N_3672,N_3538,N_3590);
xnor U3673 (N_3673,N_3518,N_3519);
nand U3674 (N_3674,N_3570,N_3532);
or U3675 (N_3675,N_3510,N_3558);
xor U3676 (N_3676,N_3555,N_3516);
or U3677 (N_3677,N_3529,N_3589);
nor U3678 (N_3678,N_3597,N_3576);
or U3679 (N_3679,N_3574,N_3500);
nor U3680 (N_3680,N_3518,N_3578);
nand U3681 (N_3681,N_3565,N_3587);
nand U3682 (N_3682,N_3584,N_3572);
and U3683 (N_3683,N_3577,N_3575);
or U3684 (N_3684,N_3564,N_3554);
nor U3685 (N_3685,N_3567,N_3522);
or U3686 (N_3686,N_3588,N_3534);
and U3687 (N_3687,N_3541,N_3515);
nand U3688 (N_3688,N_3538,N_3527);
nand U3689 (N_3689,N_3502,N_3543);
nand U3690 (N_3690,N_3559,N_3526);
xnor U3691 (N_3691,N_3582,N_3502);
and U3692 (N_3692,N_3559,N_3595);
nand U3693 (N_3693,N_3500,N_3510);
or U3694 (N_3694,N_3598,N_3582);
and U3695 (N_3695,N_3527,N_3556);
nor U3696 (N_3696,N_3594,N_3516);
and U3697 (N_3697,N_3534,N_3507);
or U3698 (N_3698,N_3539,N_3533);
xor U3699 (N_3699,N_3580,N_3532);
or U3700 (N_3700,N_3633,N_3608);
nand U3701 (N_3701,N_3660,N_3698);
nor U3702 (N_3702,N_3640,N_3602);
nor U3703 (N_3703,N_3661,N_3695);
nor U3704 (N_3704,N_3690,N_3629);
nand U3705 (N_3705,N_3677,N_3625);
nand U3706 (N_3706,N_3649,N_3616);
nand U3707 (N_3707,N_3664,N_3663);
or U3708 (N_3708,N_3600,N_3680);
nand U3709 (N_3709,N_3693,N_3606);
xor U3710 (N_3710,N_3669,N_3638);
and U3711 (N_3711,N_3665,N_3627);
and U3712 (N_3712,N_3654,N_3682);
and U3713 (N_3713,N_3697,N_3676);
nand U3714 (N_3714,N_3668,N_3672);
and U3715 (N_3715,N_3605,N_3617);
and U3716 (N_3716,N_3652,N_3637);
and U3717 (N_3717,N_3655,N_3611);
or U3718 (N_3718,N_3613,N_3688);
nand U3719 (N_3719,N_3647,N_3670);
or U3720 (N_3720,N_3662,N_3687);
nor U3721 (N_3721,N_3644,N_3634);
nor U3722 (N_3722,N_3692,N_3679);
nand U3723 (N_3723,N_3642,N_3684);
and U3724 (N_3724,N_3673,N_3603);
nand U3725 (N_3725,N_3632,N_3681);
and U3726 (N_3726,N_3648,N_3620);
and U3727 (N_3727,N_3619,N_3689);
xnor U3728 (N_3728,N_3604,N_3691);
nand U3729 (N_3729,N_3653,N_3643);
and U3730 (N_3730,N_3696,N_3614);
or U3731 (N_3731,N_3657,N_3631);
nand U3732 (N_3732,N_3667,N_3645);
or U3733 (N_3733,N_3686,N_3630);
nand U3734 (N_3734,N_3658,N_3612);
xor U3735 (N_3735,N_3666,N_3621);
nor U3736 (N_3736,N_3615,N_3622);
nand U3737 (N_3737,N_3618,N_3601);
and U3738 (N_3738,N_3675,N_3639);
nand U3739 (N_3739,N_3623,N_3609);
nor U3740 (N_3740,N_3641,N_3671);
nand U3741 (N_3741,N_3624,N_3636);
or U3742 (N_3742,N_3685,N_3699);
xor U3743 (N_3743,N_3646,N_3694);
or U3744 (N_3744,N_3678,N_3659);
and U3745 (N_3745,N_3651,N_3683);
or U3746 (N_3746,N_3650,N_3610);
and U3747 (N_3747,N_3635,N_3674);
xnor U3748 (N_3748,N_3626,N_3607);
nor U3749 (N_3749,N_3628,N_3656);
nand U3750 (N_3750,N_3683,N_3628);
nor U3751 (N_3751,N_3652,N_3636);
nor U3752 (N_3752,N_3614,N_3680);
or U3753 (N_3753,N_3655,N_3656);
nand U3754 (N_3754,N_3626,N_3618);
and U3755 (N_3755,N_3673,N_3678);
nor U3756 (N_3756,N_3657,N_3655);
nor U3757 (N_3757,N_3625,N_3693);
xor U3758 (N_3758,N_3690,N_3636);
and U3759 (N_3759,N_3656,N_3696);
xor U3760 (N_3760,N_3647,N_3622);
xor U3761 (N_3761,N_3673,N_3662);
and U3762 (N_3762,N_3690,N_3665);
nor U3763 (N_3763,N_3658,N_3695);
nor U3764 (N_3764,N_3660,N_3608);
nand U3765 (N_3765,N_3699,N_3631);
nor U3766 (N_3766,N_3688,N_3618);
nand U3767 (N_3767,N_3693,N_3655);
xor U3768 (N_3768,N_3618,N_3641);
nand U3769 (N_3769,N_3678,N_3677);
nor U3770 (N_3770,N_3663,N_3692);
and U3771 (N_3771,N_3632,N_3637);
nand U3772 (N_3772,N_3647,N_3654);
and U3773 (N_3773,N_3676,N_3680);
xnor U3774 (N_3774,N_3697,N_3632);
and U3775 (N_3775,N_3625,N_3690);
nand U3776 (N_3776,N_3695,N_3604);
nand U3777 (N_3777,N_3639,N_3679);
or U3778 (N_3778,N_3631,N_3677);
nor U3779 (N_3779,N_3645,N_3686);
nand U3780 (N_3780,N_3661,N_3647);
nand U3781 (N_3781,N_3635,N_3677);
and U3782 (N_3782,N_3687,N_3659);
nand U3783 (N_3783,N_3696,N_3686);
nor U3784 (N_3784,N_3639,N_3665);
or U3785 (N_3785,N_3668,N_3644);
or U3786 (N_3786,N_3686,N_3688);
or U3787 (N_3787,N_3639,N_3676);
or U3788 (N_3788,N_3662,N_3683);
or U3789 (N_3789,N_3619,N_3679);
or U3790 (N_3790,N_3668,N_3646);
nor U3791 (N_3791,N_3673,N_3643);
or U3792 (N_3792,N_3670,N_3637);
nor U3793 (N_3793,N_3675,N_3614);
and U3794 (N_3794,N_3618,N_3670);
or U3795 (N_3795,N_3639,N_3626);
nand U3796 (N_3796,N_3617,N_3650);
or U3797 (N_3797,N_3639,N_3668);
or U3798 (N_3798,N_3621,N_3674);
nor U3799 (N_3799,N_3646,N_3626);
xnor U3800 (N_3800,N_3788,N_3748);
or U3801 (N_3801,N_3753,N_3765);
and U3802 (N_3802,N_3795,N_3782);
and U3803 (N_3803,N_3755,N_3771);
nor U3804 (N_3804,N_3767,N_3721);
and U3805 (N_3805,N_3796,N_3734);
nand U3806 (N_3806,N_3713,N_3764);
nand U3807 (N_3807,N_3789,N_3793);
xor U3808 (N_3808,N_3733,N_3714);
nand U3809 (N_3809,N_3783,N_3719);
and U3810 (N_3810,N_3738,N_3790);
and U3811 (N_3811,N_3736,N_3772);
and U3812 (N_3812,N_3705,N_3784);
nand U3813 (N_3813,N_3739,N_3766);
or U3814 (N_3814,N_3716,N_3785);
and U3815 (N_3815,N_3750,N_3778);
nand U3816 (N_3816,N_3769,N_3777);
or U3817 (N_3817,N_3720,N_3745);
and U3818 (N_3818,N_3707,N_3762);
nand U3819 (N_3819,N_3799,N_3732);
nor U3820 (N_3820,N_3763,N_3749);
nor U3821 (N_3821,N_3725,N_3756);
and U3822 (N_3822,N_3746,N_3779);
or U3823 (N_3823,N_3724,N_3758);
nor U3824 (N_3824,N_3787,N_3715);
and U3825 (N_3825,N_3727,N_3781);
nor U3826 (N_3826,N_3794,N_3770);
nor U3827 (N_3827,N_3706,N_3775);
nand U3828 (N_3828,N_3740,N_3726);
nand U3829 (N_3829,N_3718,N_3752);
nor U3830 (N_3830,N_3744,N_3791);
nor U3831 (N_3831,N_3722,N_3747);
or U3832 (N_3832,N_3776,N_3735);
nor U3833 (N_3833,N_3754,N_3709);
nand U3834 (N_3834,N_3757,N_3703);
nand U3835 (N_3835,N_3768,N_3751);
nor U3836 (N_3836,N_3717,N_3737);
and U3837 (N_3837,N_3774,N_3712);
nor U3838 (N_3838,N_3700,N_3741);
and U3839 (N_3839,N_3711,N_3701);
or U3840 (N_3840,N_3731,N_3761);
nand U3841 (N_3841,N_3780,N_3708);
and U3842 (N_3842,N_3792,N_3760);
and U3843 (N_3843,N_3786,N_3730);
and U3844 (N_3844,N_3710,N_3702);
and U3845 (N_3845,N_3728,N_3798);
nor U3846 (N_3846,N_3743,N_3704);
or U3847 (N_3847,N_3773,N_3723);
nor U3848 (N_3848,N_3742,N_3759);
nor U3849 (N_3849,N_3729,N_3797);
or U3850 (N_3850,N_3777,N_3745);
or U3851 (N_3851,N_3755,N_3780);
nand U3852 (N_3852,N_3701,N_3764);
or U3853 (N_3853,N_3716,N_3702);
and U3854 (N_3854,N_3754,N_3757);
nor U3855 (N_3855,N_3776,N_3786);
xor U3856 (N_3856,N_3723,N_3730);
nor U3857 (N_3857,N_3703,N_3709);
nor U3858 (N_3858,N_3770,N_3716);
xor U3859 (N_3859,N_3797,N_3720);
xnor U3860 (N_3860,N_3787,N_3780);
nor U3861 (N_3861,N_3747,N_3771);
nand U3862 (N_3862,N_3778,N_3777);
nor U3863 (N_3863,N_3716,N_3727);
nor U3864 (N_3864,N_3745,N_3786);
nor U3865 (N_3865,N_3732,N_3734);
and U3866 (N_3866,N_3796,N_3787);
or U3867 (N_3867,N_3703,N_3740);
nor U3868 (N_3868,N_3731,N_3759);
nor U3869 (N_3869,N_3780,N_3752);
nor U3870 (N_3870,N_3738,N_3729);
or U3871 (N_3871,N_3761,N_3750);
nor U3872 (N_3872,N_3739,N_3788);
and U3873 (N_3873,N_3781,N_3797);
nand U3874 (N_3874,N_3765,N_3710);
and U3875 (N_3875,N_3781,N_3755);
nor U3876 (N_3876,N_3789,N_3706);
and U3877 (N_3877,N_3714,N_3773);
or U3878 (N_3878,N_3758,N_3746);
and U3879 (N_3879,N_3782,N_3716);
xnor U3880 (N_3880,N_3717,N_3781);
or U3881 (N_3881,N_3751,N_3731);
and U3882 (N_3882,N_3755,N_3794);
or U3883 (N_3883,N_3791,N_3796);
xnor U3884 (N_3884,N_3724,N_3757);
nand U3885 (N_3885,N_3725,N_3796);
xor U3886 (N_3886,N_3752,N_3779);
nand U3887 (N_3887,N_3774,N_3725);
or U3888 (N_3888,N_3703,N_3768);
or U3889 (N_3889,N_3750,N_3717);
or U3890 (N_3890,N_3700,N_3773);
or U3891 (N_3891,N_3766,N_3732);
or U3892 (N_3892,N_3714,N_3760);
and U3893 (N_3893,N_3797,N_3791);
nor U3894 (N_3894,N_3785,N_3754);
nor U3895 (N_3895,N_3755,N_3702);
and U3896 (N_3896,N_3772,N_3794);
nor U3897 (N_3897,N_3722,N_3789);
nor U3898 (N_3898,N_3768,N_3774);
xor U3899 (N_3899,N_3781,N_3725);
nand U3900 (N_3900,N_3844,N_3822);
nand U3901 (N_3901,N_3841,N_3859);
and U3902 (N_3902,N_3801,N_3862);
or U3903 (N_3903,N_3870,N_3803);
or U3904 (N_3904,N_3836,N_3827);
or U3905 (N_3905,N_3808,N_3860);
or U3906 (N_3906,N_3878,N_3838);
or U3907 (N_3907,N_3818,N_3833);
nand U3908 (N_3908,N_3842,N_3881);
nand U3909 (N_3909,N_3821,N_3897);
nand U3910 (N_3910,N_3892,N_3899);
or U3911 (N_3911,N_3856,N_3887);
nand U3912 (N_3912,N_3884,N_3815);
nor U3913 (N_3913,N_3871,N_3858);
or U3914 (N_3914,N_3855,N_3813);
nand U3915 (N_3915,N_3820,N_3890);
and U3916 (N_3916,N_3882,N_3850);
nand U3917 (N_3917,N_3811,N_3879);
nor U3918 (N_3918,N_3873,N_3861);
nand U3919 (N_3919,N_3823,N_3805);
and U3920 (N_3920,N_3800,N_3830);
or U3921 (N_3921,N_3849,N_3852);
nand U3922 (N_3922,N_3857,N_3847);
and U3923 (N_3923,N_3875,N_3877);
nor U3924 (N_3924,N_3831,N_3869);
and U3925 (N_3925,N_3835,N_3834);
nand U3926 (N_3926,N_3865,N_3874);
or U3927 (N_3927,N_3825,N_3880);
nor U3928 (N_3928,N_3817,N_3863);
or U3929 (N_3929,N_3851,N_3848);
nand U3930 (N_3930,N_3885,N_3819);
nor U3931 (N_3931,N_3845,N_3893);
nor U3932 (N_3932,N_3812,N_3816);
nor U3933 (N_3933,N_3895,N_3872);
xnor U3934 (N_3934,N_3809,N_3889);
nor U3935 (N_3935,N_3868,N_3864);
or U3936 (N_3936,N_3814,N_3826);
and U3937 (N_3937,N_3886,N_3806);
xnor U3938 (N_3938,N_3840,N_3828);
and U3939 (N_3939,N_3807,N_3894);
or U3940 (N_3940,N_3891,N_3843);
or U3941 (N_3941,N_3824,N_3837);
or U3942 (N_3942,N_3888,N_3883);
nor U3943 (N_3943,N_3829,N_3839);
or U3944 (N_3944,N_3804,N_3866);
nand U3945 (N_3945,N_3846,N_3854);
xor U3946 (N_3946,N_3896,N_3810);
nor U3947 (N_3947,N_3867,N_3832);
and U3948 (N_3948,N_3802,N_3898);
nor U3949 (N_3949,N_3876,N_3853);
nor U3950 (N_3950,N_3809,N_3867);
and U3951 (N_3951,N_3826,N_3875);
nor U3952 (N_3952,N_3817,N_3843);
and U3953 (N_3953,N_3826,N_3804);
nand U3954 (N_3954,N_3821,N_3803);
and U3955 (N_3955,N_3830,N_3818);
or U3956 (N_3956,N_3814,N_3805);
and U3957 (N_3957,N_3825,N_3891);
nor U3958 (N_3958,N_3805,N_3896);
nand U3959 (N_3959,N_3808,N_3874);
xor U3960 (N_3960,N_3861,N_3811);
nor U3961 (N_3961,N_3873,N_3853);
or U3962 (N_3962,N_3825,N_3828);
and U3963 (N_3963,N_3892,N_3875);
or U3964 (N_3964,N_3850,N_3868);
or U3965 (N_3965,N_3841,N_3813);
or U3966 (N_3966,N_3838,N_3851);
and U3967 (N_3967,N_3817,N_3854);
nor U3968 (N_3968,N_3806,N_3851);
xor U3969 (N_3969,N_3824,N_3892);
or U3970 (N_3970,N_3808,N_3830);
nand U3971 (N_3971,N_3869,N_3881);
nor U3972 (N_3972,N_3856,N_3806);
nor U3973 (N_3973,N_3845,N_3805);
nor U3974 (N_3974,N_3840,N_3877);
xor U3975 (N_3975,N_3841,N_3831);
or U3976 (N_3976,N_3816,N_3830);
nand U3977 (N_3977,N_3819,N_3825);
and U3978 (N_3978,N_3899,N_3876);
or U3979 (N_3979,N_3858,N_3864);
and U3980 (N_3980,N_3843,N_3871);
nor U3981 (N_3981,N_3894,N_3820);
or U3982 (N_3982,N_3851,N_3849);
or U3983 (N_3983,N_3801,N_3838);
and U3984 (N_3984,N_3803,N_3828);
nor U3985 (N_3985,N_3880,N_3847);
nor U3986 (N_3986,N_3869,N_3882);
nor U3987 (N_3987,N_3870,N_3860);
and U3988 (N_3988,N_3827,N_3819);
and U3989 (N_3989,N_3875,N_3847);
or U3990 (N_3990,N_3891,N_3877);
or U3991 (N_3991,N_3849,N_3832);
or U3992 (N_3992,N_3837,N_3870);
nor U3993 (N_3993,N_3870,N_3830);
nand U3994 (N_3994,N_3897,N_3891);
or U3995 (N_3995,N_3891,N_3853);
nand U3996 (N_3996,N_3843,N_3859);
or U3997 (N_3997,N_3804,N_3891);
nand U3998 (N_3998,N_3836,N_3813);
nor U3999 (N_3999,N_3894,N_3855);
xor U4000 (N_4000,N_3935,N_3955);
nand U4001 (N_4001,N_3984,N_3978);
or U4002 (N_4002,N_3920,N_3904);
nor U4003 (N_4003,N_3946,N_3954);
nor U4004 (N_4004,N_3994,N_3906);
nand U4005 (N_4005,N_3991,N_3971);
and U4006 (N_4006,N_3938,N_3905);
nor U4007 (N_4007,N_3914,N_3963);
and U4008 (N_4008,N_3944,N_3975);
and U4009 (N_4009,N_3972,N_3930);
nor U4010 (N_4010,N_3924,N_3986);
and U4011 (N_4011,N_3940,N_3959);
and U4012 (N_4012,N_3907,N_3925);
nor U4013 (N_4013,N_3912,N_3993);
or U4014 (N_4014,N_3970,N_3903);
nor U4015 (N_4015,N_3937,N_3992);
and U4016 (N_4016,N_3958,N_3941);
or U4017 (N_4017,N_3969,N_3948);
and U4018 (N_4018,N_3956,N_3965);
xor U4019 (N_4019,N_3901,N_3934);
or U4020 (N_4020,N_3982,N_3943);
nand U4021 (N_4021,N_3996,N_3918);
and U4022 (N_4022,N_3915,N_3977);
or U4023 (N_4023,N_3917,N_3913);
and U4024 (N_4024,N_3931,N_3995);
and U4025 (N_4025,N_3942,N_3964);
and U4026 (N_4026,N_3939,N_3987);
nor U4027 (N_4027,N_3957,N_3976);
xnor U4028 (N_4028,N_3902,N_3999);
nor U4029 (N_4029,N_3952,N_3967);
nor U4030 (N_4030,N_3947,N_3927);
or U4031 (N_4031,N_3989,N_3908);
or U4032 (N_4032,N_3936,N_3966);
or U4033 (N_4033,N_3911,N_3933);
nand U4034 (N_4034,N_3900,N_3949);
or U4035 (N_4035,N_3953,N_3968);
nand U4036 (N_4036,N_3962,N_3980);
nand U4037 (N_4037,N_3928,N_3973);
nor U4038 (N_4038,N_3950,N_3979);
or U4039 (N_4039,N_3988,N_3916);
nor U4040 (N_4040,N_3961,N_3951);
nor U4041 (N_4041,N_3910,N_3922);
or U4042 (N_4042,N_3981,N_3985);
nand U4043 (N_4043,N_3919,N_3983);
and U4044 (N_4044,N_3974,N_3909);
nor U4045 (N_4045,N_3926,N_3960);
and U4046 (N_4046,N_3990,N_3998);
or U4047 (N_4047,N_3923,N_3929);
nand U4048 (N_4048,N_3921,N_3997);
and U4049 (N_4049,N_3932,N_3945);
nor U4050 (N_4050,N_3915,N_3994);
nor U4051 (N_4051,N_3976,N_3942);
or U4052 (N_4052,N_3943,N_3916);
nand U4053 (N_4053,N_3962,N_3959);
nand U4054 (N_4054,N_3920,N_3982);
nand U4055 (N_4055,N_3934,N_3924);
nand U4056 (N_4056,N_3981,N_3963);
nor U4057 (N_4057,N_3973,N_3996);
or U4058 (N_4058,N_3942,N_3949);
nor U4059 (N_4059,N_3911,N_3954);
or U4060 (N_4060,N_3924,N_3983);
nand U4061 (N_4061,N_3959,N_3999);
and U4062 (N_4062,N_3914,N_3903);
or U4063 (N_4063,N_3902,N_3913);
and U4064 (N_4064,N_3998,N_3934);
or U4065 (N_4065,N_3903,N_3984);
nor U4066 (N_4066,N_3927,N_3996);
or U4067 (N_4067,N_3941,N_3924);
or U4068 (N_4068,N_3921,N_3904);
xor U4069 (N_4069,N_3982,N_3931);
and U4070 (N_4070,N_3944,N_3922);
and U4071 (N_4071,N_3942,N_3938);
or U4072 (N_4072,N_3980,N_3942);
or U4073 (N_4073,N_3929,N_3956);
nand U4074 (N_4074,N_3912,N_3986);
nor U4075 (N_4075,N_3919,N_3900);
xor U4076 (N_4076,N_3916,N_3935);
or U4077 (N_4077,N_3923,N_3991);
nor U4078 (N_4078,N_3925,N_3920);
or U4079 (N_4079,N_3913,N_3934);
xnor U4080 (N_4080,N_3910,N_3969);
or U4081 (N_4081,N_3957,N_3962);
or U4082 (N_4082,N_3945,N_3935);
xnor U4083 (N_4083,N_3993,N_3936);
or U4084 (N_4084,N_3976,N_3918);
nand U4085 (N_4085,N_3912,N_3939);
nand U4086 (N_4086,N_3912,N_3982);
or U4087 (N_4087,N_3911,N_3992);
and U4088 (N_4088,N_3948,N_3999);
or U4089 (N_4089,N_3955,N_3924);
nand U4090 (N_4090,N_3958,N_3955);
or U4091 (N_4091,N_3986,N_3918);
nand U4092 (N_4092,N_3953,N_3940);
nor U4093 (N_4093,N_3947,N_3983);
and U4094 (N_4094,N_3977,N_3996);
and U4095 (N_4095,N_3950,N_3908);
nand U4096 (N_4096,N_3940,N_3971);
or U4097 (N_4097,N_3972,N_3957);
nand U4098 (N_4098,N_3977,N_3965);
nor U4099 (N_4099,N_3918,N_3973);
nand U4100 (N_4100,N_4082,N_4089);
nand U4101 (N_4101,N_4026,N_4054);
and U4102 (N_4102,N_4069,N_4033);
and U4103 (N_4103,N_4024,N_4057);
and U4104 (N_4104,N_4064,N_4083);
nor U4105 (N_4105,N_4053,N_4012);
nand U4106 (N_4106,N_4097,N_4008);
nand U4107 (N_4107,N_4000,N_4065);
xnor U4108 (N_4108,N_4027,N_4093);
and U4109 (N_4109,N_4092,N_4014);
nor U4110 (N_4110,N_4063,N_4020);
xor U4111 (N_4111,N_4087,N_4032);
nor U4112 (N_4112,N_4043,N_4015);
nand U4113 (N_4113,N_4007,N_4029);
or U4114 (N_4114,N_4058,N_4051);
or U4115 (N_4115,N_4055,N_4011);
nand U4116 (N_4116,N_4005,N_4028);
nor U4117 (N_4117,N_4047,N_4001);
nor U4118 (N_4118,N_4038,N_4074);
nand U4119 (N_4119,N_4077,N_4078);
nand U4120 (N_4120,N_4059,N_4060);
or U4121 (N_4121,N_4018,N_4031);
nand U4122 (N_4122,N_4091,N_4002);
or U4123 (N_4123,N_4090,N_4006);
and U4124 (N_4124,N_4034,N_4049);
nor U4125 (N_4125,N_4076,N_4071);
nand U4126 (N_4126,N_4080,N_4062);
and U4127 (N_4127,N_4085,N_4075);
nand U4128 (N_4128,N_4094,N_4048);
nand U4129 (N_4129,N_4095,N_4098);
or U4130 (N_4130,N_4086,N_4021);
nor U4131 (N_4131,N_4010,N_4066);
nand U4132 (N_4132,N_4099,N_4070);
xor U4133 (N_4133,N_4036,N_4045);
or U4134 (N_4134,N_4004,N_4041);
xor U4135 (N_4135,N_4023,N_4052);
or U4136 (N_4136,N_4030,N_4096);
or U4137 (N_4137,N_4037,N_4046);
nand U4138 (N_4138,N_4061,N_4009);
nor U4139 (N_4139,N_4025,N_4084);
xnor U4140 (N_4140,N_4068,N_4081);
nor U4141 (N_4141,N_4022,N_4035);
or U4142 (N_4142,N_4039,N_4003);
and U4143 (N_4143,N_4079,N_4042);
or U4144 (N_4144,N_4073,N_4072);
nand U4145 (N_4145,N_4013,N_4044);
or U4146 (N_4146,N_4017,N_4019);
and U4147 (N_4147,N_4067,N_4016);
nor U4148 (N_4148,N_4088,N_4056);
xor U4149 (N_4149,N_4040,N_4050);
nand U4150 (N_4150,N_4015,N_4050);
nand U4151 (N_4151,N_4085,N_4031);
nor U4152 (N_4152,N_4058,N_4018);
nand U4153 (N_4153,N_4061,N_4070);
and U4154 (N_4154,N_4075,N_4025);
xnor U4155 (N_4155,N_4059,N_4025);
nor U4156 (N_4156,N_4016,N_4046);
nor U4157 (N_4157,N_4011,N_4029);
nand U4158 (N_4158,N_4085,N_4048);
nand U4159 (N_4159,N_4078,N_4000);
nand U4160 (N_4160,N_4085,N_4060);
nand U4161 (N_4161,N_4094,N_4006);
xnor U4162 (N_4162,N_4096,N_4029);
or U4163 (N_4163,N_4040,N_4041);
and U4164 (N_4164,N_4004,N_4017);
xor U4165 (N_4165,N_4015,N_4066);
nor U4166 (N_4166,N_4037,N_4069);
nand U4167 (N_4167,N_4090,N_4068);
nor U4168 (N_4168,N_4092,N_4019);
or U4169 (N_4169,N_4084,N_4058);
nor U4170 (N_4170,N_4021,N_4008);
nor U4171 (N_4171,N_4027,N_4049);
nor U4172 (N_4172,N_4058,N_4007);
or U4173 (N_4173,N_4069,N_4015);
nor U4174 (N_4174,N_4065,N_4021);
nand U4175 (N_4175,N_4081,N_4035);
nor U4176 (N_4176,N_4094,N_4014);
or U4177 (N_4177,N_4050,N_4028);
nor U4178 (N_4178,N_4033,N_4031);
xnor U4179 (N_4179,N_4011,N_4080);
xor U4180 (N_4180,N_4082,N_4059);
nand U4181 (N_4181,N_4029,N_4076);
nor U4182 (N_4182,N_4083,N_4071);
and U4183 (N_4183,N_4084,N_4027);
nor U4184 (N_4184,N_4091,N_4029);
and U4185 (N_4185,N_4085,N_4022);
nor U4186 (N_4186,N_4023,N_4022);
or U4187 (N_4187,N_4069,N_4022);
or U4188 (N_4188,N_4001,N_4076);
xnor U4189 (N_4189,N_4047,N_4059);
and U4190 (N_4190,N_4050,N_4001);
nor U4191 (N_4191,N_4068,N_4079);
nor U4192 (N_4192,N_4009,N_4086);
nor U4193 (N_4193,N_4084,N_4003);
and U4194 (N_4194,N_4034,N_4074);
and U4195 (N_4195,N_4002,N_4095);
or U4196 (N_4196,N_4046,N_4074);
and U4197 (N_4197,N_4008,N_4085);
nand U4198 (N_4198,N_4025,N_4002);
and U4199 (N_4199,N_4096,N_4098);
and U4200 (N_4200,N_4118,N_4142);
or U4201 (N_4201,N_4179,N_4149);
or U4202 (N_4202,N_4195,N_4132);
xor U4203 (N_4203,N_4163,N_4170);
xor U4204 (N_4204,N_4111,N_4108);
and U4205 (N_4205,N_4190,N_4166);
nor U4206 (N_4206,N_4151,N_4167);
nor U4207 (N_4207,N_4110,N_4172);
nor U4208 (N_4208,N_4169,N_4140);
nand U4209 (N_4209,N_4180,N_4103);
or U4210 (N_4210,N_4138,N_4192);
or U4211 (N_4211,N_4174,N_4143);
nand U4212 (N_4212,N_4148,N_4158);
nand U4213 (N_4213,N_4145,N_4187);
and U4214 (N_4214,N_4193,N_4109);
nand U4215 (N_4215,N_4135,N_4124);
xnor U4216 (N_4216,N_4128,N_4165);
and U4217 (N_4217,N_4183,N_4136);
nor U4218 (N_4218,N_4122,N_4178);
and U4219 (N_4219,N_4120,N_4134);
nand U4220 (N_4220,N_4127,N_4159);
nor U4221 (N_4221,N_4101,N_4177);
nand U4222 (N_4222,N_4100,N_4154);
or U4223 (N_4223,N_4130,N_4146);
nand U4224 (N_4224,N_4162,N_4114);
nor U4225 (N_4225,N_4197,N_4161);
nand U4226 (N_4226,N_4156,N_4144);
nor U4227 (N_4227,N_4117,N_4164);
and U4228 (N_4228,N_4131,N_4139);
or U4229 (N_4229,N_4186,N_4173);
nand U4230 (N_4230,N_4171,N_4121);
nand U4231 (N_4231,N_4185,N_4194);
nand U4232 (N_4232,N_4113,N_4125);
or U4233 (N_4233,N_4182,N_4175);
nand U4234 (N_4234,N_4106,N_4152);
and U4235 (N_4235,N_4168,N_4160);
xor U4236 (N_4236,N_4191,N_4123);
nand U4237 (N_4237,N_4198,N_4116);
or U4238 (N_4238,N_4189,N_4119);
or U4239 (N_4239,N_4157,N_4181);
xor U4240 (N_4240,N_4107,N_4196);
xor U4241 (N_4241,N_4115,N_4199);
and U4242 (N_4242,N_4153,N_4129);
nor U4243 (N_4243,N_4105,N_4184);
nand U4244 (N_4244,N_4150,N_4147);
nand U4245 (N_4245,N_4188,N_4141);
or U4246 (N_4246,N_4112,N_4137);
or U4247 (N_4247,N_4104,N_4126);
xor U4248 (N_4248,N_4155,N_4133);
or U4249 (N_4249,N_4102,N_4176);
or U4250 (N_4250,N_4119,N_4166);
nand U4251 (N_4251,N_4114,N_4182);
or U4252 (N_4252,N_4195,N_4123);
and U4253 (N_4253,N_4188,N_4171);
nor U4254 (N_4254,N_4190,N_4103);
nor U4255 (N_4255,N_4138,N_4108);
nand U4256 (N_4256,N_4157,N_4105);
nor U4257 (N_4257,N_4122,N_4123);
and U4258 (N_4258,N_4124,N_4185);
or U4259 (N_4259,N_4191,N_4188);
and U4260 (N_4260,N_4108,N_4106);
nand U4261 (N_4261,N_4136,N_4103);
nand U4262 (N_4262,N_4172,N_4119);
nor U4263 (N_4263,N_4192,N_4129);
nor U4264 (N_4264,N_4149,N_4168);
xnor U4265 (N_4265,N_4140,N_4196);
nand U4266 (N_4266,N_4107,N_4150);
nor U4267 (N_4267,N_4103,N_4115);
xnor U4268 (N_4268,N_4185,N_4166);
and U4269 (N_4269,N_4143,N_4172);
or U4270 (N_4270,N_4162,N_4157);
nand U4271 (N_4271,N_4120,N_4193);
xnor U4272 (N_4272,N_4153,N_4109);
or U4273 (N_4273,N_4139,N_4185);
xor U4274 (N_4274,N_4103,N_4159);
or U4275 (N_4275,N_4123,N_4193);
or U4276 (N_4276,N_4155,N_4184);
nand U4277 (N_4277,N_4183,N_4190);
nor U4278 (N_4278,N_4119,N_4185);
nand U4279 (N_4279,N_4182,N_4177);
nor U4280 (N_4280,N_4190,N_4119);
and U4281 (N_4281,N_4178,N_4181);
nor U4282 (N_4282,N_4198,N_4140);
or U4283 (N_4283,N_4133,N_4141);
and U4284 (N_4284,N_4160,N_4171);
and U4285 (N_4285,N_4159,N_4167);
or U4286 (N_4286,N_4181,N_4107);
nor U4287 (N_4287,N_4170,N_4142);
or U4288 (N_4288,N_4149,N_4182);
nand U4289 (N_4289,N_4191,N_4118);
nor U4290 (N_4290,N_4159,N_4151);
and U4291 (N_4291,N_4180,N_4104);
nor U4292 (N_4292,N_4131,N_4181);
and U4293 (N_4293,N_4146,N_4105);
or U4294 (N_4294,N_4111,N_4103);
or U4295 (N_4295,N_4156,N_4157);
and U4296 (N_4296,N_4185,N_4153);
and U4297 (N_4297,N_4183,N_4182);
nor U4298 (N_4298,N_4122,N_4177);
and U4299 (N_4299,N_4103,N_4177);
nor U4300 (N_4300,N_4208,N_4239);
nand U4301 (N_4301,N_4290,N_4284);
nor U4302 (N_4302,N_4298,N_4222);
nor U4303 (N_4303,N_4228,N_4218);
and U4304 (N_4304,N_4285,N_4232);
and U4305 (N_4305,N_4216,N_4240);
nor U4306 (N_4306,N_4279,N_4233);
nor U4307 (N_4307,N_4277,N_4206);
nand U4308 (N_4308,N_4231,N_4274);
nand U4309 (N_4309,N_4254,N_4283);
or U4310 (N_4310,N_4207,N_4289);
or U4311 (N_4311,N_4264,N_4201);
or U4312 (N_4312,N_4253,N_4286);
and U4313 (N_4313,N_4225,N_4257);
xnor U4314 (N_4314,N_4237,N_4209);
and U4315 (N_4315,N_4297,N_4213);
and U4316 (N_4316,N_4288,N_4275);
and U4317 (N_4317,N_4203,N_4210);
or U4318 (N_4318,N_4217,N_4265);
and U4319 (N_4319,N_4221,N_4202);
or U4320 (N_4320,N_4261,N_4259);
nor U4321 (N_4321,N_4242,N_4214);
nand U4322 (N_4322,N_4241,N_4273);
xnor U4323 (N_4323,N_4267,N_4252);
nor U4324 (N_4324,N_4211,N_4299);
and U4325 (N_4325,N_4272,N_4238);
nor U4326 (N_4326,N_4255,N_4244);
or U4327 (N_4327,N_4235,N_4247);
or U4328 (N_4328,N_4200,N_4266);
or U4329 (N_4329,N_4246,N_4248);
and U4330 (N_4330,N_4280,N_4234);
and U4331 (N_4331,N_4295,N_4224);
nand U4332 (N_4332,N_4260,N_4204);
and U4333 (N_4333,N_4263,N_4219);
or U4334 (N_4334,N_4291,N_4269);
nor U4335 (N_4335,N_4293,N_4281);
nand U4336 (N_4336,N_4227,N_4230);
nand U4337 (N_4337,N_4268,N_4243);
or U4338 (N_4338,N_4229,N_4236);
xnor U4339 (N_4339,N_4215,N_4271);
nand U4340 (N_4340,N_4223,N_4250);
and U4341 (N_4341,N_4256,N_4270);
nor U4342 (N_4342,N_4212,N_4296);
and U4343 (N_4343,N_4262,N_4294);
or U4344 (N_4344,N_4276,N_4251);
nand U4345 (N_4345,N_4287,N_4220);
nand U4346 (N_4346,N_4278,N_4282);
and U4347 (N_4347,N_4249,N_4226);
nand U4348 (N_4348,N_4258,N_4205);
xor U4349 (N_4349,N_4292,N_4245);
and U4350 (N_4350,N_4263,N_4226);
and U4351 (N_4351,N_4277,N_4214);
and U4352 (N_4352,N_4269,N_4286);
nand U4353 (N_4353,N_4237,N_4205);
and U4354 (N_4354,N_4255,N_4280);
and U4355 (N_4355,N_4217,N_4288);
and U4356 (N_4356,N_4216,N_4222);
and U4357 (N_4357,N_4232,N_4249);
and U4358 (N_4358,N_4232,N_4273);
or U4359 (N_4359,N_4260,N_4268);
xnor U4360 (N_4360,N_4284,N_4285);
nor U4361 (N_4361,N_4206,N_4210);
nand U4362 (N_4362,N_4273,N_4270);
or U4363 (N_4363,N_4278,N_4270);
nor U4364 (N_4364,N_4291,N_4259);
nor U4365 (N_4365,N_4261,N_4267);
nor U4366 (N_4366,N_4235,N_4287);
nor U4367 (N_4367,N_4217,N_4291);
nand U4368 (N_4368,N_4228,N_4287);
nor U4369 (N_4369,N_4290,N_4208);
xor U4370 (N_4370,N_4266,N_4263);
nor U4371 (N_4371,N_4207,N_4299);
or U4372 (N_4372,N_4262,N_4293);
and U4373 (N_4373,N_4265,N_4223);
nor U4374 (N_4374,N_4255,N_4266);
nor U4375 (N_4375,N_4298,N_4290);
nand U4376 (N_4376,N_4252,N_4290);
xnor U4377 (N_4377,N_4270,N_4252);
nand U4378 (N_4378,N_4257,N_4274);
xor U4379 (N_4379,N_4260,N_4277);
or U4380 (N_4380,N_4269,N_4279);
or U4381 (N_4381,N_4294,N_4206);
or U4382 (N_4382,N_4214,N_4291);
or U4383 (N_4383,N_4268,N_4233);
and U4384 (N_4384,N_4274,N_4276);
xnor U4385 (N_4385,N_4244,N_4227);
or U4386 (N_4386,N_4238,N_4282);
nor U4387 (N_4387,N_4282,N_4202);
or U4388 (N_4388,N_4221,N_4237);
or U4389 (N_4389,N_4236,N_4241);
or U4390 (N_4390,N_4288,N_4269);
or U4391 (N_4391,N_4203,N_4293);
nor U4392 (N_4392,N_4246,N_4241);
nor U4393 (N_4393,N_4243,N_4246);
nand U4394 (N_4394,N_4258,N_4274);
nand U4395 (N_4395,N_4226,N_4299);
or U4396 (N_4396,N_4293,N_4299);
xor U4397 (N_4397,N_4273,N_4295);
nor U4398 (N_4398,N_4219,N_4287);
nand U4399 (N_4399,N_4242,N_4269);
and U4400 (N_4400,N_4304,N_4384);
or U4401 (N_4401,N_4356,N_4397);
nor U4402 (N_4402,N_4315,N_4367);
and U4403 (N_4403,N_4343,N_4369);
nor U4404 (N_4404,N_4395,N_4380);
nand U4405 (N_4405,N_4319,N_4328);
and U4406 (N_4406,N_4307,N_4364);
nor U4407 (N_4407,N_4378,N_4352);
and U4408 (N_4408,N_4398,N_4382);
and U4409 (N_4409,N_4316,N_4300);
nand U4410 (N_4410,N_4326,N_4322);
or U4411 (N_4411,N_4391,N_4337);
xor U4412 (N_4412,N_4365,N_4361);
xnor U4413 (N_4413,N_4387,N_4306);
or U4414 (N_4414,N_4396,N_4335);
nor U4415 (N_4415,N_4388,N_4341);
or U4416 (N_4416,N_4325,N_4331);
xnor U4417 (N_4417,N_4363,N_4324);
nand U4418 (N_4418,N_4357,N_4393);
or U4419 (N_4419,N_4314,N_4381);
nand U4420 (N_4420,N_4338,N_4372);
or U4421 (N_4421,N_4386,N_4344);
nand U4422 (N_4422,N_4370,N_4329);
and U4423 (N_4423,N_4373,N_4345);
nor U4424 (N_4424,N_4318,N_4336);
nand U4425 (N_4425,N_4303,N_4311);
and U4426 (N_4426,N_4392,N_4321);
nor U4427 (N_4427,N_4371,N_4376);
and U4428 (N_4428,N_4302,N_4362);
nor U4429 (N_4429,N_4312,N_4385);
or U4430 (N_4430,N_4342,N_4339);
nand U4431 (N_4431,N_4346,N_4379);
or U4432 (N_4432,N_4368,N_4390);
nand U4433 (N_4433,N_4347,N_4309);
nor U4434 (N_4434,N_4353,N_4360);
nor U4435 (N_4435,N_4375,N_4334);
or U4436 (N_4436,N_4355,N_4332);
nor U4437 (N_4437,N_4333,N_4389);
xnor U4438 (N_4438,N_4320,N_4323);
or U4439 (N_4439,N_4308,N_4340);
nor U4440 (N_4440,N_4350,N_4383);
and U4441 (N_4441,N_4349,N_4374);
nand U4442 (N_4442,N_4301,N_4348);
xor U4443 (N_4443,N_4358,N_4305);
nor U4444 (N_4444,N_4313,N_4310);
nand U4445 (N_4445,N_4327,N_4399);
or U4446 (N_4446,N_4354,N_4317);
nand U4447 (N_4447,N_4394,N_4351);
nand U4448 (N_4448,N_4330,N_4366);
and U4449 (N_4449,N_4377,N_4359);
and U4450 (N_4450,N_4331,N_4337);
or U4451 (N_4451,N_4370,N_4367);
and U4452 (N_4452,N_4359,N_4398);
nand U4453 (N_4453,N_4314,N_4319);
nor U4454 (N_4454,N_4380,N_4370);
and U4455 (N_4455,N_4359,N_4322);
nand U4456 (N_4456,N_4381,N_4367);
nor U4457 (N_4457,N_4394,N_4314);
nor U4458 (N_4458,N_4309,N_4311);
nor U4459 (N_4459,N_4377,N_4349);
and U4460 (N_4460,N_4366,N_4377);
and U4461 (N_4461,N_4391,N_4375);
or U4462 (N_4462,N_4307,N_4344);
and U4463 (N_4463,N_4374,N_4388);
nor U4464 (N_4464,N_4398,N_4331);
nor U4465 (N_4465,N_4382,N_4326);
and U4466 (N_4466,N_4341,N_4367);
or U4467 (N_4467,N_4375,N_4308);
nand U4468 (N_4468,N_4321,N_4323);
or U4469 (N_4469,N_4315,N_4360);
and U4470 (N_4470,N_4300,N_4320);
xnor U4471 (N_4471,N_4343,N_4338);
xnor U4472 (N_4472,N_4349,N_4332);
xnor U4473 (N_4473,N_4353,N_4388);
and U4474 (N_4474,N_4362,N_4333);
nor U4475 (N_4475,N_4371,N_4353);
and U4476 (N_4476,N_4350,N_4367);
or U4477 (N_4477,N_4307,N_4350);
and U4478 (N_4478,N_4380,N_4326);
or U4479 (N_4479,N_4344,N_4352);
and U4480 (N_4480,N_4367,N_4308);
and U4481 (N_4481,N_4366,N_4335);
nor U4482 (N_4482,N_4368,N_4341);
and U4483 (N_4483,N_4373,N_4301);
nor U4484 (N_4484,N_4327,N_4350);
nand U4485 (N_4485,N_4331,N_4339);
xor U4486 (N_4486,N_4385,N_4341);
and U4487 (N_4487,N_4395,N_4363);
nor U4488 (N_4488,N_4315,N_4390);
and U4489 (N_4489,N_4339,N_4388);
and U4490 (N_4490,N_4371,N_4318);
and U4491 (N_4491,N_4305,N_4318);
nand U4492 (N_4492,N_4332,N_4324);
nand U4493 (N_4493,N_4384,N_4333);
and U4494 (N_4494,N_4311,N_4397);
and U4495 (N_4495,N_4357,N_4309);
nand U4496 (N_4496,N_4332,N_4304);
and U4497 (N_4497,N_4320,N_4399);
and U4498 (N_4498,N_4379,N_4332);
and U4499 (N_4499,N_4399,N_4338);
and U4500 (N_4500,N_4454,N_4400);
nand U4501 (N_4501,N_4412,N_4497);
and U4502 (N_4502,N_4492,N_4419);
nand U4503 (N_4503,N_4466,N_4479);
xor U4504 (N_4504,N_4417,N_4423);
or U4505 (N_4505,N_4420,N_4467);
xor U4506 (N_4506,N_4456,N_4442);
and U4507 (N_4507,N_4469,N_4490);
and U4508 (N_4508,N_4440,N_4408);
or U4509 (N_4509,N_4485,N_4451);
xor U4510 (N_4510,N_4444,N_4434);
or U4511 (N_4511,N_4428,N_4425);
or U4512 (N_4512,N_4443,N_4427);
nand U4513 (N_4513,N_4495,N_4445);
or U4514 (N_4514,N_4415,N_4410);
xnor U4515 (N_4515,N_4426,N_4463);
or U4516 (N_4516,N_4437,N_4450);
nand U4517 (N_4517,N_4435,N_4459);
and U4518 (N_4518,N_4432,N_4438);
and U4519 (N_4519,N_4402,N_4422);
xor U4520 (N_4520,N_4489,N_4481);
nand U4521 (N_4521,N_4455,N_4447);
or U4522 (N_4522,N_4474,N_4430);
nor U4523 (N_4523,N_4449,N_4418);
nor U4524 (N_4524,N_4452,N_4404);
nor U4525 (N_4525,N_4403,N_4436);
and U4526 (N_4526,N_4486,N_4407);
xnor U4527 (N_4527,N_4480,N_4457);
xnor U4528 (N_4528,N_4409,N_4484);
nor U4529 (N_4529,N_4491,N_4472);
and U4530 (N_4530,N_4462,N_4478);
or U4531 (N_4531,N_4493,N_4487);
nor U4532 (N_4532,N_4458,N_4498);
or U4533 (N_4533,N_4483,N_4475);
and U4534 (N_4534,N_4470,N_4405);
xnor U4535 (N_4535,N_4499,N_4406);
nand U4536 (N_4536,N_4488,N_4482);
nand U4537 (N_4537,N_4494,N_4461);
nor U4538 (N_4538,N_4411,N_4468);
and U4539 (N_4539,N_4433,N_4476);
and U4540 (N_4540,N_4424,N_4465);
nand U4541 (N_4541,N_4473,N_4414);
xor U4542 (N_4542,N_4421,N_4413);
nor U4543 (N_4543,N_4416,N_4431);
nand U4544 (N_4544,N_4448,N_4464);
nor U4545 (N_4545,N_4401,N_4446);
and U4546 (N_4546,N_4453,N_4460);
nand U4547 (N_4547,N_4441,N_4439);
nor U4548 (N_4548,N_4477,N_4429);
nand U4549 (N_4549,N_4496,N_4471);
and U4550 (N_4550,N_4443,N_4431);
and U4551 (N_4551,N_4461,N_4402);
and U4552 (N_4552,N_4442,N_4407);
nand U4553 (N_4553,N_4409,N_4456);
or U4554 (N_4554,N_4487,N_4489);
nand U4555 (N_4555,N_4490,N_4451);
nand U4556 (N_4556,N_4401,N_4423);
nor U4557 (N_4557,N_4404,N_4434);
nor U4558 (N_4558,N_4414,N_4468);
and U4559 (N_4559,N_4479,N_4434);
and U4560 (N_4560,N_4482,N_4435);
and U4561 (N_4561,N_4464,N_4446);
or U4562 (N_4562,N_4480,N_4481);
or U4563 (N_4563,N_4427,N_4477);
nand U4564 (N_4564,N_4472,N_4407);
or U4565 (N_4565,N_4493,N_4481);
nor U4566 (N_4566,N_4403,N_4450);
xor U4567 (N_4567,N_4467,N_4449);
nor U4568 (N_4568,N_4420,N_4421);
nor U4569 (N_4569,N_4414,N_4437);
or U4570 (N_4570,N_4493,N_4412);
nand U4571 (N_4571,N_4492,N_4493);
nor U4572 (N_4572,N_4452,N_4405);
nand U4573 (N_4573,N_4407,N_4476);
nor U4574 (N_4574,N_4447,N_4475);
or U4575 (N_4575,N_4464,N_4499);
and U4576 (N_4576,N_4472,N_4489);
nand U4577 (N_4577,N_4427,N_4464);
nand U4578 (N_4578,N_4462,N_4460);
nor U4579 (N_4579,N_4484,N_4447);
nand U4580 (N_4580,N_4426,N_4497);
and U4581 (N_4581,N_4496,N_4449);
or U4582 (N_4582,N_4469,N_4482);
nor U4583 (N_4583,N_4446,N_4494);
or U4584 (N_4584,N_4420,N_4435);
and U4585 (N_4585,N_4461,N_4433);
or U4586 (N_4586,N_4476,N_4405);
nor U4587 (N_4587,N_4473,N_4453);
xor U4588 (N_4588,N_4489,N_4488);
nor U4589 (N_4589,N_4482,N_4476);
or U4590 (N_4590,N_4407,N_4457);
nand U4591 (N_4591,N_4498,N_4452);
nor U4592 (N_4592,N_4462,N_4461);
nand U4593 (N_4593,N_4447,N_4490);
nand U4594 (N_4594,N_4477,N_4459);
and U4595 (N_4595,N_4443,N_4409);
or U4596 (N_4596,N_4429,N_4409);
nor U4597 (N_4597,N_4490,N_4492);
xor U4598 (N_4598,N_4426,N_4498);
nor U4599 (N_4599,N_4481,N_4495);
nor U4600 (N_4600,N_4558,N_4561);
nor U4601 (N_4601,N_4516,N_4533);
nand U4602 (N_4602,N_4585,N_4520);
nor U4603 (N_4603,N_4580,N_4502);
nor U4604 (N_4604,N_4587,N_4550);
nor U4605 (N_4605,N_4507,N_4510);
nor U4606 (N_4606,N_4517,N_4509);
nor U4607 (N_4607,N_4506,N_4592);
nor U4608 (N_4608,N_4504,N_4501);
nor U4609 (N_4609,N_4519,N_4596);
nand U4610 (N_4610,N_4583,N_4575);
nand U4611 (N_4611,N_4546,N_4505);
nand U4612 (N_4612,N_4528,N_4562);
nor U4613 (N_4613,N_4572,N_4541);
and U4614 (N_4614,N_4588,N_4570);
or U4615 (N_4615,N_4543,N_4593);
or U4616 (N_4616,N_4591,N_4566);
xor U4617 (N_4617,N_4511,N_4595);
nand U4618 (N_4618,N_4524,N_4534);
or U4619 (N_4619,N_4579,N_4597);
nand U4620 (N_4620,N_4529,N_4557);
and U4621 (N_4621,N_4553,N_4599);
and U4622 (N_4622,N_4576,N_4552);
or U4623 (N_4623,N_4554,N_4582);
nand U4624 (N_4624,N_4563,N_4532);
nor U4625 (N_4625,N_4598,N_4551);
nor U4626 (N_4626,N_4560,N_4514);
or U4627 (N_4627,N_4537,N_4503);
nor U4628 (N_4628,N_4549,N_4590);
and U4629 (N_4629,N_4565,N_4539);
nor U4630 (N_4630,N_4559,N_4508);
nor U4631 (N_4631,N_4531,N_4538);
nor U4632 (N_4632,N_4525,N_4544);
and U4633 (N_4633,N_4564,N_4574);
and U4634 (N_4634,N_4584,N_4548);
and U4635 (N_4635,N_4569,N_4515);
or U4636 (N_4636,N_4542,N_4513);
and U4637 (N_4637,N_4568,N_4540);
nor U4638 (N_4638,N_4571,N_4521);
nand U4639 (N_4639,N_4523,N_4586);
nor U4640 (N_4640,N_4512,N_4527);
or U4641 (N_4641,N_4535,N_4577);
and U4642 (N_4642,N_4581,N_4556);
xnor U4643 (N_4643,N_4573,N_4526);
xor U4644 (N_4644,N_4500,N_4547);
and U4645 (N_4645,N_4594,N_4589);
nor U4646 (N_4646,N_4567,N_4518);
nand U4647 (N_4647,N_4522,N_4536);
nand U4648 (N_4648,N_4555,N_4530);
nand U4649 (N_4649,N_4578,N_4545);
xor U4650 (N_4650,N_4547,N_4544);
or U4651 (N_4651,N_4541,N_4525);
or U4652 (N_4652,N_4540,N_4596);
or U4653 (N_4653,N_4556,N_4572);
nor U4654 (N_4654,N_4568,N_4511);
and U4655 (N_4655,N_4573,N_4542);
nand U4656 (N_4656,N_4556,N_4574);
and U4657 (N_4657,N_4533,N_4547);
or U4658 (N_4658,N_4557,N_4502);
nor U4659 (N_4659,N_4588,N_4512);
and U4660 (N_4660,N_4594,N_4567);
nand U4661 (N_4661,N_4559,N_4521);
or U4662 (N_4662,N_4531,N_4532);
nor U4663 (N_4663,N_4555,N_4575);
nor U4664 (N_4664,N_4523,N_4576);
nor U4665 (N_4665,N_4542,N_4599);
xnor U4666 (N_4666,N_4566,N_4501);
and U4667 (N_4667,N_4575,N_4537);
and U4668 (N_4668,N_4516,N_4571);
nand U4669 (N_4669,N_4536,N_4599);
nor U4670 (N_4670,N_4573,N_4597);
and U4671 (N_4671,N_4544,N_4531);
xor U4672 (N_4672,N_4536,N_4565);
nor U4673 (N_4673,N_4569,N_4591);
nand U4674 (N_4674,N_4578,N_4557);
nand U4675 (N_4675,N_4553,N_4580);
nor U4676 (N_4676,N_4586,N_4543);
nor U4677 (N_4677,N_4565,N_4526);
and U4678 (N_4678,N_4597,N_4583);
or U4679 (N_4679,N_4588,N_4551);
nand U4680 (N_4680,N_4560,N_4588);
nand U4681 (N_4681,N_4554,N_4551);
nand U4682 (N_4682,N_4527,N_4581);
nand U4683 (N_4683,N_4584,N_4569);
or U4684 (N_4684,N_4507,N_4521);
nor U4685 (N_4685,N_4547,N_4595);
nand U4686 (N_4686,N_4561,N_4584);
or U4687 (N_4687,N_4588,N_4595);
or U4688 (N_4688,N_4578,N_4588);
or U4689 (N_4689,N_4507,N_4575);
nand U4690 (N_4690,N_4523,N_4567);
or U4691 (N_4691,N_4537,N_4586);
or U4692 (N_4692,N_4541,N_4524);
or U4693 (N_4693,N_4545,N_4557);
nand U4694 (N_4694,N_4583,N_4513);
nor U4695 (N_4695,N_4515,N_4572);
nor U4696 (N_4696,N_4541,N_4508);
or U4697 (N_4697,N_4516,N_4528);
xor U4698 (N_4698,N_4587,N_4575);
xnor U4699 (N_4699,N_4558,N_4516);
nand U4700 (N_4700,N_4612,N_4613);
xor U4701 (N_4701,N_4601,N_4615);
or U4702 (N_4702,N_4642,N_4685);
and U4703 (N_4703,N_4603,N_4665);
nand U4704 (N_4704,N_4646,N_4655);
or U4705 (N_4705,N_4664,N_4658);
xor U4706 (N_4706,N_4654,N_4686);
xnor U4707 (N_4707,N_4614,N_4689);
nor U4708 (N_4708,N_4680,N_4650);
nand U4709 (N_4709,N_4620,N_4630);
nand U4710 (N_4710,N_4622,N_4628);
nor U4711 (N_4711,N_4671,N_4611);
and U4712 (N_4712,N_4660,N_4673);
nor U4713 (N_4713,N_4623,N_4634);
nand U4714 (N_4714,N_4675,N_4688);
and U4715 (N_4715,N_4617,N_4653);
nor U4716 (N_4716,N_4697,N_4661);
nand U4717 (N_4717,N_4631,N_4698);
or U4718 (N_4718,N_4692,N_4657);
or U4719 (N_4719,N_4677,N_4668);
or U4720 (N_4720,N_4600,N_4670);
nand U4721 (N_4721,N_4632,N_4621);
xnor U4722 (N_4722,N_4666,N_4699);
and U4723 (N_4723,N_4609,N_4669);
nor U4724 (N_4724,N_4695,N_4684);
and U4725 (N_4725,N_4656,N_4639);
and U4726 (N_4726,N_4635,N_4648);
or U4727 (N_4727,N_4678,N_4633);
and U4728 (N_4728,N_4651,N_4682);
or U4729 (N_4729,N_4659,N_4693);
nand U4730 (N_4730,N_4643,N_4687);
or U4731 (N_4731,N_4608,N_4637);
nand U4732 (N_4732,N_4676,N_4606);
nor U4733 (N_4733,N_4674,N_4691);
nor U4734 (N_4734,N_4681,N_4663);
or U4735 (N_4735,N_4604,N_4624);
and U4736 (N_4736,N_4645,N_4647);
or U4737 (N_4737,N_4683,N_4644);
and U4738 (N_4738,N_4626,N_4679);
xor U4739 (N_4739,N_4610,N_4638);
and U4740 (N_4740,N_4636,N_4696);
xor U4741 (N_4741,N_4605,N_4629);
nand U4742 (N_4742,N_4627,N_4602);
and U4743 (N_4743,N_4662,N_4607);
nand U4744 (N_4744,N_4690,N_4667);
and U4745 (N_4745,N_4618,N_4649);
nand U4746 (N_4746,N_4672,N_4640);
nand U4747 (N_4747,N_4641,N_4694);
or U4748 (N_4748,N_4619,N_4625);
nor U4749 (N_4749,N_4652,N_4616);
or U4750 (N_4750,N_4678,N_4648);
or U4751 (N_4751,N_4661,N_4693);
and U4752 (N_4752,N_4669,N_4626);
or U4753 (N_4753,N_4633,N_4640);
nor U4754 (N_4754,N_4676,N_4616);
or U4755 (N_4755,N_4679,N_4632);
nor U4756 (N_4756,N_4658,N_4612);
xnor U4757 (N_4757,N_4689,N_4694);
and U4758 (N_4758,N_4664,N_4678);
and U4759 (N_4759,N_4639,N_4627);
and U4760 (N_4760,N_4649,N_4660);
and U4761 (N_4761,N_4667,N_4671);
and U4762 (N_4762,N_4666,N_4600);
nand U4763 (N_4763,N_4617,N_4637);
and U4764 (N_4764,N_4683,N_4610);
or U4765 (N_4765,N_4604,N_4639);
nand U4766 (N_4766,N_4611,N_4625);
nor U4767 (N_4767,N_4629,N_4646);
nor U4768 (N_4768,N_4676,N_4614);
nor U4769 (N_4769,N_4668,N_4698);
xor U4770 (N_4770,N_4674,N_4696);
or U4771 (N_4771,N_4608,N_4600);
nor U4772 (N_4772,N_4605,N_4666);
nand U4773 (N_4773,N_4641,N_4619);
nand U4774 (N_4774,N_4651,N_4641);
nand U4775 (N_4775,N_4668,N_4690);
nor U4776 (N_4776,N_4602,N_4605);
nor U4777 (N_4777,N_4604,N_4608);
nand U4778 (N_4778,N_4600,N_4674);
nor U4779 (N_4779,N_4635,N_4643);
or U4780 (N_4780,N_4663,N_4689);
nand U4781 (N_4781,N_4672,N_4610);
or U4782 (N_4782,N_4676,N_4686);
or U4783 (N_4783,N_4601,N_4610);
nand U4784 (N_4784,N_4696,N_4695);
nor U4785 (N_4785,N_4621,N_4611);
and U4786 (N_4786,N_4615,N_4671);
xnor U4787 (N_4787,N_4684,N_4698);
and U4788 (N_4788,N_4656,N_4649);
and U4789 (N_4789,N_4629,N_4696);
nand U4790 (N_4790,N_4673,N_4619);
nor U4791 (N_4791,N_4642,N_4620);
nand U4792 (N_4792,N_4682,N_4604);
nand U4793 (N_4793,N_4671,N_4662);
xnor U4794 (N_4794,N_4677,N_4621);
nand U4795 (N_4795,N_4643,N_4652);
nand U4796 (N_4796,N_4614,N_4678);
nor U4797 (N_4797,N_4663,N_4677);
and U4798 (N_4798,N_4683,N_4692);
nor U4799 (N_4799,N_4668,N_4622);
or U4800 (N_4800,N_4794,N_4784);
nand U4801 (N_4801,N_4703,N_4778);
and U4802 (N_4802,N_4788,N_4713);
and U4803 (N_4803,N_4761,N_4777);
nand U4804 (N_4804,N_4747,N_4744);
nand U4805 (N_4805,N_4715,N_4755);
and U4806 (N_4806,N_4740,N_4782);
and U4807 (N_4807,N_4760,N_4756);
xnor U4808 (N_4808,N_4733,N_4736);
or U4809 (N_4809,N_4720,N_4732);
or U4810 (N_4810,N_4743,N_4741);
nor U4811 (N_4811,N_4759,N_4712);
and U4812 (N_4812,N_4769,N_4796);
and U4813 (N_4813,N_4791,N_4718);
and U4814 (N_4814,N_4792,N_4771);
nand U4815 (N_4815,N_4780,N_4724);
xnor U4816 (N_4816,N_4797,N_4783);
and U4817 (N_4817,N_4773,N_4795);
nand U4818 (N_4818,N_4708,N_4738);
or U4819 (N_4819,N_4774,N_4757);
xor U4820 (N_4820,N_4730,N_4719);
xor U4821 (N_4821,N_4781,N_4745);
xor U4822 (N_4822,N_4731,N_4750);
xor U4823 (N_4823,N_4751,N_4704);
and U4824 (N_4824,N_4779,N_4716);
and U4825 (N_4825,N_4776,N_4793);
nand U4826 (N_4826,N_4787,N_4725);
and U4827 (N_4827,N_4701,N_4742);
nand U4828 (N_4828,N_4706,N_4702);
nor U4829 (N_4829,N_4749,N_4799);
or U4830 (N_4830,N_4737,N_4775);
nor U4831 (N_4831,N_4766,N_4735);
or U4832 (N_4832,N_4728,N_4726);
nand U4833 (N_4833,N_4752,N_4770);
xor U4834 (N_4834,N_4727,N_4754);
and U4835 (N_4835,N_4798,N_4765);
and U4836 (N_4836,N_4767,N_4723);
and U4837 (N_4837,N_4739,N_4729);
and U4838 (N_4838,N_4700,N_4711);
nand U4839 (N_4839,N_4758,N_4714);
and U4840 (N_4840,N_4763,N_4709);
nor U4841 (N_4841,N_4717,N_4786);
or U4842 (N_4842,N_4762,N_4705);
and U4843 (N_4843,N_4785,N_4789);
and U4844 (N_4844,N_4790,N_4734);
xor U4845 (N_4845,N_4746,N_4768);
and U4846 (N_4846,N_4722,N_4748);
nor U4847 (N_4847,N_4721,N_4753);
nor U4848 (N_4848,N_4772,N_4707);
nand U4849 (N_4849,N_4764,N_4710);
or U4850 (N_4850,N_4794,N_4756);
nor U4851 (N_4851,N_4720,N_4784);
xor U4852 (N_4852,N_4742,N_4715);
nand U4853 (N_4853,N_4752,N_4787);
nor U4854 (N_4854,N_4777,N_4726);
nand U4855 (N_4855,N_4760,N_4772);
and U4856 (N_4856,N_4719,N_4761);
nand U4857 (N_4857,N_4702,N_4780);
nor U4858 (N_4858,N_4717,N_4787);
nand U4859 (N_4859,N_4733,N_4707);
xor U4860 (N_4860,N_4715,N_4706);
or U4861 (N_4861,N_4749,N_4794);
or U4862 (N_4862,N_4793,N_4791);
nor U4863 (N_4863,N_4759,N_4737);
and U4864 (N_4864,N_4729,N_4774);
and U4865 (N_4865,N_4734,N_4726);
xor U4866 (N_4866,N_4776,N_4794);
and U4867 (N_4867,N_4720,N_4779);
or U4868 (N_4868,N_4796,N_4711);
and U4869 (N_4869,N_4733,N_4755);
or U4870 (N_4870,N_4706,N_4754);
and U4871 (N_4871,N_4723,N_4762);
nand U4872 (N_4872,N_4798,N_4781);
xor U4873 (N_4873,N_4764,N_4706);
xor U4874 (N_4874,N_4705,N_4770);
nand U4875 (N_4875,N_4779,N_4765);
nor U4876 (N_4876,N_4728,N_4797);
xnor U4877 (N_4877,N_4717,N_4731);
nor U4878 (N_4878,N_4743,N_4777);
and U4879 (N_4879,N_4772,N_4730);
or U4880 (N_4880,N_4718,N_4770);
nand U4881 (N_4881,N_4779,N_4733);
and U4882 (N_4882,N_4724,N_4748);
or U4883 (N_4883,N_4701,N_4739);
nor U4884 (N_4884,N_4740,N_4722);
xor U4885 (N_4885,N_4784,N_4735);
xor U4886 (N_4886,N_4730,N_4788);
nor U4887 (N_4887,N_4708,N_4789);
and U4888 (N_4888,N_4783,N_4718);
nand U4889 (N_4889,N_4713,N_4708);
nand U4890 (N_4890,N_4736,N_4721);
or U4891 (N_4891,N_4725,N_4730);
nor U4892 (N_4892,N_4722,N_4703);
xor U4893 (N_4893,N_4707,N_4768);
or U4894 (N_4894,N_4793,N_4787);
and U4895 (N_4895,N_4798,N_4793);
nor U4896 (N_4896,N_4773,N_4747);
nand U4897 (N_4897,N_4746,N_4717);
and U4898 (N_4898,N_4794,N_4780);
xnor U4899 (N_4899,N_4723,N_4787);
nand U4900 (N_4900,N_4872,N_4838);
or U4901 (N_4901,N_4832,N_4800);
nand U4902 (N_4902,N_4840,N_4868);
nand U4903 (N_4903,N_4877,N_4829);
nand U4904 (N_4904,N_4864,N_4806);
nor U4905 (N_4905,N_4815,N_4801);
or U4906 (N_4906,N_4802,N_4845);
nor U4907 (N_4907,N_4878,N_4894);
nor U4908 (N_4908,N_4826,N_4875);
or U4909 (N_4909,N_4870,N_4884);
nor U4910 (N_4910,N_4836,N_4816);
and U4911 (N_4911,N_4859,N_4813);
and U4912 (N_4912,N_4862,N_4881);
nand U4913 (N_4913,N_4892,N_4837);
xor U4914 (N_4914,N_4866,N_4849);
or U4915 (N_4915,N_4839,N_4850);
xnor U4916 (N_4916,N_4822,N_4804);
nand U4917 (N_4917,N_4873,N_4809);
nor U4918 (N_4918,N_4851,N_4887);
and U4919 (N_4919,N_4821,N_4834);
or U4920 (N_4920,N_4876,N_4812);
xnor U4921 (N_4921,N_4860,N_4853);
nor U4922 (N_4922,N_4805,N_4895);
or U4923 (N_4923,N_4811,N_4899);
nor U4924 (N_4924,N_4848,N_4886);
xor U4925 (N_4925,N_4810,N_4841);
or U4926 (N_4926,N_4818,N_4861);
and U4927 (N_4927,N_4817,N_4898);
nand U4928 (N_4928,N_4865,N_4803);
nand U4929 (N_4929,N_4824,N_4880);
or U4930 (N_4930,N_4844,N_4835);
xor U4931 (N_4931,N_4883,N_4820);
nor U4932 (N_4932,N_4833,N_4847);
nor U4933 (N_4933,N_4896,N_4846);
nor U4934 (N_4934,N_4857,N_4874);
xor U4935 (N_4935,N_4819,N_4856);
or U4936 (N_4936,N_4825,N_4855);
nor U4937 (N_4937,N_4882,N_4897);
nor U4938 (N_4938,N_4807,N_4858);
nand U4939 (N_4939,N_4854,N_4885);
or U4940 (N_4940,N_4814,N_4889);
nand U4941 (N_4941,N_4830,N_4842);
nor U4942 (N_4942,N_4823,N_4827);
nor U4943 (N_4943,N_4831,N_4869);
and U4944 (N_4944,N_4890,N_4888);
or U4945 (N_4945,N_4808,N_4843);
and U4946 (N_4946,N_4852,N_4879);
nand U4947 (N_4947,N_4867,N_4893);
or U4948 (N_4948,N_4891,N_4871);
or U4949 (N_4949,N_4863,N_4828);
xnor U4950 (N_4950,N_4815,N_4830);
or U4951 (N_4951,N_4842,N_4854);
xor U4952 (N_4952,N_4825,N_4850);
nand U4953 (N_4953,N_4836,N_4841);
nor U4954 (N_4954,N_4826,N_4836);
nand U4955 (N_4955,N_4891,N_4802);
and U4956 (N_4956,N_4804,N_4864);
nor U4957 (N_4957,N_4810,N_4857);
and U4958 (N_4958,N_4846,N_4844);
nand U4959 (N_4959,N_4893,N_4851);
nand U4960 (N_4960,N_4893,N_4868);
nand U4961 (N_4961,N_4813,N_4811);
nor U4962 (N_4962,N_4864,N_4892);
xnor U4963 (N_4963,N_4899,N_4835);
and U4964 (N_4964,N_4809,N_4868);
and U4965 (N_4965,N_4856,N_4892);
nor U4966 (N_4966,N_4858,N_4874);
nand U4967 (N_4967,N_4825,N_4838);
and U4968 (N_4968,N_4872,N_4823);
xnor U4969 (N_4969,N_4889,N_4845);
xor U4970 (N_4970,N_4815,N_4811);
nand U4971 (N_4971,N_4839,N_4896);
nor U4972 (N_4972,N_4867,N_4815);
nand U4973 (N_4973,N_4874,N_4851);
or U4974 (N_4974,N_4871,N_4803);
nor U4975 (N_4975,N_4822,N_4818);
xor U4976 (N_4976,N_4816,N_4802);
or U4977 (N_4977,N_4814,N_4896);
nor U4978 (N_4978,N_4813,N_4829);
nand U4979 (N_4979,N_4839,N_4860);
or U4980 (N_4980,N_4899,N_4834);
nand U4981 (N_4981,N_4841,N_4858);
or U4982 (N_4982,N_4876,N_4859);
nand U4983 (N_4983,N_4868,N_4820);
or U4984 (N_4984,N_4801,N_4834);
nand U4985 (N_4985,N_4824,N_4839);
and U4986 (N_4986,N_4858,N_4849);
xor U4987 (N_4987,N_4883,N_4857);
nor U4988 (N_4988,N_4854,N_4860);
or U4989 (N_4989,N_4837,N_4843);
nor U4990 (N_4990,N_4860,N_4836);
nand U4991 (N_4991,N_4862,N_4863);
or U4992 (N_4992,N_4840,N_4828);
and U4993 (N_4993,N_4832,N_4833);
nor U4994 (N_4994,N_4852,N_4800);
xor U4995 (N_4995,N_4859,N_4870);
and U4996 (N_4996,N_4888,N_4872);
nand U4997 (N_4997,N_4839,N_4880);
nor U4998 (N_4998,N_4818,N_4863);
xor U4999 (N_4999,N_4814,N_4839);
or U5000 (N_5000,N_4970,N_4959);
or U5001 (N_5001,N_4962,N_4932);
and U5002 (N_5002,N_4966,N_4979);
nand U5003 (N_5003,N_4934,N_4928);
nand U5004 (N_5004,N_4999,N_4910);
and U5005 (N_5005,N_4946,N_4954);
nand U5006 (N_5006,N_4987,N_4929);
nand U5007 (N_5007,N_4920,N_4955);
xor U5008 (N_5008,N_4936,N_4939);
and U5009 (N_5009,N_4912,N_4996);
and U5010 (N_5010,N_4942,N_4958);
and U5011 (N_5011,N_4973,N_4991);
nand U5012 (N_5012,N_4989,N_4924);
nor U5013 (N_5013,N_4976,N_4919);
nor U5014 (N_5014,N_4963,N_4944);
xnor U5015 (N_5015,N_4974,N_4904);
nor U5016 (N_5016,N_4993,N_4906);
xor U5017 (N_5017,N_4941,N_4978);
nor U5018 (N_5018,N_4983,N_4950);
and U5019 (N_5019,N_4923,N_4971);
and U5020 (N_5020,N_4988,N_4949);
nand U5021 (N_5021,N_4933,N_4960);
nand U5022 (N_5022,N_4972,N_4922);
or U5023 (N_5023,N_4969,N_4965);
and U5024 (N_5024,N_4930,N_4994);
nor U5025 (N_5025,N_4967,N_4916);
nor U5026 (N_5026,N_4931,N_4926);
nor U5027 (N_5027,N_4913,N_4992);
xor U5028 (N_5028,N_4956,N_4945);
xnor U5029 (N_5029,N_4938,N_4902);
or U5030 (N_5030,N_4921,N_4903);
or U5031 (N_5031,N_4961,N_4935);
nor U5032 (N_5032,N_4900,N_4975);
or U5033 (N_5033,N_4943,N_4937);
nand U5034 (N_5034,N_4915,N_4901);
or U5035 (N_5035,N_4968,N_4948);
or U5036 (N_5036,N_4981,N_4947);
nor U5037 (N_5037,N_4917,N_4998);
nand U5038 (N_5038,N_4905,N_4927);
nand U5039 (N_5039,N_4995,N_4977);
nor U5040 (N_5040,N_4908,N_4985);
or U5041 (N_5041,N_4911,N_4952);
or U5042 (N_5042,N_4980,N_4997);
or U5043 (N_5043,N_4951,N_4907);
nor U5044 (N_5044,N_4940,N_4984);
or U5045 (N_5045,N_4990,N_4914);
nand U5046 (N_5046,N_4964,N_4909);
xor U5047 (N_5047,N_4957,N_4925);
nor U5048 (N_5048,N_4918,N_4986);
nand U5049 (N_5049,N_4982,N_4953);
or U5050 (N_5050,N_4949,N_4993);
xnor U5051 (N_5051,N_4978,N_4909);
or U5052 (N_5052,N_4902,N_4971);
xnor U5053 (N_5053,N_4909,N_4958);
and U5054 (N_5054,N_4911,N_4969);
xnor U5055 (N_5055,N_4958,N_4979);
nor U5056 (N_5056,N_4996,N_4998);
nor U5057 (N_5057,N_4940,N_4971);
nand U5058 (N_5058,N_4926,N_4924);
nor U5059 (N_5059,N_4949,N_4965);
nand U5060 (N_5060,N_4977,N_4974);
xnor U5061 (N_5061,N_4932,N_4969);
or U5062 (N_5062,N_4956,N_4994);
and U5063 (N_5063,N_4973,N_4916);
xnor U5064 (N_5064,N_4934,N_4925);
xor U5065 (N_5065,N_4917,N_4914);
or U5066 (N_5066,N_4980,N_4938);
nand U5067 (N_5067,N_4987,N_4933);
and U5068 (N_5068,N_4982,N_4925);
nand U5069 (N_5069,N_4937,N_4971);
or U5070 (N_5070,N_4928,N_4956);
and U5071 (N_5071,N_4908,N_4938);
and U5072 (N_5072,N_4922,N_4949);
nand U5073 (N_5073,N_4979,N_4943);
or U5074 (N_5074,N_4922,N_4955);
or U5075 (N_5075,N_4955,N_4990);
or U5076 (N_5076,N_4942,N_4947);
nand U5077 (N_5077,N_4913,N_4990);
or U5078 (N_5078,N_4910,N_4977);
and U5079 (N_5079,N_4911,N_4957);
nand U5080 (N_5080,N_4952,N_4988);
nand U5081 (N_5081,N_4931,N_4925);
xor U5082 (N_5082,N_4998,N_4923);
nor U5083 (N_5083,N_4956,N_4908);
and U5084 (N_5084,N_4952,N_4987);
and U5085 (N_5085,N_4954,N_4989);
xnor U5086 (N_5086,N_4938,N_4949);
or U5087 (N_5087,N_4912,N_4952);
nand U5088 (N_5088,N_4989,N_4918);
xor U5089 (N_5089,N_4912,N_4950);
nor U5090 (N_5090,N_4961,N_4971);
and U5091 (N_5091,N_4914,N_4935);
and U5092 (N_5092,N_4938,N_4907);
nor U5093 (N_5093,N_4969,N_4937);
nor U5094 (N_5094,N_4907,N_4968);
and U5095 (N_5095,N_4940,N_4916);
nand U5096 (N_5096,N_4934,N_4981);
nand U5097 (N_5097,N_4915,N_4983);
nor U5098 (N_5098,N_4921,N_4940);
and U5099 (N_5099,N_4924,N_4941);
nand U5100 (N_5100,N_5012,N_5035);
nor U5101 (N_5101,N_5064,N_5029);
nor U5102 (N_5102,N_5015,N_5051);
nor U5103 (N_5103,N_5037,N_5008);
and U5104 (N_5104,N_5007,N_5014);
or U5105 (N_5105,N_5092,N_5016);
or U5106 (N_5106,N_5020,N_5003);
nand U5107 (N_5107,N_5060,N_5077);
and U5108 (N_5108,N_5033,N_5063);
nand U5109 (N_5109,N_5040,N_5099);
nor U5110 (N_5110,N_5091,N_5072);
and U5111 (N_5111,N_5093,N_5088);
or U5112 (N_5112,N_5022,N_5076);
nand U5113 (N_5113,N_5041,N_5073);
nor U5114 (N_5114,N_5021,N_5011);
nor U5115 (N_5115,N_5081,N_5046);
nor U5116 (N_5116,N_5071,N_5098);
xnor U5117 (N_5117,N_5036,N_5004);
nand U5118 (N_5118,N_5026,N_5000);
xor U5119 (N_5119,N_5009,N_5048);
or U5120 (N_5120,N_5066,N_5018);
nor U5121 (N_5121,N_5034,N_5028);
nand U5122 (N_5122,N_5085,N_5049);
or U5123 (N_5123,N_5042,N_5094);
nand U5124 (N_5124,N_5044,N_5031);
nand U5125 (N_5125,N_5059,N_5079);
and U5126 (N_5126,N_5054,N_5083);
nand U5127 (N_5127,N_5017,N_5068);
or U5128 (N_5128,N_5043,N_5052);
nand U5129 (N_5129,N_5090,N_5013);
nor U5130 (N_5130,N_5010,N_5005);
or U5131 (N_5131,N_5070,N_5062);
nand U5132 (N_5132,N_5074,N_5024);
nor U5133 (N_5133,N_5058,N_5023);
nor U5134 (N_5134,N_5030,N_5089);
nor U5135 (N_5135,N_5084,N_5050);
and U5136 (N_5136,N_5047,N_5069);
nand U5137 (N_5137,N_5096,N_5075);
nor U5138 (N_5138,N_5025,N_5097);
or U5139 (N_5139,N_5080,N_5032);
nand U5140 (N_5140,N_5056,N_5086);
or U5141 (N_5141,N_5038,N_5039);
nand U5142 (N_5142,N_5082,N_5053);
nand U5143 (N_5143,N_5078,N_5006);
or U5144 (N_5144,N_5019,N_5002);
nor U5145 (N_5145,N_5095,N_5045);
and U5146 (N_5146,N_5027,N_5001);
or U5147 (N_5147,N_5061,N_5067);
nor U5148 (N_5148,N_5065,N_5055);
nor U5149 (N_5149,N_5087,N_5057);
and U5150 (N_5150,N_5052,N_5048);
nor U5151 (N_5151,N_5040,N_5080);
nand U5152 (N_5152,N_5038,N_5037);
nor U5153 (N_5153,N_5089,N_5051);
or U5154 (N_5154,N_5049,N_5001);
nand U5155 (N_5155,N_5070,N_5031);
or U5156 (N_5156,N_5028,N_5088);
or U5157 (N_5157,N_5019,N_5037);
nand U5158 (N_5158,N_5041,N_5011);
nand U5159 (N_5159,N_5033,N_5005);
and U5160 (N_5160,N_5026,N_5072);
nand U5161 (N_5161,N_5024,N_5009);
nand U5162 (N_5162,N_5062,N_5048);
nor U5163 (N_5163,N_5049,N_5007);
and U5164 (N_5164,N_5068,N_5083);
nor U5165 (N_5165,N_5027,N_5026);
or U5166 (N_5166,N_5025,N_5088);
nand U5167 (N_5167,N_5004,N_5097);
and U5168 (N_5168,N_5057,N_5044);
and U5169 (N_5169,N_5074,N_5038);
and U5170 (N_5170,N_5045,N_5072);
nor U5171 (N_5171,N_5090,N_5062);
nand U5172 (N_5172,N_5072,N_5046);
nand U5173 (N_5173,N_5045,N_5059);
nor U5174 (N_5174,N_5040,N_5007);
nand U5175 (N_5175,N_5026,N_5087);
xor U5176 (N_5176,N_5008,N_5061);
nand U5177 (N_5177,N_5017,N_5023);
or U5178 (N_5178,N_5021,N_5036);
and U5179 (N_5179,N_5049,N_5058);
nor U5180 (N_5180,N_5062,N_5059);
or U5181 (N_5181,N_5055,N_5033);
and U5182 (N_5182,N_5054,N_5007);
nor U5183 (N_5183,N_5029,N_5018);
nor U5184 (N_5184,N_5006,N_5033);
nor U5185 (N_5185,N_5099,N_5021);
nand U5186 (N_5186,N_5005,N_5053);
or U5187 (N_5187,N_5030,N_5016);
xor U5188 (N_5188,N_5095,N_5004);
and U5189 (N_5189,N_5018,N_5058);
xnor U5190 (N_5190,N_5056,N_5032);
or U5191 (N_5191,N_5050,N_5075);
nand U5192 (N_5192,N_5059,N_5017);
nor U5193 (N_5193,N_5006,N_5052);
nand U5194 (N_5194,N_5074,N_5011);
nand U5195 (N_5195,N_5082,N_5080);
xor U5196 (N_5196,N_5048,N_5008);
nand U5197 (N_5197,N_5022,N_5052);
xnor U5198 (N_5198,N_5082,N_5091);
or U5199 (N_5199,N_5077,N_5082);
and U5200 (N_5200,N_5158,N_5185);
and U5201 (N_5201,N_5155,N_5181);
or U5202 (N_5202,N_5145,N_5100);
nand U5203 (N_5203,N_5178,N_5135);
and U5204 (N_5204,N_5180,N_5121);
and U5205 (N_5205,N_5140,N_5183);
and U5206 (N_5206,N_5136,N_5137);
nor U5207 (N_5207,N_5191,N_5119);
or U5208 (N_5208,N_5130,N_5133);
nand U5209 (N_5209,N_5126,N_5115);
and U5210 (N_5210,N_5192,N_5188);
and U5211 (N_5211,N_5189,N_5176);
and U5212 (N_5212,N_5195,N_5156);
and U5213 (N_5213,N_5109,N_5184);
nand U5214 (N_5214,N_5108,N_5179);
nand U5215 (N_5215,N_5163,N_5177);
and U5216 (N_5216,N_5152,N_5132);
and U5217 (N_5217,N_5101,N_5138);
nor U5218 (N_5218,N_5154,N_5199);
and U5219 (N_5219,N_5141,N_5198);
nor U5220 (N_5220,N_5175,N_5165);
and U5221 (N_5221,N_5187,N_5167);
nor U5222 (N_5222,N_5116,N_5129);
and U5223 (N_5223,N_5131,N_5194);
nand U5224 (N_5224,N_5147,N_5146);
xor U5225 (N_5225,N_5150,N_5151);
or U5226 (N_5226,N_5190,N_5124);
nor U5227 (N_5227,N_5114,N_5159);
xor U5228 (N_5228,N_5197,N_5127);
nand U5229 (N_5229,N_5161,N_5144);
nor U5230 (N_5230,N_5166,N_5106);
xnor U5231 (N_5231,N_5170,N_5193);
nand U5232 (N_5232,N_5168,N_5157);
nand U5233 (N_5233,N_5196,N_5111);
and U5234 (N_5234,N_5186,N_5103);
nand U5235 (N_5235,N_5107,N_5118);
nor U5236 (N_5236,N_5153,N_5122);
nor U5237 (N_5237,N_5105,N_5160);
or U5238 (N_5238,N_5174,N_5169);
nor U5239 (N_5239,N_5123,N_5112);
nand U5240 (N_5240,N_5143,N_5149);
and U5241 (N_5241,N_5128,N_5162);
and U5242 (N_5242,N_5139,N_5182);
and U5243 (N_5243,N_5120,N_5117);
nand U5244 (N_5244,N_5113,N_5102);
nor U5245 (N_5245,N_5171,N_5142);
or U5246 (N_5246,N_5134,N_5173);
or U5247 (N_5247,N_5172,N_5104);
and U5248 (N_5248,N_5125,N_5164);
or U5249 (N_5249,N_5148,N_5110);
nand U5250 (N_5250,N_5194,N_5137);
nand U5251 (N_5251,N_5147,N_5188);
nand U5252 (N_5252,N_5126,N_5186);
nor U5253 (N_5253,N_5167,N_5193);
and U5254 (N_5254,N_5158,N_5111);
nor U5255 (N_5255,N_5141,N_5112);
or U5256 (N_5256,N_5136,N_5162);
nor U5257 (N_5257,N_5104,N_5183);
nor U5258 (N_5258,N_5175,N_5162);
and U5259 (N_5259,N_5110,N_5177);
or U5260 (N_5260,N_5133,N_5189);
or U5261 (N_5261,N_5165,N_5147);
nor U5262 (N_5262,N_5180,N_5161);
nor U5263 (N_5263,N_5173,N_5146);
nor U5264 (N_5264,N_5177,N_5157);
or U5265 (N_5265,N_5152,N_5194);
and U5266 (N_5266,N_5149,N_5127);
and U5267 (N_5267,N_5117,N_5138);
nor U5268 (N_5268,N_5169,N_5102);
or U5269 (N_5269,N_5127,N_5159);
nor U5270 (N_5270,N_5149,N_5138);
nand U5271 (N_5271,N_5118,N_5125);
and U5272 (N_5272,N_5168,N_5131);
xor U5273 (N_5273,N_5199,N_5123);
nor U5274 (N_5274,N_5164,N_5185);
nand U5275 (N_5275,N_5123,N_5107);
and U5276 (N_5276,N_5143,N_5168);
or U5277 (N_5277,N_5156,N_5146);
and U5278 (N_5278,N_5196,N_5113);
nand U5279 (N_5279,N_5113,N_5197);
nor U5280 (N_5280,N_5162,N_5146);
nand U5281 (N_5281,N_5153,N_5176);
or U5282 (N_5282,N_5116,N_5132);
nand U5283 (N_5283,N_5179,N_5119);
nand U5284 (N_5284,N_5169,N_5164);
and U5285 (N_5285,N_5148,N_5105);
nand U5286 (N_5286,N_5164,N_5186);
nand U5287 (N_5287,N_5144,N_5183);
xnor U5288 (N_5288,N_5194,N_5101);
xnor U5289 (N_5289,N_5104,N_5126);
and U5290 (N_5290,N_5197,N_5169);
and U5291 (N_5291,N_5179,N_5185);
nand U5292 (N_5292,N_5116,N_5177);
or U5293 (N_5293,N_5126,N_5114);
nand U5294 (N_5294,N_5172,N_5115);
or U5295 (N_5295,N_5124,N_5110);
nand U5296 (N_5296,N_5158,N_5183);
xnor U5297 (N_5297,N_5127,N_5105);
and U5298 (N_5298,N_5163,N_5183);
nand U5299 (N_5299,N_5170,N_5124);
nand U5300 (N_5300,N_5240,N_5205);
or U5301 (N_5301,N_5202,N_5220);
or U5302 (N_5302,N_5216,N_5254);
and U5303 (N_5303,N_5292,N_5289);
nor U5304 (N_5304,N_5239,N_5219);
or U5305 (N_5305,N_5266,N_5253);
and U5306 (N_5306,N_5234,N_5256);
and U5307 (N_5307,N_5291,N_5246);
and U5308 (N_5308,N_5248,N_5238);
and U5309 (N_5309,N_5299,N_5257);
nand U5310 (N_5310,N_5213,N_5290);
nor U5311 (N_5311,N_5277,N_5222);
nand U5312 (N_5312,N_5286,N_5279);
or U5313 (N_5313,N_5288,N_5227);
and U5314 (N_5314,N_5261,N_5235);
nand U5315 (N_5315,N_5224,N_5226);
nor U5316 (N_5316,N_5260,N_5287);
and U5317 (N_5317,N_5280,N_5236);
nor U5318 (N_5318,N_5283,N_5278);
nand U5319 (N_5319,N_5200,N_5263);
or U5320 (N_5320,N_5217,N_5255);
and U5321 (N_5321,N_5230,N_5237);
nand U5322 (N_5322,N_5271,N_5242);
nor U5323 (N_5323,N_5294,N_5259);
nor U5324 (N_5324,N_5282,N_5214);
nor U5325 (N_5325,N_5251,N_5258);
xor U5326 (N_5326,N_5252,N_5250);
and U5327 (N_5327,N_5229,N_5274);
nor U5328 (N_5328,N_5262,N_5233);
nand U5329 (N_5329,N_5296,N_5204);
nand U5330 (N_5330,N_5209,N_5211);
or U5331 (N_5331,N_5212,N_5245);
nand U5332 (N_5332,N_5223,N_5297);
and U5333 (N_5333,N_5218,N_5243);
nand U5334 (N_5334,N_5293,N_5281);
nor U5335 (N_5335,N_5270,N_5208);
xnor U5336 (N_5336,N_5249,N_5269);
and U5337 (N_5337,N_5265,N_5225);
and U5338 (N_5338,N_5215,N_5268);
nor U5339 (N_5339,N_5201,N_5206);
and U5340 (N_5340,N_5275,N_5221);
nor U5341 (N_5341,N_5207,N_5231);
and U5342 (N_5342,N_5264,N_5232);
nor U5343 (N_5343,N_5247,N_5284);
nor U5344 (N_5344,N_5267,N_5244);
nand U5345 (N_5345,N_5276,N_5241);
nand U5346 (N_5346,N_5298,N_5210);
or U5347 (N_5347,N_5285,N_5228);
or U5348 (N_5348,N_5272,N_5273);
or U5349 (N_5349,N_5295,N_5203);
nor U5350 (N_5350,N_5227,N_5274);
nor U5351 (N_5351,N_5248,N_5274);
nor U5352 (N_5352,N_5258,N_5209);
nand U5353 (N_5353,N_5212,N_5228);
nand U5354 (N_5354,N_5267,N_5200);
nor U5355 (N_5355,N_5236,N_5229);
nor U5356 (N_5356,N_5241,N_5278);
nor U5357 (N_5357,N_5200,N_5221);
and U5358 (N_5358,N_5271,N_5244);
or U5359 (N_5359,N_5269,N_5243);
nand U5360 (N_5360,N_5294,N_5222);
or U5361 (N_5361,N_5298,N_5261);
and U5362 (N_5362,N_5244,N_5277);
nand U5363 (N_5363,N_5210,N_5231);
or U5364 (N_5364,N_5233,N_5247);
nand U5365 (N_5365,N_5276,N_5260);
nand U5366 (N_5366,N_5274,N_5270);
and U5367 (N_5367,N_5296,N_5213);
nor U5368 (N_5368,N_5295,N_5241);
and U5369 (N_5369,N_5281,N_5296);
or U5370 (N_5370,N_5282,N_5226);
or U5371 (N_5371,N_5242,N_5273);
and U5372 (N_5372,N_5206,N_5226);
nor U5373 (N_5373,N_5273,N_5276);
nand U5374 (N_5374,N_5204,N_5268);
or U5375 (N_5375,N_5226,N_5213);
nand U5376 (N_5376,N_5203,N_5278);
and U5377 (N_5377,N_5290,N_5208);
or U5378 (N_5378,N_5258,N_5205);
and U5379 (N_5379,N_5299,N_5281);
or U5380 (N_5380,N_5298,N_5209);
and U5381 (N_5381,N_5293,N_5282);
nand U5382 (N_5382,N_5202,N_5246);
nor U5383 (N_5383,N_5235,N_5214);
and U5384 (N_5384,N_5227,N_5248);
xnor U5385 (N_5385,N_5279,N_5262);
or U5386 (N_5386,N_5260,N_5277);
or U5387 (N_5387,N_5288,N_5237);
nand U5388 (N_5388,N_5220,N_5212);
nor U5389 (N_5389,N_5286,N_5267);
and U5390 (N_5390,N_5261,N_5249);
nor U5391 (N_5391,N_5282,N_5218);
and U5392 (N_5392,N_5261,N_5226);
or U5393 (N_5393,N_5245,N_5213);
or U5394 (N_5394,N_5279,N_5255);
and U5395 (N_5395,N_5271,N_5275);
and U5396 (N_5396,N_5235,N_5255);
and U5397 (N_5397,N_5232,N_5293);
and U5398 (N_5398,N_5226,N_5203);
nand U5399 (N_5399,N_5296,N_5295);
or U5400 (N_5400,N_5352,N_5382);
nor U5401 (N_5401,N_5355,N_5376);
nand U5402 (N_5402,N_5305,N_5307);
nand U5403 (N_5403,N_5322,N_5351);
nor U5404 (N_5404,N_5385,N_5344);
or U5405 (N_5405,N_5340,N_5363);
or U5406 (N_5406,N_5362,N_5333);
and U5407 (N_5407,N_5336,N_5373);
or U5408 (N_5408,N_5330,N_5323);
nor U5409 (N_5409,N_5306,N_5301);
nor U5410 (N_5410,N_5315,N_5387);
xnor U5411 (N_5411,N_5347,N_5337);
or U5412 (N_5412,N_5316,N_5318);
nor U5413 (N_5413,N_5331,N_5324);
and U5414 (N_5414,N_5356,N_5369);
or U5415 (N_5415,N_5320,N_5358);
xnor U5416 (N_5416,N_5371,N_5321);
nand U5417 (N_5417,N_5364,N_5309);
nor U5418 (N_5418,N_5393,N_5370);
and U5419 (N_5419,N_5326,N_5327);
nand U5420 (N_5420,N_5391,N_5346);
xnor U5421 (N_5421,N_5317,N_5349);
nand U5422 (N_5422,N_5394,N_5313);
and U5423 (N_5423,N_5314,N_5392);
nand U5424 (N_5424,N_5374,N_5396);
nor U5425 (N_5425,N_5341,N_5357);
and U5426 (N_5426,N_5365,N_5380);
and U5427 (N_5427,N_5384,N_5367);
nand U5428 (N_5428,N_5303,N_5383);
xor U5429 (N_5429,N_5348,N_5353);
and U5430 (N_5430,N_5312,N_5311);
nor U5431 (N_5431,N_5381,N_5388);
nand U5432 (N_5432,N_5354,N_5310);
nor U5433 (N_5433,N_5338,N_5372);
or U5434 (N_5434,N_5304,N_5345);
or U5435 (N_5435,N_5377,N_5334);
or U5436 (N_5436,N_5332,N_5359);
nor U5437 (N_5437,N_5343,N_5389);
and U5438 (N_5438,N_5325,N_5366);
nor U5439 (N_5439,N_5379,N_5375);
or U5440 (N_5440,N_5361,N_5378);
and U5441 (N_5441,N_5386,N_5397);
nand U5442 (N_5442,N_5398,N_5342);
nor U5443 (N_5443,N_5368,N_5302);
and U5444 (N_5444,N_5300,N_5350);
nor U5445 (N_5445,N_5329,N_5335);
or U5446 (N_5446,N_5339,N_5390);
xnor U5447 (N_5447,N_5399,N_5395);
nand U5448 (N_5448,N_5328,N_5308);
and U5449 (N_5449,N_5319,N_5360);
or U5450 (N_5450,N_5383,N_5367);
xor U5451 (N_5451,N_5355,N_5325);
or U5452 (N_5452,N_5375,N_5333);
nand U5453 (N_5453,N_5366,N_5321);
nor U5454 (N_5454,N_5318,N_5304);
or U5455 (N_5455,N_5328,N_5336);
nand U5456 (N_5456,N_5383,N_5397);
nand U5457 (N_5457,N_5325,N_5345);
nor U5458 (N_5458,N_5395,N_5397);
and U5459 (N_5459,N_5319,N_5378);
or U5460 (N_5460,N_5375,N_5382);
nand U5461 (N_5461,N_5345,N_5314);
nor U5462 (N_5462,N_5365,N_5378);
nand U5463 (N_5463,N_5357,N_5301);
nor U5464 (N_5464,N_5399,N_5315);
nand U5465 (N_5465,N_5376,N_5319);
nand U5466 (N_5466,N_5345,N_5319);
xnor U5467 (N_5467,N_5302,N_5374);
and U5468 (N_5468,N_5343,N_5312);
or U5469 (N_5469,N_5306,N_5379);
xnor U5470 (N_5470,N_5371,N_5301);
or U5471 (N_5471,N_5382,N_5398);
nand U5472 (N_5472,N_5392,N_5374);
and U5473 (N_5473,N_5346,N_5324);
xnor U5474 (N_5474,N_5378,N_5362);
or U5475 (N_5475,N_5348,N_5318);
and U5476 (N_5476,N_5357,N_5302);
nand U5477 (N_5477,N_5356,N_5335);
nor U5478 (N_5478,N_5363,N_5385);
nand U5479 (N_5479,N_5324,N_5348);
and U5480 (N_5480,N_5333,N_5376);
nor U5481 (N_5481,N_5391,N_5392);
and U5482 (N_5482,N_5341,N_5325);
or U5483 (N_5483,N_5315,N_5329);
and U5484 (N_5484,N_5307,N_5333);
and U5485 (N_5485,N_5342,N_5355);
and U5486 (N_5486,N_5317,N_5338);
nand U5487 (N_5487,N_5304,N_5320);
or U5488 (N_5488,N_5317,N_5303);
nor U5489 (N_5489,N_5386,N_5341);
or U5490 (N_5490,N_5336,N_5358);
nor U5491 (N_5491,N_5317,N_5322);
and U5492 (N_5492,N_5388,N_5399);
xnor U5493 (N_5493,N_5365,N_5341);
xor U5494 (N_5494,N_5353,N_5380);
and U5495 (N_5495,N_5307,N_5337);
nand U5496 (N_5496,N_5346,N_5348);
nand U5497 (N_5497,N_5373,N_5308);
and U5498 (N_5498,N_5369,N_5383);
and U5499 (N_5499,N_5379,N_5359);
or U5500 (N_5500,N_5441,N_5460);
nand U5501 (N_5501,N_5450,N_5415);
nand U5502 (N_5502,N_5459,N_5428);
nor U5503 (N_5503,N_5482,N_5463);
and U5504 (N_5504,N_5418,N_5453);
nand U5505 (N_5505,N_5483,N_5477);
or U5506 (N_5506,N_5436,N_5402);
or U5507 (N_5507,N_5461,N_5403);
nand U5508 (N_5508,N_5433,N_5478);
or U5509 (N_5509,N_5407,N_5490);
or U5510 (N_5510,N_5462,N_5493);
xor U5511 (N_5511,N_5476,N_5409);
nand U5512 (N_5512,N_5425,N_5467);
nand U5513 (N_5513,N_5455,N_5444);
xor U5514 (N_5514,N_5429,N_5439);
nor U5515 (N_5515,N_5473,N_5468);
nand U5516 (N_5516,N_5454,N_5445);
nor U5517 (N_5517,N_5422,N_5497);
or U5518 (N_5518,N_5481,N_5452);
xor U5519 (N_5519,N_5484,N_5492);
nor U5520 (N_5520,N_5432,N_5440);
and U5521 (N_5521,N_5491,N_5437);
xor U5522 (N_5522,N_5417,N_5430);
or U5523 (N_5523,N_5400,N_5413);
and U5524 (N_5524,N_5485,N_5488);
and U5525 (N_5525,N_5495,N_5466);
and U5526 (N_5526,N_5426,N_5470);
nand U5527 (N_5527,N_5465,N_5406);
nand U5528 (N_5528,N_5457,N_5448);
or U5529 (N_5529,N_5486,N_5414);
or U5530 (N_5530,N_5411,N_5410);
or U5531 (N_5531,N_5449,N_5489);
nand U5532 (N_5532,N_5472,N_5464);
and U5533 (N_5533,N_5442,N_5401);
or U5534 (N_5534,N_5458,N_5435);
and U5535 (N_5535,N_5479,N_5420);
nor U5536 (N_5536,N_5456,N_5416);
or U5537 (N_5537,N_5405,N_5424);
xnor U5538 (N_5538,N_5427,N_5431);
or U5539 (N_5539,N_5471,N_5412);
nand U5540 (N_5540,N_5404,N_5408);
xnor U5541 (N_5541,N_5480,N_5446);
xnor U5542 (N_5542,N_5421,N_5434);
nor U5543 (N_5543,N_5494,N_5474);
nand U5544 (N_5544,N_5499,N_5469);
and U5545 (N_5545,N_5419,N_5487);
xnor U5546 (N_5546,N_5475,N_5423);
xor U5547 (N_5547,N_5498,N_5447);
nor U5548 (N_5548,N_5496,N_5443);
nor U5549 (N_5549,N_5438,N_5451);
xor U5550 (N_5550,N_5428,N_5448);
nand U5551 (N_5551,N_5440,N_5485);
or U5552 (N_5552,N_5459,N_5498);
nor U5553 (N_5553,N_5451,N_5406);
or U5554 (N_5554,N_5420,N_5451);
nand U5555 (N_5555,N_5412,N_5480);
and U5556 (N_5556,N_5473,N_5484);
and U5557 (N_5557,N_5477,N_5450);
or U5558 (N_5558,N_5426,N_5493);
nand U5559 (N_5559,N_5428,N_5419);
nand U5560 (N_5560,N_5403,N_5479);
nor U5561 (N_5561,N_5459,N_5468);
or U5562 (N_5562,N_5453,N_5490);
nand U5563 (N_5563,N_5467,N_5483);
or U5564 (N_5564,N_5471,N_5470);
nand U5565 (N_5565,N_5419,N_5468);
xnor U5566 (N_5566,N_5473,N_5410);
nand U5567 (N_5567,N_5467,N_5419);
nand U5568 (N_5568,N_5498,N_5481);
nor U5569 (N_5569,N_5490,N_5479);
or U5570 (N_5570,N_5430,N_5450);
or U5571 (N_5571,N_5452,N_5464);
or U5572 (N_5572,N_5498,N_5451);
nor U5573 (N_5573,N_5480,N_5401);
or U5574 (N_5574,N_5458,N_5447);
nor U5575 (N_5575,N_5493,N_5499);
xnor U5576 (N_5576,N_5423,N_5415);
nand U5577 (N_5577,N_5472,N_5431);
nand U5578 (N_5578,N_5473,N_5442);
and U5579 (N_5579,N_5440,N_5489);
or U5580 (N_5580,N_5450,N_5465);
nand U5581 (N_5581,N_5461,N_5404);
or U5582 (N_5582,N_5425,N_5468);
xnor U5583 (N_5583,N_5450,N_5443);
nand U5584 (N_5584,N_5401,N_5444);
nor U5585 (N_5585,N_5402,N_5447);
xor U5586 (N_5586,N_5434,N_5451);
and U5587 (N_5587,N_5480,N_5439);
nor U5588 (N_5588,N_5496,N_5454);
or U5589 (N_5589,N_5419,N_5426);
nand U5590 (N_5590,N_5484,N_5434);
or U5591 (N_5591,N_5449,N_5436);
or U5592 (N_5592,N_5497,N_5485);
nor U5593 (N_5593,N_5417,N_5487);
or U5594 (N_5594,N_5467,N_5430);
or U5595 (N_5595,N_5473,N_5446);
nand U5596 (N_5596,N_5438,N_5452);
nor U5597 (N_5597,N_5407,N_5435);
nor U5598 (N_5598,N_5494,N_5406);
nand U5599 (N_5599,N_5482,N_5412);
and U5600 (N_5600,N_5565,N_5538);
or U5601 (N_5601,N_5580,N_5573);
xor U5602 (N_5602,N_5570,N_5562);
and U5603 (N_5603,N_5589,N_5514);
and U5604 (N_5604,N_5586,N_5579);
nor U5605 (N_5605,N_5509,N_5571);
and U5606 (N_5606,N_5569,N_5581);
or U5607 (N_5607,N_5525,N_5556);
and U5608 (N_5608,N_5541,N_5521);
nand U5609 (N_5609,N_5552,N_5540);
and U5610 (N_5610,N_5504,N_5575);
or U5611 (N_5611,N_5577,N_5587);
nor U5612 (N_5612,N_5548,N_5537);
and U5613 (N_5613,N_5501,N_5524);
or U5614 (N_5614,N_5584,N_5512);
and U5615 (N_5615,N_5555,N_5561);
and U5616 (N_5616,N_5545,N_5516);
nand U5617 (N_5617,N_5526,N_5593);
nor U5618 (N_5618,N_5583,N_5544);
nor U5619 (N_5619,N_5542,N_5513);
nor U5620 (N_5620,N_5506,N_5592);
and U5621 (N_5621,N_5595,N_5527);
xor U5622 (N_5622,N_5567,N_5528);
and U5623 (N_5623,N_5517,N_5503);
and U5624 (N_5624,N_5563,N_5550);
xnor U5625 (N_5625,N_5549,N_5536);
nor U5626 (N_5626,N_5520,N_5554);
nor U5627 (N_5627,N_5560,N_5599);
or U5628 (N_5628,N_5574,N_5553);
or U5629 (N_5629,N_5551,N_5529);
nor U5630 (N_5630,N_5511,N_5547);
nor U5631 (N_5631,N_5585,N_5535);
or U5632 (N_5632,N_5558,N_5596);
xor U5633 (N_5633,N_5588,N_5543);
and U5634 (N_5634,N_5572,N_5559);
or U5635 (N_5635,N_5576,N_5507);
nor U5636 (N_5636,N_5598,N_5531);
or U5637 (N_5637,N_5568,N_5539);
xor U5638 (N_5638,N_5508,N_5523);
nor U5639 (N_5639,N_5502,N_5522);
nor U5640 (N_5640,N_5505,N_5566);
and U5641 (N_5641,N_5557,N_5530);
nor U5642 (N_5642,N_5519,N_5597);
nor U5643 (N_5643,N_5515,N_5532);
nor U5644 (N_5644,N_5591,N_5518);
xnor U5645 (N_5645,N_5533,N_5546);
or U5646 (N_5646,N_5590,N_5594);
nand U5647 (N_5647,N_5578,N_5564);
and U5648 (N_5648,N_5534,N_5500);
or U5649 (N_5649,N_5582,N_5510);
xnor U5650 (N_5650,N_5579,N_5551);
and U5651 (N_5651,N_5526,N_5523);
or U5652 (N_5652,N_5589,N_5585);
nand U5653 (N_5653,N_5520,N_5533);
or U5654 (N_5654,N_5520,N_5555);
xor U5655 (N_5655,N_5527,N_5537);
nand U5656 (N_5656,N_5579,N_5567);
nor U5657 (N_5657,N_5587,N_5523);
xor U5658 (N_5658,N_5572,N_5592);
or U5659 (N_5659,N_5586,N_5519);
and U5660 (N_5660,N_5535,N_5520);
nor U5661 (N_5661,N_5524,N_5555);
or U5662 (N_5662,N_5571,N_5525);
nand U5663 (N_5663,N_5548,N_5594);
nor U5664 (N_5664,N_5580,N_5595);
nand U5665 (N_5665,N_5519,N_5549);
nand U5666 (N_5666,N_5595,N_5544);
nor U5667 (N_5667,N_5569,N_5562);
or U5668 (N_5668,N_5521,N_5576);
and U5669 (N_5669,N_5500,N_5517);
and U5670 (N_5670,N_5584,N_5583);
and U5671 (N_5671,N_5577,N_5500);
and U5672 (N_5672,N_5514,N_5556);
xnor U5673 (N_5673,N_5547,N_5579);
nor U5674 (N_5674,N_5516,N_5503);
nand U5675 (N_5675,N_5567,N_5565);
nor U5676 (N_5676,N_5569,N_5559);
and U5677 (N_5677,N_5547,N_5598);
and U5678 (N_5678,N_5530,N_5512);
nor U5679 (N_5679,N_5528,N_5561);
or U5680 (N_5680,N_5588,N_5533);
nand U5681 (N_5681,N_5520,N_5567);
nor U5682 (N_5682,N_5512,N_5533);
nor U5683 (N_5683,N_5552,N_5597);
nor U5684 (N_5684,N_5559,N_5534);
nand U5685 (N_5685,N_5503,N_5559);
nand U5686 (N_5686,N_5595,N_5532);
nor U5687 (N_5687,N_5522,N_5557);
nand U5688 (N_5688,N_5533,N_5553);
nor U5689 (N_5689,N_5560,N_5526);
and U5690 (N_5690,N_5529,N_5537);
and U5691 (N_5691,N_5593,N_5506);
and U5692 (N_5692,N_5590,N_5550);
nand U5693 (N_5693,N_5591,N_5540);
xnor U5694 (N_5694,N_5544,N_5525);
nand U5695 (N_5695,N_5500,N_5556);
and U5696 (N_5696,N_5501,N_5526);
nor U5697 (N_5697,N_5533,N_5593);
nand U5698 (N_5698,N_5544,N_5533);
nand U5699 (N_5699,N_5596,N_5518);
nor U5700 (N_5700,N_5645,N_5661);
and U5701 (N_5701,N_5604,N_5664);
xnor U5702 (N_5702,N_5668,N_5606);
nor U5703 (N_5703,N_5696,N_5638);
or U5704 (N_5704,N_5609,N_5680);
and U5705 (N_5705,N_5683,N_5621);
and U5706 (N_5706,N_5630,N_5692);
and U5707 (N_5707,N_5602,N_5667);
xor U5708 (N_5708,N_5626,N_5611);
nor U5709 (N_5709,N_5655,N_5649);
and U5710 (N_5710,N_5628,N_5601);
nor U5711 (N_5711,N_5669,N_5637);
nor U5712 (N_5712,N_5625,N_5691);
or U5713 (N_5713,N_5616,N_5644);
nor U5714 (N_5714,N_5643,N_5663);
or U5715 (N_5715,N_5660,N_5627);
nor U5716 (N_5716,N_5646,N_5685);
and U5717 (N_5717,N_5613,N_5658);
and U5718 (N_5718,N_5670,N_5615);
and U5719 (N_5719,N_5686,N_5673);
nand U5720 (N_5720,N_5687,N_5652);
xor U5721 (N_5721,N_5694,N_5607);
and U5722 (N_5722,N_5647,N_5682);
nor U5723 (N_5723,N_5632,N_5600);
nor U5724 (N_5724,N_5642,N_5614);
or U5725 (N_5725,N_5612,N_5698);
nor U5726 (N_5726,N_5631,N_5674);
or U5727 (N_5727,N_5623,N_5666);
nor U5728 (N_5728,N_5617,N_5639);
and U5729 (N_5729,N_5681,N_5605);
nand U5730 (N_5730,N_5689,N_5672);
nor U5731 (N_5731,N_5690,N_5640);
and U5732 (N_5732,N_5679,N_5656);
or U5733 (N_5733,N_5675,N_5618);
xnor U5734 (N_5734,N_5654,N_5678);
and U5735 (N_5735,N_5695,N_5629);
nand U5736 (N_5736,N_5619,N_5651);
nor U5737 (N_5737,N_5662,N_5653);
and U5738 (N_5738,N_5699,N_5624);
nand U5739 (N_5739,N_5603,N_5677);
nor U5740 (N_5740,N_5610,N_5671);
or U5741 (N_5741,N_5608,N_5665);
nand U5742 (N_5742,N_5620,N_5650);
xor U5743 (N_5743,N_5622,N_5636);
xor U5744 (N_5744,N_5684,N_5633);
xor U5745 (N_5745,N_5676,N_5659);
and U5746 (N_5746,N_5697,N_5648);
xor U5747 (N_5747,N_5688,N_5635);
or U5748 (N_5748,N_5693,N_5657);
or U5749 (N_5749,N_5641,N_5634);
nor U5750 (N_5750,N_5674,N_5694);
and U5751 (N_5751,N_5686,N_5636);
and U5752 (N_5752,N_5619,N_5653);
nor U5753 (N_5753,N_5644,N_5605);
nor U5754 (N_5754,N_5661,N_5696);
xor U5755 (N_5755,N_5634,N_5671);
nand U5756 (N_5756,N_5615,N_5618);
and U5757 (N_5757,N_5658,N_5657);
and U5758 (N_5758,N_5635,N_5623);
or U5759 (N_5759,N_5660,N_5614);
nor U5760 (N_5760,N_5620,N_5691);
and U5761 (N_5761,N_5618,N_5653);
nor U5762 (N_5762,N_5659,N_5674);
or U5763 (N_5763,N_5679,N_5653);
nand U5764 (N_5764,N_5628,N_5624);
and U5765 (N_5765,N_5689,N_5680);
nand U5766 (N_5766,N_5603,N_5611);
nand U5767 (N_5767,N_5608,N_5650);
and U5768 (N_5768,N_5651,N_5695);
or U5769 (N_5769,N_5674,N_5690);
xnor U5770 (N_5770,N_5646,N_5689);
xnor U5771 (N_5771,N_5636,N_5613);
nand U5772 (N_5772,N_5674,N_5688);
or U5773 (N_5773,N_5611,N_5621);
xnor U5774 (N_5774,N_5662,N_5618);
nor U5775 (N_5775,N_5674,N_5661);
xor U5776 (N_5776,N_5624,N_5679);
xor U5777 (N_5777,N_5671,N_5679);
nor U5778 (N_5778,N_5657,N_5672);
or U5779 (N_5779,N_5692,N_5625);
nand U5780 (N_5780,N_5684,N_5631);
nand U5781 (N_5781,N_5686,N_5690);
or U5782 (N_5782,N_5686,N_5613);
nand U5783 (N_5783,N_5647,N_5680);
or U5784 (N_5784,N_5624,N_5636);
nand U5785 (N_5785,N_5659,N_5623);
and U5786 (N_5786,N_5621,N_5629);
or U5787 (N_5787,N_5659,N_5608);
xnor U5788 (N_5788,N_5617,N_5687);
and U5789 (N_5789,N_5680,N_5602);
and U5790 (N_5790,N_5699,N_5664);
nor U5791 (N_5791,N_5613,N_5632);
nor U5792 (N_5792,N_5694,N_5633);
nand U5793 (N_5793,N_5650,N_5659);
and U5794 (N_5794,N_5690,N_5644);
nand U5795 (N_5795,N_5629,N_5691);
and U5796 (N_5796,N_5644,N_5631);
and U5797 (N_5797,N_5664,N_5612);
nand U5798 (N_5798,N_5627,N_5606);
nor U5799 (N_5799,N_5646,N_5630);
xor U5800 (N_5800,N_5755,N_5717);
nor U5801 (N_5801,N_5792,N_5732);
nand U5802 (N_5802,N_5791,N_5761);
nor U5803 (N_5803,N_5733,N_5746);
xor U5804 (N_5804,N_5745,N_5797);
and U5805 (N_5805,N_5780,N_5721);
and U5806 (N_5806,N_5757,N_5712);
nor U5807 (N_5807,N_5771,N_5747);
nand U5808 (N_5808,N_5726,N_5783);
nand U5809 (N_5809,N_5725,N_5795);
xnor U5810 (N_5810,N_5704,N_5716);
nand U5811 (N_5811,N_5772,N_5768);
or U5812 (N_5812,N_5765,N_5727);
nor U5813 (N_5813,N_5754,N_5782);
or U5814 (N_5814,N_5731,N_5713);
or U5815 (N_5815,N_5769,N_5784);
and U5816 (N_5816,N_5734,N_5705);
xnor U5817 (N_5817,N_5711,N_5728);
or U5818 (N_5818,N_5750,N_5796);
xor U5819 (N_5819,N_5789,N_5798);
or U5820 (N_5820,N_5703,N_5777);
nand U5821 (N_5821,N_5785,N_5781);
nand U5822 (N_5822,N_5762,N_5756);
nand U5823 (N_5823,N_5707,N_5776);
and U5824 (N_5824,N_5770,N_5706);
or U5825 (N_5825,N_5786,N_5758);
and U5826 (N_5826,N_5775,N_5740);
nand U5827 (N_5827,N_5719,N_5752);
and U5828 (N_5828,N_5701,N_5736);
xnor U5829 (N_5829,N_5709,N_5738);
xnor U5830 (N_5830,N_5766,N_5723);
nand U5831 (N_5831,N_5773,N_5729);
nor U5832 (N_5832,N_5735,N_5759);
or U5833 (N_5833,N_5799,N_5751);
nor U5834 (N_5834,N_5708,N_5737);
nor U5835 (N_5835,N_5767,N_5718);
xnor U5836 (N_5836,N_5720,N_5787);
nand U5837 (N_5837,N_5744,N_5715);
nor U5838 (N_5838,N_5774,N_5730);
nor U5839 (N_5839,N_5743,N_5700);
and U5840 (N_5840,N_5749,N_5778);
nor U5841 (N_5841,N_5779,N_5753);
nor U5842 (N_5842,N_5722,N_5760);
or U5843 (N_5843,N_5794,N_5748);
or U5844 (N_5844,N_5710,N_5763);
or U5845 (N_5845,N_5793,N_5724);
or U5846 (N_5846,N_5742,N_5739);
nor U5847 (N_5847,N_5702,N_5790);
or U5848 (N_5848,N_5788,N_5714);
nor U5849 (N_5849,N_5741,N_5764);
nor U5850 (N_5850,N_5780,N_5717);
nor U5851 (N_5851,N_5773,N_5732);
nand U5852 (N_5852,N_5740,N_5707);
nand U5853 (N_5853,N_5759,N_5703);
or U5854 (N_5854,N_5767,N_5740);
nor U5855 (N_5855,N_5725,N_5782);
nand U5856 (N_5856,N_5704,N_5796);
or U5857 (N_5857,N_5792,N_5723);
or U5858 (N_5858,N_5794,N_5761);
or U5859 (N_5859,N_5727,N_5758);
nand U5860 (N_5860,N_5733,N_5762);
xor U5861 (N_5861,N_5725,N_5747);
and U5862 (N_5862,N_5770,N_5747);
and U5863 (N_5863,N_5742,N_5717);
xor U5864 (N_5864,N_5703,N_5789);
nor U5865 (N_5865,N_5748,N_5769);
or U5866 (N_5866,N_5775,N_5760);
nor U5867 (N_5867,N_5737,N_5794);
nand U5868 (N_5868,N_5777,N_5733);
nand U5869 (N_5869,N_5716,N_5723);
and U5870 (N_5870,N_5730,N_5711);
and U5871 (N_5871,N_5755,N_5773);
or U5872 (N_5872,N_5769,N_5703);
nor U5873 (N_5873,N_5711,N_5797);
nand U5874 (N_5874,N_5718,N_5794);
and U5875 (N_5875,N_5743,N_5765);
or U5876 (N_5876,N_5733,N_5716);
and U5877 (N_5877,N_5702,N_5737);
or U5878 (N_5878,N_5784,N_5776);
or U5879 (N_5879,N_5779,N_5744);
and U5880 (N_5880,N_5721,N_5775);
and U5881 (N_5881,N_5703,N_5774);
and U5882 (N_5882,N_5758,N_5797);
xor U5883 (N_5883,N_5751,N_5710);
nor U5884 (N_5884,N_5728,N_5731);
or U5885 (N_5885,N_5721,N_5708);
nor U5886 (N_5886,N_5779,N_5708);
nor U5887 (N_5887,N_5769,N_5770);
nand U5888 (N_5888,N_5720,N_5736);
nor U5889 (N_5889,N_5781,N_5745);
and U5890 (N_5890,N_5749,N_5727);
or U5891 (N_5891,N_5721,N_5764);
or U5892 (N_5892,N_5735,N_5795);
nor U5893 (N_5893,N_5742,N_5732);
nand U5894 (N_5894,N_5774,N_5731);
and U5895 (N_5895,N_5731,N_5717);
xnor U5896 (N_5896,N_5729,N_5730);
xor U5897 (N_5897,N_5791,N_5705);
nor U5898 (N_5898,N_5738,N_5754);
and U5899 (N_5899,N_5775,N_5788);
nor U5900 (N_5900,N_5867,N_5852);
nand U5901 (N_5901,N_5864,N_5866);
nand U5902 (N_5902,N_5856,N_5812);
or U5903 (N_5903,N_5826,N_5815);
or U5904 (N_5904,N_5829,N_5898);
and U5905 (N_5905,N_5806,N_5828);
and U5906 (N_5906,N_5827,N_5801);
and U5907 (N_5907,N_5842,N_5868);
xnor U5908 (N_5908,N_5835,N_5854);
or U5909 (N_5909,N_5840,N_5846);
nand U5910 (N_5910,N_5831,N_5837);
or U5911 (N_5911,N_5816,N_5838);
nor U5912 (N_5912,N_5873,N_5821);
nand U5913 (N_5913,N_5802,N_5853);
nor U5914 (N_5914,N_5884,N_5890);
nand U5915 (N_5915,N_5876,N_5810);
nand U5916 (N_5916,N_5817,N_5885);
or U5917 (N_5917,N_5841,N_5825);
or U5918 (N_5918,N_5836,N_5886);
nor U5919 (N_5919,N_5819,N_5845);
nand U5920 (N_5920,N_5814,N_5896);
or U5921 (N_5921,N_5824,N_5857);
xnor U5922 (N_5922,N_5800,N_5809);
and U5923 (N_5923,N_5820,N_5839);
nor U5924 (N_5924,N_5892,N_5878);
or U5925 (N_5925,N_5805,N_5875);
nand U5926 (N_5926,N_5843,N_5871);
and U5927 (N_5927,N_5813,N_5818);
nor U5928 (N_5928,N_5858,N_5877);
and U5929 (N_5929,N_5833,N_5822);
or U5930 (N_5930,N_5899,N_5808);
xor U5931 (N_5931,N_5834,N_5882);
nand U5932 (N_5932,N_5863,N_5851);
nor U5933 (N_5933,N_5850,N_5870);
nor U5934 (N_5934,N_5811,N_5807);
xor U5935 (N_5935,N_5861,N_5803);
nor U5936 (N_5936,N_5847,N_5844);
nor U5937 (N_5937,N_5855,N_5859);
nor U5938 (N_5938,N_5881,N_5860);
xor U5939 (N_5939,N_5848,N_5889);
and U5940 (N_5940,N_5849,N_5830);
nor U5941 (N_5941,N_5879,N_5897);
nor U5942 (N_5942,N_5832,N_5893);
and U5943 (N_5943,N_5888,N_5874);
xnor U5944 (N_5944,N_5872,N_5823);
nand U5945 (N_5945,N_5865,N_5869);
or U5946 (N_5946,N_5895,N_5862);
and U5947 (N_5947,N_5880,N_5804);
nor U5948 (N_5948,N_5894,N_5883);
nor U5949 (N_5949,N_5891,N_5887);
and U5950 (N_5950,N_5876,N_5832);
nor U5951 (N_5951,N_5820,N_5856);
or U5952 (N_5952,N_5811,N_5878);
and U5953 (N_5953,N_5884,N_5857);
or U5954 (N_5954,N_5881,N_5898);
xor U5955 (N_5955,N_5827,N_5880);
nor U5956 (N_5956,N_5890,N_5819);
and U5957 (N_5957,N_5864,N_5873);
and U5958 (N_5958,N_5865,N_5817);
or U5959 (N_5959,N_5818,N_5825);
xnor U5960 (N_5960,N_5807,N_5820);
or U5961 (N_5961,N_5898,N_5857);
or U5962 (N_5962,N_5890,N_5880);
and U5963 (N_5963,N_5853,N_5805);
or U5964 (N_5964,N_5838,N_5840);
and U5965 (N_5965,N_5838,N_5817);
or U5966 (N_5966,N_5812,N_5859);
nor U5967 (N_5967,N_5878,N_5853);
xnor U5968 (N_5968,N_5846,N_5802);
or U5969 (N_5969,N_5823,N_5875);
and U5970 (N_5970,N_5859,N_5814);
nand U5971 (N_5971,N_5854,N_5849);
nor U5972 (N_5972,N_5845,N_5898);
and U5973 (N_5973,N_5863,N_5891);
and U5974 (N_5974,N_5873,N_5882);
nand U5975 (N_5975,N_5804,N_5887);
nand U5976 (N_5976,N_5826,N_5894);
nor U5977 (N_5977,N_5811,N_5819);
and U5978 (N_5978,N_5859,N_5821);
nor U5979 (N_5979,N_5817,N_5812);
nor U5980 (N_5980,N_5848,N_5865);
and U5981 (N_5981,N_5828,N_5871);
nand U5982 (N_5982,N_5831,N_5867);
and U5983 (N_5983,N_5874,N_5841);
nand U5984 (N_5984,N_5860,N_5816);
and U5985 (N_5985,N_5832,N_5873);
xor U5986 (N_5986,N_5894,N_5899);
nor U5987 (N_5987,N_5824,N_5826);
nand U5988 (N_5988,N_5859,N_5833);
or U5989 (N_5989,N_5818,N_5833);
or U5990 (N_5990,N_5832,N_5851);
nand U5991 (N_5991,N_5806,N_5841);
nand U5992 (N_5992,N_5845,N_5811);
nand U5993 (N_5993,N_5863,N_5830);
nand U5994 (N_5994,N_5818,N_5856);
xor U5995 (N_5995,N_5811,N_5825);
nor U5996 (N_5996,N_5800,N_5816);
or U5997 (N_5997,N_5819,N_5817);
xnor U5998 (N_5998,N_5863,N_5899);
or U5999 (N_5999,N_5847,N_5870);
nor U6000 (N_6000,N_5957,N_5976);
nand U6001 (N_6001,N_5982,N_5986);
nor U6002 (N_6002,N_5981,N_5968);
nor U6003 (N_6003,N_5989,N_5939);
or U6004 (N_6004,N_5916,N_5945);
and U6005 (N_6005,N_5987,N_5993);
xnor U6006 (N_6006,N_5983,N_5912);
and U6007 (N_6007,N_5900,N_5932);
nor U6008 (N_6008,N_5995,N_5938);
nand U6009 (N_6009,N_5965,N_5906);
and U6010 (N_6010,N_5964,N_5919);
or U6011 (N_6011,N_5955,N_5941);
nor U6012 (N_6012,N_5940,N_5901);
nor U6013 (N_6013,N_5979,N_5970);
nand U6014 (N_6014,N_5948,N_5931);
nor U6015 (N_6015,N_5997,N_5963);
xnor U6016 (N_6016,N_5933,N_5913);
nor U6017 (N_6017,N_5918,N_5996);
or U6018 (N_6018,N_5973,N_5937);
or U6019 (N_6019,N_5991,N_5917);
nand U6020 (N_6020,N_5951,N_5960);
nor U6021 (N_6021,N_5962,N_5923);
nand U6022 (N_6022,N_5966,N_5946);
nor U6023 (N_6023,N_5953,N_5947);
xor U6024 (N_6024,N_5952,N_5922);
nand U6025 (N_6025,N_5984,N_5935);
and U6026 (N_6026,N_5929,N_5999);
and U6027 (N_6027,N_5908,N_5914);
nand U6028 (N_6028,N_5975,N_5927);
nand U6029 (N_6029,N_5992,N_5902);
and U6030 (N_6030,N_5903,N_5958);
and U6031 (N_6031,N_5926,N_5949);
and U6032 (N_6032,N_5980,N_5977);
nor U6033 (N_6033,N_5990,N_5978);
nor U6034 (N_6034,N_5959,N_5905);
and U6035 (N_6035,N_5928,N_5936);
nor U6036 (N_6036,N_5934,N_5954);
or U6037 (N_6037,N_5972,N_5943);
nor U6038 (N_6038,N_5998,N_5969);
or U6039 (N_6039,N_5921,N_5924);
nand U6040 (N_6040,N_5911,N_5915);
and U6041 (N_6041,N_5910,N_5967);
or U6042 (N_6042,N_5971,N_5909);
nor U6043 (N_6043,N_5904,N_5944);
nand U6044 (N_6044,N_5994,N_5907);
nand U6045 (N_6045,N_5930,N_5920);
or U6046 (N_6046,N_5988,N_5961);
and U6047 (N_6047,N_5985,N_5942);
or U6048 (N_6048,N_5974,N_5950);
xnor U6049 (N_6049,N_5925,N_5956);
and U6050 (N_6050,N_5905,N_5933);
or U6051 (N_6051,N_5919,N_5947);
nand U6052 (N_6052,N_5950,N_5923);
and U6053 (N_6053,N_5968,N_5916);
xor U6054 (N_6054,N_5921,N_5945);
nor U6055 (N_6055,N_5952,N_5984);
nor U6056 (N_6056,N_5920,N_5938);
nor U6057 (N_6057,N_5900,N_5930);
xor U6058 (N_6058,N_5972,N_5971);
nand U6059 (N_6059,N_5901,N_5904);
nand U6060 (N_6060,N_5937,N_5971);
and U6061 (N_6061,N_5903,N_5999);
or U6062 (N_6062,N_5989,N_5931);
nor U6063 (N_6063,N_5912,N_5966);
or U6064 (N_6064,N_5917,N_5942);
nand U6065 (N_6065,N_5908,N_5962);
and U6066 (N_6066,N_5954,N_5936);
nand U6067 (N_6067,N_5987,N_5924);
nand U6068 (N_6068,N_5910,N_5906);
nand U6069 (N_6069,N_5991,N_5911);
nor U6070 (N_6070,N_5970,N_5948);
nor U6071 (N_6071,N_5961,N_5991);
nor U6072 (N_6072,N_5948,N_5997);
and U6073 (N_6073,N_5930,N_5963);
nor U6074 (N_6074,N_5966,N_5928);
or U6075 (N_6075,N_5937,N_5940);
and U6076 (N_6076,N_5949,N_5988);
and U6077 (N_6077,N_5970,N_5977);
nand U6078 (N_6078,N_5979,N_5920);
xnor U6079 (N_6079,N_5907,N_5920);
nor U6080 (N_6080,N_5927,N_5981);
nor U6081 (N_6081,N_5961,N_5928);
nor U6082 (N_6082,N_5903,N_5978);
xor U6083 (N_6083,N_5985,N_5911);
and U6084 (N_6084,N_5974,N_5990);
or U6085 (N_6085,N_5937,N_5946);
or U6086 (N_6086,N_5972,N_5925);
and U6087 (N_6087,N_5997,N_5919);
and U6088 (N_6088,N_5946,N_5989);
nor U6089 (N_6089,N_5952,N_5943);
and U6090 (N_6090,N_5968,N_5970);
nand U6091 (N_6091,N_5905,N_5939);
nor U6092 (N_6092,N_5921,N_5958);
or U6093 (N_6093,N_5974,N_5972);
or U6094 (N_6094,N_5952,N_5977);
nand U6095 (N_6095,N_5956,N_5978);
or U6096 (N_6096,N_5952,N_5906);
or U6097 (N_6097,N_5956,N_5941);
xnor U6098 (N_6098,N_5952,N_5900);
nand U6099 (N_6099,N_5965,N_5938);
nor U6100 (N_6100,N_6059,N_6017);
nand U6101 (N_6101,N_6051,N_6069);
nor U6102 (N_6102,N_6022,N_6054);
or U6103 (N_6103,N_6033,N_6046);
and U6104 (N_6104,N_6048,N_6079);
nand U6105 (N_6105,N_6010,N_6074);
or U6106 (N_6106,N_6073,N_6009);
and U6107 (N_6107,N_6001,N_6091);
nand U6108 (N_6108,N_6025,N_6068);
nand U6109 (N_6109,N_6098,N_6023);
or U6110 (N_6110,N_6028,N_6049);
xnor U6111 (N_6111,N_6099,N_6097);
nor U6112 (N_6112,N_6072,N_6070);
nand U6113 (N_6113,N_6057,N_6052);
nand U6114 (N_6114,N_6032,N_6031);
xnor U6115 (N_6115,N_6064,N_6002);
or U6116 (N_6116,N_6078,N_6086);
or U6117 (N_6117,N_6084,N_6034);
and U6118 (N_6118,N_6085,N_6088);
or U6119 (N_6119,N_6062,N_6044);
nor U6120 (N_6120,N_6080,N_6030);
and U6121 (N_6121,N_6015,N_6063);
and U6122 (N_6122,N_6089,N_6055);
nor U6123 (N_6123,N_6019,N_6047);
nor U6124 (N_6124,N_6008,N_6020);
nand U6125 (N_6125,N_6007,N_6065);
or U6126 (N_6126,N_6000,N_6005);
and U6127 (N_6127,N_6036,N_6081);
and U6128 (N_6128,N_6092,N_6026);
or U6129 (N_6129,N_6024,N_6058);
or U6130 (N_6130,N_6061,N_6087);
xor U6131 (N_6131,N_6014,N_6040);
or U6132 (N_6132,N_6029,N_6021);
xor U6133 (N_6133,N_6039,N_6011);
or U6134 (N_6134,N_6012,N_6096);
nor U6135 (N_6135,N_6037,N_6027);
nor U6136 (N_6136,N_6042,N_6041);
or U6137 (N_6137,N_6006,N_6060);
nor U6138 (N_6138,N_6056,N_6083);
or U6139 (N_6139,N_6035,N_6053);
or U6140 (N_6140,N_6090,N_6075);
and U6141 (N_6141,N_6066,N_6004);
or U6142 (N_6142,N_6071,N_6013);
nor U6143 (N_6143,N_6082,N_6018);
nor U6144 (N_6144,N_6067,N_6038);
nor U6145 (N_6145,N_6043,N_6003);
nand U6146 (N_6146,N_6094,N_6076);
and U6147 (N_6147,N_6093,N_6016);
and U6148 (N_6148,N_6077,N_6095);
nand U6149 (N_6149,N_6045,N_6050);
or U6150 (N_6150,N_6064,N_6004);
and U6151 (N_6151,N_6029,N_6037);
or U6152 (N_6152,N_6005,N_6026);
or U6153 (N_6153,N_6071,N_6086);
xnor U6154 (N_6154,N_6048,N_6032);
or U6155 (N_6155,N_6086,N_6064);
or U6156 (N_6156,N_6071,N_6031);
nand U6157 (N_6157,N_6075,N_6048);
and U6158 (N_6158,N_6091,N_6038);
nand U6159 (N_6159,N_6099,N_6033);
nand U6160 (N_6160,N_6072,N_6004);
nand U6161 (N_6161,N_6030,N_6061);
nor U6162 (N_6162,N_6054,N_6052);
nand U6163 (N_6163,N_6012,N_6003);
and U6164 (N_6164,N_6008,N_6003);
and U6165 (N_6165,N_6027,N_6026);
or U6166 (N_6166,N_6051,N_6016);
nand U6167 (N_6167,N_6050,N_6081);
nand U6168 (N_6168,N_6086,N_6044);
nor U6169 (N_6169,N_6003,N_6021);
nor U6170 (N_6170,N_6042,N_6026);
and U6171 (N_6171,N_6048,N_6045);
nor U6172 (N_6172,N_6035,N_6003);
nor U6173 (N_6173,N_6062,N_6061);
and U6174 (N_6174,N_6021,N_6069);
or U6175 (N_6175,N_6060,N_6015);
nor U6176 (N_6176,N_6089,N_6007);
and U6177 (N_6177,N_6072,N_6011);
xor U6178 (N_6178,N_6010,N_6024);
or U6179 (N_6179,N_6084,N_6040);
nand U6180 (N_6180,N_6087,N_6076);
and U6181 (N_6181,N_6087,N_6011);
or U6182 (N_6182,N_6098,N_6060);
xor U6183 (N_6183,N_6046,N_6098);
or U6184 (N_6184,N_6006,N_6019);
nor U6185 (N_6185,N_6013,N_6041);
nand U6186 (N_6186,N_6082,N_6088);
or U6187 (N_6187,N_6044,N_6048);
nor U6188 (N_6188,N_6043,N_6008);
and U6189 (N_6189,N_6049,N_6081);
nand U6190 (N_6190,N_6042,N_6000);
nand U6191 (N_6191,N_6041,N_6012);
xnor U6192 (N_6192,N_6014,N_6058);
or U6193 (N_6193,N_6020,N_6026);
or U6194 (N_6194,N_6068,N_6061);
nand U6195 (N_6195,N_6008,N_6032);
and U6196 (N_6196,N_6038,N_6042);
nand U6197 (N_6197,N_6094,N_6011);
and U6198 (N_6198,N_6008,N_6030);
nor U6199 (N_6199,N_6074,N_6030);
and U6200 (N_6200,N_6127,N_6152);
nor U6201 (N_6201,N_6183,N_6191);
and U6202 (N_6202,N_6125,N_6189);
nor U6203 (N_6203,N_6151,N_6161);
nor U6204 (N_6204,N_6199,N_6148);
or U6205 (N_6205,N_6132,N_6134);
nand U6206 (N_6206,N_6115,N_6186);
and U6207 (N_6207,N_6128,N_6171);
or U6208 (N_6208,N_6109,N_6122);
nand U6209 (N_6209,N_6182,N_6164);
or U6210 (N_6210,N_6178,N_6184);
nor U6211 (N_6211,N_6153,N_6147);
or U6212 (N_6212,N_6102,N_6124);
nor U6213 (N_6213,N_6103,N_6110);
and U6214 (N_6214,N_6106,N_6158);
nand U6215 (N_6215,N_6104,N_6140);
and U6216 (N_6216,N_6118,N_6119);
and U6217 (N_6217,N_6120,N_6170);
nor U6218 (N_6218,N_6105,N_6130);
nor U6219 (N_6219,N_6146,N_6181);
nand U6220 (N_6220,N_6107,N_6155);
or U6221 (N_6221,N_6169,N_6177);
nor U6222 (N_6222,N_6172,N_6117);
nor U6223 (N_6223,N_6111,N_6136);
or U6224 (N_6224,N_6145,N_6143);
nor U6225 (N_6225,N_6173,N_6187);
or U6226 (N_6226,N_6133,N_6129);
or U6227 (N_6227,N_6149,N_6162);
and U6228 (N_6228,N_6139,N_6160);
and U6229 (N_6229,N_6141,N_6188);
nand U6230 (N_6230,N_6135,N_6131);
nand U6231 (N_6231,N_6165,N_6166);
and U6232 (N_6232,N_6138,N_6112);
or U6233 (N_6233,N_6156,N_6100);
nor U6234 (N_6234,N_6116,N_6150);
or U6235 (N_6235,N_6179,N_6195);
nand U6236 (N_6236,N_6193,N_6198);
xor U6237 (N_6237,N_6101,N_6137);
nand U6238 (N_6238,N_6180,N_6194);
nand U6239 (N_6239,N_6114,N_6175);
nand U6240 (N_6240,N_6123,N_6192);
nor U6241 (N_6241,N_6185,N_6197);
or U6242 (N_6242,N_6126,N_6196);
nor U6243 (N_6243,N_6167,N_6113);
nor U6244 (N_6244,N_6154,N_6142);
or U6245 (N_6245,N_6176,N_6163);
xor U6246 (N_6246,N_6121,N_6190);
or U6247 (N_6247,N_6159,N_6108);
nand U6248 (N_6248,N_6144,N_6174);
or U6249 (N_6249,N_6168,N_6157);
nor U6250 (N_6250,N_6153,N_6191);
or U6251 (N_6251,N_6184,N_6187);
nand U6252 (N_6252,N_6114,N_6113);
xnor U6253 (N_6253,N_6192,N_6169);
xnor U6254 (N_6254,N_6196,N_6194);
or U6255 (N_6255,N_6181,N_6179);
nor U6256 (N_6256,N_6144,N_6167);
or U6257 (N_6257,N_6113,N_6128);
and U6258 (N_6258,N_6178,N_6126);
nor U6259 (N_6259,N_6105,N_6157);
and U6260 (N_6260,N_6144,N_6161);
and U6261 (N_6261,N_6135,N_6116);
and U6262 (N_6262,N_6136,N_6117);
or U6263 (N_6263,N_6111,N_6180);
or U6264 (N_6264,N_6165,N_6136);
or U6265 (N_6265,N_6103,N_6191);
nor U6266 (N_6266,N_6103,N_6137);
xnor U6267 (N_6267,N_6144,N_6135);
or U6268 (N_6268,N_6177,N_6183);
and U6269 (N_6269,N_6154,N_6158);
nor U6270 (N_6270,N_6148,N_6194);
and U6271 (N_6271,N_6164,N_6168);
nor U6272 (N_6272,N_6169,N_6128);
nand U6273 (N_6273,N_6130,N_6137);
and U6274 (N_6274,N_6135,N_6132);
or U6275 (N_6275,N_6141,N_6103);
or U6276 (N_6276,N_6139,N_6187);
nor U6277 (N_6277,N_6144,N_6148);
or U6278 (N_6278,N_6116,N_6111);
nor U6279 (N_6279,N_6109,N_6137);
or U6280 (N_6280,N_6141,N_6113);
nor U6281 (N_6281,N_6150,N_6196);
and U6282 (N_6282,N_6139,N_6175);
nor U6283 (N_6283,N_6108,N_6152);
xor U6284 (N_6284,N_6107,N_6128);
and U6285 (N_6285,N_6104,N_6125);
or U6286 (N_6286,N_6198,N_6106);
and U6287 (N_6287,N_6153,N_6137);
or U6288 (N_6288,N_6108,N_6151);
nand U6289 (N_6289,N_6143,N_6188);
nor U6290 (N_6290,N_6152,N_6198);
nand U6291 (N_6291,N_6166,N_6171);
and U6292 (N_6292,N_6184,N_6117);
nand U6293 (N_6293,N_6135,N_6185);
nor U6294 (N_6294,N_6189,N_6167);
and U6295 (N_6295,N_6159,N_6191);
and U6296 (N_6296,N_6110,N_6144);
and U6297 (N_6297,N_6134,N_6106);
or U6298 (N_6298,N_6164,N_6154);
or U6299 (N_6299,N_6113,N_6125);
and U6300 (N_6300,N_6266,N_6279);
and U6301 (N_6301,N_6296,N_6268);
nor U6302 (N_6302,N_6258,N_6293);
nand U6303 (N_6303,N_6255,N_6283);
and U6304 (N_6304,N_6252,N_6270);
xor U6305 (N_6305,N_6206,N_6230);
and U6306 (N_6306,N_6251,N_6201);
or U6307 (N_6307,N_6257,N_6234);
or U6308 (N_6308,N_6242,N_6210);
or U6309 (N_6309,N_6219,N_6236);
and U6310 (N_6310,N_6204,N_6282);
nor U6311 (N_6311,N_6290,N_6278);
nand U6312 (N_6312,N_6287,N_6213);
nand U6313 (N_6313,N_6256,N_6291);
nor U6314 (N_6314,N_6272,N_6254);
or U6315 (N_6315,N_6221,N_6262);
and U6316 (N_6316,N_6241,N_6228);
and U6317 (N_6317,N_6260,N_6240);
nand U6318 (N_6318,N_6203,N_6248);
xnor U6319 (N_6319,N_6284,N_6249);
and U6320 (N_6320,N_6267,N_6238);
nand U6321 (N_6321,N_6229,N_6285);
and U6322 (N_6322,N_6274,N_6223);
nand U6323 (N_6323,N_6200,N_6298);
nor U6324 (N_6324,N_6276,N_6295);
xnor U6325 (N_6325,N_6232,N_6247);
or U6326 (N_6326,N_6235,N_6231);
nand U6327 (N_6327,N_6273,N_6222);
nor U6328 (N_6328,N_6205,N_6277);
nor U6329 (N_6329,N_6288,N_6246);
xor U6330 (N_6330,N_6211,N_6226);
nand U6331 (N_6331,N_6239,N_6265);
or U6332 (N_6332,N_6297,N_6216);
nor U6333 (N_6333,N_6218,N_6259);
nor U6334 (N_6334,N_6237,N_6286);
xor U6335 (N_6335,N_6227,N_6250);
nor U6336 (N_6336,N_6208,N_6224);
and U6337 (N_6337,N_6253,N_6220);
nor U6338 (N_6338,N_6292,N_6263);
nor U6339 (N_6339,N_6212,N_6217);
nand U6340 (N_6340,N_6271,N_6207);
or U6341 (N_6341,N_6275,N_6233);
and U6342 (N_6342,N_6245,N_6289);
and U6343 (N_6343,N_6261,N_6202);
nand U6344 (N_6344,N_6209,N_6280);
or U6345 (N_6345,N_6299,N_6281);
or U6346 (N_6346,N_6214,N_6243);
or U6347 (N_6347,N_6294,N_6225);
nor U6348 (N_6348,N_6264,N_6269);
nand U6349 (N_6349,N_6244,N_6215);
xnor U6350 (N_6350,N_6224,N_6258);
nor U6351 (N_6351,N_6250,N_6246);
nand U6352 (N_6352,N_6288,N_6278);
nand U6353 (N_6353,N_6261,N_6236);
and U6354 (N_6354,N_6230,N_6280);
nand U6355 (N_6355,N_6284,N_6292);
nor U6356 (N_6356,N_6271,N_6256);
nand U6357 (N_6357,N_6263,N_6201);
nor U6358 (N_6358,N_6251,N_6277);
nand U6359 (N_6359,N_6202,N_6276);
or U6360 (N_6360,N_6285,N_6296);
nand U6361 (N_6361,N_6253,N_6276);
xnor U6362 (N_6362,N_6250,N_6254);
xor U6363 (N_6363,N_6226,N_6201);
and U6364 (N_6364,N_6270,N_6207);
and U6365 (N_6365,N_6219,N_6234);
nand U6366 (N_6366,N_6247,N_6265);
xnor U6367 (N_6367,N_6246,N_6281);
and U6368 (N_6368,N_6229,N_6220);
nand U6369 (N_6369,N_6218,N_6261);
or U6370 (N_6370,N_6278,N_6254);
or U6371 (N_6371,N_6269,N_6275);
nand U6372 (N_6372,N_6281,N_6295);
nand U6373 (N_6373,N_6240,N_6255);
or U6374 (N_6374,N_6287,N_6246);
or U6375 (N_6375,N_6286,N_6287);
and U6376 (N_6376,N_6264,N_6232);
nand U6377 (N_6377,N_6231,N_6253);
nor U6378 (N_6378,N_6229,N_6200);
and U6379 (N_6379,N_6246,N_6225);
or U6380 (N_6380,N_6210,N_6205);
nor U6381 (N_6381,N_6281,N_6200);
xor U6382 (N_6382,N_6287,N_6275);
nor U6383 (N_6383,N_6253,N_6206);
or U6384 (N_6384,N_6263,N_6244);
or U6385 (N_6385,N_6288,N_6296);
nand U6386 (N_6386,N_6208,N_6256);
and U6387 (N_6387,N_6295,N_6280);
nand U6388 (N_6388,N_6283,N_6269);
nand U6389 (N_6389,N_6215,N_6270);
xor U6390 (N_6390,N_6240,N_6271);
nand U6391 (N_6391,N_6250,N_6259);
or U6392 (N_6392,N_6204,N_6229);
and U6393 (N_6393,N_6269,N_6285);
or U6394 (N_6394,N_6232,N_6298);
nand U6395 (N_6395,N_6216,N_6285);
and U6396 (N_6396,N_6224,N_6298);
nand U6397 (N_6397,N_6277,N_6209);
or U6398 (N_6398,N_6214,N_6298);
or U6399 (N_6399,N_6221,N_6287);
nand U6400 (N_6400,N_6300,N_6383);
nand U6401 (N_6401,N_6397,N_6373);
nor U6402 (N_6402,N_6362,N_6390);
or U6403 (N_6403,N_6379,N_6371);
and U6404 (N_6404,N_6385,N_6333);
nor U6405 (N_6405,N_6346,N_6381);
xnor U6406 (N_6406,N_6321,N_6378);
nor U6407 (N_6407,N_6301,N_6364);
nand U6408 (N_6408,N_6388,N_6304);
xnor U6409 (N_6409,N_6337,N_6359);
nor U6410 (N_6410,N_6322,N_6335);
and U6411 (N_6411,N_6357,N_6328);
and U6412 (N_6412,N_6355,N_6365);
nor U6413 (N_6413,N_6377,N_6303);
nand U6414 (N_6414,N_6341,N_6354);
nor U6415 (N_6415,N_6319,N_6352);
nand U6416 (N_6416,N_6324,N_6351);
or U6417 (N_6417,N_6396,N_6361);
and U6418 (N_6418,N_6336,N_6316);
or U6419 (N_6419,N_6311,N_6310);
nand U6420 (N_6420,N_6389,N_6393);
nor U6421 (N_6421,N_6363,N_6387);
nor U6422 (N_6422,N_6334,N_6339);
nor U6423 (N_6423,N_6369,N_6320);
or U6424 (N_6424,N_6326,N_6302);
or U6425 (N_6425,N_6384,N_6350);
or U6426 (N_6426,N_6349,N_6318);
nor U6427 (N_6427,N_6360,N_6313);
nor U6428 (N_6428,N_6317,N_6391);
xnor U6429 (N_6429,N_6330,N_6380);
or U6430 (N_6430,N_6375,N_6398);
xor U6431 (N_6431,N_6323,N_6372);
and U6432 (N_6432,N_6392,N_6367);
and U6433 (N_6433,N_6347,N_6395);
nand U6434 (N_6434,N_6307,N_6332);
nand U6435 (N_6435,N_6342,N_6306);
or U6436 (N_6436,N_6348,N_6329);
or U6437 (N_6437,N_6305,N_6312);
nor U6438 (N_6438,N_6353,N_6358);
nor U6439 (N_6439,N_6343,N_6370);
nand U6440 (N_6440,N_6309,N_6314);
nand U6441 (N_6441,N_6394,N_6368);
or U6442 (N_6442,N_6325,N_6356);
and U6443 (N_6443,N_6308,N_6376);
or U6444 (N_6444,N_6382,N_6374);
nand U6445 (N_6445,N_6344,N_6331);
and U6446 (N_6446,N_6315,N_6340);
nor U6447 (N_6447,N_6345,N_6338);
xnor U6448 (N_6448,N_6399,N_6327);
xor U6449 (N_6449,N_6386,N_6366);
nor U6450 (N_6450,N_6356,N_6333);
nor U6451 (N_6451,N_6319,N_6335);
and U6452 (N_6452,N_6375,N_6347);
nor U6453 (N_6453,N_6361,N_6308);
nand U6454 (N_6454,N_6377,N_6324);
or U6455 (N_6455,N_6387,N_6377);
and U6456 (N_6456,N_6306,N_6364);
nor U6457 (N_6457,N_6319,N_6385);
nand U6458 (N_6458,N_6354,N_6386);
nor U6459 (N_6459,N_6336,N_6391);
or U6460 (N_6460,N_6308,N_6340);
nor U6461 (N_6461,N_6352,N_6354);
or U6462 (N_6462,N_6384,N_6342);
or U6463 (N_6463,N_6384,N_6325);
and U6464 (N_6464,N_6306,N_6370);
xor U6465 (N_6465,N_6345,N_6392);
and U6466 (N_6466,N_6396,N_6381);
or U6467 (N_6467,N_6304,N_6357);
or U6468 (N_6468,N_6327,N_6315);
and U6469 (N_6469,N_6393,N_6373);
or U6470 (N_6470,N_6356,N_6399);
xnor U6471 (N_6471,N_6311,N_6355);
or U6472 (N_6472,N_6312,N_6306);
and U6473 (N_6473,N_6311,N_6398);
nand U6474 (N_6474,N_6374,N_6314);
nor U6475 (N_6475,N_6321,N_6314);
nor U6476 (N_6476,N_6308,N_6302);
and U6477 (N_6477,N_6365,N_6318);
nand U6478 (N_6478,N_6327,N_6312);
xnor U6479 (N_6479,N_6324,N_6350);
and U6480 (N_6480,N_6355,N_6379);
and U6481 (N_6481,N_6382,N_6366);
nand U6482 (N_6482,N_6308,N_6305);
nand U6483 (N_6483,N_6391,N_6322);
or U6484 (N_6484,N_6330,N_6321);
or U6485 (N_6485,N_6338,N_6381);
nand U6486 (N_6486,N_6306,N_6368);
nand U6487 (N_6487,N_6307,N_6397);
or U6488 (N_6488,N_6348,N_6300);
and U6489 (N_6489,N_6380,N_6399);
or U6490 (N_6490,N_6345,N_6352);
nand U6491 (N_6491,N_6365,N_6357);
and U6492 (N_6492,N_6399,N_6359);
nor U6493 (N_6493,N_6324,N_6304);
and U6494 (N_6494,N_6356,N_6352);
or U6495 (N_6495,N_6394,N_6367);
xnor U6496 (N_6496,N_6355,N_6326);
nor U6497 (N_6497,N_6340,N_6300);
and U6498 (N_6498,N_6380,N_6390);
nand U6499 (N_6499,N_6397,N_6308);
and U6500 (N_6500,N_6403,N_6444);
nor U6501 (N_6501,N_6446,N_6440);
xor U6502 (N_6502,N_6469,N_6459);
or U6503 (N_6503,N_6414,N_6473);
nor U6504 (N_6504,N_6479,N_6453);
or U6505 (N_6505,N_6443,N_6461);
and U6506 (N_6506,N_6435,N_6498);
and U6507 (N_6507,N_6412,N_6402);
and U6508 (N_6508,N_6491,N_6475);
nand U6509 (N_6509,N_6465,N_6437);
nor U6510 (N_6510,N_6497,N_6474);
nand U6511 (N_6511,N_6417,N_6404);
and U6512 (N_6512,N_6481,N_6434);
nor U6513 (N_6513,N_6472,N_6438);
nand U6514 (N_6514,N_6462,N_6406);
xnor U6515 (N_6515,N_6470,N_6439);
and U6516 (N_6516,N_6496,N_6415);
and U6517 (N_6517,N_6456,N_6489);
or U6518 (N_6518,N_6447,N_6418);
and U6519 (N_6519,N_6448,N_6467);
and U6520 (N_6520,N_6408,N_6445);
and U6521 (N_6521,N_6484,N_6454);
nand U6522 (N_6522,N_6430,N_6458);
nor U6523 (N_6523,N_6490,N_6488);
xnor U6524 (N_6524,N_6492,N_6441);
nand U6525 (N_6525,N_6486,N_6450);
xor U6526 (N_6526,N_6429,N_6468);
nand U6527 (N_6527,N_6485,N_6433);
nor U6528 (N_6528,N_6466,N_6455);
nand U6529 (N_6529,N_6436,N_6422);
and U6530 (N_6530,N_6457,N_6400);
nor U6531 (N_6531,N_6428,N_6477);
or U6532 (N_6532,N_6449,N_6423);
nor U6533 (N_6533,N_6478,N_6420);
nand U6534 (N_6534,N_6407,N_6494);
nand U6535 (N_6535,N_6476,N_6409);
or U6536 (N_6536,N_6480,N_6421);
nor U6537 (N_6537,N_6426,N_6401);
nand U6538 (N_6538,N_6411,N_6493);
nand U6539 (N_6539,N_6451,N_6427);
and U6540 (N_6540,N_6410,N_6482);
nor U6541 (N_6541,N_6463,N_6432);
nor U6542 (N_6542,N_6431,N_6483);
and U6543 (N_6543,N_6460,N_6413);
nand U6544 (N_6544,N_6487,N_6495);
xnor U6545 (N_6545,N_6464,N_6419);
and U6546 (N_6546,N_6416,N_6452);
xnor U6547 (N_6547,N_6405,N_6425);
xnor U6548 (N_6548,N_6424,N_6471);
or U6549 (N_6549,N_6499,N_6442);
and U6550 (N_6550,N_6414,N_6492);
or U6551 (N_6551,N_6482,N_6461);
and U6552 (N_6552,N_6472,N_6430);
nand U6553 (N_6553,N_6437,N_6486);
nor U6554 (N_6554,N_6484,N_6417);
or U6555 (N_6555,N_6407,N_6466);
nor U6556 (N_6556,N_6466,N_6467);
nor U6557 (N_6557,N_6497,N_6411);
and U6558 (N_6558,N_6400,N_6480);
nor U6559 (N_6559,N_6481,N_6468);
nor U6560 (N_6560,N_6449,N_6415);
or U6561 (N_6561,N_6466,N_6432);
nand U6562 (N_6562,N_6413,N_6496);
nor U6563 (N_6563,N_6401,N_6416);
xnor U6564 (N_6564,N_6465,N_6496);
nor U6565 (N_6565,N_6416,N_6474);
nor U6566 (N_6566,N_6478,N_6455);
and U6567 (N_6567,N_6428,N_6437);
xnor U6568 (N_6568,N_6432,N_6440);
nand U6569 (N_6569,N_6431,N_6459);
nor U6570 (N_6570,N_6420,N_6445);
or U6571 (N_6571,N_6449,N_6425);
and U6572 (N_6572,N_6438,N_6427);
nor U6573 (N_6573,N_6422,N_6476);
or U6574 (N_6574,N_6438,N_6457);
and U6575 (N_6575,N_6440,N_6404);
or U6576 (N_6576,N_6491,N_6458);
xnor U6577 (N_6577,N_6403,N_6481);
nor U6578 (N_6578,N_6489,N_6486);
and U6579 (N_6579,N_6497,N_6459);
and U6580 (N_6580,N_6406,N_6475);
nand U6581 (N_6581,N_6426,N_6403);
nor U6582 (N_6582,N_6408,N_6440);
xnor U6583 (N_6583,N_6452,N_6486);
xor U6584 (N_6584,N_6434,N_6442);
nand U6585 (N_6585,N_6473,N_6485);
nand U6586 (N_6586,N_6422,N_6411);
or U6587 (N_6587,N_6426,N_6425);
nand U6588 (N_6588,N_6407,N_6461);
nor U6589 (N_6589,N_6408,N_6473);
nand U6590 (N_6590,N_6492,N_6469);
xnor U6591 (N_6591,N_6490,N_6473);
nand U6592 (N_6592,N_6440,N_6492);
nand U6593 (N_6593,N_6407,N_6450);
nor U6594 (N_6594,N_6416,N_6431);
or U6595 (N_6595,N_6443,N_6493);
nor U6596 (N_6596,N_6466,N_6454);
nand U6597 (N_6597,N_6402,N_6499);
nor U6598 (N_6598,N_6494,N_6405);
or U6599 (N_6599,N_6488,N_6468);
or U6600 (N_6600,N_6576,N_6563);
xor U6601 (N_6601,N_6530,N_6586);
nor U6602 (N_6602,N_6516,N_6592);
nand U6603 (N_6603,N_6578,N_6511);
and U6604 (N_6604,N_6559,N_6540);
nor U6605 (N_6605,N_6509,N_6557);
and U6606 (N_6606,N_6566,N_6580);
and U6607 (N_6607,N_6597,N_6517);
nor U6608 (N_6608,N_6572,N_6505);
or U6609 (N_6609,N_6541,N_6550);
nand U6610 (N_6610,N_6545,N_6599);
nand U6611 (N_6611,N_6538,N_6573);
nor U6612 (N_6612,N_6508,N_6569);
and U6613 (N_6613,N_6513,N_6504);
nand U6614 (N_6614,N_6594,N_6591);
or U6615 (N_6615,N_6565,N_6531);
nand U6616 (N_6616,N_6548,N_6528);
and U6617 (N_6617,N_6524,N_6575);
nor U6618 (N_6618,N_6544,N_6577);
nand U6619 (N_6619,N_6525,N_6543);
and U6620 (N_6620,N_6518,N_6590);
and U6621 (N_6621,N_6561,N_6585);
xor U6622 (N_6622,N_6598,N_6546);
or U6623 (N_6623,N_6501,N_6571);
nor U6624 (N_6624,N_6515,N_6579);
or U6625 (N_6625,N_6536,N_6535);
nand U6626 (N_6626,N_6558,N_6584);
nor U6627 (N_6627,N_6502,N_6587);
nor U6628 (N_6628,N_6593,N_6564);
or U6629 (N_6629,N_6512,N_6568);
nor U6630 (N_6630,N_6519,N_6551);
nand U6631 (N_6631,N_6562,N_6555);
or U6632 (N_6632,N_6500,N_6581);
nand U6633 (N_6633,N_6503,N_6549);
nand U6634 (N_6634,N_6547,N_6556);
nand U6635 (N_6635,N_6510,N_6527);
nand U6636 (N_6636,N_6537,N_6570);
nor U6637 (N_6637,N_6532,N_6588);
nor U6638 (N_6638,N_6534,N_6583);
and U6639 (N_6639,N_6553,N_6507);
or U6640 (N_6640,N_6560,N_6552);
or U6641 (N_6641,N_6539,N_6523);
or U6642 (N_6642,N_6514,N_6521);
and U6643 (N_6643,N_6520,N_6554);
nand U6644 (N_6644,N_6595,N_6582);
and U6645 (N_6645,N_6567,N_6506);
and U6646 (N_6646,N_6542,N_6533);
nor U6647 (N_6647,N_6574,N_6526);
and U6648 (N_6648,N_6589,N_6596);
or U6649 (N_6649,N_6522,N_6529);
and U6650 (N_6650,N_6513,N_6581);
and U6651 (N_6651,N_6502,N_6572);
nor U6652 (N_6652,N_6592,N_6514);
nor U6653 (N_6653,N_6574,N_6553);
nand U6654 (N_6654,N_6590,N_6515);
and U6655 (N_6655,N_6585,N_6587);
xor U6656 (N_6656,N_6511,N_6565);
xnor U6657 (N_6657,N_6576,N_6524);
nor U6658 (N_6658,N_6597,N_6512);
and U6659 (N_6659,N_6593,N_6569);
xor U6660 (N_6660,N_6523,N_6589);
or U6661 (N_6661,N_6513,N_6500);
and U6662 (N_6662,N_6531,N_6500);
nor U6663 (N_6663,N_6533,N_6599);
nor U6664 (N_6664,N_6575,N_6556);
nand U6665 (N_6665,N_6504,N_6545);
nand U6666 (N_6666,N_6577,N_6518);
nor U6667 (N_6667,N_6565,N_6553);
nor U6668 (N_6668,N_6543,N_6548);
nor U6669 (N_6669,N_6518,N_6529);
xnor U6670 (N_6670,N_6583,N_6528);
nand U6671 (N_6671,N_6593,N_6520);
or U6672 (N_6672,N_6564,N_6513);
or U6673 (N_6673,N_6594,N_6519);
nand U6674 (N_6674,N_6549,N_6573);
and U6675 (N_6675,N_6552,N_6561);
nor U6676 (N_6676,N_6513,N_6573);
or U6677 (N_6677,N_6567,N_6545);
nand U6678 (N_6678,N_6540,N_6563);
and U6679 (N_6679,N_6533,N_6532);
xnor U6680 (N_6680,N_6519,N_6575);
and U6681 (N_6681,N_6511,N_6544);
nor U6682 (N_6682,N_6547,N_6519);
xnor U6683 (N_6683,N_6549,N_6502);
and U6684 (N_6684,N_6515,N_6585);
xor U6685 (N_6685,N_6508,N_6567);
nand U6686 (N_6686,N_6524,N_6533);
nor U6687 (N_6687,N_6505,N_6546);
and U6688 (N_6688,N_6559,N_6576);
and U6689 (N_6689,N_6563,N_6529);
or U6690 (N_6690,N_6542,N_6575);
xnor U6691 (N_6691,N_6563,N_6573);
or U6692 (N_6692,N_6558,N_6524);
xnor U6693 (N_6693,N_6589,N_6547);
xnor U6694 (N_6694,N_6526,N_6549);
nand U6695 (N_6695,N_6505,N_6555);
xnor U6696 (N_6696,N_6513,N_6561);
and U6697 (N_6697,N_6552,N_6507);
nor U6698 (N_6698,N_6584,N_6576);
nor U6699 (N_6699,N_6515,N_6571);
and U6700 (N_6700,N_6695,N_6688);
or U6701 (N_6701,N_6617,N_6665);
nor U6702 (N_6702,N_6625,N_6621);
or U6703 (N_6703,N_6658,N_6600);
nor U6704 (N_6704,N_6614,N_6652);
and U6705 (N_6705,N_6689,N_6641);
nor U6706 (N_6706,N_6673,N_6699);
nand U6707 (N_6707,N_6683,N_6622);
nor U6708 (N_6708,N_6675,N_6606);
nor U6709 (N_6709,N_6601,N_6627);
and U6710 (N_6710,N_6632,N_6678);
nor U6711 (N_6711,N_6647,N_6679);
nand U6712 (N_6712,N_6643,N_6649);
nor U6713 (N_6713,N_6680,N_6618);
or U6714 (N_6714,N_6623,N_6616);
nand U6715 (N_6715,N_6655,N_6659);
nand U6716 (N_6716,N_6687,N_6639);
nand U6717 (N_6717,N_6697,N_6646);
nor U6718 (N_6718,N_6671,N_6609);
nor U6719 (N_6719,N_6611,N_6696);
nand U6720 (N_6720,N_6619,N_6691);
xor U6721 (N_6721,N_6610,N_6638);
nor U6722 (N_6722,N_6612,N_6660);
or U6723 (N_6723,N_6651,N_6620);
nand U6724 (N_6724,N_6613,N_6657);
or U6725 (N_6725,N_6634,N_6667);
nor U6726 (N_6726,N_6624,N_6677);
xor U6727 (N_6727,N_6693,N_6653);
and U6728 (N_6728,N_6605,N_6690);
xnor U6729 (N_6729,N_6668,N_6650);
nand U6730 (N_6730,N_6692,N_6637);
or U6731 (N_6731,N_6698,N_6664);
nand U6732 (N_6732,N_6661,N_6682);
and U6733 (N_6733,N_6654,N_6607);
nand U6734 (N_6734,N_6674,N_6672);
and U6735 (N_6735,N_6629,N_6644);
nand U6736 (N_6736,N_6630,N_6684);
and U6737 (N_6737,N_6676,N_6633);
and U6738 (N_6738,N_6635,N_6694);
or U6739 (N_6739,N_6656,N_6670);
nor U6740 (N_6740,N_6685,N_6662);
nand U6741 (N_6741,N_6603,N_6615);
nand U6742 (N_6742,N_6642,N_6648);
xor U6743 (N_6743,N_6681,N_6631);
nor U6744 (N_6744,N_6645,N_6663);
nor U6745 (N_6745,N_6666,N_6604);
and U6746 (N_6746,N_6628,N_6608);
nand U6747 (N_6747,N_6602,N_6626);
nor U6748 (N_6748,N_6640,N_6686);
xnor U6749 (N_6749,N_6636,N_6669);
nor U6750 (N_6750,N_6671,N_6647);
or U6751 (N_6751,N_6604,N_6615);
nand U6752 (N_6752,N_6643,N_6667);
nor U6753 (N_6753,N_6662,N_6606);
and U6754 (N_6754,N_6670,N_6627);
and U6755 (N_6755,N_6635,N_6670);
xnor U6756 (N_6756,N_6658,N_6684);
or U6757 (N_6757,N_6618,N_6631);
nand U6758 (N_6758,N_6611,N_6689);
nor U6759 (N_6759,N_6670,N_6600);
and U6760 (N_6760,N_6657,N_6665);
nor U6761 (N_6761,N_6684,N_6621);
xor U6762 (N_6762,N_6603,N_6609);
nor U6763 (N_6763,N_6645,N_6636);
nand U6764 (N_6764,N_6602,N_6650);
or U6765 (N_6765,N_6636,N_6691);
nor U6766 (N_6766,N_6641,N_6620);
or U6767 (N_6767,N_6661,N_6697);
nor U6768 (N_6768,N_6651,N_6632);
nor U6769 (N_6769,N_6662,N_6622);
nor U6770 (N_6770,N_6684,N_6653);
nor U6771 (N_6771,N_6652,N_6666);
nor U6772 (N_6772,N_6691,N_6687);
nor U6773 (N_6773,N_6661,N_6664);
or U6774 (N_6774,N_6603,N_6611);
xor U6775 (N_6775,N_6615,N_6691);
nand U6776 (N_6776,N_6612,N_6640);
nor U6777 (N_6777,N_6608,N_6639);
and U6778 (N_6778,N_6665,N_6651);
or U6779 (N_6779,N_6692,N_6691);
and U6780 (N_6780,N_6607,N_6678);
nor U6781 (N_6781,N_6636,N_6624);
and U6782 (N_6782,N_6630,N_6680);
and U6783 (N_6783,N_6633,N_6694);
nor U6784 (N_6784,N_6666,N_6684);
nand U6785 (N_6785,N_6669,N_6615);
nor U6786 (N_6786,N_6615,N_6699);
and U6787 (N_6787,N_6674,N_6651);
nand U6788 (N_6788,N_6662,N_6669);
nor U6789 (N_6789,N_6659,N_6605);
and U6790 (N_6790,N_6634,N_6651);
or U6791 (N_6791,N_6650,N_6631);
and U6792 (N_6792,N_6647,N_6661);
or U6793 (N_6793,N_6615,N_6654);
or U6794 (N_6794,N_6608,N_6621);
nand U6795 (N_6795,N_6632,N_6653);
nand U6796 (N_6796,N_6602,N_6696);
and U6797 (N_6797,N_6617,N_6637);
nand U6798 (N_6798,N_6662,N_6688);
and U6799 (N_6799,N_6640,N_6613);
xnor U6800 (N_6800,N_6783,N_6715);
or U6801 (N_6801,N_6781,N_6765);
nor U6802 (N_6802,N_6752,N_6799);
or U6803 (N_6803,N_6757,N_6777);
nor U6804 (N_6804,N_6725,N_6776);
nor U6805 (N_6805,N_6712,N_6736);
and U6806 (N_6806,N_6740,N_6741);
or U6807 (N_6807,N_6762,N_6787);
and U6808 (N_6808,N_6709,N_6796);
and U6809 (N_6809,N_6728,N_6731);
nor U6810 (N_6810,N_6779,N_6778);
or U6811 (N_6811,N_6742,N_6753);
nand U6812 (N_6812,N_6747,N_6797);
or U6813 (N_6813,N_6700,N_6758);
nand U6814 (N_6814,N_6724,N_6721);
nand U6815 (N_6815,N_6719,N_6743);
nand U6816 (N_6816,N_6795,N_6716);
nand U6817 (N_6817,N_6794,N_6703);
and U6818 (N_6818,N_6766,N_6734);
xnor U6819 (N_6819,N_6791,N_6702);
nor U6820 (N_6820,N_6722,N_6789);
xor U6821 (N_6821,N_6763,N_6744);
nand U6822 (N_6822,N_6723,N_6775);
nand U6823 (N_6823,N_6755,N_6717);
or U6824 (N_6824,N_6748,N_6714);
nor U6825 (N_6825,N_6730,N_6739);
nor U6826 (N_6826,N_6704,N_6750);
xor U6827 (N_6827,N_6720,N_6745);
nand U6828 (N_6828,N_6780,N_6746);
xor U6829 (N_6829,N_6782,N_6760);
xnor U6830 (N_6830,N_6754,N_6772);
and U6831 (N_6831,N_6764,N_6759);
and U6832 (N_6832,N_6732,N_6733);
nand U6833 (N_6833,N_6729,N_6711);
nor U6834 (N_6834,N_6756,N_6710);
and U6835 (N_6835,N_6751,N_6708);
or U6836 (N_6836,N_6713,N_6767);
and U6837 (N_6837,N_6788,N_6737);
nand U6838 (N_6838,N_6701,N_6749);
or U6839 (N_6839,N_6790,N_6774);
and U6840 (N_6840,N_6706,N_6773);
and U6841 (N_6841,N_6718,N_6771);
and U6842 (N_6842,N_6726,N_6793);
or U6843 (N_6843,N_6707,N_6761);
xnor U6844 (N_6844,N_6798,N_6769);
or U6845 (N_6845,N_6705,N_6727);
nand U6846 (N_6846,N_6784,N_6768);
or U6847 (N_6847,N_6792,N_6770);
or U6848 (N_6848,N_6735,N_6738);
and U6849 (N_6849,N_6786,N_6785);
or U6850 (N_6850,N_6750,N_6778);
xor U6851 (N_6851,N_6780,N_6777);
nand U6852 (N_6852,N_6714,N_6794);
and U6853 (N_6853,N_6772,N_6745);
or U6854 (N_6854,N_6749,N_6739);
nand U6855 (N_6855,N_6738,N_6702);
nand U6856 (N_6856,N_6750,N_6734);
nand U6857 (N_6857,N_6766,N_6746);
or U6858 (N_6858,N_6704,N_6745);
xor U6859 (N_6859,N_6721,N_6776);
xnor U6860 (N_6860,N_6793,N_6763);
or U6861 (N_6861,N_6722,N_6701);
or U6862 (N_6862,N_6790,N_6795);
nor U6863 (N_6863,N_6765,N_6788);
xnor U6864 (N_6864,N_6772,N_6706);
nor U6865 (N_6865,N_6788,N_6701);
or U6866 (N_6866,N_6756,N_6746);
xor U6867 (N_6867,N_6783,N_6728);
and U6868 (N_6868,N_6788,N_6795);
nand U6869 (N_6869,N_6792,N_6797);
nand U6870 (N_6870,N_6750,N_6774);
and U6871 (N_6871,N_6760,N_6779);
xnor U6872 (N_6872,N_6709,N_6750);
nand U6873 (N_6873,N_6728,N_6751);
xnor U6874 (N_6874,N_6707,N_6754);
and U6875 (N_6875,N_6784,N_6708);
nand U6876 (N_6876,N_6749,N_6768);
and U6877 (N_6877,N_6724,N_6793);
nor U6878 (N_6878,N_6799,N_6775);
or U6879 (N_6879,N_6746,N_6753);
and U6880 (N_6880,N_6758,N_6727);
or U6881 (N_6881,N_6763,N_6717);
xnor U6882 (N_6882,N_6772,N_6775);
and U6883 (N_6883,N_6713,N_6783);
nor U6884 (N_6884,N_6774,N_6745);
nor U6885 (N_6885,N_6786,N_6720);
xor U6886 (N_6886,N_6771,N_6702);
or U6887 (N_6887,N_6778,N_6711);
nor U6888 (N_6888,N_6781,N_6716);
xor U6889 (N_6889,N_6721,N_6787);
nand U6890 (N_6890,N_6740,N_6701);
or U6891 (N_6891,N_6795,N_6705);
or U6892 (N_6892,N_6769,N_6740);
nand U6893 (N_6893,N_6710,N_6750);
nand U6894 (N_6894,N_6738,N_6743);
nand U6895 (N_6895,N_6764,N_6710);
and U6896 (N_6896,N_6749,N_6771);
and U6897 (N_6897,N_6714,N_6700);
xnor U6898 (N_6898,N_6790,N_6763);
nor U6899 (N_6899,N_6795,N_6709);
nor U6900 (N_6900,N_6812,N_6814);
xnor U6901 (N_6901,N_6835,N_6839);
or U6902 (N_6902,N_6837,N_6853);
and U6903 (N_6903,N_6820,N_6824);
or U6904 (N_6904,N_6881,N_6851);
nor U6905 (N_6905,N_6846,N_6882);
and U6906 (N_6906,N_6815,N_6878);
nor U6907 (N_6907,N_6821,N_6834);
nor U6908 (N_6908,N_6807,N_6849);
and U6909 (N_6909,N_6875,N_6861);
xor U6910 (N_6910,N_6864,N_6802);
and U6911 (N_6911,N_6801,N_6866);
nor U6912 (N_6912,N_6850,N_6894);
nand U6913 (N_6913,N_6877,N_6845);
nor U6914 (N_6914,N_6819,N_6813);
nor U6915 (N_6915,N_6887,N_6872);
and U6916 (N_6916,N_6859,N_6822);
and U6917 (N_6917,N_6862,N_6867);
or U6918 (N_6918,N_6869,N_6855);
xor U6919 (N_6919,N_6874,N_6830);
nor U6920 (N_6920,N_6896,N_6827);
nand U6921 (N_6921,N_6829,N_6826);
nand U6922 (N_6922,N_6876,N_6809);
nand U6923 (N_6923,N_6805,N_6884);
and U6924 (N_6924,N_6868,N_6880);
nand U6925 (N_6925,N_6865,N_6825);
nand U6926 (N_6926,N_6897,N_6836);
nor U6927 (N_6927,N_6842,N_6854);
nor U6928 (N_6928,N_6890,N_6810);
and U6929 (N_6929,N_6816,N_6870);
or U6930 (N_6930,N_6883,N_6899);
and U6931 (N_6931,N_6857,N_6817);
xnor U6932 (N_6932,N_6898,N_6804);
or U6933 (N_6933,N_6847,N_6871);
or U6934 (N_6934,N_6879,N_6811);
and U6935 (N_6935,N_6885,N_6840);
and U6936 (N_6936,N_6828,N_6873);
or U6937 (N_6937,N_6803,N_6856);
nor U6938 (N_6938,N_6808,N_6831);
nand U6939 (N_6939,N_6886,N_6844);
and U6940 (N_6940,N_6806,N_6858);
xnor U6941 (N_6941,N_6893,N_6889);
xor U6942 (N_6942,N_6833,N_6891);
nor U6943 (N_6943,N_6832,N_6860);
and U6944 (N_6944,N_6895,N_6852);
nand U6945 (N_6945,N_6841,N_6863);
nand U6946 (N_6946,N_6848,N_6843);
nor U6947 (N_6947,N_6888,N_6800);
nand U6948 (N_6948,N_6838,N_6892);
xor U6949 (N_6949,N_6823,N_6818);
and U6950 (N_6950,N_6841,N_6865);
or U6951 (N_6951,N_6897,N_6863);
and U6952 (N_6952,N_6826,N_6840);
xnor U6953 (N_6953,N_6889,N_6891);
and U6954 (N_6954,N_6871,N_6814);
xnor U6955 (N_6955,N_6804,N_6809);
xnor U6956 (N_6956,N_6872,N_6837);
or U6957 (N_6957,N_6898,N_6841);
or U6958 (N_6958,N_6827,N_6858);
xor U6959 (N_6959,N_6897,N_6850);
and U6960 (N_6960,N_6830,N_6816);
or U6961 (N_6961,N_6807,N_6828);
nand U6962 (N_6962,N_6823,N_6864);
nor U6963 (N_6963,N_6880,N_6847);
nand U6964 (N_6964,N_6844,N_6873);
and U6965 (N_6965,N_6885,N_6850);
nor U6966 (N_6966,N_6877,N_6862);
and U6967 (N_6967,N_6803,N_6897);
or U6968 (N_6968,N_6812,N_6820);
xor U6969 (N_6969,N_6826,N_6893);
or U6970 (N_6970,N_6816,N_6876);
and U6971 (N_6971,N_6876,N_6849);
or U6972 (N_6972,N_6856,N_6835);
or U6973 (N_6973,N_6860,N_6835);
nor U6974 (N_6974,N_6866,N_6817);
nand U6975 (N_6975,N_6824,N_6850);
nand U6976 (N_6976,N_6874,N_6850);
and U6977 (N_6977,N_6873,N_6829);
or U6978 (N_6978,N_6898,N_6843);
nor U6979 (N_6979,N_6822,N_6872);
nor U6980 (N_6980,N_6832,N_6858);
nand U6981 (N_6981,N_6836,N_6813);
and U6982 (N_6982,N_6820,N_6838);
and U6983 (N_6983,N_6851,N_6894);
nor U6984 (N_6984,N_6838,N_6896);
and U6985 (N_6985,N_6828,N_6809);
nand U6986 (N_6986,N_6806,N_6800);
or U6987 (N_6987,N_6856,N_6864);
nand U6988 (N_6988,N_6823,N_6872);
or U6989 (N_6989,N_6831,N_6804);
nand U6990 (N_6990,N_6856,N_6828);
xnor U6991 (N_6991,N_6852,N_6858);
nand U6992 (N_6992,N_6801,N_6863);
nand U6993 (N_6993,N_6855,N_6861);
and U6994 (N_6994,N_6842,N_6806);
nor U6995 (N_6995,N_6884,N_6836);
or U6996 (N_6996,N_6896,N_6811);
nand U6997 (N_6997,N_6845,N_6872);
or U6998 (N_6998,N_6850,N_6811);
nor U6999 (N_6999,N_6837,N_6814);
xor U7000 (N_7000,N_6908,N_6935);
nand U7001 (N_7001,N_6934,N_6912);
or U7002 (N_7002,N_6996,N_6961);
or U7003 (N_7003,N_6973,N_6907);
or U7004 (N_7004,N_6901,N_6986);
nor U7005 (N_7005,N_6999,N_6978);
nand U7006 (N_7006,N_6982,N_6958);
nand U7007 (N_7007,N_6947,N_6926);
nor U7008 (N_7008,N_6976,N_6954);
nor U7009 (N_7009,N_6930,N_6992);
nand U7010 (N_7010,N_6922,N_6914);
or U7011 (N_7011,N_6949,N_6940);
nor U7012 (N_7012,N_6968,N_6987);
and U7013 (N_7013,N_6988,N_6969);
or U7014 (N_7014,N_6933,N_6905);
nor U7015 (N_7015,N_6945,N_6917);
or U7016 (N_7016,N_6989,N_6937);
or U7017 (N_7017,N_6927,N_6995);
nand U7018 (N_7018,N_6963,N_6913);
nand U7019 (N_7019,N_6967,N_6943);
and U7020 (N_7020,N_6964,N_6932);
or U7021 (N_7021,N_6960,N_6974);
and U7022 (N_7022,N_6915,N_6991);
and U7023 (N_7023,N_6924,N_6971);
and U7024 (N_7024,N_6925,N_6980);
and U7025 (N_7025,N_6910,N_6950);
and U7026 (N_7026,N_6966,N_6942);
and U7027 (N_7027,N_6948,N_6998);
nand U7028 (N_7028,N_6993,N_6939);
nor U7029 (N_7029,N_6981,N_6959);
xor U7030 (N_7030,N_6975,N_6962);
and U7031 (N_7031,N_6972,N_6928);
nand U7032 (N_7032,N_6931,N_6918);
and U7033 (N_7033,N_6994,N_6956);
xnor U7034 (N_7034,N_6900,N_6929);
nand U7035 (N_7035,N_6936,N_6902);
xnor U7036 (N_7036,N_6923,N_6965);
or U7037 (N_7037,N_6955,N_6903);
nand U7038 (N_7038,N_6953,N_6920);
xor U7039 (N_7039,N_6979,N_6906);
and U7040 (N_7040,N_6957,N_6919);
nand U7041 (N_7041,N_6983,N_6970);
nor U7042 (N_7042,N_6997,N_6916);
nand U7043 (N_7043,N_6952,N_6944);
or U7044 (N_7044,N_6911,N_6921);
or U7045 (N_7045,N_6990,N_6938);
or U7046 (N_7046,N_6946,N_6984);
nor U7047 (N_7047,N_6904,N_6951);
nor U7048 (N_7048,N_6941,N_6909);
nor U7049 (N_7049,N_6977,N_6985);
or U7050 (N_7050,N_6918,N_6939);
nand U7051 (N_7051,N_6988,N_6918);
nand U7052 (N_7052,N_6933,N_6939);
nand U7053 (N_7053,N_6977,N_6955);
nor U7054 (N_7054,N_6996,N_6921);
nor U7055 (N_7055,N_6987,N_6996);
or U7056 (N_7056,N_6908,N_6930);
nor U7057 (N_7057,N_6932,N_6976);
nand U7058 (N_7058,N_6981,N_6986);
or U7059 (N_7059,N_6963,N_6951);
nand U7060 (N_7060,N_6927,N_6913);
and U7061 (N_7061,N_6961,N_6902);
and U7062 (N_7062,N_6954,N_6963);
nor U7063 (N_7063,N_6984,N_6907);
and U7064 (N_7064,N_6946,N_6971);
xor U7065 (N_7065,N_6976,N_6925);
and U7066 (N_7066,N_6945,N_6993);
or U7067 (N_7067,N_6919,N_6916);
nand U7068 (N_7068,N_6904,N_6970);
nand U7069 (N_7069,N_6966,N_6974);
or U7070 (N_7070,N_6952,N_6932);
xnor U7071 (N_7071,N_6990,N_6940);
or U7072 (N_7072,N_6926,N_6941);
or U7073 (N_7073,N_6954,N_6991);
and U7074 (N_7074,N_6958,N_6961);
nand U7075 (N_7075,N_6948,N_6990);
and U7076 (N_7076,N_6972,N_6977);
and U7077 (N_7077,N_6978,N_6913);
nor U7078 (N_7078,N_6990,N_6973);
xor U7079 (N_7079,N_6932,N_6900);
or U7080 (N_7080,N_6999,N_6958);
and U7081 (N_7081,N_6939,N_6970);
nand U7082 (N_7082,N_6978,N_6986);
nor U7083 (N_7083,N_6956,N_6912);
nor U7084 (N_7084,N_6938,N_6922);
nand U7085 (N_7085,N_6908,N_6902);
nor U7086 (N_7086,N_6940,N_6946);
xnor U7087 (N_7087,N_6948,N_6912);
xnor U7088 (N_7088,N_6910,N_6956);
and U7089 (N_7089,N_6918,N_6969);
nand U7090 (N_7090,N_6966,N_6996);
nor U7091 (N_7091,N_6914,N_6974);
nor U7092 (N_7092,N_6912,N_6987);
nor U7093 (N_7093,N_6992,N_6990);
or U7094 (N_7094,N_6984,N_6975);
or U7095 (N_7095,N_6922,N_6962);
nor U7096 (N_7096,N_6959,N_6917);
and U7097 (N_7097,N_6942,N_6948);
nand U7098 (N_7098,N_6973,N_6950);
nand U7099 (N_7099,N_6935,N_6998);
nor U7100 (N_7100,N_7009,N_7067);
nand U7101 (N_7101,N_7094,N_7001);
nor U7102 (N_7102,N_7028,N_7082);
or U7103 (N_7103,N_7092,N_7016);
nor U7104 (N_7104,N_7098,N_7021);
xnor U7105 (N_7105,N_7079,N_7091);
nand U7106 (N_7106,N_7069,N_7010);
or U7107 (N_7107,N_7057,N_7034);
or U7108 (N_7108,N_7078,N_7035);
nor U7109 (N_7109,N_7083,N_7051);
nor U7110 (N_7110,N_7025,N_7058);
nand U7111 (N_7111,N_7075,N_7086);
nand U7112 (N_7112,N_7041,N_7073);
nand U7113 (N_7113,N_7071,N_7022);
or U7114 (N_7114,N_7093,N_7011);
and U7115 (N_7115,N_7030,N_7039);
nand U7116 (N_7116,N_7059,N_7070);
xnor U7117 (N_7117,N_7049,N_7026);
nand U7118 (N_7118,N_7090,N_7089);
nor U7119 (N_7119,N_7024,N_7096);
nor U7120 (N_7120,N_7076,N_7023);
nor U7121 (N_7121,N_7020,N_7074);
nand U7122 (N_7122,N_7014,N_7085);
nand U7123 (N_7123,N_7072,N_7048);
or U7124 (N_7124,N_7003,N_7013);
and U7125 (N_7125,N_7012,N_7015);
and U7126 (N_7126,N_7064,N_7068);
and U7127 (N_7127,N_7046,N_7033);
nor U7128 (N_7128,N_7077,N_7042);
or U7129 (N_7129,N_7027,N_7088);
nor U7130 (N_7130,N_7005,N_7029);
nor U7131 (N_7131,N_7008,N_7043);
nor U7132 (N_7132,N_7080,N_7097);
or U7133 (N_7133,N_7081,N_7063);
and U7134 (N_7134,N_7017,N_7084);
xor U7135 (N_7135,N_7031,N_7047);
nand U7136 (N_7136,N_7018,N_7045);
and U7137 (N_7137,N_7040,N_7095);
nand U7138 (N_7138,N_7036,N_7062);
and U7139 (N_7139,N_7061,N_7056);
xor U7140 (N_7140,N_7006,N_7065);
xnor U7141 (N_7141,N_7066,N_7050);
xor U7142 (N_7142,N_7052,N_7099);
and U7143 (N_7143,N_7032,N_7037);
or U7144 (N_7144,N_7087,N_7044);
nor U7145 (N_7145,N_7002,N_7055);
or U7146 (N_7146,N_7060,N_7038);
and U7147 (N_7147,N_7019,N_7007);
and U7148 (N_7148,N_7004,N_7054);
or U7149 (N_7149,N_7000,N_7053);
or U7150 (N_7150,N_7046,N_7018);
and U7151 (N_7151,N_7085,N_7026);
and U7152 (N_7152,N_7014,N_7058);
and U7153 (N_7153,N_7013,N_7035);
and U7154 (N_7154,N_7063,N_7042);
and U7155 (N_7155,N_7029,N_7084);
and U7156 (N_7156,N_7023,N_7019);
or U7157 (N_7157,N_7062,N_7020);
nor U7158 (N_7158,N_7007,N_7018);
nand U7159 (N_7159,N_7075,N_7037);
or U7160 (N_7160,N_7044,N_7034);
nor U7161 (N_7161,N_7036,N_7023);
and U7162 (N_7162,N_7029,N_7023);
or U7163 (N_7163,N_7046,N_7063);
nor U7164 (N_7164,N_7026,N_7035);
nor U7165 (N_7165,N_7065,N_7023);
xor U7166 (N_7166,N_7082,N_7095);
nand U7167 (N_7167,N_7064,N_7085);
or U7168 (N_7168,N_7078,N_7036);
nand U7169 (N_7169,N_7044,N_7024);
and U7170 (N_7170,N_7016,N_7073);
nor U7171 (N_7171,N_7047,N_7094);
and U7172 (N_7172,N_7031,N_7095);
nor U7173 (N_7173,N_7020,N_7032);
and U7174 (N_7174,N_7049,N_7080);
or U7175 (N_7175,N_7052,N_7042);
or U7176 (N_7176,N_7018,N_7082);
and U7177 (N_7177,N_7008,N_7026);
or U7178 (N_7178,N_7089,N_7040);
and U7179 (N_7179,N_7089,N_7062);
and U7180 (N_7180,N_7022,N_7095);
or U7181 (N_7181,N_7022,N_7026);
and U7182 (N_7182,N_7096,N_7029);
and U7183 (N_7183,N_7012,N_7010);
and U7184 (N_7184,N_7065,N_7084);
or U7185 (N_7185,N_7054,N_7076);
nor U7186 (N_7186,N_7057,N_7077);
or U7187 (N_7187,N_7067,N_7045);
or U7188 (N_7188,N_7099,N_7077);
nor U7189 (N_7189,N_7093,N_7091);
or U7190 (N_7190,N_7044,N_7042);
and U7191 (N_7191,N_7046,N_7000);
or U7192 (N_7192,N_7030,N_7063);
nand U7193 (N_7193,N_7003,N_7067);
or U7194 (N_7194,N_7047,N_7044);
nand U7195 (N_7195,N_7074,N_7024);
xnor U7196 (N_7196,N_7045,N_7040);
and U7197 (N_7197,N_7009,N_7037);
and U7198 (N_7198,N_7094,N_7043);
or U7199 (N_7199,N_7036,N_7046);
xnor U7200 (N_7200,N_7186,N_7115);
nand U7201 (N_7201,N_7131,N_7168);
nor U7202 (N_7202,N_7193,N_7185);
nand U7203 (N_7203,N_7172,N_7108);
nand U7204 (N_7204,N_7167,N_7104);
or U7205 (N_7205,N_7177,N_7147);
nand U7206 (N_7206,N_7179,N_7190);
or U7207 (N_7207,N_7126,N_7103);
nand U7208 (N_7208,N_7140,N_7109);
nor U7209 (N_7209,N_7137,N_7112);
nor U7210 (N_7210,N_7142,N_7165);
xor U7211 (N_7211,N_7124,N_7133);
and U7212 (N_7212,N_7163,N_7136);
nand U7213 (N_7213,N_7102,N_7150);
and U7214 (N_7214,N_7188,N_7107);
nand U7215 (N_7215,N_7143,N_7141);
nor U7216 (N_7216,N_7132,N_7139);
or U7217 (N_7217,N_7160,N_7183);
or U7218 (N_7218,N_7182,N_7197);
nor U7219 (N_7219,N_7128,N_7116);
nor U7220 (N_7220,N_7156,N_7152);
nor U7221 (N_7221,N_7191,N_7170);
nand U7222 (N_7222,N_7151,N_7175);
and U7223 (N_7223,N_7161,N_7145);
nand U7224 (N_7224,N_7149,N_7125);
and U7225 (N_7225,N_7144,N_7181);
nor U7226 (N_7226,N_7194,N_7158);
nand U7227 (N_7227,N_7153,N_7180);
xor U7228 (N_7228,N_7110,N_7127);
nand U7229 (N_7229,N_7148,N_7157);
nor U7230 (N_7230,N_7118,N_7187);
and U7231 (N_7231,N_7173,N_7176);
nor U7232 (N_7232,N_7113,N_7192);
nand U7233 (N_7233,N_7171,N_7122);
and U7234 (N_7234,N_7178,N_7184);
nand U7235 (N_7235,N_7162,N_7199);
xnor U7236 (N_7236,N_7134,N_7106);
nor U7237 (N_7237,N_7166,N_7111);
or U7238 (N_7238,N_7169,N_7189);
nor U7239 (N_7239,N_7155,N_7174);
nand U7240 (N_7240,N_7164,N_7119);
and U7241 (N_7241,N_7195,N_7105);
and U7242 (N_7242,N_7159,N_7121);
or U7243 (N_7243,N_7135,N_7146);
and U7244 (N_7244,N_7138,N_7130);
or U7245 (N_7245,N_7100,N_7198);
or U7246 (N_7246,N_7123,N_7129);
nor U7247 (N_7247,N_7117,N_7114);
xor U7248 (N_7248,N_7154,N_7120);
nor U7249 (N_7249,N_7196,N_7101);
or U7250 (N_7250,N_7134,N_7140);
and U7251 (N_7251,N_7191,N_7115);
or U7252 (N_7252,N_7185,N_7176);
or U7253 (N_7253,N_7154,N_7197);
and U7254 (N_7254,N_7197,N_7140);
and U7255 (N_7255,N_7196,N_7124);
xnor U7256 (N_7256,N_7197,N_7113);
nor U7257 (N_7257,N_7157,N_7186);
or U7258 (N_7258,N_7125,N_7111);
or U7259 (N_7259,N_7176,N_7183);
xor U7260 (N_7260,N_7158,N_7175);
and U7261 (N_7261,N_7172,N_7197);
nor U7262 (N_7262,N_7153,N_7168);
nor U7263 (N_7263,N_7102,N_7152);
nand U7264 (N_7264,N_7142,N_7177);
nand U7265 (N_7265,N_7162,N_7115);
xnor U7266 (N_7266,N_7197,N_7132);
nand U7267 (N_7267,N_7181,N_7162);
nor U7268 (N_7268,N_7142,N_7194);
nor U7269 (N_7269,N_7160,N_7104);
nor U7270 (N_7270,N_7130,N_7143);
or U7271 (N_7271,N_7189,N_7135);
or U7272 (N_7272,N_7155,N_7121);
nor U7273 (N_7273,N_7143,N_7124);
nor U7274 (N_7274,N_7195,N_7165);
nand U7275 (N_7275,N_7162,N_7182);
or U7276 (N_7276,N_7194,N_7135);
nor U7277 (N_7277,N_7109,N_7157);
or U7278 (N_7278,N_7165,N_7184);
nor U7279 (N_7279,N_7199,N_7170);
or U7280 (N_7280,N_7103,N_7163);
or U7281 (N_7281,N_7135,N_7183);
nor U7282 (N_7282,N_7102,N_7137);
and U7283 (N_7283,N_7107,N_7149);
nor U7284 (N_7284,N_7181,N_7174);
or U7285 (N_7285,N_7177,N_7171);
nor U7286 (N_7286,N_7118,N_7131);
or U7287 (N_7287,N_7112,N_7165);
and U7288 (N_7288,N_7122,N_7163);
nand U7289 (N_7289,N_7130,N_7185);
or U7290 (N_7290,N_7162,N_7160);
or U7291 (N_7291,N_7158,N_7137);
nand U7292 (N_7292,N_7164,N_7182);
and U7293 (N_7293,N_7192,N_7165);
and U7294 (N_7294,N_7181,N_7139);
and U7295 (N_7295,N_7176,N_7151);
or U7296 (N_7296,N_7104,N_7132);
nand U7297 (N_7297,N_7164,N_7121);
or U7298 (N_7298,N_7132,N_7179);
nand U7299 (N_7299,N_7113,N_7137);
and U7300 (N_7300,N_7222,N_7289);
or U7301 (N_7301,N_7215,N_7224);
nand U7302 (N_7302,N_7225,N_7219);
nor U7303 (N_7303,N_7292,N_7295);
xnor U7304 (N_7304,N_7284,N_7230);
and U7305 (N_7305,N_7255,N_7266);
and U7306 (N_7306,N_7273,N_7210);
and U7307 (N_7307,N_7226,N_7204);
or U7308 (N_7308,N_7296,N_7205);
nor U7309 (N_7309,N_7269,N_7293);
nand U7310 (N_7310,N_7288,N_7246);
and U7311 (N_7311,N_7252,N_7207);
nand U7312 (N_7312,N_7238,N_7299);
xor U7313 (N_7313,N_7249,N_7217);
xor U7314 (N_7314,N_7270,N_7240);
nand U7315 (N_7315,N_7277,N_7298);
nor U7316 (N_7316,N_7254,N_7274);
nor U7317 (N_7317,N_7221,N_7237);
or U7318 (N_7318,N_7235,N_7228);
nor U7319 (N_7319,N_7234,N_7247);
and U7320 (N_7320,N_7264,N_7257);
xnor U7321 (N_7321,N_7256,N_7211);
nand U7322 (N_7322,N_7276,N_7212);
and U7323 (N_7323,N_7253,N_7287);
and U7324 (N_7324,N_7268,N_7206);
nor U7325 (N_7325,N_7259,N_7286);
and U7326 (N_7326,N_7223,N_7250);
and U7327 (N_7327,N_7282,N_7231);
nor U7328 (N_7328,N_7281,N_7260);
nand U7329 (N_7329,N_7233,N_7200);
and U7330 (N_7330,N_7244,N_7278);
or U7331 (N_7331,N_7220,N_7232);
xor U7332 (N_7332,N_7229,N_7272);
or U7333 (N_7333,N_7261,N_7209);
nand U7334 (N_7334,N_7241,N_7265);
or U7335 (N_7335,N_7294,N_7267);
nand U7336 (N_7336,N_7218,N_7297);
nor U7337 (N_7337,N_7242,N_7262);
nand U7338 (N_7338,N_7202,N_7291);
and U7339 (N_7339,N_7214,N_7275);
and U7340 (N_7340,N_7290,N_7203);
nand U7341 (N_7341,N_7251,N_7280);
and U7342 (N_7342,N_7285,N_7239);
nand U7343 (N_7343,N_7271,N_7258);
xor U7344 (N_7344,N_7216,N_7201);
nor U7345 (N_7345,N_7279,N_7243);
and U7346 (N_7346,N_7263,N_7245);
and U7347 (N_7347,N_7236,N_7283);
nand U7348 (N_7348,N_7208,N_7248);
nand U7349 (N_7349,N_7213,N_7227);
nor U7350 (N_7350,N_7245,N_7211);
nand U7351 (N_7351,N_7257,N_7252);
xnor U7352 (N_7352,N_7242,N_7204);
xnor U7353 (N_7353,N_7231,N_7243);
and U7354 (N_7354,N_7218,N_7211);
nand U7355 (N_7355,N_7218,N_7228);
xor U7356 (N_7356,N_7245,N_7229);
nand U7357 (N_7357,N_7298,N_7232);
or U7358 (N_7358,N_7211,N_7232);
and U7359 (N_7359,N_7268,N_7291);
nand U7360 (N_7360,N_7271,N_7242);
nand U7361 (N_7361,N_7232,N_7283);
nand U7362 (N_7362,N_7217,N_7224);
nor U7363 (N_7363,N_7263,N_7202);
or U7364 (N_7364,N_7251,N_7272);
nand U7365 (N_7365,N_7244,N_7296);
nor U7366 (N_7366,N_7224,N_7260);
xnor U7367 (N_7367,N_7291,N_7249);
nand U7368 (N_7368,N_7261,N_7269);
and U7369 (N_7369,N_7232,N_7231);
and U7370 (N_7370,N_7293,N_7209);
nor U7371 (N_7371,N_7232,N_7284);
or U7372 (N_7372,N_7236,N_7256);
or U7373 (N_7373,N_7248,N_7278);
nand U7374 (N_7374,N_7203,N_7261);
or U7375 (N_7375,N_7228,N_7210);
nor U7376 (N_7376,N_7256,N_7247);
or U7377 (N_7377,N_7220,N_7270);
nand U7378 (N_7378,N_7228,N_7229);
nor U7379 (N_7379,N_7206,N_7299);
nor U7380 (N_7380,N_7235,N_7297);
nor U7381 (N_7381,N_7226,N_7254);
nor U7382 (N_7382,N_7222,N_7247);
nor U7383 (N_7383,N_7274,N_7241);
nor U7384 (N_7384,N_7243,N_7268);
or U7385 (N_7385,N_7286,N_7299);
and U7386 (N_7386,N_7238,N_7200);
nand U7387 (N_7387,N_7228,N_7257);
nor U7388 (N_7388,N_7258,N_7200);
and U7389 (N_7389,N_7255,N_7214);
or U7390 (N_7390,N_7265,N_7258);
nand U7391 (N_7391,N_7224,N_7291);
or U7392 (N_7392,N_7203,N_7245);
nand U7393 (N_7393,N_7242,N_7283);
nand U7394 (N_7394,N_7231,N_7244);
nand U7395 (N_7395,N_7246,N_7205);
and U7396 (N_7396,N_7251,N_7239);
or U7397 (N_7397,N_7252,N_7271);
and U7398 (N_7398,N_7295,N_7222);
nor U7399 (N_7399,N_7251,N_7258);
or U7400 (N_7400,N_7399,N_7374);
nor U7401 (N_7401,N_7324,N_7340);
nand U7402 (N_7402,N_7378,N_7384);
nor U7403 (N_7403,N_7361,N_7356);
or U7404 (N_7404,N_7389,N_7321);
and U7405 (N_7405,N_7322,N_7372);
nor U7406 (N_7406,N_7327,N_7307);
or U7407 (N_7407,N_7366,N_7338);
nor U7408 (N_7408,N_7391,N_7373);
nand U7409 (N_7409,N_7376,N_7308);
nand U7410 (N_7410,N_7354,N_7362);
and U7411 (N_7411,N_7326,N_7346);
or U7412 (N_7412,N_7318,N_7347);
or U7413 (N_7413,N_7353,N_7335);
nor U7414 (N_7414,N_7320,N_7368);
nor U7415 (N_7415,N_7314,N_7383);
nand U7416 (N_7416,N_7312,N_7377);
or U7417 (N_7417,N_7375,N_7363);
nand U7418 (N_7418,N_7398,N_7325);
and U7419 (N_7419,N_7385,N_7339);
or U7420 (N_7420,N_7355,N_7360);
nor U7421 (N_7421,N_7388,N_7309);
and U7422 (N_7422,N_7344,N_7319);
nor U7423 (N_7423,N_7333,N_7393);
and U7424 (N_7424,N_7305,N_7387);
or U7425 (N_7425,N_7345,N_7301);
xnor U7426 (N_7426,N_7367,N_7328);
or U7427 (N_7427,N_7390,N_7332);
or U7428 (N_7428,N_7330,N_7342);
or U7429 (N_7429,N_7371,N_7382);
or U7430 (N_7430,N_7317,N_7336);
nor U7431 (N_7431,N_7351,N_7310);
nand U7432 (N_7432,N_7364,N_7365);
or U7433 (N_7433,N_7381,N_7316);
nand U7434 (N_7434,N_7313,N_7311);
or U7435 (N_7435,N_7331,N_7380);
or U7436 (N_7436,N_7352,N_7357);
or U7437 (N_7437,N_7359,N_7386);
nor U7438 (N_7438,N_7329,N_7306);
nor U7439 (N_7439,N_7303,N_7350);
or U7440 (N_7440,N_7379,N_7392);
and U7441 (N_7441,N_7358,N_7394);
and U7442 (N_7442,N_7348,N_7315);
xnor U7443 (N_7443,N_7302,N_7341);
nand U7444 (N_7444,N_7395,N_7323);
or U7445 (N_7445,N_7334,N_7349);
or U7446 (N_7446,N_7397,N_7337);
or U7447 (N_7447,N_7369,N_7370);
nor U7448 (N_7448,N_7300,N_7343);
nand U7449 (N_7449,N_7396,N_7304);
or U7450 (N_7450,N_7355,N_7323);
or U7451 (N_7451,N_7390,N_7395);
nor U7452 (N_7452,N_7339,N_7396);
nand U7453 (N_7453,N_7305,N_7316);
and U7454 (N_7454,N_7322,N_7304);
or U7455 (N_7455,N_7347,N_7398);
or U7456 (N_7456,N_7375,N_7347);
nor U7457 (N_7457,N_7322,N_7392);
nor U7458 (N_7458,N_7379,N_7337);
nand U7459 (N_7459,N_7332,N_7365);
nand U7460 (N_7460,N_7381,N_7397);
nor U7461 (N_7461,N_7379,N_7361);
nand U7462 (N_7462,N_7367,N_7344);
nor U7463 (N_7463,N_7378,N_7367);
and U7464 (N_7464,N_7347,N_7327);
xor U7465 (N_7465,N_7348,N_7343);
and U7466 (N_7466,N_7320,N_7332);
xor U7467 (N_7467,N_7313,N_7334);
nor U7468 (N_7468,N_7334,N_7358);
xnor U7469 (N_7469,N_7366,N_7343);
nand U7470 (N_7470,N_7321,N_7304);
or U7471 (N_7471,N_7335,N_7364);
xor U7472 (N_7472,N_7370,N_7327);
nand U7473 (N_7473,N_7380,N_7302);
nand U7474 (N_7474,N_7305,N_7370);
or U7475 (N_7475,N_7316,N_7353);
nor U7476 (N_7476,N_7317,N_7306);
nor U7477 (N_7477,N_7336,N_7361);
nand U7478 (N_7478,N_7345,N_7367);
and U7479 (N_7479,N_7354,N_7347);
and U7480 (N_7480,N_7300,N_7397);
and U7481 (N_7481,N_7322,N_7349);
xor U7482 (N_7482,N_7333,N_7372);
and U7483 (N_7483,N_7343,N_7339);
nor U7484 (N_7484,N_7386,N_7345);
or U7485 (N_7485,N_7357,N_7346);
or U7486 (N_7486,N_7357,N_7381);
and U7487 (N_7487,N_7378,N_7388);
and U7488 (N_7488,N_7329,N_7369);
or U7489 (N_7489,N_7332,N_7329);
nor U7490 (N_7490,N_7363,N_7305);
nand U7491 (N_7491,N_7399,N_7376);
nor U7492 (N_7492,N_7351,N_7348);
nand U7493 (N_7493,N_7387,N_7325);
xnor U7494 (N_7494,N_7394,N_7364);
xnor U7495 (N_7495,N_7333,N_7381);
nor U7496 (N_7496,N_7367,N_7359);
or U7497 (N_7497,N_7383,N_7318);
or U7498 (N_7498,N_7372,N_7320);
and U7499 (N_7499,N_7387,N_7385);
nor U7500 (N_7500,N_7458,N_7450);
nor U7501 (N_7501,N_7432,N_7449);
xnor U7502 (N_7502,N_7417,N_7407);
xnor U7503 (N_7503,N_7488,N_7431);
and U7504 (N_7504,N_7456,N_7494);
nor U7505 (N_7505,N_7405,N_7473);
xnor U7506 (N_7506,N_7442,N_7408);
nor U7507 (N_7507,N_7401,N_7423);
xnor U7508 (N_7508,N_7459,N_7498);
nand U7509 (N_7509,N_7471,N_7411);
nand U7510 (N_7510,N_7416,N_7491);
nand U7511 (N_7511,N_7454,N_7418);
nand U7512 (N_7512,N_7447,N_7410);
nor U7513 (N_7513,N_7451,N_7472);
nand U7514 (N_7514,N_7457,N_7439);
nand U7515 (N_7515,N_7435,N_7430);
and U7516 (N_7516,N_7461,N_7484);
nor U7517 (N_7517,N_7441,N_7470);
xor U7518 (N_7518,N_7424,N_7420);
and U7519 (N_7519,N_7404,N_7468);
nand U7520 (N_7520,N_7434,N_7436);
nor U7521 (N_7521,N_7497,N_7426);
nand U7522 (N_7522,N_7452,N_7462);
and U7523 (N_7523,N_7469,N_7480);
or U7524 (N_7524,N_7440,N_7421);
or U7525 (N_7525,N_7412,N_7478);
nand U7526 (N_7526,N_7448,N_7406);
nand U7527 (N_7527,N_7409,N_7433);
or U7528 (N_7528,N_7479,N_7482);
or U7529 (N_7529,N_7403,N_7445);
nor U7530 (N_7530,N_7475,N_7493);
xnor U7531 (N_7531,N_7443,N_7413);
and U7532 (N_7532,N_7446,N_7490);
nor U7533 (N_7533,N_7428,N_7437);
or U7534 (N_7534,N_7465,N_7438);
nor U7535 (N_7535,N_7489,N_7422);
nand U7536 (N_7536,N_7400,N_7477);
nand U7537 (N_7537,N_7453,N_7499);
nand U7538 (N_7538,N_7474,N_7419);
or U7539 (N_7539,N_7460,N_7466);
nor U7540 (N_7540,N_7429,N_7495);
xor U7541 (N_7541,N_7487,N_7415);
xnor U7542 (N_7542,N_7485,N_7486);
nor U7543 (N_7543,N_7496,N_7492);
nor U7544 (N_7544,N_7467,N_7414);
and U7545 (N_7545,N_7444,N_7455);
nor U7546 (N_7546,N_7464,N_7481);
or U7547 (N_7547,N_7463,N_7425);
and U7548 (N_7548,N_7476,N_7483);
and U7549 (N_7549,N_7427,N_7402);
nand U7550 (N_7550,N_7458,N_7415);
or U7551 (N_7551,N_7408,N_7426);
nor U7552 (N_7552,N_7485,N_7440);
and U7553 (N_7553,N_7496,N_7475);
or U7554 (N_7554,N_7463,N_7445);
nor U7555 (N_7555,N_7428,N_7491);
xor U7556 (N_7556,N_7445,N_7409);
xor U7557 (N_7557,N_7495,N_7462);
and U7558 (N_7558,N_7462,N_7414);
nor U7559 (N_7559,N_7474,N_7486);
or U7560 (N_7560,N_7408,N_7493);
and U7561 (N_7561,N_7485,N_7409);
nand U7562 (N_7562,N_7437,N_7478);
and U7563 (N_7563,N_7420,N_7419);
or U7564 (N_7564,N_7430,N_7442);
and U7565 (N_7565,N_7463,N_7438);
nand U7566 (N_7566,N_7474,N_7490);
xnor U7567 (N_7567,N_7411,N_7484);
nand U7568 (N_7568,N_7424,N_7409);
nand U7569 (N_7569,N_7495,N_7469);
or U7570 (N_7570,N_7497,N_7446);
and U7571 (N_7571,N_7468,N_7442);
nand U7572 (N_7572,N_7477,N_7470);
and U7573 (N_7573,N_7476,N_7425);
nand U7574 (N_7574,N_7451,N_7456);
xor U7575 (N_7575,N_7415,N_7449);
or U7576 (N_7576,N_7476,N_7426);
xnor U7577 (N_7577,N_7434,N_7433);
xnor U7578 (N_7578,N_7434,N_7447);
nand U7579 (N_7579,N_7468,N_7412);
nor U7580 (N_7580,N_7409,N_7481);
nor U7581 (N_7581,N_7447,N_7416);
or U7582 (N_7582,N_7459,N_7409);
nor U7583 (N_7583,N_7475,N_7470);
or U7584 (N_7584,N_7477,N_7484);
nand U7585 (N_7585,N_7416,N_7492);
nor U7586 (N_7586,N_7415,N_7439);
nand U7587 (N_7587,N_7479,N_7458);
or U7588 (N_7588,N_7456,N_7421);
and U7589 (N_7589,N_7482,N_7469);
nand U7590 (N_7590,N_7495,N_7458);
nor U7591 (N_7591,N_7424,N_7474);
or U7592 (N_7592,N_7477,N_7429);
and U7593 (N_7593,N_7479,N_7474);
nand U7594 (N_7594,N_7489,N_7498);
xnor U7595 (N_7595,N_7448,N_7436);
or U7596 (N_7596,N_7490,N_7495);
and U7597 (N_7597,N_7479,N_7497);
and U7598 (N_7598,N_7472,N_7482);
nand U7599 (N_7599,N_7416,N_7404);
or U7600 (N_7600,N_7578,N_7527);
and U7601 (N_7601,N_7568,N_7597);
xor U7602 (N_7602,N_7575,N_7520);
nand U7603 (N_7603,N_7501,N_7592);
nand U7604 (N_7604,N_7594,N_7564);
xor U7605 (N_7605,N_7505,N_7551);
and U7606 (N_7606,N_7595,N_7523);
nand U7607 (N_7607,N_7524,N_7553);
or U7608 (N_7608,N_7515,N_7565);
and U7609 (N_7609,N_7579,N_7566);
xor U7610 (N_7610,N_7580,N_7509);
nor U7611 (N_7611,N_7546,N_7587);
and U7612 (N_7612,N_7517,N_7503);
nand U7613 (N_7613,N_7532,N_7576);
nor U7614 (N_7614,N_7571,N_7557);
nand U7615 (N_7615,N_7561,N_7525);
and U7616 (N_7616,N_7540,N_7544);
nand U7617 (N_7617,N_7534,N_7530);
nor U7618 (N_7618,N_7591,N_7513);
and U7619 (N_7619,N_7533,N_7593);
or U7620 (N_7620,N_7529,N_7586);
nand U7621 (N_7621,N_7521,N_7536);
nor U7622 (N_7622,N_7598,N_7542);
nor U7623 (N_7623,N_7569,N_7506);
nor U7624 (N_7624,N_7562,N_7574);
nand U7625 (N_7625,N_7507,N_7589);
or U7626 (N_7626,N_7545,N_7502);
and U7627 (N_7627,N_7584,N_7573);
nor U7628 (N_7628,N_7547,N_7554);
and U7629 (N_7629,N_7550,N_7583);
nand U7630 (N_7630,N_7516,N_7590);
or U7631 (N_7631,N_7522,N_7596);
xnor U7632 (N_7632,N_7526,N_7512);
xor U7633 (N_7633,N_7560,N_7500);
nand U7634 (N_7634,N_7537,N_7563);
nor U7635 (N_7635,N_7572,N_7582);
nand U7636 (N_7636,N_7539,N_7552);
or U7637 (N_7637,N_7581,N_7511);
xor U7638 (N_7638,N_7543,N_7556);
or U7639 (N_7639,N_7519,N_7535);
xnor U7640 (N_7640,N_7531,N_7555);
nor U7641 (N_7641,N_7570,N_7585);
or U7642 (N_7642,N_7567,N_7559);
or U7643 (N_7643,N_7518,N_7558);
and U7644 (N_7644,N_7599,N_7528);
xnor U7645 (N_7645,N_7514,N_7538);
nand U7646 (N_7646,N_7549,N_7504);
or U7647 (N_7647,N_7588,N_7577);
nor U7648 (N_7648,N_7541,N_7510);
and U7649 (N_7649,N_7548,N_7508);
nor U7650 (N_7650,N_7533,N_7560);
nor U7651 (N_7651,N_7555,N_7595);
nand U7652 (N_7652,N_7576,N_7570);
or U7653 (N_7653,N_7568,N_7563);
nand U7654 (N_7654,N_7565,N_7521);
or U7655 (N_7655,N_7586,N_7519);
or U7656 (N_7656,N_7524,N_7510);
nor U7657 (N_7657,N_7592,N_7534);
and U7658 (N_7658,N_7531,N_7509);
nand U7659 (N_7659,N_7576,N_7531);
nand U7660 (N_7660,N_7522,N_7513);
and U7661 (N_7661,N_7562,N_7596);
nor U7662 (N_7662,N_7555,N_7511);
and U7663 (N_7663,N_7531,N_7522);
and U7664 (N_7664,N_7534,N_7582);
nor U7665 (N_7665,N_7577,N_7551);
or U7666 (N_7666,N_7555,N_7550);
nand U7667 (N_7667,N_7557,N_7553);
nor U7668 (N_7668,N_7597,N_7542);
nor U7669 (N_7669,N_7572,N_7528);
or U7670 (N_7670,N_7569,N_7576);
and U7671 (N_7671,N_7579,N_7569);
nand U7672 (N_7672,N_7559,N_7563);
or U7673 (N_7673,N_7539,N_7562);
or U7674 (N_7674,N_7510,N_7598);
xnor U7675 (N_7675,N_7553,N_7589);
nor U7676 (N_7676,N_7505,N_7557);
nand U7677 (N_7677,N_7585,N_7526);
or U7678 (N_7678,N_7530,N_7593);
nand U7679 (N_7679,N_7568,N_7507);
nand U7680 (N_7680,N_7595,N_7560);
nor U7681 (N_7681,N_7551,N_7501);
nor U7682 (N_7682,N_7549,N_7518);
nor U7683 (N_7683,N_7590,N_7542);
nand U7684 (N_7684,N_7578,N_7554);
or U7685 (N_7685,N_7578,N_7547);
xnor U7686 (N_7686,N_7535,N_7539);
or U7687 (N_7687,N_7511,N_7521);
nor U7688 (N_7688,N_7503,N_7567);
nand U7689 (N_7689,N_7536,N_7523);
and U7690 (N_7690,N_7582,N_7505);
nor U7691 (N_7691,N_7509,N_7516);
nor U7692 (N_7692,N_7526,N_7503);
nand U7693 (N_7693,N_7576,N_7581);
xnor U7694 (N_7694,N_7565,N_7542);
nor U7695 (N_7695,N_7575,N_7510);
or U7696 (N_7696,N_7553,N_7509);
and U7697 (N_7697,N_7558,N_7525);
or U7698 (N_7698,N_7586,N_7559);
nand U7699 (N_7699,N_7582,N_7526);
or U7700 (N_7700,N_7629,N_7652);
and U7701 (N_7701,N_7678,N_7686);
nor U7702 (N_7702,N_7653,N_7675);
nand U7703 (N_7703,N_7687,N_7627);
nand U7704 (N_7704,N_7626,N_7611);
and U7705 (N_7705,N_7669,N_7680);
or U7706 (N_7706,N_7688,N_7695);
nand U7707 (N_7707,N_7681,N_7600);
nor U7708 (N_7708,N_7633,N_7632);
or U7709 (N_7709,N_7685,N_7620);
xnor U7710 (N_7710,N_7651,N_7608);
and U7711 (N_7711,N_7658,N_7676);
nor U7712 (N_7712,N_7618,N_7637);
or U7713 (N_7713,N_7677,N_7689);
xor U7714 (N_7714,N_7671,N_7667);
xnor U7715 (N_7715,N_7660,N_7648);
nor U7716 (N_7716,N_7661,N_7684);
or U7717 (N_7717,N_7664,N_7673);
or U7718 (N_7718,N_7603,N_7672);
nor U7719 (N_7719,N_7692,N_7649);
or U7720 (N_7720,N_7612,N_7691);
or U7721 (N_7721,N_7614,N_7698);
and U7722 (N_7722,N_7696,N_7656);
nor U7723 (N_7723,N_7679,N_7639);
nor U7724 (N_7724,N_7615,N_7647);
nand U7725 (N_7725,N_7636,N_7662);
or U7726 (N_7726,N_7613,N_7619);
nor U7727 (N_7727,N_7694,N_7606);
and U7728 (N_7728,N_7674,N_7642);
or U7729 (N_7729,N_7690,N_7670);
or U7730 (N_7730,N_7641,N_7699);
and U7731 (N_7731,N_7638,N_7605);
nand U7732 (N_7732,N_7644,N_7655);
or U7733 (N_7733,N_7630,N_7624);
nor U7734 (N_7734,N_7610,N_7666);
and U7735 (N_7735,N_7622,N_7659);
nor U7736 (N_7736,N_7631,N_7634);
nand U7737 (N_7737,N_7682,N_7654);
xnor U7738 (N_7738,N_7668,N_7609);
or U7739 (N_7739,N_7665,N_7645);
and U7740 (N_7740,N_7693,N_7616);
or U7741 (N_7741,N_7601,N_7650);
or U7742 (N_7742,N_7663,N_7643);
and U7743 (N_7743,N_7635,N_7697);
and U7744 (N_7744,N_7646,N_7640);
nor U7745 (N_7745,N_7604,N_7683);
or U7746 (N_7746,N_7625,N_7617);
nand U7747 (N_7747,N_7623,N_7602);
or U7748 (N_7748,N_7607,N_7657);
nand U7749 (N_7749,N_7628,N_7621);
and U7750 (N_7750,N_7618,N_7694);
nor U7751 (N_7751,N_7657,N_7650);
nor U7752 (N_7752,N_7675,N_7684);
xnor U7753 (N_7753,N_7602,N_7656);
and U7754 (N_7754,N_7686,N_7615);
or U7755 (N_7755,N_7623,N_7665);
or U7756 (N_7756,N_7676,N_7637);
and U7757 (N_7757,N_7610,N_7660);
nand U7758 (N_7758,N_7687,N_7638);
or U7759 (N_7759,N_7686,N_7628);
and U7760 (N_7760,N_7637,N_7651);
and U7761 (N_7761,N_7677,N_7687);
nor U7762 (N_7762,N_7678,N_7604);
and U7763 (N_7763,N_7684,N_7613);
or U7764 (N_7764,N_7605,N_7602);
and U7765 (N_7765,N_7671,N_7691);
and U7766 (N_7766,N_7693,N_7688);
or U7767 (N_7767,N_7667,N_7608);
or U7768 (N_7768,N_7693,N_7603);
or U7769 (N_7769,N_7654,N_7611);
and U7770 (N_7770,N_7687,N_7610);
and U7771 (N_7771,N_7653,N_7657);
and U7772 (N_7772,N_7659,N_7697);
and U7773 (N_7773,N_7606,N_7643);
and U7774 (N_7774,N_7634,N_7607);
nor U7775 (N_7775,N_7634,N_7637);
nand U7776 (N_7776,N_7676,N_7669);
and U7777 (N_7777,N_7616,N_7607);
nor U7778 (N_7778,N_7612,N_7628);
and U7779 (N_7779,N_7673,N_7608);
xor U7780 (N_7780,N_7605,N_7612);
or U7781 (N_7781,N_7607,N_7677);
nor U7782 (N_7782,N_7603,N_7602);
nand U7783 (N_7783,N_7642,N_7652);
nor U7784 (N_7784,N_7697,N_7653);
or U7785 (N_7785,N_7647,N_7683);
nand U7786 (N_7786,N_7655,N_7686);
or U7787 (N_7787,N_7688,N_7630);
nor U7788 (N_7788,N_7619,N_7680);
and U7789 (N_7789,N_7669,N_7622);
nand U7790 (N_7790,N_7659,N_7615);
and U7791 (N_7791,N_7668,N_7697);
or U7792 (N_7792,N_7696,N_7688);
or U7793 (N_7793,N_7626,N_7662);
nor U7794 (N_7794,N_7670,N_7685);
or U7795 (N_7795,N_7659,N_7658);
nand U7796 (N_7796,N_7626,N_7644);
nand U7797 (N_7797,N_7638,N_7671);
or U7798 (N_7798,N_7640,N_7684);
nand U7799 (N_7799,N_7676,N_7660);
nand U7800 (N_7800,N_7784,N_7779);
nand U7801 (N_7801,N_7767,N_7797);
nor U7802 (N_7802,N_7703,N_7772);
nand U7803 (N_7803,N_7759,N_7775);
or U7804 (N_7804,N_7701,N_7726);
or U7805 (N_7805,N_7764,N_7776);
nand U7806 (N_7806,N_7798,N_7731);
and U7807 (N_7807,N_7755,N_7733);
and U7808 (N_7808,N_7774,N_7783);
and U7809 (N_7809,N_7751,N_7734);
nor U7810 (N_7810,N_7781,N_7787);
nand U7811 (N_7811,N_7782,N_7732);
nor U7812 (N_7812,N_7741,N_7702);
and U7813 (N_7813,N_7745,N_7752);
xor U7814 (N_7814,N_7716,N_7771);
and U7815 (N_7815,N_7765,N_7736);
xor U7816 (N_7816,N_7711,N_7746);
or U7817 (N_7817,N_7794,N_7737);
and U7818 (N_7818,N_7740,N_7770);
nand U7819 (N_7819,N_7721,N_7748);
nand U7820 (N_7820,N_7753,N_7743);
or U7821 (N_7821,N_7778,N_7724);
and U7822 (N_7822,N_7799,N_7704);
nor U7823 (N_7823,N_7756,N_7712);
or U7824 (N_7824,N_7728,N_7727);
and U7825 (N_7825,N_7713,N_7786);
and U7826 (N_7826,N_7738,N_7768);
and U7827 (N_7827,N_7762,N_7723);
nor U7828 (N_7828,N_7769,N_7700);
nor U7829 (N_7829,N_7777,N_7761);
nor U7830 (N_7830,N_7717,N_7715);
or U7831 (N_7831,N_7735,N_7730);
nand U7832 (N_7832,N_7742,N_7722);
or U7833 (N_7833,N_7719,N_7792);
nor U7834 (N_7834,N_7785,N_7754);
and U7835 (N_7835,N_7766,N_7706);
nor U7836 (N_7836,N_7791,N_7744);
xnor U7837 (N_7837,N_7710,N_7729);
nor U7838 (N_7838,N_7705,N_7747);
nand U7839 (N_7839,N_7714,N_7749);
and U7840 (N_7840,N_7709,N_7708);
nand U7841 (N_7841,N_7718,N_7720);
and U7842 (N_7842,N_7796,N_7757);
and U7843 (N_7843,N_7707,N_7750);
or U7844 (N_7844,N_7795,N_7758);
or U7845 (N_7845,N_7789,N_7790);
and U7846 (N_7846,N_7793,N_7773);
or U7847 (N_7847,N_7788,N_7739);
xnor U7848 (N_7848,N_7725,N_7780);
nand U7849 (N_7849,N_7760,N_7763);
and U7850 (N_7850,N_7719,N_7732);
nor U7851 (N_7851,N_7774,N_7789);
nor U7852 (N_7852,N_7799,N_7770);
xnor U7853 (N_7853,N_7732,N_7706);
nand U7854 (N_7854,N_7792,N_7736);
nor U7855 (N_7855,N_7756,N_7732);
nand U7856 (N_7856,N_7784,N_7797);
xor U7857 (N_7857,N_7721,N_7787);
nand U7858 (N_7858,N_7706,N_7755);
xnor U7859 (N_7859,N_7752,N_7738);
nand U7860 (N_7860,N_7711,N_7715);
xor U7861 (N_7861,N_7732,N_7742);
nand U7862 (N_7862,N_7755,N_7750);
nor U7863 (N_7863,N_7721,N_7799);
nand U7864 (N_7864,N_7710,N_7734);
or U7865 (N_7865,N_7713,N_7737);
and U7866 (N_7866,N_7776,N_7768);
nand U7867 (N_7867,N_7748,N_7762);
nand U7868 (N_7868,N_7763,N_7712);
nand U7869 (N_7869,N_7750,N_7731);
nand U7870 (N_7870,N_7769,N_7778);
xnor U7871 (N_7871,N_7700,N_7790);
or U7872 (N_7872,N_7764,N_7759);
or U7873 (N_7873,N_7783,N_7730);
and U7874 (N_7874,N_7702,N_7793);
and U7875 (N_7875,N_7732,N_7746);
nand U7876 (N_7876,N_7729,N_7728);
nand U7877 (N_7877,N_7761,N_7722);
and U7878 (N_7878,N_7730,N_7756);
and U7879 (N_7879,N_7706,N_7777);
nand U7880 (N_7880,N_7797,N_7759);
or U7881 (N_7881,N_7734,N_7754);
and U7882 (N_7882,N_7701,N_7748);
nor U7883 (N_7883,N_7714,N_7747);
nand U7884 (N_7884,N_7714,N_7756);
or U7885 (N_7885,N_7784,N_7770);
nor U7886 (N_7886,N_7730,N_7790);
nand U7887 (N_7887,N_7793,N_7763);
or U7888 (N_7888,N_7757,N_7732);
nand U7889 (N_7889,N_7716,N_7769);
or U7890 (N_7890,N_7716,N_7778);
nor U7891 (N_7891,N_7739,N_7718);
and U7892 (N_7892,N_7710,N_7763);
and U7893 (N_7893,N_7777,N_7790);
or U7894 (N_7894,N_7755,N_7754);
nor U7895 (N_7895,N_7769,N_7730);
nor U7896 (N_7896,N_7729,N_7765);
nand U7897 (N_7897,N_7771,N_7777);
and U7898 (N_7898,N_7752,N_7709);
nand U7899 (N_7899,N_7754,N_7726);
nand U7900 (N_7900,N_7876,N_7846);
and U7901 (N_7901,N_7843,N_7844);
or U7902 (N_7902,N_7802,N_7823);
nand U7903 (N_7903,N_7881,N_7812);
nor U7904 (N_7904,N_7815,N_7864);
and U7905 (N_7905,N_7871,N_7877);
nor U7906 (N_7906,N_7891,N_7879);
nand U7907 (N_7907,N_7810,N_7856);
or U7908 (N_7908,N_7837,N_7808);
nand U7909 (N_7909,N_7872,N_7890);
nor U7910 (N_7910,N_7829,N_7800);
nor U7911 (N_7911,N_7801,N_7826);
nor U7912 (N_7912,N_7878,N_7817);
nor U7913 (N_7913,N_7886,N_7888);
or U7914 (N_7914,N_7894,N_7805);
nor U7915 (N_7915,N_7813,N_7867);
nand U7916 (N_7916,N_7873,N_7820);
nor U7917 (N_7917,N_7852,N_7822);
and U7918 (N_7918,N_7818,N_7897);
nand U7919 (N_7919,N_7869,N_7845);
nand U7920 (N_7920,N_7865,N_7847);
or U7921 (N_7921,N_7803,N_7816);
or U7922 (N_7922,N_7870,N_7884);
xor U7923 (N_7923,N_7831,N_7828);
and U7924 (N_7924,N_7898,N_7889);
nand U7925 (N_7925,N_7866,N_7859);
or U7926 (N_7926,N_7861,N_7835);
xor U7927 (N_7927,N_7858,N_7830);
or U7928 (N_7928,N_7853,N_7807);
or U7929 (N_7929,N_7887,N_7860);
or U7930 (N_7930,N_7825,N_7868);
or U7931 (N_7931,N_7863,N_7842);
nor U7932 (N_7932,N_7814,N_7840);
or U7933 (N_7933,N_7841,N_7819);
and U7934 (N_7934,N_7833,N_7855);
or U7935 (N_7935,N_7821,N_7854);
or U7936 (N_7936,N_7896,N_7895);
nor U7937 (N_7937,N_7893,N_7804);
nand U7938 (N_7938,N_7809,N_7849);
nor U7939 (N_7939,N_7851,N_7850);
or U7940 (N_7940,N_7836,N_7857);
xor U7941 (N_7941,N_7824,N_7834);
or U7942 (N_7942,N_7848,N_7875);
xnor U7943 (N_7943,N_7806,N_7832);
xor U7944 (N_7944,N_7827,N_7880);
or U7945 (N_7945,N_7883,N_7885);
xor U7946 (N_7946,N_7899,N_7862);
nor U7947 (N_7947,N_7892,N_7838);
nand U7948 (N_7948,N_7874,N_7839);
nand U7949 (N_7949,N_7811,N_7882);
nor U7950 (N_7950,N_7845,N_7873);
or U7951 (N_7951,N_7841,N_7860);
or U7952 (N_7952,N_7835,N_7880);
or U7953 (N_7953,N_7858,N_7851);
nand U7954 (N_7954,N_7841,N_7863);
nor U7955 (N_7955,N_7803,N_7818);
nor U7956 (N_7956,N_7887,N_7846);
nand U7957 (N_7957,N_7865,N_7823);
nand U7958 (N_7958,N_7854,N_7807);
or U7959 (N_7959,N_7848,N_7857);
and U7960 (N_7960,N_7879,N_7805);
nor U7961 (N_7961,N_7887,N_7850);
nand U7962 (N_7962,N_7897,N_7816);
or U7963 (N_7963,N_7808,N_7877);
and U7964 (N_7964,N_7855,N_7844);
xnor U7965 (N_7965,N_7874,N_7848);
and U7966 (N_7966,N_7857,N_7899);
or U7967 (N_7967,N_7879,N_7846);
nor U7968 (N_7968,N_7897,N_7840);
and U7969 (N_7969,N_7819,N_7848);
or U7970 (N_7970,N_7820,N_7818);
or U7971 (N_7971,N_7879,N_7813);
nor U7972 (N_7972,N_7835,N_7850);
and U7973 (N_7973,N_7808,N_7803);
or U7974 (N_7974,N_7887,N_7854);
nor U7975 (N_7975,N_7859,N_7867);
nand U7976 (N_7976,N_7899,N_7822);
nor U7977 (N_7977,N_7880,N_7800);
or U7978 (N_7978,N_7814,N_7894);
nor U7979 (N_7979,N_7843,N_7835);
or U7980 (N_7980,N_7860,N_7875);
or U7981 (N_7981,N_7806,N_7853);
and U7982 (N_7982,N_7860,N_7840);
or U7983 (N_7983,N_7844,N_7828);
and U7984 (N_7984,N_7849,N_7839);
nand U7985 (N_7985,N_7837,N_7870);
or U7986 (N_7986,N_7814,N_7831);
nand U7987 (N_7987,N_7866,N_7824);
or U7988 (N_7988,N_7846,N_7800);
or U7989 (N_7989,N_7847,N_7884);
or U7990 (N_7990,N_7896,N_7866);
and U7991 (N_7991,N_7833,N_7893);
nand U7992 (N_7992,N_7814,N_7852);
nand U7993 (N_7993,N_7808,N_7871);
and U7994 (N_7994,N_7893,N_7844);
and U7995 (N_7995,N_7845,N_7846);
nand U7996 (N_7996,N_7823,N_7803);
nor U7997 (N_7997,N_7895,N_7822);
or U7998 (N_7998,N_7835,N_7858);
and U7999 (N_7999,N_7819,N_7887);
or U8000 (N_8000,N_7981,N_7972);
nand U8001 (N_8001,N_7997,N_7951);
nand U8002 (N_8002,N_7947,N_7928);
nand U8003 (N_8003,N_7989,N_7923);
xnor U8004 (N_8004,N_7960,N_7994);
or U8005 (N_8005,N_7967,N_7945);
nor U8006 (N_8006,N_7946,N_7992);
and U8007 (N_8007,N_7966,N_7958);
or U8008 (N_8008,N_7930,N_7927);
nor U8009 (N_8009,N_7907,N_7983);
nand U8010 (N_8010,N_7934,N_7933);
xor U8011 (N_8011,N_7948,N_7971);
and U8012 (N_8012,N_7993,N_7943);
nand U8013 (N_8013,N_7939,N_7908);
nand U8014 (N_8014,N_7999,N_7941);
nor U8015 (N_8015,N_7926,N_7902);
or U8016 (N_8016,N_7986,N_7932);
or U8017 (N_8017,N_7906,N_7952);
nor U8018 (N_8018,N_7919,N_7909);
and U8019 (N_8019,N_7970,N_7988);
or U8020 (N_8020,N_7904,N_7921);
nand U8021 (N_8021,N_7962,N_7977);
nor U8022 (N_8022,N_7931,N_7991);
nor U8023 (N_8023,N_7910,N_7990);
nor U8024 (N_8024,N_7979,N_7922);
xnor U8025 (N_8025,N_7918,N_7903);
or U8026 (N_8026,N_7995,N_7949);
or U8027 (N_8027,N_7950,N_7912);
or U8028 (N_8028,N_7937,N_7953);
nand U8029 (N_8029,N_7900,N_7956);
nand U8030 (N_8030,N_7929,N_7913);
nor U8031 (N_8031,N_7968,N_7969);
or U8032 (N_8032,N_7975,N_7961);
nand U8033 (N_8033,N_7917,N_7963);
and U8034 (N_8034,N_7978,N_7911);
nor U8035 (N_8035,N_7924,N_7935);
nor U8036 (N_8036,N_7936,N_7914);
nand U8037 (N_8037,N_7955,N_7985);
or U8038 (N_8038,N_7998,N_7974);
or U8039 (N_8039,N_7957,N_7944);
nor U8040 (N_8040,N_7940,N_7973);
nor U8041 (N_8041,N_7942,N_7954);
and U8042 (N_8042,N_7905,N_7901);
xnor U8043 (N_8043,N_7984,N_7925);
nor U8044 (N_8044,N_7996,N_7920);
nand U8045 (N_8045,N_7980,N_7916);
nand U8046 (N_8046,N_7987,N_7915);
or U8047 (N_8047,N_7938,N_7976);
or U8048 (N_8048,N_7964,N_7982);
nor U8049 (N_8049,N_7965,N_7959);
or U8050 (N_8050,N_7987,N_7921);
or U8051 (N_8051,N_7931,N_7922);
nand U8052 (N_8052,N_7991,N_7945);
xor U8053 (N_8053,N_7906,N_7922);
nor U8054 (N_8054,N_7936,N_7956);
and U8055 (N_8055,N_7951,N_7947);
nand U8056 (N_8056,N_7927,N_7911);
nor U8057 (N_8057,N_7941,N_7984);
xnor U8058 (N_8058,N_7928,N_7929);
or U8059 (N_8059,N_7956,N_7934);
or U8060 (N_8060,N_7933,N_7947);
and U8061 (N_8061,N_7945,N_7994);
and U8062 (N_8062,N_7965,N_7953);
xor U8063 (N_8063,N_7993,N_7969);
nor U8064 (N_8064,N_7941,N_7930);
xnor U8065 (N_8065,N_7949,N_7979);
nand U8066 (N_8066,N_7971,N_7932);
and U8067 (N_8067,N_7989,N_7942);
nand U8068 (N_8068,N_7964,N_7957);
or U8069 (N_8069,N_7967,N_7926);
nor U8070 (N_8070,N_7904,N_7963);
and U8071 (N_8071,N_7996,N_7936);
and U8072 (N_8072,N_7905,N_7916);
or U8073 (N_8073,N_7933,N_7937);
nand U8074 (N_8074,N_7941,N_7997);
nor U8075 (N_8075,N_7926,N_7993);
or U8076 (N_8076,N_7990,N_7982);
xnor U8077 (N_8077,N_7932,N_7942);
nor U8078 (N_8078,N_7956,N_7997);
xnor U8079 (N_8079,N_7980,N_7965);
and U8080 (N_8080,N_7911,N_7975);
nor U8081 (N_8081,N_7903,N_7978);
nor U8082 (N_8082,N_7996,N_7964);
or U8083 (N_8083,N_7984,N_7954);
nor U8084 (N_8084,N_7913,N_7910);
nor U8085 (N_8085,N_7957,N_7988);
or U8086 (N_8086,N_7983,N_7948);
or U8087 (N_8087,N_7910,N_7963);
nand U8088 (N_8088,N_7974,N_7947);
nand U8089 (N_8089,N_7977,N_7947);
and U8090 (N_8090,N_7984,N_7999);
nand U8091 (N_8091,N_7990,N_7986);
or U8092 (N_8092,N_7909,N_7913);
xnor U8093 (N_8093,N_7964,N_7969);
nand U8094 (N_8094,N_7965,N_7940);
and U8095 (N_8095,N_7988,N_7964);
or U8096 (N_8096,N_7913,N_7967);
xnor U8097 (N_8097,N_7925,N_7954);
nor U8098 (N_8098,N_7994,N_7921);
and U8099 (N_8099,N_7919,N_7983);
nand U8100 (N_8100,N_8026,N_8028);
or U8101 (N_8101,N_8078,N_8012);
nor U8102 (N_8102,N_8045,N_8080);
nor U8103 (N_8103,N_8004,N_8094);
xnor U8104 (N_8104,N_8092,N_8031);
nor U8105 (N_8105,N_8032,N_8091);
nand U8106 (N_8106,N_8006,N_8019);
xnor U8107 (N_8107,N_8054,N_8062);
nor U8108 (N_8108,N_8003,N_8014);
and U8109 (N_8109,N_8041,N_8095);
xor U8110 (N_8110,N_8077,N_8097);
nor U8111 (N_8111,N_8033,N_8061);
or U8112 (N_8112,N_8027,N_8064);
nand U8113 (N_8113,N_8052,N_8039);
nand U8114 (N_8114,N_8007,N_8058);
and U8115 (N_8115,N_8085,N_8036);
and U8116 (N_8116,N_8022,N_8086);
nand U8117 (N_8117,N_8021,N_8005);
and U8118 (N_8118,N_8008,N_8046);
nand U8119 (N_8119,N_8079,N_8020);
xor U8120 (N_8120,N_8082,N_8055);
and U8121 (N_8121,N_8044,N_8065);
and U8122 (N_8122,N_8000,N_8075);
nand U8123 (N_8123,N_8068,N_8048);
nor U8124 (N_8124,N_8024,N_8047);
and U8125 (N_8125,N_8018,N_8017);
nor U8126 (N_8126,N_8074,N_8090);
and U8127 (N_8127,N_8038,N_8050);
or U8128 (N_8128,N_8084,N_8037);
nor U8129 (N_8129,N_8099,N_8060);
and U8130 (N_8130,N_8069,N_8072);
or U8131 (N_8131,N_8043,N_8035);
and U8132 (N_8132,N_8087,N_8093);
and U8133 (N_8133,N_8034,N_8040);
or U8134 (N_8134,N_8063,N_8089);
and U8135 (N_8135,N_8076,N_8096);
or U8136 (N_8136,N_8067,N_8011);
and U8137 (N_8137,N_8053,N_8098);
nand U8138 (N_8138,N_8010,N_8066);
and U8139 (N_8139,N_8001,N_8051);
and U8140 (N_8140,N_8083,N_8025);
xor U8141 (N_8141,N_8059,N_8049);
nor U8142 (N_8142,N_8023,N_8042);
and U8143 (N_8143,N_8081,N_8071);
and U8144 (N_8144,N_8013,N_8070);
or U8145 (N_8145,N_8002,N_8073);
nand U8146 (N_8146,N_8088,N_8016);
nor U8147 (N_8147,N_8056,N_8009);
and U8148 (N_8148,N_8030,N_8029);
nand U8149 (N_8149,N_8015,N_8057);
nor U8150 (N_8150,N_8054,N_8097);
nand U8151 (N_8151,N_8084,N_8043);
or U8152 (N_8152,N_8063,N_8033);
nand U8153 (N_8153,N_8036,N_8081);
or U8154 (N_8154,N_8017,N_8064);
and U8155 (N_8155,N_8009,N_8014);
nor U8156 (N_8156,N_8025,N_8044);
or U8157 (N_8157,N_8062,N_8045);
or U8158 (N_8158,N_8091,N_8059);
nor U8159 (N_8159,N_8010,N_8017);
or U8160 (N_8160,N_8057,N_8034);
or U8161 (N_8161,N_8077,N_8029);
and U8162 (N_8162,N_8006,N_8093);
nor U8163 (N_8163,N_8034,N_8065);
xnor U8164 (N_8164,N_8081,N_8010);
nor U8165 (N_8165,N_8043,N_8081);
nor U8166 (N_8166,N_8007,N_8063);
and U8167 (N_8167,N_8079,N_8004);
and U8168 (N_8168,N_8070,N_8008);
and U8169 (N_8169,N_8019,N_8032);
nand U8170 (N_8170,N_8081,N_8079);
xor U8171 (N_8171,N_8061,N_8088);
nand U8172 (N_8172,N_8077,N_8047);
or U8173 (N_8173,N_8044,N_8050);
or U8174 (N_8174,N_8006,N_8076);
nand U8175 (N_8175,N_8092,N_8078);
and U8176 (N_8176,N_8038,N_8082);
nand U8177 (N_8177,N_8023,N_8049);
nor U8178 (N_8178,N_8039,N_8056);
or U8179 (N_8179,N_8004,N_8029);
nor U8180 (N_8180,N_8059,N_8054);
nor U8181 (N_8181,N_8036,N_8005);
or U8182 (N_8182,N_8085,N_8093);
or U8183 (N_8183,N_8037,N_8009);
xor U8184 (N_8184,N_8047,N_8025);
nand U8185 (N_8185,N_8091,N_8090);
nor U8186 (N_8186,N_8080,N_8041);
nand U8187 (N_8187,N_8014,N_8015);
nor U8188 (N_8188,N_8018,N_8026);
xor U8189 (N_8189,N_8040,N_8064);
nor U8190 (N_8190,N_8044,N_8023);
nand U8191 (N_8191,N_8008,N_8037);
nor U8192 (N_8192,N_8002,N_8064);
nor U8193 (N_8193,N_8066,N_8080);
or U8194 (N_8194,N_8006,N_8042);
and U8195 (N_8195,N_8052,N_8091);
nand U8196 (N_8196,N_8026,N_8074);
and U8197 (N_8197,N_8052,N_8016);
nor U8198 (N_8198,N_8098,N_8036);
or U8199 (N_8199,N_8047,N_8076);
nand U8200 (N_8200,N_8185,N_8129);
and U8201 (N_8201,N_8158,N_8137);
and U8202 (N_8202,N_8162,N_8155);
or U8203 (N_8203,N_8103,N_8146);
or U8204 (N_8204,N_8134,N_8163);
and U8205 (N_8205,N_8194,N_8177);
and U8206 (N_8206,N_8165,N_8161);
and U8207 (N_8207,N_8191,N_8190);
and U8208 (N_8208,N_8151,N_8169);
or U8209 (N_8209,N_8143,N_8189);
or U8210 (N_8210,N_8152,N_8187);
and U8211 (N_8211,N_8118,N_8116);
and U8212 (N_8212,N_8193,N_8131);
or U8213 (N_8213,N_8106,N_8184);
or U8214 (N_8214,N_8173,N_8154);
and U8215 (N_8215,N_8156,N_8178);
nand U8216 (N_8216,N_8168,N_8139);
xor U8217 (N_8217,N_8108,N_8144);
and U8218 (N_8218,N_8142,N_8113);
xnor U8219 (N_8219,N_8104,N_8145);
and U8220 (N_8220,N_8140,N_8181);
xor U8221 (N_8221,N_8186,N_8171);
and U8222 (N_8222,N_8105,N_8141);
nand U8223 (N_8223,N_8115,N_8121);
xnor U8224 (N_8224,N_8195,N_8174);
and U8225 (N_8225,N_8182,N_8107);
nor U8226 (N_8226,N_8160,N_8188);
nand U8227 (N_8227,N_8147,N_8175);
or U8228 (N_8228,N_8180,N_8148);
nand U8229 (N_8229,N_8179,N_8135);
nor U8230 (N_8230,N_8157,N_8159);
nand U8231 (N_8231,N_8149,N_8122);
nor U8232 (N_8232,N_8176,N_8123);
nor U8233 (N_8233,N_8153,N_8124);
nand U8234 (N_8234,N_8119,N_8138);
and U8235 (N_8235,N_8167,N_8198);
nand U8236 (N_8236,N_8133,N_8132);
xor U8237 (N_8237,N_8127,N_8128);
nand U8238 (N_8238,N_8164,N_8109);
nand U8239 (N_8239,N_8120,N_8172);
nand U8240 (N_8240,N_8125,N_8126);
and U8241 (N_8241,N_8111,N_8199);
and U8242 (N_8242,N_8170,N_8110);
xor U8243 (N_8243,N_8100,N_8166);
nand U8244 (N_8244,N_8196,N_8183);
and U8245 (N_8245,N_8192,N_8136);
nand U8246 (N_8246,N_8117,N_8130);
or U8247 (N_8247,N_8101,N_8102);
nand U8248 (N_8248,N_8114,N_8150);
nand U8249 (N_8249,N_8112,N_8197);
nor U8250 (N_8250,N_8142,N_8103);
nor U8251 (N_8251,N_8142,N_8121);
or U8252 (N_8252,N_8136,N_8195);
nand U8253 (N_8253,N_8107,N_8101);
and U8254 (N_8254,N_8115,N_8170);
and U8255 (N_8255,N_8154,N_8158);
nand U8256 (N_8256,N_8152,N_8151);
and U8257 (N_8257,N_8109,N_8157);
and U8258 (N_8258,N_8111,N_8150);
or U8259 (N_8259,N_8155,N_8102);
nand U8260 (N_8260,N_8177,N_8169);
xnor U8261 (N_8261,N_8105,N_8149);
and U8262 (N_8262,N_8122,N_8124);
or U8263 (N_8263,N_8184,N_8170);
nor U8264 (N_8264,N_8113,N_8183);
nand U8265 (N_8265,N_8156,N_8150);
or U8266 (N_8266,N_8172,N_8152);
or U8267 (N_8267,N_8120,N_8176);
and U8268 (N_8268,N_8198,N_8136);
nand U8269 (N_8269,N_8112,N_8114);
and U8270 (N_8270,N_8152,N_8145);
nor U8271 (N_8271,N_8152,N_8133);
or U8272 (N_8272,N_8157,N_8156);
nand U8273 (N_8273,N_8101,N_8119);
or U8274 (N_8274,N_8199,N_8185);
or U8275 (N_8275,N_8137,N_8157);
or U8276 (N_8276,N_8172,N_8122);
nor U8277 (N_8277,N_8147,N_8139);
nor U8278 (N_8278,N_8151,N_8157);
xnor U8279 (N_8279,N_8156,N_8169);
or U8280 (N_8280,N_8175,N_8148);
or U8281 (N_8281,N_8101,N_8193);
and U8282 (N_8282,N_8192,N_8197);
nand U8283 (N_8283,N_8132,N_8178);
nand U8284 (N_8284,N_8193,N_8106);
nor U8285 (N_8285,N_8118,N_8164);
or U8286 (N_8286,N_8183,N_8126);
and U8287 (N_8287,N_8120,N_8113);
nor U8288 (N_8288,N_8179,N_8162);
nand U8289 (N_8289,N_8146,N_8129);
nand U8290 (N_8290,N_8189,N_8183);
or U8291 (N_8291,N_8162,N_8127);
or U8292 (N_8292,N_8195,N_8149);
nand U8293 (N_8293,N_8115,N_8145);
nor U8294 (N_8294,N_8110,N_8197);
and U8295 (N_8295,N_8150,N_8119);
nor U8296 (N_8296,N_8128,N_8180);
or U8297 (N_8297,N_8127,N_8151);
or U8298 (N_8298,N_8126,N_8113);
nor U8299 (N_8299,N_8139,N_8141);
nor U8300 (N_8300,N_8236,N_8202);
nand U8301 (N_8301,N_8295,N_8273);
nand U8302 (N_8302,N_8209,N_8267);
nand U8303 (N_8303,N_8220,N_8213);
xnor U8304 (N_8304,N_8247,N_8203);
or U8305 (N_8305,N_8227,N_8243);
nor U8306 (N_8306,N_8255,N_8268);
xnor U8307 (N_8307,N_8285,N_8206);
or U8308 (N_8308,N_8208,N_8201);
or U8309 (N_8309,N_8290,N_8216);
and U8310 (N_8310,N_8292,N_8274);
and U8311 (N_8311,N_8284,N_8293);
nand U8312 (N_8312,N_8269,N_8204);
or U8313 (N_8313,N_8210,N_8259);
nor U8314 (N_8314,N_8280,N_8254);
and U8315 (N_8315,N_8270,N_8249);
and U8316 (N_8316,N_8257,N_8215);
xnor U8317 (N_8317,N_8218,N_8224);
and U8318 (N_8318,N_8261,N_8244);
xnor U8319 (N_8319,N_8294,N_8266);
and U8320 (N_8320,N_8238,N_8252);
nand U8321 (N_8321,N_8233,N_8297);
and U8322 (N_8322,N_8291,N_8228);
xor U8323 (N_8323,N_8296,N_8214);
and U8324 (N_8324,N_8223,N_8289);
nand U8325 (N_8325,N_8253,N_8240);
nand U8326 (N_8326,N_8225,N_8200);
nor U8327 (N_8327,N_8278,N_8248);
or U8328 (N_8328,N_8205,N_8246);
nor U8329 (N_8329,N_8229,N_8272);
or U8330 (N_8330,N_8242,N_8281);
and U8331 (N_8331,N_8279,N_8282);
nor U8332 (N_8332,N_8221,N_8212);
or U8333 (N_8333,N_8230,N_8241);
nand U8334 (N_8334,N_8231,N_8264);
or U8335 (N_8335,N_8262,N_8276);
nor U8336 (N_8336,N_8234,N_8211);
and U8337 (N_8337,N_8222,N_8288);
nor U8338 (N_8338,N_8235,N_8271);
and U8339 (N_8339,N_8239,N_8250);
and U8340 (N_8340,N_8283,N_8275);
and U8341 (N_8341,N_8287,N_8277);
and U8342 (N_8342,N_8219,N_8217);
nand U8343 (N_8343,N_8263,N_8299);
or U8344 (N_8344,N_8207,N_8265);
xnor U8345 (N_8345,N_8298,N_8260);
nand U8346 (N_8346,N_8237,N_8232);
and U8347 (N_8347,N_8286,N_8251);
xnor U8348 (N_8348,N_8256,N_8258);
and U8349 (N_8349,N_8226,N_8245);
or U8350 (N_8350,N_8242,N_8271);
and U8351 (N_8351,N_8218,N_8242);
and U8352 (N_8352,N_8299,N_8283);
nand U8353 (N_8353,N_8233,N_8250);
nand U8354 (N_8354,N_8286,N_8226);
or U8355 (N_8355,N_8220,N_8266);
nand U8356 (N_8356,N_8252,N_8214);
nor U8357 (N_8357,N_8209,N_8235);
nand U8358 (N_8358,N_8293,N_8276);
xor U8359 (N_8359,N_8297,N_8252);
and U8360 (N_8360,N_8205,N_8265);
nand U8361 (N_8361,N_8204,N_8257);
nand U8362 (N_8362,N_8219,N_8276);
or U8363 (N_8363,N_8233,N_8276);
nand U8364 (N_8364,N_8241,N_8286);
nand U8365 (N_8365,N_8257,N_8266);
and U8366 (N_8366,N_8227,N_8255);
nor U8367 (N_8367,N_8213,N_8215);
and U8368 (N_8368,N_8218,N_8281);
nand U8369 (N_8369,N_8209,N_8254);
or U8370 (N_8370,N_8279,N_8247);
nor U8371 (N_8371,N_8264,N_8232);
or U8372 (N_8372,N_8221,N_8224);
and U8373 (N_8373,N_8280,N_8252);
nand U8374 (N_8374,N_8264,N_8240);
nand U8375 (N_8375,N_8270,N_8219);
nor U8376 (N_8376,N_8248,N_8204);
nor U8377 (N_8377,N_8254,N_8205);
or U8378 (N_8378,N_8233,N_8205);
nand U8379 (N_8379,N_8211,N_8223);
nor U8380 (N_8380,N_8217,N_8259);
or U8381 (N_8381,N_8203,N_8211);
or U8382 (N_8382,N_8265,N_8217);
xor U8383 (N_8383,N_8228,N_8242);
and U8384 (N_8384,N_8262,N_8209);
nor U8385 (N_8385,N_8224,N_8296);
or U8386 (N_8386,N_8249,N_8286);
nand U8387 (N_8387,N_8241,N_8204);
or U8388 (N_8388,N_8273,N_8258);
or U8389 (N_8389,N_8283,N_8217);
nand U8390 (N_8390,N_8291,N_8289);
and U8391 (N_8391,N_8225,N_8260);
nor U8392 (N_8392,N_8259,N_8256);
xnor U8393 (N_8393,N_8231,N_8236);
and U8394 (N_8394,N_8228,N_8276);
and U8395 (N_8395,N_8210,N_8217);
or U8396 (N_8396,N_8203,N_8249);
xor U8397 (N_8397,N_8265,N_8240);
and U8398 (N_8398,N_8212,N_8228);
or U8399 (N_8399,N_8204,N_8215);
xor U8400 (N_8400,N_8397,N_8373);
nor U8401 (N_8401,N_8393,N_8352);
and U8402 (N_8402,N_8376,N_8379);
nand U8403 (N_8403,N_8313,N_8395);
and U8404 (N_8404,N_8381,N_8331);
nor U8405 (N_8405,N_8339,N_8324);
or U8406 (N_8406,N_8380,N_8326);
nor U8407 (N_8407,N_8348,N_8332);
and U8408 (N_8408,N_8355,N_8362);
and U8409 (N_8409,N_8300,N_8378);
or U8410 (N_8410,N_8368,N_8347);
or U8411 (N_8411,N_8342,N_8308);
nand U8412 (N_8412,N_8346,N_8318);
or U8413 (N_8413,N_8398,N_8323);
and U8414 (N_8414,N_8343,N_8329);
nand U8415 (N_8415,N_8314,N_8330);
and U8416 (N_8416,N_8333,N_8336);
and U8417 (N_8417,N_8304,N_8351);
and U8418 (N_8418,N_8307,N_8325);
nand U8419 (N_8419,N_8345,N_8302);
or U8420 (N_8420,N_8361,N_8370);
nand U8421 (N_8421,N_8360,N_8310);
or U8422 (N_8422,N_8383,N_8350);
nand U8423 (N_8423,N_8389,N_8388);
and U8424 (N_8424,N_8334,N_8306);
or U8425 (N_8425,N_8364,N_8319);
nor U8426 (N_8426,N_8356,N_8385);
and U8427 (N_8427,N_8374,N_8322);
and U8428 (N_8428,N_8303,N_8320);
and U8429 (N_8429,N_8392,N_8354);
nand U8430 (N_8430,N_8312,N_8371);
or U8431 (N_8431,N_8317,N_8321);
nand U8432 (N_8432,N_8344,N_8399);
and U8433 (N_8433,N_8340,N_8372);
or U8434 (N_8434,N_8386,N_8301);
nand U8435 (N_8435,N_8341,N_8309);
or U8436 (N_8436,N_8363,N_8394);
nor U8437 (N_8437,N_8338,N_8382);
nand U8438 (N_8438,N_8377,N_8366);
nand U8439 (N_8439,N_8375,N_8311);
and U8440 (N_8440,N_8390,N_8391);
and U8441 (N_8441,N_8387,N_8369);
nor U8442 (N_8442,N_8316,N_8349);
and U8443 (N_8443,N_8335,N_8327);
or U8444 (N_8444,N_8337,N_8315);
or U8445 (N_8445,N_8365,N_8384);
or U8446 (N_8446,N_8396,N_8359);
or U8447 (N_8447,N_8328,N_8305);
nand U8448 (N_8448,N_8353,N_8358);
or U8449 (N_8449,N_8357,N_8367);
or U8450 (N_8450,N_8399,N_8308);
nor U8451 (N_8451,N_8393,N_8385);
or U8452 (N_8452,N_8315,N_8330);
or U8453 (N_8453,N_8387,N_8324);
and U8454 (N_8454,N_8328,N_8307);
and U8455 (N_8455,N_8315,N_8355);
and U8456 (N_8456,N_8382,N_8313);
or U8457 (N_8457,N_8309,N_8336);
and U8458 (N_8458,N_8383,N_8330);
and U8459 (N_8459,N_8395,N_8360);
and U8460 (N_8460,N_8318,N_8375);
xor U8461 (N_8461,N_8393,N_8307);
nand U8462 (N_8462,N_8389,N_8321);
nand U8463 (N_8463,N_8323,N_8327);
and U8464 (N_8464,N_8389,N_8304);
and U8465 (N_8465,N_8319,N_8393);
or U8466 (N_8466,N_8329,N_8384);
and U8467 (N_8467,N_8354,N_8382);
nor U8468 (N_8468,N_8325,N_8392);
or U8469 (N_8469,N_8351,N_8318);
and U8470 (N_8470,N_8395,N_8317);
or U8471 (N_8471,N_8328,N_8334);
and U8472 (N_8472,N_8369,N_8364);
and U8473 (N_8473,N_8320,N_8326);
and U8474 (N_8474,N_8324,N_8398);
nor U8475 (N_8475,N_8369,N_8391);
nand U8476 (N_8476,N_8349,N_8338);
or U8477 (N_8477,N_8384,N_8322);
nand U8478 (N_8478,N_8382,N_8309);
xor U8479 (N_8479,N_8351,N_8361);
and U8480 (N_8480,N_8301,N_8373);
nor U8481 (N_8481,N_8312,N_8322);
nand U8482 (N_8482,N_8367,N_8326);
nor U8483 (N_8483,N_8326,N_8357);
and U8484 (N_8484,N_8396,N_8336);
and U8485 (N_8485,N_8344,N_8302);
nand U8486 (N_8486,N_8332,N_8376);
nand U8487 (N_8487,N_8378,N_8316);
nor U8488 (N_8488,N_8356,N_8397);
and U8489 (N_8489,N_8355,N_8323);
or U8490 (N_8490,N_8381,N_8305);
xnor U8491 (N_8491,N_8315,N_8332);
nand U8492 (N_8492,N_8327,N_8379);
nand U8493 (N_8493,N_8378,N_8344);
or U8494 (N_8494,N_8316,N_8301);
and U8495 (N_8495,N_8374,N_8334);
and U8496 (N_8496,N_8391,N_8374);
and U8497 (N_8497,N_8369,N_8388);
and U8498 (N_8498,N_8317,N_8328);
xor U8499 (N_8499,N_8308,N_8366);
nand U8500 (N_8500,N_8451,N_8436);
xor U8501 (N_8501,N_8431,N_8432);
nand U8502 (N_8502,N_8434,N_8468);
and U8503 (N_8503,N_8499,N_8408);
nand U8504 (N_8504,N_8448,N_8493);
nand U8505 (N_8505,N_8421,N_8464);
nand U8506 (N_8506,N_8424,N_8495);
and U8507 (N_8507,N_8400,N_8443);
nor U8508 (N_8508,N_8480,N_8459);
or U8509 (N_8509,N_8469,N_8465);
nand U8510 (N_8510,N_8497,N_8454);
nor U8511 (N_8511,N_8490,N_8456);
xor U8512 (N_8512,N_8494,N_8478);
nor U8513 (N_8513,N_8471,N_8415);
nor U8514 (N_8514,N_8492,N_8470);
and U8515 (N_8515,N_8477,N_8439);
or U8516 (N_8516,N_8461,N_8472);
nor U8517 (N_8517,N_8476,N_8473);
nand U8518 (N_8518,N_8407,N_8425);
nand U8519 (N_8519,N_8403,N_8466);
nor U8520 (N_8520,N_8402,N_8442);
nor U8521 (N_8521,N_8449,N_8487);
nor U8522 (N_8522,N_8405,N_8410);
nor U8523 (N_8523,N_8441,N_8450);
and U8524 (N_8524,N_8475,N_8452);
and U8525 (N_8525,N_8462,N_8457);
and U8526 (N_8526,N_8467,N_8489);
xor U8527 (N_8527,N_8453,N_8438);
nand U8528 (N_8528,N_8430,N_8481);
nand U8529 (N_8529,N_8435,N_8416);
or U8530 (N_8530,N_8447,N_8433);
xnor U8531 (N_8531,N_8455,N_8491);
or U8532 (N_8532,N_8412,N_8404);
xor U8533 (N_8533,N_8460,N_8426);
nand U8534 (N_8534,N_8401,N_8428);
or U8535 (N_8535,N_8446,N_8419);
or U8536 (N_8536,N_8429,N_8422);
and U8537 (N_8537,N_8485,N_8458);
nand U8538 (N_8538,N_8418,N_8486);
nand U8539 (N_8539,N_8479,N_8444);
nand U8540 (N_8540,N_8427,N_8420);
and U8541 (N_8541,N_8445,N_8406);
nor U8542 (N_8542,N_8409,N_8484);
nor U8543 (N_8543,N_8414,N_8496);
xnor U8544 (N_8544,N_8413,N_8411);
nand U8545 (N_8545,N_8488,N_8463);
xnor U8546 (N_8546,N_8474,N_8437);
and U8547 (N_8547,N_8417,N_8483);
or U8548 (N_8548,N_8482,N_8423);
or U8549 (N_8549,N_8498,N_8440);
nand U8550 (N_8550,N_8409,N_8455);
or U8551 (N_8551,N_8424,N_8430);
and U8552 (N_8552,N_8414,N_8453);
and U8553 (N_8553,N_8401,N_8482);
xor U8554 (N_8554,N_8429,N_8481);
nor U8555 (N_8555,N_8419,N_8472);
or U8556 (N_8556,N_8426,N_8445);
or U8557 (N_8557,N_8415,N_8439);
nor U8558 (N_8558,N_8484,N_8411);
xnor U8559 (N_8559,N_8483,N_8412);
xor U8560 (N_8560,N_8453,N_8464);
xnor U8561 (N_8561,N_8439,N_8451);
and U8562 (N_8562,N_8451,N_8429);
nand U8563 (N_8563,N_8499,N_8452);
or U8564 (N_8564,N_8468,N_8473);
nand U8565 (N_8565,N_8462,N_8492);
nand U8566 (N_8566,N_8429,N_8456);
and U8567 (N_8567,N_8491,N_8411);
and U8568 (N_8568,N_8455,N_8419);
nand U8569 (N_8569,N_8468,N_8443);
nand U8570 (N_8570,N_8473,N_8448);
nand U8571 (N_8571,N_8442,N_8496);
nand U8572 (N_8572,N_8495,N_8452);
and U8573 (N_8573,N_8457,N_8477);
and U8574 (N_8574,N_8440,N_8401);
nand U8575 (N_8575,N_8442,N_8439);
nor U8576 (N_8576,N_8460,N_8440);
and U8577 (N_8577,N_8414,N_8450);
and U8578 (N_8578,N_8452,N_8403);
or U8579 (N_8579,N_8456,N_8414);
nor U8580 (N_8580,N_8446,N_8491);
and U8581 (N_8581,N_8448,N_8433);
or U8582 (N_8582,N_8456,N_8461);
nor U8583 (N_8583,N_8497,N_8444);
and U8584 (N_8584,N_8418,N_8458);
and U8585 (N_8585,N_8461,N_8469);
and U8586 (N_8586,N_8412,N_8488);
nor U8587 (N_8587,N_8457,N_8424);
nand U8588 (N_8588,N_8401,N_8467);
xor U8589 (N_8589,N_8421,N_8445);
or U8590 (N_8590,N_8432,N_8481);
nor U8591 (N_8591,N_8459,N_8406);
nor U8592 (N_8592,N_8489,N_8448);
or U8593 (N_8593,N_8482,N_8408);
or U8594 (N_8594,N_8432,N_8416);
nand U8595 (N_8595,N_8458,N_8421);
nor U8596 (N_8596,N_8438,N_8476);
nand U8597 (N_8597,N_8457,N_8439);
and U8598 (N_8598,N_8484,N_8474);
xnor U8599 (N_8599,N_8431,N_8409);
nand U8600 (N_8600,N_8555,N_8574);
and U8601 (N_8601,N_8589,N_8587);
or U8602 (N_8602,N_8529,N_8536);
nor U8603 (N_8603,N_8558,N_8508);
or U8604 (N_8604,N_8581,N_8583);
or U8605 (N_8605,N_8577,N_8531);
nand U8606 (N_8606,N_8526,N_8505);
nand U8607 (N_8607,N_8596,N_8593);
or U8608 (N_8608,N_8534,N_8569);
nand U8609 (N_8609,N_8562,N_8538);
nand U8610 (N_8610,N_8549,N_8530);
nor U8611 (N_8611,N_8580,N_8500);
xnor U8612 (N_8612,N_8563,N_8588);
and U8613 (N_8613,N_8503,N_8546);
nand U8614 (N_8614,N_8515,N_8502);
or U8615 (N_8615,N_8584,N_8533);
or U8616 (N_8616,N_8553,N_8599);
nand U8617 (N_8617,N_8592,N_8551);
and U8618 (N_8618,N_8597,N_8572);
and U8619 (N_8619,N_8528,N_8579);
or U8620 (N_8620,N_8594,N_8509);
or U8621 (N_8621,N_8511,N_8578);
xnor U8622 (N_8622,N_8554,N_8552);
nor U8623 (N_8623,N_8566,N_8527);
nor U8624 (N_8624,N_8541,N_8506);
xnor U8625 (N_8625,N_8573,N_8514);
or U8626 (N_8626,N_8586,N_8564);
nor U8627 (N_8627,N_8550,N_8595);
and U8628 (N_8628,N_8510,N_8517);
and U8629 (N_8629,N_8537,N_8560);
or U8630 (N_8630,N_8525,N_8561);
and U8631 (N_8631,N_8504,N_8585);
nand U8632 (N_8632,N_8575,N_8556);
and U8633 (N_8633,N_8568,N_8559);
and U8634 (N_8634,N_8512,N_8576);
nand U8635 (N_8635,N_8571,N_8591);
or U8636 (N_8636,N_8522,N_8520);
or U8637 (N_8637,N_8501,N_8535);
or U8638 (N_8638,N_8513,N_8565);
or U8639 (N_8639,N_8516,N_8557);
or U8640 (N_8640,N_8547,N_8582);
nand U8641 (N_8641,N_8521,N_8544);
nor U8642 (N_8642,N_8524,N_8543);
and U8643 (N_8643,N_8532,N_8523);
and U8644 (N_8644,N_8567,N_8545);
and U8645 (N_8645,N_8548,N_8540);
and U8646 (N_8646,N_8598,N_8507);
nor U8647 (N_8647,N_8539,N_8590);
and U8648 (N_8648,N_8542,N_8519);
and U8649 (N_8649,N_8518,N_8570);
or U8650 (N_8650,N_8534,N_8525);
or U8651 (N_8651,N_8551,N_8587);
or U8652 (N_8652,N_8505,N_8582);
nand U8653 (N_8653,N_8523,N_8565);
or U8654 (N_8654,N_8512,N_8567);
xor U8655 (N_8655,N_8548,N_8509);
nor U8656 (N_8656,N_8543,N_8538);
nand U8657 (N_8657,N_8578,N_8524);
or U8658 (N_8658,N_8510,N_8560);
xor U8659 (N_8659,N_8500,N_8592);
and U8660 (N_8660,N_8517,N_8593);
nand U8661 (N_8661,N_8514,N_8588);
xor U8662 (N_8662,N_8548,N_8598);
nor U8663 (N_8663,N_8525,N_8540);
nor U8664 (N_8664,N_8500,N_8574);
xor U8665 (N_8665,N_8527,N_8567);
nor U8666 (N_8666,N_8594,N_8598);
and U8667 (N_8667,N_8530,N_8504);
and U8668 (N_8668,N_8501,N_8599);
and U8669 (N_8669,N_8582,N_8567);
or U8670 (N_8670,N_8588,N_8500);
nor U8671 (N_8671,N_8587,N_8502);
nand U8672 (N_8672,N_8511,N_8554);
nor U8673 (N_8673,N_8558,N_8577);
nand U8674 (N_8674,N_8540,N_8510);
nand U8675 (N_8675,N_8597,N_8509);
and U8676 (N_8676,N_8552,N_8519);
or U8677 (N_8677,N_8570,N_8526);
or U8678 (N_8678,N_8564,N_8505);
or U8679 (N_8679,N_8569,N_8570);
and U8680 (N_8680,N_8585,N_8528);
nor U8681 (N_8681,N_8560,N_8569);
and U8682 (N_8682,N_8542,N_8553);
or U8683 (N_8683,N_8528,N_8595);
nand U8684 (N_8684,N_8569,N_8573);
and U8685 (N_8685,N_8529,N_8504);
and U8686 (N_8686,N_8583,N_8506);
and U8687 (N_8687,N_8511,N_8516);
nand U8688 (N_8688,N_8542,N_8550);
nand U8689 (N_8689,N_8585,N_8546);
and U8690 (N_8690,N_8516,N_8582);
and U8691 (N_8691,N_8589,N_8586);
or U8692 (N_8692,N_8538,N_8589);
or U8693 (N_8693,N_8540,N_8574);
or U8694 (N_8694,N_8514,N_8541);
nand U8695 (N_8695,N_8504,N_8573);
xnor U8696 (N_8696,N_8596,N_8590);
nand U8697 (N_8697,N_8516,N_8589);
and U8698 (N_8698,N_8552,N_8531);
or U8699 (N_8699,N_8542,N_8566);
xor U8700 (N_8700,N_8661,N_8628);
and U8701 (N_8701,N_8671,N_8674);
nor U8702 (N_8702,N_8603,N_8647);
xnor U8703 (N_8703,N_8651,N_8624);
and U8704 (N_8704,N_8660,N_8635);
nor U8705 (N_8705,N_8664,N_8666);
xnor U8706 (N_8706,N_8652,N_8680);
nor U8707 (N_8707,N_8699,N_8618);
or U8708 (N_8708,N_8644,N_8695);
or U8709 (N_8709,N_8645,N_8639);
and U8710 (N_8710,N_8646,N_8689);
xor U8711 (N_8711,N_8662,N_8614);
and U8712 (N_8712,N_8625,N_8610);
and U8713 (N_8713,N_8611,N_8678);
and U8714 (N_8714,N_8672,N_8691);
and U8715 (N_8715,N_8600,N_8658);
and U8716 (N_8716,N_8620,N_8637);
xor U8717 (N_8717,N_8632,N_8668);
and U8718 (N_8718,N_8609,N_8675);
or U8719 (N_8719,N_8636,N_8643);
and U8720 (N_8720,N_8601,N_8605);
nand U8721 (N_8721,N_8682,N_8638);
nand U8722 (N_8722,N_8627,N_8655);
nor U8723 (N_8723,N_8612,N_8667);
xor U8724 (N_8724,N_8608,N_8654);
nand U8725 (N_8725,N_8626,N_8623);
nand U8726 (N_8726,N_8656,N_8673);
or U8727 (N_8727,N_8683,N_8653);
or U8728 (N_8728,N_8615,N_8665);
nand U8729 (N_8729,N_8686,N_8613);
nor U8730 (N_8730,N_8684,N_8621);
or U8731 (N_8731,N_8687,N_8663);
nand U8732 (N_8732,N_8634,N_8607);
and U8733 (N_8733,N_8630,N_8685);
xnor U8734 (N_8734,N_8648,N_8604);
and U8735 (N_8735,N_8692,N_8640);
and U8736 (N_8736,N_8669,N_8693);
nand U8737 (N_8737,N_8677,N_8606);
nand U8738 (N_8738,N_8616,N_8657);
or U8739 (N_8739,N_8617,N_8619);
nand U8740 (N_8740,N_8642,N_8688);
nand U8741 (N_8741,N_8697,N_8641);
or U8742 (N_8742,N_8670,N_8681);
and U8743 (N_8743,N_8631,N_8679);
nand U8744 (N_8744,N_8622,N_8698);
and U8745 (N_8745,N_8629,N_8694);
nand U8746 (N_8746,N_8659,N_8633);
xor U8747 (N_8747,N_8690,N_8696);
nor U8748 (N_8748,N_8649,N_8676);
nand U8749 (N_8749,N_8650,N_8602);
and U8750 (N_8750,N_8674,N_8647);
or U8751 (N_8751,N_8651,N_8642);
or U8752 (N_8752,N_8608,N_8659);
nand U8753 (N_8753,N_8638,N_8657);
and U8754 (N_8754,N_8695,N_8633);
nor U8755 (N_8755,N_8699,N_8689);
xnor U8756 (N_8756,N_8600,N_8605);
nor U8757 (N_8757,N_8627,N_8674);
xnor U8758 (N_8758,N_8610,N_8679);
nand U8759 (N_8759,N_8673,N_8676);
and U8760 (N_8760,N_8612,N_8635);
nand U8761 (N_8761,N_8633,N_8697);
nor U8762 (N_8762,N_8652,N_8643);
or U8763 (N_8763,N_8623,N_8608);
and U8764 (N_8764,N_8642,N_8661);
nand U8765 (N_8765,N_8663,N_8675);
nand U8766 (N_8766,N_8649,N_8632);
nor U8767 (N_8767,N_8602,N_8644);
or U8768 (N_8768,N_8630,N_8663);
nor U8769 (N_8769,N_8678,N_8672);
nand U8770 (N_8770,N_8669,N_8648);
and U8771 (N_8771,N_8636,N_8694);
nand U8772 (N_8772,N_8632,N_8620);
xor U8773 (N_8773,N_8616,N_8613);
or U8774 (N_8774,N_8697,N_8608);
nor U8775 (N_8775,N_8651,N_8630);
xnor U8776 (N_8776,N_8613,N_8646);
and U8777 (N_8777,N_8691,N_8620);
or U8778 (N_8778,N_8688,N_8654);
and U8779 (N_8779,N_8648,N_8623);
nand U8780 (N_8780,N_8628,N_8643);
nand U8781 (N_8781,N_8663,N_8695);
and U8782 (N_8782,N_8623,N_8682);
nand U8783 (N_8783,N_8655,N_8658);
nand U8784 (N_8784,N_8649,N_8698);
and U8785 (N_8785,N_8697,N_8665);
xor U8786 (N_8786,N_8682,N_8685);
xnor U8787 (N_8787,N_8616,N_8668);
or U8788 (N_8788,N_8603,N_8671);
or U8789 (N_8789,N_8670,N_8637);
xnor U8790 (N_8790,N_8626,N_8678);
or U8791 (N_8791,N_8661,N_8646);
and U8792 (N_8792,N_8690,N_8637);
or U8793 (N_8793,N_8619,N_8663);
and U8794 (N_8794,N_8691,N_8632);
and U8795 (N_8795,N_8660,N_8619);
and U8796 (N_8796,N_8686,N_8664);
or U8797 (N_8797,N_8649,N_8620);
and U8798 (N_8798,N_8677,N_8616);
and U8799 (N_8799,N_8656,N_8690);
or U8800 (N_8800,N_8750,N_8731);
nand U8801 (N_8801,N_8783,N_8740);
nand U8802 (N_8802,N_8798,N_8730);
xor U8803 (N_8803,N_8765,N_8775);
and U8804 (N_8804,N_8782,N_8754);
xnor U8805 (N_8805,N_8702,N_8764);
nand U8806 (N_8806,N_8759,N_8790);
or U8807 (N_8807,N_8768,N_8792);
and U8808 (N_8808,N_8752,N_8763);
nor U8809 (N_8809,N_8743,N_8729);
or U8810 (N_8810,N_8758,N_8781);
and U8811 (N_8811,N_8799,N_8795);
or U8812 (N_8812,N_8709,N_8724);
xor U8813 (N_8813,N_8797,N_8760);
nand U8814 (N_8814,N_8769,N_8748);
nor U8815 (N_8815,N_8786,N_8789);
nand U8816 (N_8816,N_8700,N_8756);
xnor U8817 (N_8817,N_8733,N_8727);
xor U8818 (N_8818,N_8717,N_8725);
xnor U8819 (N_8819,N_8746,N_8737);
nor U8820 (N_8820,N_8757,N_8723);
nand U8821 (N_8821,N_8780,N_8706);
or U8822 (N_8822,N_8785,N_8715);
and U8823 (N_8823,N_8744,N_8776);
nor U8824 (N_8824,N_8774,N_8716);
nor U8825 (N_8825,N_8738,N_8751);
xnor U8826 (N_8826,N_8704,N_8734);
nor U8827 (N_8827,N_8705,N_8710);
nor U8828 (N_8828,N_8722,N_8726);
nand U8829 (N_8829,N_8773,N_8793);
nand U8830 (N_8830,N_8732,N_8794);
or U8831 (N_8831,N_8766,N_8711);
nor U8832 (N_8832,N_8714,N_8728);
xnor U8833 (N_8833,N_8772,N_8777);
and U8834 (N_8834,N_8771,N_8707);
and U8835 (N_8835,N_8761,N_8762);
or U8836 (N_8836,N_8713,N_8741);
nand U8837 (N_8837,N_8779,N_8735);
or U8838 (N_8838,N_8784,N_8770);
nand U8839 (N_8839,N_8701,N_8712);
nor U8840 (N_8840,N_8742,N_8747);
or U8841 (N_8841,N_8721,N_8708);
nand U8842 (N_8842,N_8736,N_8787);
nor U8843 (N_8843,N_8753,N_8739);
and U8844 (N_8844,N_8755,N_8791);
nand U8845 (N_8845,N_8703,N_8720);
and U8846 (N_8846,N_8778,N_8719);
nor U8847 (N_8847,N_8718,N_8749);
xnor U8848 (N_8848,N_8767,N_8745);
or U8849 (N_8849,N_8796,N_8788);
xor U8850 (N_8850,N_8715,N_8719);
nand U8851 (N_8851,N_8701,N_8707);
and U8852 (N_8852,N_8796,N_8777);
nor U8853 (N_8853,N_8704,N_8736);
and U8854 (N_8854,N_8798,N_8788);
nand U8855 (N_8855,N_8788,N_8707);
nand U8856 (N_8856,N_8786,N_8797);
and U8857 (N_8857,N_8779,N_8717);
nor U8858 (N_8858,N_8781,N_8716);
nand U8859 (N_8859,N_8704,N_8707);
nand U8860 (N_8860,N_8737,N_8722);
nor U8861 (N_8861,N_8721,N_8787);
nand U8862 (N_8862,N_8775,N_8736);
and U8863 (N_8863,N_8794,N_8727);
and U8864 (N_8864,N_8797,N_8714);
and U8865 (N_8865,N_8766,N_8790);
nand U8866 (N_8866,N_8780,N_8775);
and U8867 (N_8867,N_8755,N_8747);
nor U8868 (N_8868,N_8799,N_8771);
and U8869 (N_8869,N_8739,N_8747);
or U8870 (N_8870,N_8710,N_8781);
or U8871 (N_8871,N_8792,N_8779);
nand U8872 (N_8872,N_8795,N_8734);
or U8873 (N_8873,N_8749,N_8761);
nor U8874 (N_8874,N_8737,N_8779);
and U8875 (N_8875,N_8716,N_8739);
or U8876 (N_8876,N_8752,N_8734);
nor U8877 (N_8877,N_8774,N_8748);
nor U8878 (N_8878,N_8798,N_8720);
nor U8879 (N_8879,N_8770,N_8757);
or U8880 (N_8880,N_8768,N_8761);
xnor U8881 (N_8881,N_8770,N_8783);
xor U8882 (N_8882,N_8785,N_8728);
or U8883 (N_8883,N_8729,N_8714);
or U8884 (N_8884,N_8728,N_8740);
nor U8885 (N_8885,N_8755,N_8792);
nor U8886 (N_8886,N_8706,N_8718);
and U8887 (N_8887,N_8757,N_8735);
nand U8888 (N_8888,N_8752,N_8776);
nand U8889 (N_8889,N_8705,N_8704);
nor U8890 (N_8890,N_8771,N_8736);
and U8891 (N_8891,N_8704,N_8784);
nor U8892 (N_8892,N_8705,N_8719);
nor U8893 (N_8893,N_8760,N_8768);
nor U8894 (N_8894,N_8716,N_8796);
nand U8895 (N_8895,N_8704,N_8724);
or U8896 (N_8896,N_8722,N_8769);
and U8897 (N_8897,N_8730,N_8702);
and U8898 (N_8898,N_8738,N_8725);
or U8899 (N_8899,N_8787,N_8712);
xnor U8900 (N_8900,N_8812,N_8873);
nand U8901 (N_8901,N_8887,N_8804);
and U8902 (N_8902,N_8825,N_8897);
nand U8903 (N_8903,N_8841,N_8838);
nand U8904 (N_8904,N_8880,N_8835);
and U8905 (N_8905,N_8823,N_8800);
or U8906 (N_8906,N_8858,N_8808);
nor U8907 (N_8907,N_8843,N_8831);
nand U8908 (N_8908,N_8884,N_8848);
nand U8909 (N_8909,N_8829,N_8803);
nand U8910 (N_8910,N_8802,N_8861);
and U8911 (N_8911,N_8855,N_8814);
nand U8912 (N_8912,N_8853,N_8868);
nand U8913 (N_8913,N_8866,N_8886);
and U8914 (N_8914,N_8883,N_8834);
nand U8915 (N_8915,N_8864,N_8863);
and U8916 (N_8916,N_8871,N_8879);
nor U8917 (N_8917,N_8805,N_8816);
and U8918 (N_8918,N_8822,N_8859);
nand U8919 (N_8919,N_8839,N_8870);
or U8920 (N_8920,N_8882,N_8807);
and U8921 (N_8921,N_8846,N_8847);
or U8922 (N_8922,N_8815,N_8824);
or U8923 (N_8923,N_8867,N_8872);
nor U8924 (N_8924,N_8828,N_8874);
and U8925 (N_8925,N_8850,N_8840);
nand U8926 (N_8926,N_8833,N_8827);
or U8927 (N_8927,N_8826,N_8862);
and U8928 (N_8928,N_8811,N_8898);
nor U8929 (N_8929,N_8860,N_8810);
and U8930 (N_8930,N_8801,N_8896);
or U8931 (N_8931,N_8865,N_8845);
nor U8932 (N_8932,N_8894,N_8849);
and U8933 (N_8933,N_8818,N_8809);
or U8934 (N_8934,N_8856,N_8881);
nand U8935 (N_8935,N_8891,N_8876);
and U8936 (N_8936,N_8813,N_8844);
and U8937 (N_8937,N_8852,N_8832);
nand U8938 (N_8938,N_8889,N_8819);
nand U8939 (N_8939,N_8869,N_8892);
nor U8940 (N_8940,N_8885,N_8821);
nand U8941 (N_8941,N_8878,N_8837);
nand U8942 (N_8942,N_8893,N_8820);
nor U8943 (N_8943,N_8888,N_8875);
and U8944 (N_8944,N_8851,N_8877);
or U8945 (N_8945,N_8842,N_8857);
and U8946 (N_8946,N_8899,N_8854);
or U8947 (N_8947,N_8895,N_8817);
xor U8948 (N_8948,N_8806,N_8830);
nand U8949 (N_8949,N_8890,N_8836);
or U8950 (N_8950,N_8831,N_8850);
nand U8951 (N_8951,N_8868,N_8831);
or U8952 (N_8952,N_8845,N_8894);
nand U8953 (N_8953,N_8875,N_8893);
nor U8954 (N_8954,N_8896,N_8804);
nand U8955 (N_8955,N_8887,N_8821);
nand U8956 (N_8956,N_8840,N_8802);
or U8957 (N_8957,N_8820,N_8855);
and U8958 (N_8958,N_8878,N_8870);
nand U8959 (N_8959,N_8828,N_8801);
nand U8960 (N_8960,N_8859,N_8874);
and U8961 (N_8961,N_8841,N_8864);
nor U8962 (N_8962,N_8820,N_8887);
nor U8963 (N_8963,N_8882,N_8885);
and U8964 (N_8964,N_8801,N_8872);
nand U8965 (N_8965,N_8809,N_8846);
and U8966 (N_8966,N_8874,N_8833);
or U8967 (N_8967,N_8888,N_8851);
nand U8968 (N_8968,N_8848,N_8806);
and U8969 (N_8969,N_8881,N_8873);
xnor U8970 (N_8970,N_8872,N_8893);
or U8971 (N_8971,N_8844,N_8842);
nand U8972 (N_8972,N_8818,N_8856);
or U8973 (N_8973,N_8807,N_8803);
nand U8974 (N_8974,N_8828,N_8864);
xnor U8975 (N_8975,N_8852,N_8803);
nand U8976 (N_8976,N_8800,N_8898);
nor U8977 (N_8977,N_8834,N_8844);
and U8978 (N_8978,N_8844,N_8896);
nor U8979 (N_8979,N_8882,N_8896);
or U8980 (N_8980,N_8828,N_8850);
nand U8981 (N_8981,N_8880,N_8845);
and U8982 (N_8982,N_8894,N_8897);
or U8983 (N_8983,N_8836,N_8807);
nor U8984 (N_8984,N_8879,N_8844);
nor U8985 (N_8985,N_8864,N_8851);
nand U8986 (N_8986,N_8896,N_8891);
nor U8987 (N_8987,N_8849,N_8865);
nor U8988 (N_8988,N_8852,N_8851);
nor U8989 (N_8989,N_8800,N_8841);
and U8990 (N_8990,N_8880,N_8807);
nand U8991 (N_8991,N_8827,N_8891);
nand U8992 (N_8992,N_8836,N_8847);
or U8993 (N_8993,N_8846,N_8883);
and U8994 (N_8994,N_8847,N_8885);
nor U8995 (N_8995,N_8833,N_8843);
nand U8996 (N_8996,N_8825,N_8882);
nand U8997 (N_8997,N_8832,N_8810);
or U8998 (N_8998,N_8843,N_8858);
nor U8999 (N_8999,N_8814,N_8861);
and U9000 (N_9000,N_8965,N_8959);
and U9001 (N_9001,N_8952,N_8905);
nand U9002 (N_9002,N_8931,N_8981);
or U9003 (N_9003,N_8903,N_8997);
xor U9004 (N_9004,N_8945,N_8938);
and U9005 (N_9005,N_8940,N_8999);
and U9006 (N_9006,N_8969,N_8973);
nor U9007 (N_9007,N_8910,N_8930);
nor U9008 (N_9008,N_8923,N_8942);
nand U9009 (N_9009,N_8960,N_8953);
nor U9010 (N_9010,N_8970,N_8980);
and U9011 (N_9011,N_8950,N_8967);
or U9012 (N_9012,N_8920,N_8958);
and U9013 (N_9013,N_8989,N_8909);
nor U9014 (N_9014,N_8994,N_8964);
or U9015 (N_9015,N_8904,N_8936);
and U9016 (N_9016,N_8990,N_8916);
nor U9017 (N_9017,N_8979,N_8917);
nand U9018 (N_9018,N_8961,N_8957);
and U9019 (N_9019,N_8993,N_8928);
nand U9020 (N_9020,N_8908,N_8934);
or U9021 (N_9021,N_8988,N_8985);
nor U9022 (N_9022,N_8998,N_8927);
xnor U9023 (N_9023,N_8939,N_8963);
or U9024 (N_9024,N_8983,N_8941);
or U9025 (N_9025,N_8947,N_8968);
and U9026 (N_9026,N_8951,N_8992);
xnor U9027 (N_9027,N_8919,N_8924);
nor U9028 (N_9028,N_8978,N_8918);
nand U9029 (N_9029,N_8925,N_8984);
and U9030 (N_9030,N_8954,N_8974);
or U9031 (N_9031,N_8962,N_8996);
and U9032 (N_9032,N_8913,N_8935);
and U9033 (N_9033,N_8944,N_8943);
nand U9034 (N_9034,N_8902,N_8977);
nand U9035 (N_9035,N_8982,N_8921);
nor U9036 (N_9036,N_8991,N_8933);
and U9037 (N_9037,N_8995,N_8966);
and U9038 (N_9038,N_8900,N_8948);
nand U9039 (N_9039,N_8955,N_8972);
nand U9040 (N_9040,N_8986,N_8987);
nor U9041 (N_9041,N_8911,N_8929);
nor U9042 (N_9042,N_8912,N_8932);
or U9043 (N_9043,N_8906,N_8901);
nand U9044 (N_9044,N_8956,N_8926);
nor U9045 (N_9045,N_8914,N_8922);
nor U9046 (N_9046,N_8907,N_8971);
nor U9047 (N_9047,N_8949,N_8975);
or U9048 (N_9048,N_8976,N_8915);
nand U9049 (N_9049,N_8937,N_8946);
nor U9050 (N_9050,N_8919,N_8952);
and U9051 (N_9051,N_8950,N_8952);
and U9052 (N_9052,N_8946,N_8942);
nand U9053 (N_9053,N_8925,N_8955);
and U9054 (N_9054,N_8995,N_8983);
nor U9055 (N_9055,N_8942,N_8976);
nor U9056 (N_9056,N_8992,N_8969);
nor U9057 (N_9057,N_8940,N_8969);
or U9058 (N_9058,N_8974,N_8958);
and U9059 (N_9059,N_8941,N_8910);
nor U9060 (N_9060,N_8930,N_8928);
and U9061 (N_9061,N_8956,N_8991);
and U9062 (N_9062,N_8974,N_8973);
xnor U9063 (N_9063,N_8911,N_8951);
nand U9064 (N_9064,N_8976,N_8996);
nand U9065 (N_9065,N_8920,N_8947);
and U9066 (N_9066,N_8976,N_8907);
and U9067 (N_9067,N_8949,N_8938);
nand U9068 (N_9068,N_8912,N_8974);
nand U9069 (N_9069,N_8964,N_8916);
nand U9070 (N_9070,N_8901,N_8981);
or U9071 (N_9071,N_8947,N_8959);
nor U9072 (N_9072,N_8926,N_8934);
or U9073 (N_9073,N_8985,N_8922);
nor U9074 (N_9074,N_8910,N_8947);
or U9075 (N_9075,N_8999,N_8951);
and U9076 (N_9076,N_8996,N_8951);
and U9077 (N_9077,N_8973,N_8910);
or U9078 (N_9078,N_8982,N_8930);
or U9079 (N_9079,N_8953,N_8932);
and U9080 (N_9080,N_8989,N_8900);
and U9081 (N_9081,N_8922,N_8991);
nand U9082 (N_9082,N_8976,N_8939);
or U9083 (N_9083,N_8921,N_8930);
nand U9084 (N_9084,N_8971,N_8968);
or U9085 (N_9085,N_8969,N_8963);
nand U9086 (N_9086,N_8925,N_8901);
or U9087 (N_9087,N_8948,N_8922);
and U9088 (N_9088,N_8975,N_8948);
nor U9089 (N_9089,N_8997,N_8950);
nor U9090 (N_9090,N_8909,N_8998);
or U9091 (N_9091,N_8907,N_8955);
nand U9092 (N_9092,N_8961,N_8912);
nand U9093 (N_9093,N_8965,N_8944);
nor U9094 (N_9094,N_8927,N_8978);
xnor U9095 (N_9095,N_8991,N_8932);
and U9096 (N_9096,N_8942,N_8928);
nand U9097 (N_9097,N_8925,N_8911);
nor U9098 (N_9098,N_8913,N_8954);
or U9099 (N_9099,N_8978,N_8935);
and U9100 (N_9100,N_9062,N_9008);
nand U9101 (N_9101,N_9052,N_9023);
nand U9102 (N_9102,N_9090,N_9017);
or U9103 (N_9103,N_9036,N_9012);
nand U9104 (N_9104,N_9013,N_9033);
nor U9105 (N_9105,N_9081,N_9061);
and U9106 (N_9106,N_9049,N_9074);
and U9107 (N_9107,N_9022,N_9001);
or U9108 (N_9108,N_9096,N_9046);
nor U9109 (N_9109,N_9063,N_9009);
nor U9110 (N_9110,N_9000,N_9019);
and U9111 (N_9111,N_9010,N_9016);
and U9112 (N_9112,N_9079,N_9064);
and U9113 (N_9113,N_9099,N_9055);
and U9114 (N_9114,N_9070,N_9085);
or U9115 (N_9115,N_9034,N_9069);
nand U9116 (N_9116,N_9048,N_9066);
or U9117 (N_9117,N_9005,N_9026);
nor U9118 (N_9118,N_9027,N_9043);
nand U9119 (N_9119,N_9084,N_9057);
nor U9120 (N_9120,N_9083,N_9007);
and U9121 (N_9121,N_9072,N_9025);
or U9122 (N_9122,N_9003,N_9095);
or U9123 (N_9123,N_9093,N_9056);
or U9124 (N_9124,N_9040,N_9053);
nand U9125 (N_9125,N_9089,N_9018);
and U9126 (N_9126,N_9014,N_9060);
nor U9127 (N_9127,N_9042,N_9097);
nand U9128 (N_9128,N_9030,N_9075);
xnor U9129 (N_9129,N_9091,N_9045);
and U9130 (N_9130,N_9059,N_9050);
nor U9131 (N_9131,N_9006,N_9028);
xor U9132 (N_9132,N_9002,N_9094);
nand U9133 (N_9133,N_9039,N_9021);
and U9134 (N_9134,N_9087,N_9080);
or U9135 (N_9135,N_9035,N_9031);
and U9136 (N_9136,N_9098,N_9041);
nor U9137 (N_9137,N_9020,N_9067);
nor U9138 (N_9138,N_9068,N_9073);
nor U9139 (N_9139,N_9011,N_9058);
and U9140 (N_9140,N_9076,N_9051);
or U9141 (N_9141,N_9024,N_9077);
xor U9142 (N_9142,N_9015,N_9044);
xnor U9143 (N_9143,N_9047,N_9082);
and U9144 (N_9144,N_9071,N_9037);
nor U9145 (N_9145,N_9029,N_9038);
xor U9146 (N_9146,N_9078,N_9065);
and U9147 (N_9147,N_9054,N_9032);
or U9148 (N_9148,N_9086,N_9092);
nand U9149 (N_9149,N_9004,N_9088);
nand U9150 (N_9150,N_9057,N_9053);
or U9151 (N_9151,N_9013,N_9048);
nand U9152 (N_9152,N_9038,N_9004);
nor U9153 (N_9153,N_9077,N_9044);
nor U9154 (N_9154,N_9090,N_9009);
nor U9155 (N_9155,N_9076,N_9096);
or U9156 (N_9156,N_9024,N_9022);
and U9157 (N_9157,N_9010,N_9074);
nor U9158 (N_9158,N_9082,N_9044);
and U9159 (N_9159,N_9024,N_9060);
or U9160 (N_9160,N_9092,N_9081);
and U9161 (N_9161,N_9081,N_9051);
nand U9162 (N_9162,N_9006,N_9000);
and U9163 (N_9163,N_9019,N_9042);
and U9164 (N_9164,N_9004,N_9003);
nand U9165 (N_9165,N_9021,N_9094);
or U9166 (N_9166,N_9081,N_9065);
xnor U9167 (N_9167,N_9034,N_9091);
and U9168 (N_9168,N_9063,N_9001);
nor U9169 (N_9169,N_9062,N_9073);
or U9170 (N_9170,N_9021,N_9067);
or U9171 (N_9171,N_9093,N_9013);
nor U9172 (N_9172,N_9086,N_9079);
and U9173 (N_9173,N_9026,N_9098);
or U9174 (N_9174,N_9096,N_9030);
nand U9175 (N_9175,N_9034,N_9052);
and U9176 (N_9176,N_9013,N_9022);
and U9177 (N_9177,N_9035,N_9087);
or U9178 (N_9178,N_9084,N_9033);
or U9179 (N_9179,N_9032,N_9074);
and U9180 (N_9180,N_9088,N_9076);
and U9181 (N_9181,N_9063,N_9080);
and U9182 (N_9182,N_9012,N_9007);
xnor U9183 (N_9183,N_9007,N_9076);
or U9184 (N_9184,N_9018,N_9088);
nor U9185 (N_9185,N_9087,N_9010);
nand U9186 (N_9186,N_9053,N_9068);
or U9187 (N_9187,N_9001,N_9086);
nand U9188 (N_9188,N_9039,N_9093);
or U9189 (N_9189,N_9049,N_9099);
nand U9190 (N_9190,N_9027,N_9031);
nand U9191 (N_9191,N_9082,N_9097);
and U9192 (N_9192,N_9089,N_9016);
xor U9193 (N_9193,N_9003,N_9089);
xor U9194 (N_9194,N_9067,N_9077);
nand U9195 (N_9195,N_9097,N_9062);
nor U9196 (N_9196,N_9062,N_9065);
nand U9197 (N_9197,N_9092,N_9078);
xor U9198 (N_9198,N_9015,N_9003);
xor U9199 (N_9199,N_9087,N_9090);
xor U9200 (N_9200,N_9164,N_9162);
nand U9201 (N_9201,N_9167,N_9188);
nand U9202 (N_9202,N_9148,N_9113);
xnor U9203 (N_9203,N_9158,N_9172);
xor U9204 (N_9204,N_9177,N_9144);
and U9205 (N_9205,N_9173,N_9165);
nor U9206 (N_9206,N_9191,N_9128);
nor U9207 (N_9207,N_9145,N_9124);
or U9208 (N_9208,N_9121,N_9169);
nor U9209 (N_9209,N_9175,N_9174);
nand U9210 (N_9210,N_9156,N_9107);
or U9211 (N_9211,N_9168,N_9140);
or U9212 (N_9212,N_9184,N_9163);
or U9213 (N_9213,N_9138,N_9102);
nor U9214 (N_9214,N_9131,N_9133);
nor U9215 (N_9215,N_9195,N_9100);
nand U9216 (N_9216,N_9186,N_9142);
xor U9217 (N_9217,N_9111,N_9159);
nor U9218 (N_9218,N_9176,N_9119);
xnor U9219 (N_9219,N_9105,N_9134);
or U9220 (N_9220,N_9198,N_9104);
nand U9221 (N_9221,N_9181,N_9179);
and U9222 (N_9222,N_9178,N_9190);
nand U9223 (N_9223,N_9153,N_9129);
and U9224 (N_9224,N_9171,N_9147);
nor U9225 (N_9225,N_9161,N_9106);
and U9226 (N_9226,N_9160,N_9112);
and U9227 (N_9227,N_9152,N_9136);
nand U9228 (N_9228,N_9108,N_9101);
nand U9229 (N_9229,N_9117,N_9130);
and U9230 (N_9230,N_9125,N_9137);
nand U9231 (N_9231,N_9135,N_9123);
or U9232 (N_9232,N_9116,N_9182);
and U9233 (N_9233,N_9118,N_9189);
nand U9234 (N_9234,N_9109,N_9115);
or U9235 (N_9235,N_9122,N_9143);
xnor U9236 (N_9236,N_9154,N_9192);
and U9237 (N_9237,N_9197,N_9114);
and U9238 (N_9238,N_9155,N_9132);
and U9239 (N_9239,N_9139,N_9166);
nor U9240 (N_9240,N_9194,N_9141);
nand U9241 (N_9241,N_9180,N_9187);
nand U9242 (N_9242,N_9199,N_9150);
nor U9243 (N_9243,N_9110,N_9183);
or U9244 (N_9244,N_9120,N_9127);
nor U9245 (N_9245,N_9146,N_9170);
or U9246 (N_9246,N_9193,N_9151);
nor U9247 (N_9247,N_9185,N_9103);
nand U9248 (N_9248,N_9126,N_9196);
nand U9249 (N_9249,N_9157,N_9149);
nand U9250 (N_9250,N_9167,N_9131);
nand U9251 (N_9251,N_9143,N_9153);
or U9252 (N_9252,N_9136,N_9106);
or U9253 (N_9253,N_9155,N_9101);
nand U9254 (N_9254,N_9138,N_9184);
or U9255 (N_9255,N_9120,N_9190);
nor U9256 (N_9256,N_9163,N_9183);
or U9257 (N_9257,N_9139,N_9199);
nand U9258 (N_9258,N_9160,N_9133);
nor U9259 (N_9259,N_9167,N_9103);
or U9260 (N_9260,N_9194,N_9140);
nor U9261 (N_9261,N_9157,N_9129);
nand U9262 (N_9262,N_9169,N_9135);
or U9263 (N_9263,N_9137,N_9195);
and U9264 (N_9264,N_9103,N_9151);
nor U9265 (N_9265,N_9146,N_9110);
nor U9266 (N_9266,N_9122,N_9173);
and U9267 (N_9267,N_9151,N_9134);
xor U9268 (N_9268,N_9132,N_9189);
and U9269 (N_9269,N_9155,N_9153);
or U9270 (N_9270,N_9133,N_9189);
xnor U9271 (N_9271,N_9107,N_9132);
nand U9272 (N_9272,N_9187,N_9186);
or U9273 (N_9273,N_9150,N_9128);
and U9274 (N_9274,N_9136,N_9113);
or U9275 (N_9275,N_9123,N_9157);
nor U9276 (N_9276,N_9167,N_9132);
or U9277 (N_9277,N_9174,N_9162);
or U9278 (N_9278,N_9193,N_9130);
or U9279 (N_9279,N_9152,N_9104);
and U9280 (N_9280,N_9130,N_9103);
nor U9281 (N_9281,N_9109,N_9150);
or U9282 (N_9282,N_9100,N_9135);
or U9283 (N_9283,N_9137,N_9103);
and U9284 (N_9284,N_9167,N_9166);
or U9285 (N_9285,N_9130,N_9118);
nor U9286 (N_9286,N_9175,N_9143);
nor U9287 (N_9287,N_9174,N_9148);
nor U9288 (N_9288,N_9163,N_9146);
nor U9289 (N_9289,N_9199,N_9151);
or U9290 (N_9290,N_9102,N_9185);
and U9291 (N_9291,N_9190,N_9114);
nand U9292 (N_9292,N_9164,N_9192);
nor U9293 (N_9293,N_9155,N_9103);
nor U9294 (N_9294,N_9163,N_9159);
or U9295 (N_9295,N_9199,N_9101);
xor U9296 (N_9296,N_9128,N_9160);
nand U9297 (N_9297,N_9199,N_9179);
nor U9298 (N_9298,N_9194,N_9198);
and U9299 (N_9299,N_9100,N_9145);
and U9300 (N_9300,N_9293,N_9200);
nand U9301 (N_9301,N_9248,N_9256);
nand U9302 (N_9302,N_9212,N_9239);
and U9303 (N_9303,N_9281,N_9289);
nor U9304 (N_9304,N_9273,N_9279);
xnor U9305 (N_9305,N_9250,N_9235);
nor U9306 (N_9306,N_9287,N_9265);
and U9307 (N_9307,N_9247,N_9278);
nand U9308 (N_9308,N_9263,N_9232);
and U9309 (N_9309,N_9228,N_9218);
nor U9310 (N_9310,N_9286,N_9226);
or U9311 (N_9311,N_9282,N_9277);
nor U9312 (N_9312,N_9292,N_9274);
nand U9313 (N_9313,N_9276,N_9272);
or U9314 (N_9314,N_9245,N_9259);
nor U9315 (N_9315,N_9234,N_9298);
or U9316 (N_9316,N_9219,N_9291);
nor U9317 (N_9317,N_9242,N_9211);
or U9318 (N_9318,N_9238,N_9285);
or U9319 (N_9319,N_9216,N_9251);
or U9320 (N_9320,N_9270,N_9240);
or U9321 (N_9321,N_9241,N_9201);
and U9322 (N_9322,N_9261,N_9220);
xnor U9323 (N_9323,N_9210,N_9254);
or U9324 (N_9324,N_9215,N_9266);
nor U9325 (N_9325,N_9203,N_9207);
nand U9326 (N_9326,N_9227,N_9267);
and U9327 (N_9327,N_9243,N_9224);
or U9328 (N_9328,N_9230,N_9231);
nand U9329 (N_9329,N_9284,N_9258);
xor U9330 (N_9330,N_9271,N_9217);
or U9331 (N_9331,N_9269,N_9297);
nor U9332 (N_9332,N_9262,N_9255);
and U9333 (N_9333,N_9253,N_9252);
nor U9334 (N_9334,N_9221,N_9264);
nor U9335 (N_9335,N_9288,N_9246);
and U9336 (N_9336,N_9206,N_9233);
or U9337 (N_9337,N_9236,N_9223);
and U9338 (N_9338,N_9290,N_9296);
and U9339 (N_9339,N_9299,N_9257);
xor U9340 (N_9340,N_9204,N_9208);
nand U9341 (N_9341,N_9268,N_9295);
nor U9342 (N_9342,N_9214,N_9225);
or U9343 (N_9343,N_9202,N_9222);
nor U9344 (N_9344,N_9260,N_9229);
and U9345 (N_9345,N_9294,N_9249);
and U9346 (N_9346,N_9205,N_9283);
or U9347 (N_9347,N_9280,N_9244);
nor U9348 (N_9348,N_9237,N_9275);
nand U9349 (N_9349,N_9209,N_9213);
nor U9350 (N_9350,N_9290,N_9208);
and U9351 (N_9351,N_9296,N_9277);
or U9352 (N_9352,N_9246,N_9230);
and U9353 (N_9353,N_9288,N_9220);
nand U9354 (N_9354,N_9210,N_9267);
xor U9355 (N_9355,N_9204,N_9228);
xnor U9356 (N_9356,N_9240,N_9283);
xnor U9357 (N_9357,N_9277,N_9204);
xnor U9358 (N_9358,N_9219,N_9295);
nand U9359 (N_9359,N_9234,N_9229);
nand U9360 (N_9360,N_9231,N_9270);
nand U9361 (N_9361,N_9287,N_9204);
or U9362 (N_9362,N_9232,N_9285);
xor U9363 (N_9363,N_9212,N_9271);
and U9364 (N_9364,N_9222,N_9213);
xnor U9365 (N_9365,N_9216,N_9281);
or U9366 (N_9366,N_9282,N_9210);
nor U9367 (N_9367,N_9215,N_9208);
and U9368 (N_9368,N_9234,N_9264);
and U9369 (N_9369,N_9277,N_9286);
or U9370 (N_9370,N_9205,N_9268);
nand U9371 (N_9371,N_9247,N_9245);
and U9372 (N_9372,N_9227,N_9283);
nor U9373 (N_9373,N_9225,N_9233);
nand U9374 (N_9374,N_9223,N_9218);
nand U9375 (N_9375,N_9218,N_9213);
and U9376 (N_9376,N_9295,N_9270);
or U9377 (N_9377,N_9279,N_9200);
nand U9378 (N_9378,N_9246,N_9268);
nor U9379 (N_9379,N_9225,N_9289);
nand U9380 (N_9380,N_9210,N_9205);
or U9381 (N_9381,N_9245,N_9279);
or U9382 (N_9382,N_9209,N_9265);
or U9383 (N_9383,N_9282,N_9235);
or U9384 (N_9384,N_9214,N_9221);
xor U9385 (N_9385,N_9213,N_9266);
nand U9386 (N_9386,N_9215,N_9204);
xnor U9387 (N_9387,N_9272,N_9239);
and U9388 (N_9388,N_9253,N_9260);
and U9389 (N_9389,N_9236,N_9244);
nand U9390 (N_9390,N_9215,N_9212);
xnor U9391 (N_9391,N_9206,N_9284);
and U9392 (N_9392,N_9266,N_9269);
nand U9393 (N_9393,N_9275,N_9231);
and U9394 (N_9394,N_9233,N_9216);
nor U9395 (N_9395,N_9230,N_9207);
and U9396 (N_9396,N_9284,N_9201);
xor U9397 (N_9397,N_9298,N_9262);
and U9398 (N_9398,N_9202,N_9204);
or U9399 (N_9399,N_9217,N_9292);
or U9400 (N_9400,N_9305,N_9381);
xnor U9401 (N_9401,N_9352,N_9329);
and U9402 (N_9402,N_9398,N_9373);
and U9403 (N_9403,N_9316,N_9369);
and U9404 (N_9404,N_9354,N_9383);
and U9405 (N_9405,N_9335,N_9377);
xnor U9406 (N_9406,N_9355,N_9360);
or U9407 (N_9407,N_9328,N_9389);
or U9408 (N_9408,N_9379,N_9320);
nor U9409 (N_9409,N_9333,N_9346);
and U9410 (N_9410,N_9345,N_9372);
and U9411 (N_9411,N_9388,N_9327);
xor U9412 (N_9412,N_9353,N_9348);
nor U9413 (N_9413,N_9336,N_9395);
nand U9414 (N_9414,N_9351,N_9315);
nand U9415 (N_9415,N_9358,N_9370);
and U9416 (N_9416,N_9385,N_9350);
xnor U9417 (N_9417,N_9374,N_9396);
and U9418 (N_9418,N_9380,N_9392);
nor U9419 (N_9419,N_9317,N_9397);
and U9420 (N_9420,N_9302,N_9349);
nor U9421 (N_9421,N_9324,N_9331);
and U9422 (N_9422,N_9332,N_9306);
nand U9423 (N_9423,N_9310,N_9347);
xor U9424 (N_9424,N_9341,N_9309);
xnor U9425 (N_9425,N_9344,N_9363);
nand U9426 (N_9426,N_9337,N_9319);
nand U9427 (N_9427,N_9312,N_9371);
nor U9428 (N_9428,N_9359,N_9338);
nand U9429 (N_9429,N_9342,N_9303);
and U9430 (N_9430,N_9390,N_9313);
and U9431 (N_9431,N_9393,N_9311);
or U9432 (N_9432,N_9399,N_9321);
nor U9433 (N_9433,N_9394,N_9339);
and U9434 (N_9434,N_9356,N_9367);
xnor U9435 (N_9435,N_9382,N_9378);
and U9436 (N_9436,N_9314,N_9323);
and U9437 (N_9437,N_9387,N_9361);
and U9438 (N_9438,N_9326,N_9325);
nand U9439 (N_9439,N_9368,N_9365);
or U9440 (N_9440,N_9318,N_9308);
nor U9441 (N_9441,N_9343,N_9386);
nand U9442 (N_9442,N_9366,N_9376);
nor U9443 (N_9443,N_9375,N_9391);
nand U9444 (N_9444,N_9322,N_9300);
nor U9445 (N_9445,N_9357,N_9340);
nand U9446 (N_9446,N_9384,N_9334);
or U9447 (N_9447,N_9301,N_9330);
nor U9448 (N_9448,N_9304,N_9362);
nor U9449 (N_9449,N_9307,N_9364);
nor U9450 (N_9450,N_9322,N_9328);
or U9451 (N_9451,N_9342,N_9320);
xnor U9452 (N_9452,N_9397,N_9365);
or U9453 (N_9453,N_9362,N_9308);
and U9454 (N_9454,N_9328,N_9323);
xor U9455 (N_9455,N_9314,N_9375);
and U9456 (N_9456,N_9308,N_9301);
nor U9457 (N_9457,N_9385,N_9373);
nand U9458 (N_9458,N_9375,N_9303);
nor U9459 (N_9459,N_9321,N_9390);
and U9460 (N_9460,N_9340,N_9300);
nor U9461 (N_9461,N_9328,N_9318);
xor U9462 (N_9462,N_9383,N_9376);
nand U9463 (N_9463,N_9386,N_9397);
and U9464 (N_9464,N_9319,N_9345);
xnor U9465 (N_9465,N_9344,N_9343);
nand U9466 (N_9466,N_9379,N_9370);
and U9467 (N_9467,N_9317,N_9383);
nand U9468 (N_9468,N_9305,N_9389);
nand U9469 (N_9469,N_9387,N_9393);
and U9470 (N_9470,N_9388,N_9382);
xor U9471 (N_9471,N_9377,N_9382);
nor U9472 (N_9472,N_9399,N_9333);
or U9473 (N_9473,N_9322,N_9361);
xor U9474 (N_9474,N_9310,N_9362);
and U9475 (N_9475,N_9318,N_9372);
xor U9476 (N_9476,N_9369,N_9377);
or U9477 (N_9477,N_9388,N_9385);
nand U9478 (N_9478,N_9359,N_9382);
nor U9479 (N_9479,N_9346,N_9325);
and U9480 (N_9480,N_9321,N_9317);
and U9481 (N_9481,N_9316,N_9394);
nor U9482 (N_9482,N_9370,N_9372);
nor U9483 (N_9483,N_9389,N_9395);
or U9484 (N_9484,N_9305,N_9386);
or U9485 (N_9485,N_9312,N_9321);
nor U9486 (N_9486,N_9342,N_9359);
and U9487 (N_9487,N_9301,N_9349);
and U9488 (N_9488,N_9328,N_9366);
or U9489 (N_9489,N_9318,N_9330);
nand U9490 (N_9490,N_9352,N_9394);
nor U9491 (N_9491,N_9303,N_9385);
or U9492 (N_9492,N_9301,N_9356);
or U9493 (N_9493,N_9375,N_9370);
or U9494 (N_9494,N_9381,N_9344);
or U9495 (N_9495,N_9393,N_9396);
xor U9496 (N_9496,N_9338,N_9398);
nand U9497 (N_9497,N_9365,N_9390);
or U9498 (N_9498,N_9311,N_9380);
nor U9499 (N_9499,N_9331,N_9379);
nor U9500 (N_9500,N_9469,N_9437);
nor U9501 (N_9501,N_9436,N_9407);
nand U9502 (N_9502,N_9491,N_9483);
nor U9503 (N_9503,N_9422,N_9443);
nand U9504 (N_9504,N_9497,N_9489);
and U9505 (N_9505,N_9415,N_9414);
nor U9506 (N_9506,N_9482,N_9479);
and U9507 (N_9507,N_9435,N_9484);
xnor U9508 (N_9508,N_9488,N_9474);
nor U9509 (N_9509,N_9444,N_9433);
nor U9510 (N_9510,N_9403,N_9438);
xor U9511 (N_9511,N_9411,N_9464);
nand U9512 (N_9512,N_9495,N_9463);
and U9513 (N_9513,N_9410,N_9467);
or U9514 (N_9514,N_9480,N_9409);
nand U9515 (N_9515,N_9476,N_9473);
nand U9516 (N_9516,N_9478,N_9470);
nor U9517 (N_9517,N_9453,N_9421);
xor U9518 (N_9518,N_9449,N_9458);
nor U9519 (N_9519,N_9429,N_9405);
and U9520 (N_9520,N_9448,N_9452);
and U9521 (N_9521,N_9499,N_9412);
nand U9522 (N_9522,N_9408,N_9404);
xnor U9523 (N_9523,N_9494,N_9492);
nand U9524 (N_9524,N_9401,N_9423);
xor U9525 (N_9525,N_9424,N_9426);
and U9526 (N_9526,N_9455,N_9461);
nor U9527 (N_9527,N_9472,N_9431);
and U9528 (N_9528,N_9406,N_9481);
or U9529 (N_9529,N_9418,N_9446);
and U9530 (N_9530,N_9477,N_9486);
and U9531 (N_9531,N_9413,N_9471);
and U9532 (N_9532,N_9434,N_9457);
or U9533 (N_9533,N_9428,N_9456);
or U9534 (N_9534,N_9400,N_9465);
nand U9535 (N_9535,N_9485,N_9487);
nand U9536 (N_9536,N_9402,N_9442);
and U9537 (N_9537,N_9432,N_9493);
nor U9538 (N_9538,N_9440,N_9427);
nor U9539 (N_9539,N_9460,N_9459);
nor U9540 (N_9540,N_9496,N_9439);
and U9541 (N_9541,N_9462,N_9475);
nand U9542 (N_9542,N_9441,N_9468);
or U9543 (N_9543,N_9425,N_9419);
nand U9544 (N_9544,N_9445,N_9498);
xnor U9545 (N_9545,N_9451,N_9416);
nand U9546 (N_9546,N_9466,N_9430);
nand U9547 (N_9547,N_9420,N_9454);
or U9548 (N_9548,N_9417,N_9490);
or U9549 (N_9549,N_9450,N_9447);
nor U9550 (N_9550,N_9456,N_9458);
xor U9551 (N_9551,N_9464,N_9429);
nor U9552 (N_9552,N_9489,N_9498);
nand U9553 (N_9553,N_9460,N_9409);
xnor U9554 (N_9554,N_9497,N_9418);
nand U9555 (N_9555,N_9456,N_9441);
or U9556 (N_9556,N_9474,N_9462);
or U9557 (N_9557,N_9445,N_9472);
nor U9558 (N_9558,N_9481,N_9405);
nor U9559 (N_9559,N_9403,N_9417);
nand U9560 (N_9560,N_9486,N_9450);
or U9561 (N_9561,N_9484,N_9479);
or U9562 (N_9562,N_9407,N_9484);
and U9563 (N_9563,N_9475,N_9453);
nor U9564 (N_9564,N_9454,N_9499);
xnor U9565 (N_9565,N_9426,N_9467);
nand U9566 (N_9566,N_9461,N_9445);
nor U9567 (N_9567,N_9441,N_9411);
nor U9568 (N_9568,N_9422,N_9472);
xor U9569 (N_9569,N_9448,N_9446);
nor U9570 (N_9570,N_9481,N_9423);
xor U9571 (N_9571,N_9414,N_9496);
and U9572 (N_9572,N_9466,N_9487);
xor U9573 (N_9573,N_9445,N_9412);
xnor U9574 (N_9574,N_9472,N_9401);
nand U9575 (N_9575,N_9453,N_9477);
nand U9576 (N_9576,N_9465,N_9443);
nand U9577 (N_9577,N_9479,N_9455);
xor U9578 (N_9578,N_9421,N_9438);
and U9579 (N_9579,N_9412,N_9448);
nand U9580 (N_9580,N_9440,N_9454);
nand U9581 (N_9581,N_9472,N_9454);
and U9582 (N_9582,N_9454,N_9497);
nor U9583 (N_9583,N_9445,N_9488);
or U9584 (N_9584,N_9487,N_9423);
or U9585 (N_9585,N_9458,N_9473);
nor U9586 (N_9586,N_9487,N_9405);
and U9587 (N_9587,N_9446,N_9405);
nand U9588 (N_9588,N_9464,N_9436);
nand U9589 (N_9589,N_9404,N_9473);
nand U9590 (N_9590,N_9421,N_9464);
xor U9591 (N_9591,N_9431,N_9432);
nor U9592 (N_9592,N_9401,N_9412);
nand U9593 (N_9593,N_9427,N_9467);
or U9594 (N_9594,N_9411,N_9453);
xor U9595 (N_9595,N_9443,N_9445);
nand U9596 (N_9596,N_9491,N_9438);
or U9597 (N_9597,N_9480,N_9405);
and U9598 (N_9598,N_9412,N_9426);
and U9599 (N_9599,N_9494,N_9483);
and U9600 (N_9600,N_9577,N_9581);
or U9601 (N_9601,N_9549,N_9561);
xnor U9602 (N_9602,N_9503,N_9571);
or U9603 (N_9603,N_9511,N_9584);
and U9604 (N_9604,N_9589,N_9563);
xnor U9605 (N_9605,N_9539,N_9556);
nand U9606 (N_9606,N_9505,N_9543);
and U9607 (N_9607,N_9575,N_9565);
and U9608 (N_9608,N_9597,N_9591);
nand U9609 (N_9609,N_9529,N_9533);
nor U9610 (N_9610,N_9554,N_9586);
nor U9611 (N_9611,N_9524,N_9528);
or U9612 (N_9612,N_9509,N_9596);
nand U9613 (N_9613,N_9538,N_9526);
nor U9614 (N_9614,N_9535,N_9558);
or U9615 (N_9615,N_9576,N_9568);
or U9616 (N_9616,N_9592,N_9544);
nor U9617 (N_9617,N_9569,N_9521);
xnor U9618 (N_9618,N_9574,N_9518);
xor U9619 (N_9619,N_9519,N_9507);
nand U9620 (N_9620,N_9585,N_9599);
or U9621 (N_9621,N_9560,N_9502);
and U9622 (N_9622,N_9501,N_9536);
or U9623 (N_9623,N_9525,N_9555);
and U9624 (N_9624,N_9531,N_9588);
or U9625 (N_9625,N_9517,N_9508);
nand U9626 (N_9626,N_9580,N_9530);
and U9627 (N_9627,N_9520,N_9593);
nand U9628 (N_9628,N_9567,N_9594);
or U9629 (N_9629,N_9513,N_9595);
or U9630 (N_9630,N_9504,N_9514);
nor U9631 (N_9631,N_9583,N_9510);
or U9632 (N_9632,N_9515,N_9562);
and U9633 (N_9633,N_9500,N_9522);
or U9634 (N_9634,N_9534,N_9598);
and U9635 (N_9635,N_9506,N_9537);
nor U9636 (N_9636,N_9559,N_9590);
nand U9637 (N_9637,N_9572,N_9578);
nand U9638 (N_9638,N_9542,N_9546);
nand U9639 (N_9639,N_9527,N_9516);
nand U9640 (N_9640,N_9545,N_9564);
nand U9641 (N_9641,N_9512,N_9548);
xnor U9642 (N_9642,N_9540,N_9550);
xor U9643 (N_9643,N_9541,N_9573);
and U9644 (N_9644,N_9566,N_9570);
or U9645 (N_9645,N_9532,N_9552);
nor U9646 (N_9646,N_9587,N_9553);
and U9647 (N_9647,N_9523,N_9551);
xor U9648 (N_9648,N_9557,N_9547);
and U9649 (N_9649,N_9582,N_9579);
or U9650 (N_9650,N_9545,N_9546);
and U9651 (N_9651,N_9581,N_9534);
xnor U9652 (N_9652,N_9515,N_9583);
and U9653 (N_9653,N_9523,N_9511);
nand U9654 (N_9654,N_9507,N_9516);
or U9655 (N_9655,N_9593,N_9540);
and U9656 (N_9656,N_9583,N_9593);
or U9657 (N_9657,N_9525,N_9536);
or U9658 (N_9658,N_9506,N_9587);
and U9659 (N_9659,N_9598,N_9589);
nand U9660 (N_9660,N_9542,N_9573);
and U9661 (N_9661,N_9574,N_9512);
or U9662 (N_9662,N_9573,N_9505);
and U9663 (N_9663,N_9564,N_9571);
and U9664 (N_9664,N_9516,N_9538);
or U9665 (N_9665,N_9514,N_9566);
and U9666 (N_9666,N_9583,N_9572);
nor U9667 (N_9667,N_9563,N_9540);
or U9668 (N_9668,N_9501,N_9544);
nand U9669 (N_9669,N_9543,N_9582);
or U9670 (N_9670,N_9569,N_9502);
nor U9671 (N_9671,N_9597,N_9511);
nor U9672 (N_9672,N_9530,N_9579);
and U9673 (N_9673,N_9558,N_9508);
or U9674 (N_9674,N_9513,N_9524);
nor U9675 (N_9675,N_9532,N_9592);
xnor U9676 (N_9676,N_9581,N_9585);
xor U9677 (N_9677,N_9541,N_9562);
nor U9678 (N_9678,N_9516,N_9588);
and U9679 (N_9679,N_9538,N_9568);
nor U9680 (N_9680,N_9541,N_9549);
and U9681 (N_9681,N_9516,N_9501);
nand U9682 (N_9682,N_9526,N_9575);
or U9683 (N_9683,N_9533,N_9595);
nand U9684 (N_9684,N_9576,N_9537);
or U9685 (N_9685,N_9508,N_9565);
nor U9686 (N_9686,N_9576,N_9546);
or U9687 (N_9687,N_9524,N_9539);
and U9688 (N_9688,N_9593,N_9528);
nor U9689 (N_9689,N_9543,N_9525);
nand U9690 (N_9690,N_9520,N_9516);
xor U9691 (N_9691,N_9581,N_9599);
nor U9692 (N_9692,N_9527,N_9557);
or U9693 (N_9693,N_9584,N_9503);
and U9694 (N_9694,N_9519,N_9505);
nor U9695 (N_9695,N_9585,N_9574);
and U9696 (N_9696,N_9500,N_9583);
nor U9697 (N_9697,N_9563,N_9565);
nor U9698 (N_9698,N_9509,N_9518);
and U9699 (N_9699,N_9573,N_9546);
nand U9700 (N_9700,N_9632,N_9680);
or U9701 (N_9701,N_9633,N_9676);
and U9702 (N_9702,N_9641,N_9609);
xor U9703 (N_9703,N_9616,N_9677);
nand U9704 (N_9704,N_9697,N_9652);
and U9705 (N_9705,N_9624,N_9653);
and U9706 (N_9706,N_9682,N_9671);
and U9707 (N_9707,N_9626,N_9638);
and U9708 (N_9708,N_9619,N_9651);
or U9709 (N_9709,N_9693,N_9613);
xor U9710 (N_9710,N_9644,N_9611);
or U9711 (N_9711,N_9690,N_9650);
or U9712 (N_9712,N_9674,N_9669);
nand U9713 (N_9713,N_9637,N_9666);
or U9714 (N_9714,N_9691,N_9608);
xor U9715 (N_9715,N_9678,N_9630);
xor U9716 (N_9716,N_9655,N_9687);
and U9717 (N_9717,N_9695,N_9657);
and U9718 (N_9718,N_9664,N_9647);
nor U9719 (N_9719,N_9640,N_9618);
and U9720 (N_9720,N_9658,N_9600);
nor U9721 (N_9721,N_9623,N_9689);
xnor U9722 (N_9722,N_9615,N_9659);
and U9723 (N_9723,N_9639,N_9667);
and U9724 (N_9724,N_9696,N_9614);
nor U9725 (N_9725,N_9662,N_9698);
nor U9726 (N_9726,N_9699,N_9636);
and U9727 (N_9727,N_9629,N_9681);
xnor U9728 (N_9728,N_9648,N_9603);
nand U9729 (N_9729,N_9621,N_9625);
and U9730 (N_9730,N_9688,N_9654);
nand U9731 (N_9731,N_9610,N_9602);
xnor U9732 (N_9732,N_9617,N_9679);
nor U9733 (N_9733,N_9606,N_9627);
nor U9734 (N_9734,N_9612,N_9649);
nand U9735 (N_9735,N_9694,N_9670);
nand U9736 (N_9736,N_9656,N_9661);
or U9737 (N_9737,N_9685,N_9665);
and U9738 (N_9738,N_9634,N_9628);
and U9739 (N_9739,N_9601,N_9672);
or U9740 (N_9740,N_9605,N_9673);
nor U9741 (N_9741,N_9631,N_9604);
or U9742 (N_9742,N_9643,N_9684);
nor U9743 (N_9743,N_9683,N_9607);
and U9744 (N_9744,N_9622,N_9642);
nand U9745 (N_9745,N_9692,N_9645);
nor U9746 (N_9746,N_9668,N_9635);
xnor U9747 (N_9747,N_9660,N_9686);
nand U9748 (N_9748,N_9675,N_9620);
xor U9749 (N_9749,N_9663,N_9646);
nand U9750 (N_9750,N_9648,N_9630);
nor U9751 (N_9751,N_9646,N_9618);
nor U9752 (N_9752,N_9651,N_9666);
and U9753 (N_9753,N_9630,N_9619);
nor U9754 (N_9754,N_9659,N_9626);
or U9755 (N_9755,N_9619,N_9610);
or U9756 (N_9756,N_9616,N_9696);
or U9757 (N_9757,N_9607,N_9637);
and U9758 (N_9758,N_9639,N_9613);
or U9759 (N_9759,N_9653,N_9656);
or U9760 (N_9760,N_9662,N_9692);
or U9761 (N_9761,N_9684,N_9631);
and U9762 (N_9762,N_9673,N_9684);
nor U9763 (N_9763,N_9691,N_9633);
or U9764 (N_9764,N_9693,N_9622);
or U9765 (N_9765,N_9673,N_9652);
and U9766 (N_9766,N_9680,N_9659);
and U9767 (N_9767,N_9625,N_9644);
nor U9768 (N_9768,N_9608,N_9640);
and U9769 (N_9769,N_9661,N_9673);
nor U9770 (N_9770,N_9677,N_9690);
or U9771 (N_9771,N_9639,N_9661);
or U9772 (N_9772,N_9614,N_9656);
xor U9773 (N_9773,N_9677,N_9644);
nor U9774 (N_9774,N_9670,N_9623);
or U9775 (N_9775,N_9685,N_9650);
and U9776 (N_9776,N_9675,N_9680);
or U9777 (N_9777,N_9612,N_9697);
and U9778 (N_9778,N_9619,N_9668);
nand U9779 (N_9779,N_9684,N_9652);
nor U9780 (N_9780,N_9641,N_9684);
and U9781 (N_9781,N_9612,N_9643);
or U9782 (N_9782,N_9601,N_9632);
or U9783 (N_9783,N_9659,N_9625);
and U9784 (N_9784,N_9621,N_9634);
and U9785 (N_9785,N_9679,N_9699);
or U9786 (N_9786,N_9618,N_9665);
and U9787 (N_9787,N_9618,N_9607);
nand U9788 (N_9788,N_9669,N_9694);
or U9789 (N_9789,N_9625,N_9654);
nor U9790 (N_9790,N_9637,N_9651);
and U9791 (N_9791,N_9619,N_9638);
and U9792 (N_9792,N_9677,N_9610);
nor U9793 (N_9793,N_9620,N_9689);
or U9794 (N_9794,N_9607,N_9687);
or U9795 (N_9795,N_9654,N_9636);
nor U9796 (N_9796,N_9651,N_9645);
and U9797 (N_9797,N_9698,N_9667);
xnor U9798 (N_9798,N_9685,N_9666);
nand U9799 (N_9799,N_9646,N_9656);
and U9800 (N_9800,N_9703,N_9750);
nor U9801 (N_9801,N_9732,N_9709);
xor U9802 (N_9802,N_9792,N_9738);
nand U9803 (N_9803,N_9753,N_9705);
and U9804 (N_9804,N_9779,N_9713);
and U9805 (N_9805,N_9735,N_9780);
xnor U9806 (N_9806,N_9736,N_9770);
nand U9807 (N_9807,N_9724,N_9771);
nand U9808 (N_9808,N_9783,N_9701);
or U9809 (N_9809,N_9765,N_9720);
nor U9810 (N_9810,N_9725,N_9747);
and U9811 (N_9811,N_9733,N_9723);
nand U9812 (N_9812,N_9749,N_9790);
nand U9813 (N_9813,N_9798,N_9757);
or U9814 (N_9814,N_9734,N_9730);
and U9815 (N_9815,N_9767,N_9768);
and U9816 (N_9816,N_9791,N_9789);
or U9817 (N_9817,N_9739,N_9785);
nor U9818 (N_9818,N_9706,N_9773);
nor U9819 (N_9819,N_9799,N_9710);
nand U9820 (N_9820,N_9762,N_9766);
nand U9821 (N_9821,N_9782,N_9742);
nand U9822 (N_9822,N_9774,N_9743);
nand U9823 (N_9823,N_9752,N_9775);
nand U9824 (N_9824,N_9788,N_9746);
nand U9825 (N_9825,N_9796,N_9711);
nor U9826 (N_9826,N_9721,N_9756);
nand U9827 (N_9827,N_9712,N_9714);
or U9828 (N_9828,N_9741,N_9716);
nor U9829 (N_9829,N_9776,N_9744);
xor U9830 (N_9830,N_9760,N_9795);
nor U9831 (N_9831,N_9751,N_9764);
or U9832 (N_9832,N_9763,N_9740);
nand U9833 (N_9833,N_9731,N_9726);
and U9834 (N_9834,N_9700,N_9759);
nor U9835 (N_9835,N_9781,N_9708);
nor U9836 (N_9836,N_9772,N_9797);
nand U9837 (N_9837,N_9793,N_9715);
nor U9838 (N_9838,N_9728,N_9707);
or U9839 (N_9839,N_9784,N_9787);
nor U9840 (N_9840,N_9722,N_9704);
or U9841 (N_9841,N_9737,N_9786);
nor U9842 (N_9842,N_9777,N_9769);
nor U9843 (N_9843,N_9745,N_9761);
or U9844 (N_9844,N_9717,N_9748);
or U9845 (N_9845,N_9755,N_9794);
or U9846 (N_9846,N_9778,N_9729);
and U9847 (N_9847,N_9719,N_9718);
and U9848 (N_9848,N_9754,N_9702);
xor U9849 (N_9849,N_9758,N_9727);
nand U9850 (N_9850,N_9765,N_9724);
nand U9851 (N_9851,N_9763,N_9733);
or U9852 (N_9852,N_9759,N_9707);
and U9853 (N_9853,N_9733,N_9765);
nand U9854 (N_9854,N_9778,N_9754);
nand U9855 (N_9855,N_9740,N_9788);
and U9856 (N_9856,N_9791,N_9762);
and U9857 (N_9857,N_9704,N_9706);
and U9858 (N_9858,N_9755,N_9742);
and U9859 (N_9859,N_9774,N_9790);
or U9860 (N_9860,N_9700,N_9701);
or U9861 (N_9861,N_9748,N_9769);
and U9862 (N_9862,N_9716,N_9730);
xnor U9863 (N_9863,N_9795,N_9762);
and U9864 (N_9864,N_9766,N_9780);
nor U9865 (N_9865,N_9784,N_9709);
or U9866 (N_9866,N_9704,N_9719);
and U9867 (N_9867,N_9780,N_9733);
or U9868 (N_9868,N_9758,N_9779);
or U9869 (N_9869,N_9797,N_9784);
or U9870 (N_9870,N_9714,N_9733);
or U9871 (N_9871,N_9780,N_9723);
and U9872 (N_9872,N_9782,N_9718);
and U9873 (N_9873,N_9776,N_9796);
nand U9874 (N_9874,N_9723,N_9702);
nor U9875 (N_9875,N_9793,N_9762);
or U9876 (N_9876,N_9766,N_9724);
or U9877 (N_9877,N_9717,N_9781);
nand U9878 (N_9878,N_9757,N_9716);
nand U9879 (N_9879,N_9737,N_9717);
nand U9880 (N_9880,N_9798,N_9720);
or U9881 (N_9881,N_9735,N_9701);
nand U9882 (N_9882,N_9760,N_9719);
nand U9883 (N_9883,N_9772,N_9724);
nor U9884 (N_9884,N_9768,N_9758);
nor U9885 (N_9885,N_9732,N_9723);
nor U9886 (N_9886,N_9761,N_9758);
nand U9887 (N_9887,N_9758,N_9772);
and U9888 (N_9888,N_9736,N_9717);
nand U9889 (N_9889,N_9735,N_9765);
and U9890 (N_9890,N_9760,N_9700);
nor U9891 (N_9891,N_9723,N_9710);
and U9892 (N_9892,N_9770,N_9726);
and U9893 (N_9893,N_9724,N_9726);
or U9894 (N_9894,N_9757,N_9713);
or U9895 (N_9895,N_9713,N_9705);
nor U9896 (N_9896,N_9740,N_9739);
and U9897 (N_9897,N_9741,N_9783);
xnor U9898 (N_9898,N_9711,N_9732);
nor U9899 (N_9899,N_9767,N_9700);
and U9900 (N_9900,N_9824,N_9853);
nand U9901 (N_9901,N_9877,N_9876);
and U9902 (N_9902,N_9839,N_9891);
nand U9903 (N_9903,N_9869,N_9864);
and U9904 (N_9904,N_9832,N_9859);
or U9905 (N_9905,N_9852,N_9844);
nand U9906 (N_9906,N_9802,N_9871);
and U9907 (N_9907,N_9803,N_9880);
xnor U9908 (N_9908,N_9872,N_9895);
and U9909 (N_9909,N_9834,N_9886);
and U9910 (N_9910,N_9833,N_9870);
nor U9911 (N_9911,N_9861,N_9807);
and U9912 (N_9912,N_9890,N_9816);
and U9913 (N_9913,N_9821,N_9849);
and U9914 (N_9914,N_9836,N_9801);
or U9915 (N_9915,N_9850,N_9815);
or U9916 (N_9916,N_9881,N_9843);
nand U9917 (N_9917,N_9885,N_9812);
nor U9918 (N_9918,N_9813,N_9896);
nand U9919 (N_9919,N_9826,N_9867);
or U9920 (N_9920,N_9889,N_9811);
and U9921 (N_9921,N_9800,N_9884);
or U9922 (N_9922,N_9874,N_9804);
nand U9923 (N_9923,N_9809,N_9855);
nand U9924 (N_9924,N_9847,N_9810);
nand U9925 (N_9925,N_9860,N_9888);
nor U9926 (N_9926,N_9848,N_9825);
and U9927 (N_9927,N_9878,N_9842);
nor U9928 (N_9928,N_9898,N_9806);
nor U9929 (N_9929,N_9840,N_9831);
and U9930 (N_9930,N_9835,N_9893);
and U9931 (N_9931,N_9823,N_9883);
and U9932 (N_9932,N_9838,N_9814);
and U9933 (N_9933,N_9866,N_9830);
or U9934 (N_9934,N_9873,N_9865);
nand U9935 (N_9935,N_9882,N_9856);
nand U9936 (N_9936,N_9827,N_9841);
nand U9937 (N_9937,N_9858,N_9805);
and U9938 (N_9938,N_9868,N_9845);
nand U9939 (N_9939,N_9808,N_9829);
and U9940 (N_9940,N_9879,N_9819);
and U9941 (N_9941,N_9846,N_9851);
nor U9942 (N_9942,N_9892,N_9828);
and U9943 (N_9943,N_9822,N_9820);
nand U9944 (N_9944,N_9857,N_9875);
or U9945 (N_9945,N_9837,N_9887);
and U9946 (N_9946,N_9854,N_9894);
nor U9947 (N_9947,N_9818,N_9897);
or U9948 (N_9948,N_9863,N_9862);
nand U9949 (N_9949,N_9817,N_9899);
nand U9950 (N_9950,N_9882,N_9880);
or U9951 (N_9951,N_9876,N_9868);
nor U9952 (N_9952,N_9820,N_9846);
or U9953 (N_9953,N_9875,N_9829);
and U9954 (N_9954,N_9818,N_9875);
xor U9955 (N_9955,N_9863,N_9846);
or U9956 (N_9956,N_9800,N_9803);
nor U9957 (N_9957,N_9811,N_9882);
nor U9958 (N_9958,N_9815,N_9836);
and U9959 (N_9959,N_9874,N_9893);
nand U9960 (N_9960,N_9853,N_9827);
and U9961 (N_9961,N_9852,N_9874);
and U9962 (N_9962,N_9874,N_9828);
nor U9963 (N_9963,N_9807,N_9835);
nand U9964 (N_9964,N_9867,N_9888);
or U9965 (N_9965,N_9848,N_9837);
nand U9966 (N_9966,N_9851,N_9819);
nor U9967 (N_9967,N_9862,N_9845);
and U9968 (N_9968,N_9800,N_9810);
nand U9969 (N_9969,N_9899,N_9819);
nor U9970 (N_9970,N_9814,N_9851);
xor U9971 (N_9971,N_9865,N_9856);
xor U9972 (N_9972,N_9884,N_9889);
or U9973 (N_9973,N_9800,N_9841);
nor U9974 (N_9974,N_9825,N_9875);
and U9975 (N_9975,N_9860,N_9824);
nor U9976 (N_9976,N_9856,N_9862);
nand U9977 (N_9977,N_9859,N_9891);
nand U9978 (N_9978,N_9804,N_9817);
or U9979 (N_9979,N_9819,N_9866);
nand U9980 (N_9980,N_9833,N_9830);
and U9981 (N_9981,N_9845,N_9805);
or U9982 (N_9982,N_9847,N_9891);
nor U9983 (N_9983,N_9837,N_9803);
or U9984 (N_9984,N_9839,N_9861);
nor U9985 (N_9985,N_9837,N_9826);
xnor U9986 (N_9986,N_9843,N_9816);
xnor U9987 (N_9987,N_9854,N_9824);
nor U9988 (N_9988,N_9820,N_9862);
or U9989 (N_9989,N_9811,N_9807);
and U9990 (N_9990,N_9801,N_9880);
nor U9991 (N_9991,N_9840,N_9839);
and U9992 (N_9992,N_9883,N_9824);
and U9993 (N_9993,N_9821,N_9891);
or U9994 (N_9994,N_9838,N_9815);
nand U9995 (N_9995,N_9877,N_9881);
or U9996 (N_9996,N_9804,N_9884);
nand U9997 (N_9997,N_9830,N_9870);
nor U9998 (N_9998,N_9804,N_9848);
or U9999 (N_9999,N_9800,N_9813);
nor UO_0 (O_0,N_9907,N_9909);
and UO_1 (O_1,N_9906,N_9987);
nand UO_2 (O_2,N_9939,N_9949);
and UO_3 (O_3,N_9913,N_9920);
nand UO_4 (O_4,N_9914,N_9997);
nand UO_5 (O_5,N_9960,N_9911);
or UO_6 (O_6,N_9928,N_9931);
nor UO_7 (O_7,N_9919,N_9980);
nand UO_8 (O_8,N_9902,N_9982);
xnor UO_9 (O_9,N_9983,N_9985);
or UO_10 (O_10,N_9979,N_9972);
nor UO_11 (O_11,N_9961,N_9926);
nand UO_12 (O_12,N_9970,N_9901);
nor UO_13 (O_13,N_9932,N_9973);
nand UO_14 (O_14,N_9971,N_9918);
nor UO_15 (O_15,N_9923,N_9936);
and UO_16 (O_16,N_9993,N_9946);
or UO_17 (O_17,N_9999,N_9950);
nor UO_18 (O_18,N_9976,N_9903);
nand UO_19 (O_19,N_9967,N_9958);
and UO_20 (O_20,N_9977,N_9910);
or UO_21 (O_21,N_9988,N_9996);
and UO_22 (O_22,N_9934,N_9917);
nor UO_23 (O_23,N_9915,N_9943);
nor UO_24 (O_24,N_9998,N_9992);
or UO_25 (O_25,N_9944,N_9900);
and UO_26 (O_26,N_9925,N_9904);
and UO_27 (O_27,N_9952,N_9912);
and UO_28 (O_28,N_9975,N_9922);
and UO_29 (O_29,N_9954,N_9966);
nand UO_30 (O_30,N_9984,N_9916);
nand UO_31 (O_31,N_9974,N_9968);
xnor UO_32 (O_32,N_9930,N_9959);
and UO_33 (O_33,N_9986,N_9964);
or UO_34 (O_34,N_9963,N_9935);
or UO_35 (O_35,N_9991,N_9929);
or UO_36 (O_36,N_9981,N_9941);
or UO_37 (O_37,N_9948,N_9933);
or UO_38 (O_38,N_9989,N_9955);
or UO_39 (O_39,N_9940,N_9905);
and UO_40 (O_40,N_9995,N_9945);
nor UO_41 (O_41,N_9942,N_9953);
nand UO_42 (O_42,N_9908,N_9969);
or UO_43 (O_43,N_9951,N_9921);
or UO_44 (O_44,N_9947,N_9994);
nand UO_45 (O_45,N_9924,N_9957);
and UO_46 (O_46,N_9927,N_9990);
nor UO_47 (O_47,N_9978,N_9938);
nor UO_48 (O_48,N_9962,N_9965);
and UO_49 (O_49,N_9937,N_9956);
nand UO_50 (O_50,N_9928,N_9930);
nand UO_51 (O_51,N_9945,N_9951);
xor UO_52 (O_52,N_9965,N_9900);
nand UO_53 (O_53,N_9915,N_9974);
xor UO_54 (O_54,N_9970,N_9979);
nor UO_55 (O_55,N_9963,N_9922);
or UO_56 (O_56,N_9983,N_9959);
and UO_57 (O_57,N_9951,N_9986);
nor UO_58 (O_58,N_9909,N_9951);
nand UO_59 (O_59,N_9907,N_9966);
and UO_60 (O_60,N_9957,N_9964);
nor UO_61 (O_61,N_9931,N_9991);
nor UO_62 (O_62,N_9952,N_9921);
and UO_63 (O_63,N_9994,N_9913);
and UO_64 (O_64,N_9986,N_9930);
nand UO_65 (O_65,N_9991,N_9926);
or UO_66 (O_66,N_9956,N_9930);
nand UO_67 (O_67,N_9978,N_9958);
or UO_68 (O_68,N_9978,N_9973);
nor UO_69 (O_69,N_9922,N_9964);
nor UO_70 (O_70,N_9939,N_9916);
nor UO_71 (O_71,N_9972,N_9970);
and UO_72 (O_72,N_9930,N_9987);
nand UO_73 (O_73,N_9954,N_9960);
and UO_74 (O_74,N_9987,N_9941);
nor UO_75 (O_75,N_9986,N_9974);
or UO_76 (O_76,N_9933,N_9926);
or UO_77 (O_77,N_9985,N_9960);
nand UO_78 (O_78,N_9955,N_9995);
nand UO_79 (O_79,N_9927,N_9987);
and UO_80 (O_80,N_9987,N_9911);
and UO_81 (O_81,N_9976,N_9970);
and UO_82 (O_82,N_9980,N_9992);
or UO_83 (O_83,N_9984,N_9913);
or UO_84 (O_84,N_9960,N_9992);
nor UO_85 (O_85,N_9992,N_9918);
and UO_86 (O_86,N_9916,N_9901);
xnor UO_87 (O_87,N_9925,N_9935);
nor UO_88 (O_88,N_9934,N_9971);
and UO_89 (O_89,N_9973,N_9930);
nand UO_90 (O_90,N_9955,N_9992);
nand UO_91 (O_91,N_9959,N_9995);
xnor UO_92 (O_92,N_9993,N_9943);
and UO_93 (O_93,N_9971,N_9943);
and UO_94 (O_94,N_9927,N_9986);
nand UO_95 (O_95,N_9998,N_9945);
nand UO_96 (O_96,N_9922,N_9966);
nor UO_97 (O_97,N_9908,N_9973);
nand UO_98 (O_98,N_9903,N_9926);
or UO_99 (O_99,N_9971,N_9977);
and UO_100 (O_100,N_9968,N_9939);
nor UO_101 (O_101,N_9964,N_9999);
or UO_102 (O_102,N_9910,N_9912);
and UO_103 (O_103,N_9903,N_9986);
nor UO_104 (O_104,N_9918,N_9974);
nor UO_105 (O_105,N_9987,N_9986);
nor UO_106 (O_106,N_9974,N_9929);
and UO_107 (O_107,N_9965,N_9951);
or UO_108 (O_108,N_9911,N_9980);
or UO_109 (O_109,N_9986,N_9902);
or UO_110 (O_110,N_9925,N_9960);
nand UO_111 (O_111,N_9907,N_9946);
nand UO_112 (O_112,N_9925,N_9982);
nand UO_113 (O_113,N_9945,N_9931);
nand UO_114 (O_114,N_9993,N_9986);
nor UO_115 (O_115,N_9955,N_9919);
nand UO_116 (O_116,N_9928,N_9941);
xnor UO_117 (O_117,N_9958,N_9975);
or UO_118 (O_118,N_9917,N_9914);
nor UO_119 (O_119,N_9914,N_9981);
nor UO_120 (O_120,N_9924,N_9949);
and UO_121 (O_121,N_9989,N_9915);
and UO_122 (O_122,N_9969,N_9900);
and UO_123 (O_123,N_9940,N_9913);
or UO_124 (O_124,N_9926,N_9998);
nand UO_125 (O_125,N_9950,N_9940);
and UO_126 (O_126,N_9981,N_9992);
and UO_127 (O_127,N_9941,N_9940);
nand UO_128 (O_128,N_9936,N_9967);
or UO_129 (O_129,N_9976,N_9994);
xnor UO_130 (O_130,N_9926,N_9906);
nand UO_131 (O_131,N_9997,N_9944);
nand UO_132 (O_132,N_9921,N_9986);
nand UO_133 (O_133,N_9942,N_9956);
nand UO_134 (O_134,N_9922,N_9941);
nor UO_135 (O_135,N_9982,N_9959);
xnor UO_136 (O_136,N_9929,N_9928);
and UO_137 (O_137,N_9909,N_9911);
or UO_138 (O_138,N_9967,N_9930);
and UO_139 (O_139,N_9913,N_9933);
nand UO_140 (O_140,N_9970,N_9962);
or UO_141 (O_141,N_9982,N_9927);
nand UO_142 (O_142,N_9902,N_9918);
nand UO_143 (O_143,N_9952,N_9907);
nand UO_144 (O_144,N_9900,N_9958);
nand UO_145 (O_145,N_9923,N_9986);
nor UO_146 (O_146,N_9979,N_9984);
nor UO_147 (O_147,N_9925,N_9955);
nand UO_148 (O_148,N_9933,N_9968);
or UO_149 (O_149,N_9992,N_9953);
nand UO_150 (O_150,N_9907,N_9979);
and UO_151 (O_151,N_9909,N_9953);
xor UO_152 (O_152,N_9962,N_9920);
nand UO_153 (O_153,N_9905,N_9997);
or UO_154 (O_154,N_9967,N_9931);
nand UO_155 (O_155,N_9947,N_9960);
nand UO_156 (O_156,N_9950,N_9995);
nor UO_157 (O_157,N_9904,N_9908);
or UO_158 (O_158,N_9922,N_9925);
or UO_159 (O_159,N_9904,N_9974);
nor UO_160 (O_160,N_9977,N_9985);
or UO_161 (O_161,N_9952,N_9909);
and UO_162 (O_162,N_9910,N_9971);
or UO_163 (O_163,N_9934,N_9923);
xnor UO_164 (O_164,N_9946,N_9987);
nand UO_165 (O_165,N_9995,N_9992);
and UO_166 (O_166,N_9945,N_9947);
nand UO_167 (O_167,N_9914,N_9930);
nor UO_168 (O_168,N_9936,N_9926);
nor UO_169 (O_169,N_9981,N_9996);
nand UO_170 (O_170,N_9985,N_9904);
nand UO_171 (O_171,N_9972,N_9910);
nor UO_172 (O_172,N_9954,N_9922);
or UO_173 (O_173,N_9933,N_9987);
nor UO_174 (O_174,N_9967,N_9922);
and UO_175 (O_175,N_9924,N_9993);
nand UO_176 (O_176,N_9948,N_9968);
and UO_177 (O_177,N_9960,N_9968);
and UO_178 (O_178,N_9976,N_9946);
nand UO_179 (O_179,N_9945,N_9952);
nor UO_180 (O_180,N_9999,N_9924);
nand UO_181 (O_181,N_9948,N_9991);
nand UO_182 (O_182,N_9983,N_9971);
nor UO_183 (O_183,N_9901,N_9968);
nand UO_184 (O_184,N_9963,N_9912);
or UO_185 (O_185,N_9974,N_9996);
and UO_186 (O_186,N_9934,N_9910);
and UO_187 (O_187,N_9964,N_9981);
nand UO_188 (O_188,N_9944,N_9994);
nor UO_189 (O_189,N_9921,N_9964);
nor UO_190 (O_190,N_9962,N_9972);
and UO_191 (O_191,N_9963,N_9960);
xnor UO_192 (O_192,N_9972,N_9974);
nor UO_193 (O_193,N_9906,N_9967);
or UO_194 (O_194,N_9996,N_9944);
xor UO_195 (O_195,N_9909,N_9943);
and UO_196 (O_196,N_9944,N_9937);
and UO_197 (O_197,N_9994,N_9989);
or UO_198 (O_198,N_9950,N_9979);
nor UO_199 (O_199,N_9917,N_9907);
or UO_200 (O_200,N_9915,N_9970);
or UO_201 (O_201,N_9934,N_9979);
and UO_202 (O_202,N_9999,N_9921);
and UO_203 (O_203,N_9962,N_9946);
xor UO_204 (O_204,N_9958,N_9999);
or UO_205 (O_205,N_9917,N_9943);
or UO_206 (O_206,N_9900,N_9952);
xnor UO_207 (O_207,N_9918,N_9910);
xnor UO_208 (O_208,N_9986,N_9958);
and UO_209 (O_209,N_9921,N_9994);
xor UO_210 (O_210,N_9907,N_9926);
nor UO_211 (O_211,N_9910,N_9950);
and UO_212 (O_212,N_9989,N_9924);
and UO_213 (O_213,N_9986,N_9968);
nor UO_214 (O_214,N_9998,N_9903);
nand UO_215 (O_215,N_9905,N_9951);
or UO_216 (O_216,N_9949,N_9985);
xor UO_217 (O_217,N_9912,N_9970);
nor UO_218 (O_218,N_9936,N_9916);
nand UO_219 (O_219,N_9912,N_9950);
xnor UO_220 (O_220,N_9923,N_9919);
nand UO_221 (O_221,N_9970,N_9999);
and UO_222 (O_222,N_9928,N_9939);
or UO_223 (O_223,N_9931,N_9922);
and UO_224 (O_224,N_9911,N_9950);
nor UO_225 (O_225,N_9953,N_9923);
nor UO_226 (O_226,N_9974,N_9931);
nor UO_227 (O_227,N_9985,N_9969);
and UO_228 (O_228,N_9942,N_9923);
nor UO_229 (O_229,N_9954,N_9973);
or UO_230 (O_230,N_9969,N_9914);
or UO_231 (O_231,N_9948,N_9931);
xor UO_232 (O_232,N_9956,N_9963);
nor UO_233 (O_233,N_9961,N_9907);
and UO_234 (O_234,N_9917,N_9958);
nor UO_235 (O_235,N_9928,N_9901);
and UO_236 (O_236,N_9979,N_9920);
and UO_237 (O_237,N_9931,N_9906);
nand UO_238 (O_238,N_9957,N_9958);
and UO_239 (O_239,N_9987,N_9956);
nand UO_240 (O_240,N_9912,N_9932);
or UO_241 (O_241,N_9988,N_9920);
nor UO_242 (O_242,N_9917,N_9906);
xor UO_243 (O_243,N_9991,N_9978);
or UO_244 (O_244,N_9948,N_9964);
and UO_245 (O_245,N_9977,N_9937);
nor UO_246 (O_246,N_9910,N_9941);
nand UO_247 (O_247,N_9960,N_9956);
or UO_248 (O_248,N_9935,N_9938);
nand UO_249 (O_249,N_9992,N_9999);
nor UO_250 (O_250,N_9920,N_9954);
nor UO_251 (O_251,N_9926,N_9912);
nor UO_252 (O_252,N_9964,N_9983);
xor UO_253 (O_253,N_9991,N_9985);
and UO_254 (O_254,N_9913,N_9976);
and UO_255 (O_255,N_9943,N_9905);
nor UO_256 (O_256,N_9948,N_9960);
nor UO_257 (O_257,N_9937,N_9986);
nor UO_258 (O_258,N_9920,N_9968);
xor UO_259 (O_259,N_9979,N_9942);
xnor UO_260 (O_260,N_9998,N_9985);
or UO_261 (O_261,N_9965,N_9961);
nor UO_262 (O_262,N_9992,N_9977);
nand UO_263 (O_263,N_9941,N_9948);
nor UO_264 (O_264,N_9951,N_9944);
or UO_265 (O_265,N_9981,N_9921);
nor UO_266 (O_266,N_9960,N_9976);
and UO_267 (O_267,N_9988,N_9946);
nor UO_268 (O_268,N_9952,N_9993);
nand UO_269 (O_269,N_9958,N_9904);
and UO_270 (O_270,N_9909,N_9960);
and UO_271 (O_271,N_9999,N_9930);
nor UO_272 (O_272,N_9940,N_9909);
or UO_273 (O_273,N_9931,N_9916);
nand UO_274 (O_274,N_9938,N_9961);
or UO_275 (O_275,N_9902,N_9919);
nand UO_276 (O_276,N_9937,N_9943);
and UO_277 (O_277,N_9941,N_9964);
nand UO_278 (O_278,N_9969,N_9978);
nor UO_279 (O_279,N_9994,N_9980);
or UO_280 (O_280,N_9975,N_9978);
and UO_281 (O_281,N_9989,N_9901);
nor UO_282 (O_282,N_9936,N_9947);
nor UO_283 (O_283,N_9976,N_9996);
or UO_284 (O_284,N_9908,N_9985);
nand UO_285 (O_285,N_9936,N_9998);
or UO_286 (O_286,N_9954,N_9914);
and UO_287 (O_287,N_9991,N_9909);
nand UO_288 (O_288,N_9917,N_9963);
nand UO_289 (O_289,N_9946,N_9960);
nor UO_290 (O_290,N_9933,N_9984);
or UO_291 (O_291,N_9999,N_9955);
nand UO_292 (O_292,N_9906,N_9960);
or UO_293 (O_293,N_9976,N_9925);
or UO_294 (O_294,N_9975,N_9934);
nor UO_295 (O_295,N_9927,N_9950);
nor UO_296 (O_296,N_9991,N_9927);
nor UO_297 (O_297,N_9930,N_9965);
xnor UO_298 (O_298,N_9902,N_9904);
xor UO_299 (O_299,N_9975,N_9945);
and UO_300 (O_300,N_9999,N_9982);
and UO_301 (O_301,N_9947,N_9935);
or UO_302 (O_302,N_9926,N_9951);
or UO_303 (O_303,N_9926,N_9935);
xnor UO_304 (O_304,N_9945,N_9913);
and UO_305 (O_305,N_9998,N_9927);
xnor UO_306 (O_306,N_9911,N_9989);
xnor UO_307 (O_307,N_9962,N_9942);
nand UO_308 (O_308,N_9950,N_9959);
nor UO_309 (O_309,N_9926,N_9989);
nand UO_310 (O_310,N_9922,N_9948);
nor UO_311 (O_311,N_9914,N_9922);
nand UO_312 (O_312,N_9969,N_9959);
nor UO_313 (O_313,N_9962,N_9973);
nand UO_314 (O_314,N_9968,N_9975);
xor UO_315 (O_315,N_9997,N_9930);
xnor UO_316 (O_316,N_9935,N_9957);
nor UO_317 (O_317,N_9999,N_9944);
nand UO_318 (O_318,N_9946,N_9912);
and UO_319 (O_319,N_9932,N_9985);
xor UO_320 (O_320,N_9948,N_9939);
nand UO_321 (O_321,N_9957,N_9928);
nor UO_322 (O_322,N_9980,N_9923);
and UO_323 (O_323,N_9900,N_9977);
xor UO_324 (O_324,N_9921,N_9989);
or UO_325 (O_325,N_9911,N_9964);
xnor UO_326 (O_326,N_9945,N_9976);
and UO_327 (O_327,N_9926,N_9955);
nand UO_328 (O_328,N_9903,N_9934);
nand UO_329 (O_329,N_9952,N_9927);
or UO_330 (O_330,N_9915,N_9931);
nor UO_331 (O_331,N_9958,N_9919);
nand UO_332 (O_332,N_9982,N_9961);
nor UO_333 (O_333,N_9913,N_9948);
xnor UO_334 (O_334,N_9904,N_9964);
nor UO_335 (O_335,N_9981,N_9976);
or UO_336 (O_336,N_9997,N_9909);
nand UO_337 (O_337,N_9982,N_9940);
xnor UO_338 (O_338,N_9973,N_9951);
nor UO_339 (O_339,N_9951,N_9995);
nand UO_340 (O_340,N_9999,N_9912);
or UO_341 (O_341,N_9968,N_9937);
and UO_342 (O_342,N_9934,N_9961);
nand UO_343 (O_343,N_9950,N_9918);
or UO_344 (O_344,N_9954,N_9989);
or UO_345 (O_345,N_9974,N_9982);
or UO_346 (O_346,N_9940,N_9983);
or UO_347 (O_347,N_9938,N_9995);
and UO_348 (O_348,N_9901,N_9948);
nand UO_349 (O_349,N_9950,N_9969);
or UO_350 (O_350,N_9961,N_9941);
nand UO_351 (O_351,N_9936,N_9991);
nor UO_352 (O_352,N_9901,N_9965);
and UO_353 (O_353,N_9948,N_9909);
or UO_354 (O_354,N_9905,N_9922);
or UO_355 (O_355,N_9911,N_9934);
and UO_356 (O_356,N_9902,N_9954);
or UO_357 (O_357,N_9939,N_9935);
or UO_358 (O_358,N_9993,N_9940);
nor UO_359 (O_359,N_9996,N_9908);
xor UO_360 (O_360,N_9916,N_9983);
nor UO_361 (O_361,N_9945,N_9966);
or UO_362 (O_362,N_9907,N_9991);
nor UO_363 (O_363,N_9977,N_9939);
nand UO_364 (O_364,N_9994,N_9910);
nand UO_365 (O_365,N_9977,N_9962);
and UO_366 (O_366,N_9904,N_9930);
or UO_367 (O_367,N_9953,N_9915);
or UO_368 (O_368,N_9982,N_9930);
xnor UO_369 (O_369,N_9936,N_9978);
and UO_370 (O_370,N_9945,N_9967);
xnor UO_371 (O_371,N_9907,N_9924);
or UO_372 (O_372,N_9962,N_9950);
nor UO_373 (O_373,N_9916,N_9977);
nor UO_374 (O_374,N_9916,N_9975);
or UO_375 (O_375,N_9911,N_9988);
nand UO_376 (O_376,N_9907,N_9999);
nand UO_377 (O_377,N_9960,N_9934);
or UO_378 (O_378,N_9949,N_9933);
and UO_379 (O_379,N_9920,N_9942);
or UO_380 (O_380,N_9929,N_9906);
xnor UO_381 (O_381,N_9939,N_9995);
and UO_382 (O_382,N_9972,N_9906);
and UO_383 (O_383,N_9998,N_9972);
nor UO_384 (O_384,N_9963,N_9950);
or UO_385 (O_385,N_9974,N_9940);
nor UO_386 (O_386,N_9945,N_9922);
nor UO_387 (O_387,N_9954,N_9987);
nor UO_388 (O_388,N_9947,N_9978);
nor UO_389 (O_389,N_9931,N_9935);
nor UO_390 (O_390,N_9921,N_9963);
and UO_391 (O_391,N_9956,N_9943);
or UO_392 (O_392,N_9904,N_9959);
or UO_393 (O_393,N_9910,N_9939);
xnor UO_394 (O_394,N_9979,N_9933);
nor UO_395 (O_395,N_9917,N_9983);
or UO_396 (O_396,N_9949,N_9913);
and UO_397 (O_397,N_9970,N_9973);
or UO_398 (O_398,N_9908,N_9940);
nor UO_399 (O_399,N_9952,N_9953);
nor UO_400 (O_400,N_9932,N_9937);
and UO_401 (O_401,N_9964,N_9976);
xnor UO_402 (O_402,N_9912,N_9968);
xnor UO_403 (O_403,N_9950,N_9987);
nor UO_404 (O_404,N_9975,N_9971);
or UO_405 (O_405,N_9921,N_9954);
or UO_406 (O_406,N_9970,N_9993);
or UO_407 (O_407,N_9997,N_9906);
nand UO_408 (O_408,N_9912,N_9956);
or UO_409 (O_409,N_9913,N_9961);
or UO_410 (O_410,N_9934,N_9900);
nor UO_411 (O_411,N_9913,N_9978);
nor UO_412 (O_412,N_9962,N_9985);
and UO_413 (O_413,N_9924,N_9934);
nand UO_414 (O_414,N_9985,N_9975);
nor UO_415 (O_415,N_9994,N_9968);
and UO_416 (O_416,N_9958,N_9918);
xor UO_417 (O_417,N_9914,N_9973);
and UO_418 (O_418,N_9935,N_9980);
nor UO_419 (O_419,N_9963,N_9939);
or UO_420 (O_420,N_9978,N_9993);
or UO_421 (O_421,N_9922,N_9965);
xnor UO_422 (O_422,N_9964,N_9905);
nor UO_423 (O_423,N_9929,N_9923);
xnor UO_424 (O_424,N_9990,N_9926);
xor UO_425 (O_425,N_9907,N_9932);
nand UO_426 (O_426,N_9957,N_9920);
and UO_427 (O_427,N_9925,N_9937);
nand UO_428 (O_428,N_9955,N_9903);
xnor UO_429 (O_429,N_9921,N_9960);
nand UO_430 (O_430,N_9932,N_9930);
nor UO_431 (O_431,N_9988,N_9934);
and UO_432 (O_432,N_9903,N_9919);
nor UO_433 (O_433,N_9977,N_9954);
nand UO_434 (O_434,N_9910,N_9956);
and UO_435 (O_435,N_9978,N_9967);
or UO_436 (O_436,N_9987,N_9945);
or UO_437 (O_437,N_9979,N_9945);
nand UO_438 (O_438,N_9937,N_9929);
or UO_439 (O_439,N_9939,N_9969);
nand UO_440 (O_440,N_9979,N_9978);
nand UO_441 (O_441,N_9966,N_9932);
nor UO_442 (O_442,N_9952,N_9995);
and UO_443 (O_443,N_9935,N_9978);
and UO_444 (O_444,N_9953,N_9914);
and UO_445 (O_445,N_9915,N_9944);
and UO_446 (O_446,N_9993,N_9921);
or UO_447 (O_447,N_9967,N_9980);
or UO_448 (O_448,N_9901,N_9994);
and UO_449 (O_449,N_9977,N_9911);
and UO_450 (O_450,N_9916,N_9962);
nor UO_451 (O_451,N_9973,N_9956);
nand UO_452 (O_452,N_9996,N_9921);
nand UO_453 (O_453,N_9957,N_9905);
nor UO_454 (O_454,N_9991,N_9910);
nor UO_455 (O_455,N_9942,N_9917);
or UO_456 (O_456,N_9974,N_9910);
and UO_457 (O_457,N_9987,N_9959);
or UO_458 (O_458,N_9926,N_9945);
and UO_459 (O_459,N_9975,N_9994);
nand UO_460 (O_460,N_9942,N_9965);
and UO_461 (O_461,N_9995,N_9927);
and UO_462 (O_462,N_9983,N_9946);
and UO_463 (O_463,N_9923,N_9993);
nand UO_464 (O_464,N_9995,N_9976);
nand UO_465 (O_465,N_9903,N_9950);
nor UO_466 (O_466,N_9998,N_9969);
or UO_467 (O_467,N_9990,N_9996);
nand UO_468 (O_468,N_9976,N_9910);
nor UO_469 (O_469,N_9945,N_9905);
or UO_470 (O_470,N_9983,N_9988);
nand UO_471 (O_471,N_9980,N_9906);
nand UO_472 (O_472,N_9910,N_9959);
xnor UO_473 (O_473,N_9940,N_9949);
nand UO_474 (O_474,N_9906,N_9990);
nand UO_475 (O_475,N_9908,N_9931);
nand UO_476 (O_476,N_9920,N_9929);
nor UO_477 (O_477,N_9927,N_9979);
nand UO_478 (O_478,N_9947,N_9918);
nand UO_479 (O_479,N_9917,N_9974);
nand UO_480 (O_480,N_9974,N_9911);
nor UO_481 (O_481,N_9991,N_9937);
or UO_482 (O_482,N_9911,N_9908);
nand UO_483 (O_483,N_9932,N_9999);
or UO_484 (O_484,N_9943,N_9906);
nor UO_485 (O_485,N_9977,N_9920);
or UO_486 (O_486,N_9942,N_9985);
nand UO_487 (O_487,N_9993,N_9911);
nand UO_488 (O_488,N_9917,N_9947);
nand UO_489 (O_489,N_9950,N_9993);
or UO_490 (O_490,N_9937,N_9992);
nor UO_491 (O_491,N_9984,N_9940);
or UO_492 (O_492,N_9956,N_9944);
nand UO_493 (O_493,N_9967,N_9987);
and UO_494 (O_494,N_9935,N_9913);
and UO_495 (O_495,N_9948,N_9927);
and UO_496 (O_496,N_9916,N_9909);
and UO_497 (O_497,N_9945,N_9924);
nor UO_498 (O_498,N_9954,N_9944);
or UO_499 (O_499,N_9946,N_9954);
and UO_500 (O_500,N_9984,N_9939);
nor UO_501 (O_501,N_9938,N_9931);
nor UO_502 (O_502,N_9952,N_9990);
nor UO_503 (O_503,N_9958,N_9907);
nor UO_504 (O_504,N_9900,N_9978);
xnor UO_505 (O_505,N_9900,N_9989);
nand UO_506 (O_506,N_9928,N_9967);
or UO_507 (O_507,N_9937,N_9928);
or UO_508 (O_508,N_9918,N_9907);
and UO_509 (O_509,N_9960,N_9959);
nand UO_510 (O_510,N_9932,N_9994);
nor UO_511 (O_511,N_9965,N_9996);
or UO_512 (O_512,N_9908,N_9934);
and UO_513 (O_513,N_9925,N_9978);
or UO_514 (O_514,N_9947,N_9955);
nor UO_515 (O_515,N_9928,N_9965);
nand UO_516 (O_516,N_9922,N_9926);
or UO_517 (O_517,N_9934,N_9904);
and UO_518 (O_518,N_9962,N_9974);
xnor UO_519 (O_519,N_9982,N_9920);
nor UO_520 (O_520,N_9986,N_9988);
nand UO_521 (O_521,N_9974,N_9928);
nand UO_522 (O_522,N_9999,N_9939);
nand UO_523 (O_523,N_9949,N_9946);
nand UO_524 (O_524,N_9914,N_9988);
nor UO_525 (O_525,N_9906,N_9942);
nand UO_526 (O_526,N_9989,N_9993);
or UO_527 (O_527,N_9932,N_9964);
and UO_528 (O_528,N_9919,N_9963);
or UO_529 (O_529,N_9935,N_9940);
nor UO_530 (O_530,N_9917,N_9951);
xnor UO_531 (O_531,N_9921,N_9974);
nand UO_532 (O_532,N_9961,N_9939);
and UO_533 (O_533,N_9967,N_9977);
xnor UO_534 (O_534,N_9960,N_9938);
or UO_535 (O_535,N_9918,N_9983);
nor UO_536 (O_536,N_9916,N_9904);
nand UO_537 (O_537,N_9983,N_9954);
xnor UO_538 (O_538,N_9933,N_9908);
nor UO_539 (O_539,N_9943,N_9953);
nand UO_540 (O_540,N_9984,N_9973);
nor UO_541 (O_541,N_9953,N_9954);
and UO_542 (O_542,N_9936,N_9906);
nand UO_543 (O_543,N_9986,N_9932);
nor UO_544 (O_544,N_9964,N_9918);
or UO_545 (O_545,N_9947,N_9923);
nor UO_546 (O_546,N_9948,N_9971);
nand UO_547 (O_547,N_9984,N_9927);
and UO_548 (O_548,N_9945,N_9938);
and UO_549 (O_549,N_9972,N_9964);
or UO_550 (O_550,N_9972,N_9963);
or UO_551 (O_551,N_9968,N_9927);
nor UO_552 (O_552,N_9982,N_9941);
and UO_553 (O_553,N_9951,N_9948);
and UO_554 (O_554,N_9993,N_9938);
and UO_555 (O_555,N_9995,N_9932);
nand UO_556 (O_556,N_9982,N_9946);
nand UO_557 (O_557,N_9944,N_9929);
and UO_558 (O_558,N_9990,N_9921);
and UO_559 (O_559,N_9928,N_9905);
xnor UO_560 (O_560,N_9949,N_9919);
nand UO_561 (O_561,N_9916,N_9948);
nand UO_562 (O_562,N_9945,N_9983);
nand UO_563 (O_563,N_9951,N_9999);
and UO_564 (O_564,N_9977,N_9942);
or UO_565 (O_565,N_9961,N_9923);
or UO_566 (O_566,N_9977,N_9951);
or UO_567 (O_567,N_9992,N_9913);
and UO_568 (O_568,N_9950,N_9954);
nor UO_569 (O_569,N_9977,N_9931);
and UO_570 (O_570,N_9937,N_9999);
and UO_571 (O_571,N_9982,N_9919);
nand UO_572 (O_572,N_9978,N_9957);
and UO_573 (O_573,N_9913,N_9987);
and UO_574 (O_574,N_9955,N_9952);
nand UO_575 (O_575,N_9944,N_9975);
nor UO_576 (O_576,N_9989,N_9983);
and UO_577 (O_577,N_9948,N_9978);
nand UO_578 (O_578,N_9974,N_9994);
or UO_579 (O_579,N_9978,N_9944);
or UO_580 (O_580,N_9973,N_9925);
nand UO_581 (O_581,N_9995,N_9924);
nor UO_582 (O_582,N_9926,N_9901);
nand UO_583 (O_583,N_9964,N_9954);
nor UO_584 (O_584,N_9914,N_9933);
nand UO_585 (O_585,N_9988,N_9962);
nand UO_586 (O_586,N_9952,N_9985);
nand UO_587 (O_587,N_9992,N_9957);
nor UO_588 (O_588,N_9996,N_9967);
and UO_589 (O_589,N_9944,N_9939);
nand UO_590 (O_590,N_9921,N_9943);
nand UO_591 (O_591,N_9912,N_9939);
or UO_592 (O_592,N_9929,N_9939);
or UO_593 (O_593,N_9922,N_9917);
nor UO_594 (O_594,N_9991,N_9946);
and UO_595 (O_595,N_9960,N_9908);
nand UO_596 (O_596,N_9912,N_9951);
nand UO_597 (O_597,N_9909,N_9933);
nor UO_598 (O_598,N_9932,N_9922);
xnor UO_599 (O_599,N_9920,N_9948);
and UO_600 (O_600,N_9913,N_9923);
nor UO_601 (O_601,N_9926,N_9908);
nand UO_602 (O_602,N_9991,N_9994);
and UO_603 (O_603,N_9974,N_9948);
nor UO_604 (O_604,N_9951,N_9946);
and UO_605 (O_605,N_9906,N_9914);
or UO_606 (O_606,N_9940,N_9919);
nor UO_607 (O_607,N_9928,N_9987);
nor UO_608 (O_608,N_9982,N_9995);
or UO_609 (O_609,N_9902,N_9936);
nand UO_610 (O_610,N_9915,N_9968);
or UO_611 (O_611,N_9992,N_9985);
nand UO_612 (O_612,N_9906,N_9918);
nor UO_613 (O_613,N_9944,N_9921);
and UO_614 (O_614,N_9953,N_9960);
nand UO_615 (O_615,N_9969,N_9991);
nand UO_616 (O_616,N_9977,N_9923);
and UO_617 (O_617,N_9990,N_9959);
xor UO_618 (O_618,N_9950,N_9976);
or UO_619 (O_619,N_9979,N_9919);
nand UO_620 (O_620,N_9956,N_9978);
nor UO_621 (O_621,N_9973,N_9959);
or UO_622 (O_622,N_9962,N_9982);
nand UO_623 (O_623,N_9940,N_9971);
and UO_624 (O_624,N_9977,N_9999);
or UO_625 (O_625,N_9950,N_9928);
nor UO_626 (O_626,N_9981,N_9965);
nand UO_627 (O_627,N_9984,N_9949);
or UO_628 (O_628,N_9952,N_9966);
or UO_629 (O_629,N_9973,N_9907);
nor UO_630 (O_630,N_9911,N_9945);
nand UO_631 (O_631,N_9990,N_9955);
and UO_632 (O_632,N_9982,N_9917);
and UO_633 (O_633,N_9974,N_9961);
nor UO_634 (O_634,N_9981,N_9922);
or UO_635 (O_635,N_9951,N_9975);
and UO_636 (O_636,N_9933,N_9924);
and UO_637 (O_637,N_9968,N_9987);
or UO_638 (O_638,N_9963,N_9943);
and UO_639 (O_639,N_9918,N_9932);
xor UO_640 (O_640,N_9992,N_9910);
nor UO_641 (O_641,N_9978,N_9916);
or UO_642 (O_642,N_9966,N_9928);
nand UO_643 (O_643,N_9990,N_9938);
nand UO_644 (O_644,N_9941,N_9936);
and UO_645 (O_645,N_9977,N_9986);
and UO_646 (O_646,N_9973,N_9941);
and UO_647 (O_647,N_9934,N_9916);
nor UO_648 (O_648,N_9970,N_9903);
and UO_649 (O_649,N_9993,N_9958);
nor UO_650 (O_650,N_9921,N_9980);
nand UO_651 (O_651,N_9946,N_9942);
nor UO_652 (O_652,N_9951,N_9981);
nor UO_653 (O_653,N_9900,N_9982);
nand UO_654 (O_654,N_9931,N_9943);
nor UO_655 (O_655,N_9974,N_9922);
and UO_656 (O_656,N_9991,N_9960);
and UO_657 (O_657,N_9901,N_9971);
or UO_658 (O_658,N_9915,N_9950);
and UO_659 (O_659,N_9966,N_9939);
nor UO_660 (O_660,N_9993,N_9910);
nand UO_661 (O_661,N_9971,N_9955);
nand UO_662 (O_662,N_9905,N_9938);
nand UO_663 (O_663,N_9977,N_9944);
and UO_664 (O_664,N_9908,N_9915);
nand UO_665 (O_665,N_9909,N_9957);
nand UO_666 (O_666,N_9908,N_9976);
and UO_667 (O_667,N_9919,N_9926);
nor UO_668 (O_668,N_9946,N_9999);
or UO_669 (O_669,N_9949,N_9960);
and UO_670 (O_670,N_9974,N_9988);
nor UO_671 (O_671,N_9984,N_9911);
and UO_672 (O_672,N_9988,N_9956);
and UO_673 (O_673,N_9902,N_9903);
nor UO_674 (O_674,N_9986,N_9924);
nor UO_675 (O_675,N_9995,N_9913);
nand UO_676 (O_676,N_9927,N_9969);
and UO_677 (O_677,N_9901,N_9937);
or UO_678 (O_678,N_9956,N_9949);
xor UO_679 (O_679,N_9903,N_9908);
and UO_680 (O_680,N_9928,N_9903);
nand UO_681 (O_681,N_9947,N_9929);
or UO_682 (O_682,N_9928,N_9922);
and UO_683 (O_683,N_9921,N_9931);
and UO_684 (O_684,N_9975,N_9915);
or UO_685 (O_685,N_9965,N_9972);
nand UO_686 (O_686,N_9905,N_9985);
or UO_687 (O_687,N_9975,N_9961);
or UO_688 (O_688,N_9966,N_9962);
and UO_689 (O_689,N_9960,N_9931);
nor UO_690 (O_690,N_9943,N_9925);
nor UO_691 (O_691,N_9902,N_9927);
nor UO_692 (O_692,N_9930,N_9995);
and UO_693 (O_693,N_9996,N_9968);
and UO_694 (O_694,N_9932,N_9981);
xor UO_695 (O_695,N_9931,N_9939);
nor UO_696 (O_696,N_9920,N_9927);
and UO_697 (O_697,N_9939,N_9947);
xnor UO_698 (O_698,N_9926,N_9924);
nor UO_699 (O_699,N_9915,N_9901);
nor UO_700 (O_700,N_9953,N_9935);
and UO_701 (O_701,N_9980,N_9944);
nand UO_702 (O_702,N_9933,N_9922);
or UO_703 (O_703,N_9947,N_9986);
nand UO_704 (O_704,N_9930,N_9976);
and UO_705 (O_705,N_9904,N_9978);
nand UO_706 (O_706,N_9961,N_9986);
nand UO_707 (O_707,N_9948,N_9975);
nor UO_708 (O_708,N_9916,N_9918);
xnor UO_709 (O_709,N_9996,N_9943);
or UO_710 (O_710,N_9905,N_9962);
nand UO_711 (O_711,N_9919,N_9986);
and UO_712 (O_712,N_9930,N_9943);
xnor UO_713 (O_713,N_9924,N_9921);
or UO_714 (O_714,N_9931,N_9970);
and UO_715 (O_715,N_9975,N_9998);
nor UO_716 (O_716,N_9927,N_9937);
xnor UO_717 (O_717,N_9922,N_9936);
or UO_718 (O_718,N_9943,N_9929);
nand UO_719 (O_719,N_9945,N_9944);
nand UO_720 (O_720,N_9972,N_9932);
or UO_721 (O_721,N_9994,N_9929);
or UO_722 (O_722,N_9993,N_9975);
nand UO_723 (O_723,N_9932,N_9956);
nor UO_724 (O_724,N_9905,N_9955);
nand UO_725 (O_725,N_9944,N_9928);
xnor UO_726 (O_726,N_9959,N_9923);
nand UO_727 (O_727,N_9988,N_9969);
and UO_728 (O_728,N_9928,N_9958);
and UO_729 (O_729,N_9932,N_9989);
nand UO_730 (O_730,N_9906,N_9901);
nor UO_731 (O_731,N_9954,N_9992);
or UO_732 (O_732,N_9980,N_9922);
or UO_733 (O_733,N_9926,N_9960);
or UO_734 (O_734,N_9907,N_9993);
and UO_735 (O_735,N_9956,N_9915);
xnor UO_736 (O_736,N_9974,N_9971);
or UO_737 (O_737,N_9924,N_9956);
and UO_738 (O_738,N_9922,N_9937);
or UO_739 (O_739,N_9906,N_9969);
or UO_740 (O_740,N_9934,N_9942);
or UO_741 (O_741,N_9963,N_9990);
nand UO_742 (O_742,N_9991,N_9973);
or UO_743 (O_743,N_9983,N_9902);
or UO_744 (O_744,N_9920,N_9928);
nand UO_745 (O_745,N_9992,N_9973);
and UO_746 (O_746,N_9970,N_9905);
and UO_747 (O_747,N_9971,N_9936);
nand UO_748 (O_748,N_9923,N_9908);
nor UO_749 (O_749,N_9984,N_9982);
and UO_750 (O_750,N_9959,N_9942);
nand UO_751 (O_751,N_9944,N_9955);
nand UO_752 (O_752,N_9948,N_9956);
nand UO_753 (O_753,N_9976,N_9978);
and UO_754 (O_754,N_9910,N_9962);
and UO_755 (O_755,N_9939,N_9956);
nand UO_756 (O_756,N_9946,N_9926);
nor UO_757 (O_757,N_9933,N_9932);
or UO_758 (O_758,N_9965,N_9923);
and UO_759 (O_759,N_9990,N_9975);
nand UO_760 (O_760,N_9946,N_9935);
nor UO_761 (O_761,N_9976,N_9942);
and UO_762 (O_762,N_9934,N_9918);
and UO_763 (O_763,N_9937,N_9934);
xnor UO_764 (O_764,N_9957,N_9929);
nor UO_765 (O_765,N_9949,N_9967);
and UO_766 (O_766,N_9908,N_9902);
nand UO_767 (O_767,N_9998,N_9993);
or UO_768 (O_768,N_9980,N_9952);
or UO_769 (O_769,N_9973,N_9971);
nand UO_770 (O_770,N_9902,N_9914);
and UO_771 (O_771,N_9908,N_9916);
nand UO_772 (O_772,N_9997,N_9928);
and UO_773 (O_773,N_9955,N_9939);
nor UO_774 (O_774,N_9987,N_9955);
or UO_775 (O_775,N_9951,N_9954);
or UO_776 (O_776,N_9986,N_9952);
nor UO_777 (O_777,N_9923,N_9910);
nor UO_778 (O_778,N_9976,N_9933);
nand UO_779 (O_779,N_9986,N_9990);
or UO_780 (O_780,N_9993,N_9918);
nand UO_781 (O_781,N_9947,N_9948);
and UO_782 (O_782,N_9915,N_9957);
and UO_783 (O_783,N_9934,N_9986);
or UO_784 (O_784,N_9970,N_9984);
or UO_785 (O_785,N_9995,N_9957);
or UO_786 (O_786,N_9916,N_9912);
and UO_787 (O_787,N_9979,N_9963);
or UO_788 (O_788,N_9967,N_9990);
and UO_789 (O_789,N_9957,N_9936);
or UO_790 (O_790,N_9928,N_9993);
xnor UO_791 (O_791,N_9989,N_9905);
nand UO_792 (O_792,N_9923,N_9928);
nor UO_793 (O_793,N_9980,N_9924);
nor UO_794 (O_794,N_9951,N_9969);
and UO_795 (O_795,N_9904,N_9944);
and UO_796 (O_796,N_9917,N_9990);
or UO_797 (O_797,N_9942,N_9991);
nor UO_798 (O_798,N_9938,N_9998);
and UO_799 (O_799,N_9935,N_9991);
or UO_800 (O_800,N_9984,N_9962);
nand UO_801 (O_801,N_9967,N_9984);
nand UO_802 (O_802,N_9981,N_9934);
or UO_803 (O_803,N_9996,N_9900);
nand UO_804 (O_804,N_9933,N_9937);
nand UO_805 (O_805,N_9903,N_9918);
and UO_806 (O_806,N_9903,N_9995);
and UO_807 (O_807,N_9904,N_9967);
xnor UO_808 (O_808,N_9927,N_9919);
nand UO_809 (O_809,N_9918,N_9979);
and UO_810 (O_810,N_9933,N_9921);
nand UO_811 (O_811,N_9944,N_9982);
nand UO_812 (O_812,N_9910,N_9987);
nand UO_813 (O_813,N_9967,N_9992);
or UO_814 (O_814,N_9973,N_9985);
or UO_815 (O_815,N_9991,N_9901);
and UO_816 (O_816,N_9975,N_9935);
and UO_817 (O_817,N_9909,N_9937);
or UO_818 (O_818,N_9965,N_9948);
and UO_819 (O_819,N_9936,N_9903);
and UO_820 (O_820,N_9952,N_9928);
and UO_821 (O_821,N_9955,N_9984);
or UO_822 (O_822,N_9968,N_9934);
nand UO_823 (O_823,N_9971,N_9968);
and UO_824 (O_824,N_9924,N_9987);
nand UO_825 (O_825,N_9921,N_9965);
nand UO_826 (O_826,N_9967,N_9912);
and UO_827 (O_827,N_9951,N_9960);
or UO_828 (O_828,N_9927,N_9958);
and UO_829 (O_829,N_9922,N_9999);
nor UO_830 (O_830,N_9916,N_9935);
nor UO_831 (O_831,N_9993,N_9957);
or UO_832 (O_832,N_9986,N_9914);
nand UO_833 (O_833,N_9992,N_9907);
xor UO_834 (O_834,N_9911,N_9917);
nand UO_835 (O_835,N_9997,N_9907);
and UO_836 (O_836,N_9991,N_9964);
or UO_837 (O_837,N_9975,N_9964);
nor UO_838 (O_838,N_9991,N_9924);
or UO_839 (O_839,N_9942,N_9992);
or UO_840 (O_840,N_9908,N_9944);
or UO_841 (O_841,N_9943,N_9986);
nor UO_842 (O_842,N_9965,N_9970);
or UO_843 (O_843,N_9962,N_9919);
or UO_844 (O_844,N_9936,N_9918);
nor UO_845 (O_845,N_9926,N_9913);
nor UO_846 (O_846,N_9943,N_9939);
and UO_847 (O_847,N_9956,N_9999);
xnor UO_848 (O_848,N_9997,N_9975);
and UO_849 (O_849,N_9924,N_9952);
and UO_850 (O_850,N_9935,N_9918);
or UO_851 (O_851,N_9912,N_9934);
nand UO_852 (O_852,N_9946,N_9977);
and UO_853 (O_853,N_9905,N_9963);
or UO_854 (O_854,N_9936,N_9911);
nor UO_855 (O_855,N_9946,N_9978);
xnor UO_856 (O_856,N_9929,N_9915);
nand UO_857 (O_857,N_9969,N_9910);
nor UO_858 (O_858,N_9956,N_9989);
nor UO_859 (O_859,N_9908,N_9977);
nor UO_860 (O_860,N_9925,N_9965);
nor UO_861 (O_861,N_9942,N_9969);
and UO_862 (O_862,N_9989,N_9971);
and UO_863 (O_863,N_9948,N_9904);
or UO_864 (O_864,N_9986,N_9959);
xor UO_865 (O_865,N_9913,N_9904);
xor UO_866 (O_866,N_9909,N_9998);
nor UO_867 (O_867,N_9951,N_9941);
and UO_868 (O_868,N_9935,N_9908);
and UO_869 (O_869,N_9945,N_9968);
nand UO_870 (O_870,N_9978,N_9984);
and UO_871 (O_871,N_9908,N_9986);
nor UO_872 (O_872,N_9920,N_9919);
nand UO_873 (O_873,N_9915,N_9981);
or UO_874 (O_874,N_9926,N_9921);
xnor UO_875 (O_875,N_9996,N_9963);
nor UO_876 (O_876,N_9915,N_9978);
or UO_877 (O_877,N_9993,N_9916);
and UO_878 (O_878,N_9913,N_9974);
xor UO_879 (O_879,N_9905,N_9916);
or UO_880 (O_880,N_9901,N_9988);
or UO_881 (O_881,N_9977,N_9968);
and UO_882 (O_882,N_9947,N_9931);
nand UO_883 (O_883,N_9909,N_9972);
or UO_884 (O_884,N_9935,N_9923);
and UO_885 (O_885,N_9925,N_9949);
and UO_886 (O_886,N_9979,N_9921);
nand UO_887 (O_887,N_9983,N_9948);
and UO_888 (O_888,N_9967,N_9985);
nand UO_889 (O_889,N_9921,N_9969);
and UO_890 (O_890,N_9965,N_9974);
and UO_891 (O_891,N_9943,N_9948);
xnor UO_892 (O_892,N_9936,N_9972);
xor UO_893 (O_893,N_9951,N_9996);
and UO_894 (O_894,N_9984,N_9904);
and UO_895 (O_895,N_9908,N_9942);
or UO_896 (O_896,N_9942,N_9978);
nor UO_897 (O_897,N_9960,N_9942);
xor UO_898 (O_898,N_9911,N_9902);
nand UO_899 (O_899,N_9942,N_9907);
nand UO_900 (O_900,N_9905,N_9919);
nand UO_901 (O_901,N_9963,N_9937);
nand UO_902 (O_902,N_9990,N_9962);
nor UO_903 (O_903,N_9973,N_9923);
and UO_904 (O_904,N_9976,N_9974);
nand UO_905 (O_905,N_9967,N_9910);
or UO_906 (O_906,N_9988,N_9906);
or UO_907 (O_907,N_9963,N_9959);
and UO_908 (O_908,N_9916,N_9989);
or UO_909 (O_909,N_9976,N_9979);
or UO_910 (O_910,N_9911,N_9995);
nand UO_911 (O_911,N_9901,N_9909);
nor UO_912 (O_912,N_9901,N_9953);
nand UO_913 (O_913,N_9913,N_9900);
and UO_914 (O_914,N_9922,N_9961);
xnor UO_915 (O_915,N_9920,N_9963);
and UO_916 (O_916,N_9915,N_9919);
and UO_917 (O_917,N_9996,N_9998);
and UO_918 (O_918,N_9911,N_9916);
nand UO_919 (O_919,N_9970,N_9987);
xor UO_920 (O_920,N_9919,N_9969);
nand UO_921 (O_921,N_9907,N_9915);
or UO_922 (O_922,N_9929,N_9910);
xor UO_923 (O_923,N_9946,N_9995);
or UO_924 (O_924,N_9931,N_9904);
and UO_925 (O_925,N_9991,N_9939);
nand UO_926 (O_926,N_9954,N_9901);
or UO_927 (O_927,N_9925,N_9957);
and UO_928 (O_928,N_9961,N_9929);
and UO_929 (O_929,N_9927,N_9975);
nand UO_930 (O_930,N_9968,N_9997);
nor UO_931 (O_931,N_9928,N_9959);
or UO_932 (O_932,N_9963,N_9946);
and UO_933 (O_933,N_9925,N_9946);
or UO_934 (O_934,N_9929,N_9949);
or UO_935 (O_935,N_9929,N_9925);
or UO_936 (O_936,N_9935,N_9992);
nor UO_937 (O_937,N_9907,N_9986);
nor UO_938 (O_938,N_9937,N_9998);
or UO_939 (O_939,N_9976,N_9927);
or UO_940 (O_940,N_9925,N_9951);
nand UO_941 (O_941,N_9995,N_9993);
and UO_942 (O_942,N_9918,N_9987);
and UO_943 (O_943,N_9962,N_9948);
nand UO_944 (O_944,N_9935,N_9966);
nand UO_945 (O_945,N_9944,N_9983);
nand UO_946 (O_946,N_9924,N_9983);
or UO_947 (O_947,N_9955,N_9959);
and UO_948 (O_948,N_9935,N_9915);
and UO_949 (O_949,N_9986,N_9985);
or UO_950 (O_950,N_9903,N_9956);
nor UO_951 (O_951,N_9900,N_9966);
nor UO_952 (O_952,N_9955,N_9941);
nand UO_953 (O_953,N_9965,N_9977);
nor UO_954 (O_954,N_9983,N_9961);
and UO_955 (O_955,N_9936,N_9938);
xor UO_956 (O_956,N_9955,N_9907);
and UO_957 (O_957,N_9916,N_9920);
nand UO_958 (O_958,N_9913,N_9951);
nand UO_959 (O_959,N_9955,N_9911);
xnor UO_960 (O_960,N_9987,N_9912);
or UO_961 (O_961,N_9900,N_9975);
nor UO_962 (O_962,N_9934,N_9936);
and UO_963 (O_963,N_9943,N_9968);
and UO_964 (O_964,N_9962,N_9997);
and UO_965 (O_965,N_9924,N_9912);
or UO_966 (O_966,N_9934,N_9984);
and UO_967 (O_967,N_9998,N_9941);
nor UO_968 (O_968,N_9939,N_9976);
nor UO_969 (O_969,N_9980,N_9948);
nand UO_970 (O_970,N_9921,N_9976);
nand UO_971 (O_971,N_9905,N_9968);
and UO_972 (O_972,N_9930,N_9907);
nor UO_973 (O_973,N_9929,N_9953);
nor UO_974 (O_974,N_9944,N_9987);
nor UO_975 (O_975,N_9954,N_9930);
and UO_976 (O_976,N_9960,N_9929);
xor UO_977 (O_977,N_9905,N_9944);
nand UO_978 (O_978,N_9902,N_9987);
nand UO_979 (O_979,N_9989,N_9930);
or UO_980 (O_980,N_9967,N_9948);
xor UO_981 (O_981,N_9934,N_9967);
xnor UO_982 (O_982,N_9965,N_9998);
nor UO_983 (O_983,N_9995,N_9997);
and UO_984 (O_984,N_9976,N_9986);
and UO_985 (O_985,N_9922,N_9958);
and UO_986 (O_986,N_9953,N_9980);
nand UO_987 (O_987,N_9925,N_9950);
or UO_988 (O_988,N_9997,N_9950);
and UO_989 (O_989,N_9981,N_9999);
nand UO_990 (O_990,N_9971,N_9969);
nand UO_991 (O_991,N_9942,N_9996);
and UO_992 (O_992,N_9963,N_9995);
nand UO_993 (O_993,N_9958,N_9912);
and UO_994 (O_994,N_9925,N_9970);
nor UO_995 (O_995,N_9931,N_9923);
nand UO_996 (O_996,N_9947,N_9977);
nor UO_997 (O_997,N_9916,N_9986);
or UO_998 (O_998,N_9989,N_9907);
nand UO_999 (O_999,N_9984,N_9952);
nand UO_1000 (O_1000,N_9904,N_9929);
nor UO_1001 (O_1001,N_9948,N_9995);
nor UO_1002 (O_1002,N_9996,N_9975);
xor UO_1003 (O_1003,N_9933,N_9989);
or UO_1004 (O_1004,N_9968,N_9928);
xnor UO_1005 (O_1005,N_9926,N_9992);
nor UO_1006 (O_1006,N_9983,N_9904);
nor UO_1007 (O_1007,N_9941,N_9963);
and UO_1008 (O_1008,N_9952,N_9905);
xnor UO_1009 (O_1009,N_9987,N_9964);
and UO_1010 (O_1010,N_9996,N_9995);
nand UO_1011 (O_1011,N_9993,N_9926);
nand UO_1012 (O_1012,N_9988,N_9957);
nand UO_1013 (O_1013,N_9904,N_9991);
nor UO_1014 (O_1014,N_9957,N_9980);
nand UO_1015 (O_1015,N_9952,N_9944);
and UO_1016 (O_1016,N_9972,N_9989);
or UO_1017 (O_1017,N_9921,N_9923);
nand UO_1018 (O_1018,N_9945,N_9990);
nor UO_1019 (O_1019,N_9930,N_9960);
and UO_1020 (O_1020,N_9927,N_9997);
nand UO_1021 (O_1021,N_9985,N_9928);
nor UO_1022 (O_1022,N_9901,N_9922);
nand UO_1023 (O_1023,N_9959,N_9916);
or UO_1024 (O_1024,N_9944,N_9950);
xnor UO_1025 (O_1025,N_9994,N_9946);
nand UO_1026 (O_1026,N_9969,N_9976);
or UO_1027 (O_1027,N_9972,N_9960);
nand UO_1028 (O_1028,N_9937,N_9938);
nand UO_1029 (O_1029,N_9943,N_9954);
nor UO_1030 (O_1030,N_9989,N_9980);
or UO_1031 (O_1031,N_9941,N_9912);
nand UO_1032 (O_1032,N_9956,N_9974);
nand UO_1033 (O_1033,N_9995,N_9914);
nor UO_1034 (O_1034,N_9975,N_9926);
or UO_1035 (O_1035,N_9956,N_9955);
xnor UO_1036 (O_1036,N_9973,N_9910);
and UO_1037 (O_1037,N_9931,N_9905);
nand UO_1038 (O_1038,N_9982,N_9964);
and UO_1039 (O_1039,N_9919,N_9993);
xor UO_1040 (O_1040,N_9913,N_9950);
or UO_1041 (O_1041,N_9941,N_9962);
nor UO_1042 (O_1042,N_9956,N_9951);
nor UO_1043 (O_1043,N_9934,N_9957);
or UO_1044 (O_1044,N_9980,N_9942);
xor UO_1045 (O_1045,N_9936,N_9985);
or UO_1046 (O_1046,N_9979,N_9906);
nor UO_1047 (O_1047,N_9906,N_9991);
and UO_1048 (O_1048,N_9943,N_9918);
and UO_1049 (O_1049,N_9990,N_9953);
nand UO_1050 (O_1050,N_9928,N_9933);
and UO_1051 (O_1051,N_9944,N_9968);
nand UO_1052 (O_1052,N_9994,N_9952);
nand UO_1053 (O_1053,N_9935,N_9979);
nor UO_1054 (O_1054,N_9924,N_9942);
or UO_1055 (O_1055,N_9934,N_9989);
and UO_1056 (O_1056,N_9940,N_9907);
xnor UO_1057 (O_1057,N_9994,N_9906);
nand UO_1058 (O_1058,N_9959,N_9935);
and UO_1059 (O_1059,N_9949,N_9918);
or UO_1060 (O_1060,N_9998,N_9981);
nor UO_1061 (O_1061,N_9987,N_9989);
nor UO_1062 (O_1062,N_9943,N_9965);
and UO_1063 (O_1063,N_9917,N_9977);
nor UO_1064 (O_1064,N_9962,N_9901);
nand UO_1065 (O_1065,N_9982,N_9948);
nand UO_1066 (O_1066,N_9971,N_9916);
nor UO_1067 (O_1067,N_9993,N_9967);
nor UO_1068 (O_1068,N_9906,N_9986);
nand UO_1069 (O_1069,N_9929,N_9996);
nor UO_1070 (O_1070,N_9953,N_9912);
or UO_1071 (O_1071,N_9926,N_9964);
nor UO_1072 (O_1072,N_9961,N_9953);
nand UO_1073 (O_1073,N_9934,N_9974);
and UO_1074 (O_1074,N_9911,N_9998);
and UO_1075 (O_1075,N_9947,N_9981);
nor UO_1076 (O_1076,N_9954,N_9907);
xor UO_1077 (O_1077,N_9938,N_9989);
and UO_1078 (O_1078,N_9957,N_9997);
xor UO_1079 (O_1079,N_9941,N_9934);
and UO_1080 (O_1080,N_9988,N_9943);
nand UO_1081 (O_1081,N_9997,N_9921);
xor UO_1082 (O_1082,N_9966,N_9961);
and UO_1083 (O_1083,N_9900,N_9951);
nand UO_1084 (O_1084,N_9968,N_9929);
nand UO_1085 (O_1085,N_9998,N_9902);
or UO_1086 (O_1086,N_9987,N_9926);
or UO_1087 (O_1087,N_9909,N_9996);
or UO_1088 (O_1088,N_9901,N_9923);
nand UO_1089 (O_1089,N_9963,N_9931);
and UO_1090 (O_1090,N_9980,N_9981);
or UO_1091 (O_1091,N_9912,N_9919);
and UO_1092 (O_1092,N_9934,N_9914);
and UO_1093 (O_1093,N_9952,N_9962);
nor UO_1094 (O_1094,N_9979,N_9958);
nand UO_1095 (O_1095,N_9921,N_9929);
nand UO_1096 (O_1096,N_9946,N_9904);
xor UO_1097 (O_1097,N_9914,N_9985);
or UO_1098 (O_1098,N_9982,N_9973);
and UO_1099 (O_1099,N_9981,N_9958);
nor UO_1100 (O_1100,N_9960,N_9920);
xnor UO_1101 (O_1101,N_9956,N_9901);
nand UO_1102 (O_1102,N_9926,N_9957);
and UO_1103 (O_1103,N_9931,N_9973);
nor UO_1104 (O_1104,N_9929,N_9956);
or UO_1105 (O_1105,N_9958,N_9940);
nand UO_1106 (O_1106,N_9978,N_9968);
nor UO_1107 (O_1107,N_9955,N_9942);
nor UO_1108 (O_1108,N_9923,N_9927);
nor UO_1109 (O_1109,N_9915,N_9973);
and UO_1110 (O_1110,N_9918,N_9994);
nand UO_1111 (O_1111,N_9965,N_9963);
and UO_1112 (O_1112,N_9903,N_9990);
or UO_1113 (O_1113,N_9933,N_9994);
and UO_1114 (O_1114,N_9942,N_9926);
nand UO_1115 (O_1115,N_9966,N_9983);
and UO_1116 (O_1116,N_9997,N_9945);
nor UO_1117 (O_1117,N_9967,N_9924);
xnor UO_1118 (O_1118,N_9985,N_9946);
nand UO_1119 (O_1119,N_9969,N_9987);
nand UO_1120 (O_1120,N_9954,N_9975);
nand UO_1121 (O_1121,N_9992,N_9991);
nand UO_1122 (O_1122,N_9969,N_9915);
nor UO_1123 (O_1123,N_9986,N_9972);
nand UO_1124 (O_1124,N_9950,N_9980);
nor UO_1125 (O_1125,N_9985,N_9933);
or UO_1126 (O_1126,N_9985,N_9970);
or UO_1127 (O_1127,N_9998,N_9990);
nor UO_1128 (O_1128,N_9959,N_9929);
nand UO_1129 (O_1129,N_9967,N_9991);
xnor UO_1130 (O_1130,N_9998,N_9977);
nand UO_1131 (O_1131,N_9902,N_9971);
nor UO_1132 (O_1132,N_9919,N_9917);
nor UO_1133 (O_1133,N_9944,N_9959);
and UO_1134 (O_1134,N_9942,N_9918);
xor UO_1135 (O_1135,N_9924,N_9990);
and UO_1136 (O_1136,N_9962,N_9927);
nand UO_1137 (O_1137,N_9933,N_9929);
nor UO_1138 (O_1138,N_9973,N_9961);
nor UO_1139 (O_1139,N_9998,N_9940);
or UO_1140 (O_1140,N_9925,N_9923);
or UO_1141 (O_1141,N_9955,N_9933);
or UO_1142 (O_1142,N_9901,N_9907);
and UO_1143 (O_1143,N_9945,N_9958);
xnor UO_1144 (O_1144,N_9967,N_9900);
or UO_1145 (O_1145,N_9962,N_9921);
or UO_1146 (O_1146,N_9912,N_9922);
nand UO_1147 (O_1147,N_9933,N_9938);
nor UO_1148 (O_1148,N_9939,N_9993);
nor UO_1149 (O_1149,N_9985,N_9920);
or UO_1150 (O_1150,N_9954,N_9998);
or UO_1151 (O_1151,N_9967,N_9907);
xnor UO_1152 (O_1152,N_9950,N_9965);
nor UO_1153 (O_1153,N_9913,N_9967);
nor UO_1154 (O_1154,N_9916,N_9994);
or UO_1155 (O_1155,N_9964,N_9917);
nand UO_1156 (O_1156,N_9904,N_9938);
and UO_1157 (O_1157,N_9997,N_9961);
or UO_1158 (O_1158,N_9900,N_9994);
nand UO_1159 (O_1159,N_9932,N_9936);
and UO_1160 (O_1160,N_9999,N_9972);
xnor UO_1161 (O_1161,N_9994,N_9982);
and UO_1162 (O_1162,N_9929,N_9977);
or UO_1163 (O_1163,N_9999,N_9997);
nand UO_1164 (O_1164,N_9976,N_9975);
and UO_1165 (O_1165,N_9913,N_9991);
nor UO_1166 (O_1166,N_9938,N_9980);
nor UO_1167 (O_1167,N_9965,N_9933);
xnor UO_1168 (O_1168,N_9909,N_9973);
and UO_1169 (O_1169,N_9979,N_9904);
and UO_1170 (O_1170,N_9966,N_9904);
or UO_1171 (O_1171,N_9972,N_9907);
nand UO_1172 (O_1172,N_9925,N_9908);
nand UO_1173 (O_1173,N_9982,N_9958);
xnor UO_1174 (O_1174,N_9964,N_9978);
or UO_1175 (O_1175,N_9976,N_9951);
nand UO_1176 (O_1176,N_9947,N_9974);
and UO_1177 (O_1177,N_9907,N_9928);
and UO_1178 (O_1178,N_9916,N_9926);
or UO_1179 (O_1179,N_9997,N_9974);
nor UO_1180 (O_1180,N_9966,N_9956);
nor UO_1181 (O_1181,N_9918,N_9912);
nand UO_1182 (O_1182,N_9901,N_9980);
and UO_1183 (O_1183,N_9939,N_9994);
and UO_1184 (O_1184,N_9901,N_9949);
nor UO_1185 (O_1185,N_9919,N_9968);
and UO_1186 (O_1186,N_9913,N_9988);
nor UO_1187 (O_1187,N_9982,N_9983);
or UO_1188 (O_1188,N_9986,N_9915);
nand UO_1189 (O_1189,N_9921,N_9967);
or UO_1190 (O_1190,N_9922,N_9907);
nor UO_1191 (O_1191,N_9959,N_9933);
nor UO_1192 (O_1192,N_9924,N_9911);
or UO_1193 (O_1193,N_9969,N_9957);
nor UO_1194 (O_1194,N_9994,N_9915);
or UO_1195 (O_1195,N_9971,N_9996);
nor UO_1196 (O_1196,N_9934,N_9991);
nand UO_1197 (O_1197,N_9930,N_9958);
or UO_1198 (O_1198,N_9917,N_9962);
nand UO_1199 (O_1199,N_9938,N_9971);
nand UO_1200 (O_1200,N_9988,N_9904);
nor UO_1201 (O_1201,N_9980,N_9960);
nor UO_1202 (O_1202,N_9999,N_9901);
nor UO_1203 (O_1203,N_9976,N_9982);
nand UO_1204 (O_1204,N_9964,N_9920);
nor UO_1205 (O_1205,N_9918,N_9921);
nand UO_1206 (O_1206,N_9920,N_9943);
and UO_1207 (O_1207,N_9945,N_9907);
or UO_1208 (O_1208,N_9908,N_9957);
nand UO_1209 (O_1209,N_9923,N_9932);
or UO_1210 (O_1210,N_9983,N_9986);
nand UO_1211 (O_1211,N_9946,N_9924);
and UO_1212 (O_1212,N_9992,N_9917);
nand UO_1213 (O_1213,N_9995,N_9994);
nor UO_1214 (O_1214,N_9913,N_9986);
nor UO_1215 (O_1215,N_9942,N_9902);
nand UO_1216 (O_1216,N_9915,N_9926);
xnor UO_1217 (O_1217,N_9970,N_9989);
or UO_1218 (O_1218,N_9948,N_9959);
nor UO_1219 (O_1219,N_9983,N_9922);
nand UO_1220 (O_1220,N_9950,N_9968);
and UO_1221 (O_1221,N_9918,N_9982);
or UO_1222 (O_1222,N_9978,N_9985);
and UO_1223 (O_1223,N_9992,N_9988);
and UO_1224 (O_1224,N_9904,N_9973);
nand UO_1225 (O_1225,N_9944,N_9936);
nand UO_1226 (O_1226,N_9916,N_9954);
or UO_1227 (O_1227,N_9957,N_9942);
or UO_1228 (O_1228,N_9920,N_9900);
or UO_1229 (O_1229,N_9970,N_9994);
xnor UO_1230 (O_1230,N_9907,N_9927);
nand UO_1231 (O_1231,N_9977,N_9926);
nor UO_1232 (O_1232,N_9914,N_9992);
or UO_1233 (O_1233,N_9944,N_9971);
xnor UO_1234 (O_1234,N_9905,N_9991);
nor UO_1235 (O_1235,N_9900,N_9933);
or UO_1236 (O_1236,N_9958,N_9950);
nor UO_1237 (O_1237,N_9952,N_9992);
and UO_1238 (O_1238,N_9947,N_9964);
and UO_1239 (O_1239,N_9900,N_9903);
xnor UO_1240 (O_1240,N_9969,N_9930);
and UO_1241 (O_1241,N_9983,N_9910);
nand UO_1242 (O_1242,N_9931,N_9952);
nand UO_1243 (O_1243,N_9993,N_9973);
and UO_1244 (O_1244,N_9927,N_9989);
nor UO_1245 (O_1245,N_9949,N_9983);
nand UO_1246 (O_1246,N_9909,N_9995);
xnor UO_1247 (O_1247,N_9935,N_9968);
nand UO_1248 (O_1248,N_9990,N_9976);
nand UO_1249 (O_1249,N_9986,N_9901);
or UO_1250 (O_1250,N_9945,N_9915);
or UO_1251 (O_1251,N_9979,N_9932);
or UO_1252 (O_1252,N_9913,N_9999);
xor UO_1253 (O_1253,N_9979,N_9997);
nand UO_1254 (O_1254,N_9930,N_9910);
nor UO_1255 (O_1255,N_9918,N_9913);
nor UO_1256 (O_1256,N_9923,N_9904);
nor UO_1257 (O_1257,N_9948,N_9940);
and UO_1258 (O_1258,N_9904,N_9932);
and UO_1259 (O_1259,N_9908,N_9971);
or UO_1260 (O_1260,N_9930,N_9955);
nand UO_1261 (O_1261,N_9980,N_9971);
or UO_1262 (O_1262,N_9970,N_9945);
nand UO_1263 (O_1263,N_9968,N_9967);
nor UO_1264 (O_1264,N_9987,N_9994);
xnor UO_1265 (O_1265,N_9957,N_9906);
nor UO_1266 (O_1266,N_9946,N_9921);
nand UO_1267 (O_1267,N_9999,N_9986);
or UO_1268 (O_1268,N_9948,N_9912);
xnor UO_1269 (O_1269,N_9929,N_9952);
or UO_1270 (O_1270,N_9919,N_9998);
nand UO_1271 (O_1271,N_9915,N_9949);
nor UO_1272 (O_1272,N_9903,N_9905);
xor UO_1273 (O_1273,N_9951,N_9928);
or UO_1274 (O_1274,N_9933,N_9931);
xnor UO_1275 (O_1275,N_9974,N_9966);
or UO_1276 (O_1276,N_9928,N_9963);
nand UO_1277 (O_1277,N_9968,N_9995);
nor UO_1278 (O_1278,N_9988,N_9955);
nand UO_1279 (O_1279,N_9962,N_9976);
nor UO_1280 (O_1280,N_9969,N_9977);
nor UO_1281 (O_1281,N_9908,N_9950);
nand UO_1282 (O_1282,N_9969,N_9920);
nand UO_1283 (O_1283,N_9972,N_9988);
or UO_1284 (O_1284,N_9948,N_9919);
nor UO_1285 (O_1285,N_9983,N_9972);
and UO_1286 (O_1286,N_9963,N_9969);
and UO_1287 (O_1287,N_9969,N_9925);
and UO_1288 (O_1288,N_9905,N_9993);
nand UO_1289 (O_1289,N_9952,N_9947);
or UO_1290 (O_1290,N_9944,N_9989);
nor UO_1291 (O_1291,N_9971,N_9959);
nor UO_1292 (O_1292,N_9967,N_9908);
and UO_1293 (O_1293,N_9929,N_9986);
nand UO_1294 (O_1294,N_9975,N_9917);
or UO_1295 (O_1295,N_9971,N_9963);
nor UO_1296 (O_1296,N_9974,N_9935);
or UO_1297 (O_1297,N_9919,N_9988);
or UO_1298 (O_1298,N_9923,N_9982);
or UO_1299 (O_1299,N_9939,N_9942);
or UO_1300 (O_1300,N_9990,N_9909);
nand UO_1301 (O_1301,N_9980,N_9977);
nor UO_1302 (O_1302,N_9949,N_9930);
and UO_1303 (O_1303,N_9983,N_9984);
and UO_1304 (O_1304,N_9964,N_9979);
or UO_1305 (O_1305,N_9902,N_9901);
nor UO_1306 (O_1306,N_9991,N_9990);
nor UO_1307 (O_1307,N_9930,N_9936);
nand UO_1308 (O_1308,N_9955,N_9975);
and UO_1309 (O_1309,N_9912,N_9992);
or UO_1310 (O_1310,N_9904,N_9962);
nand UO_1311 (O_1311,N_9928,N_9994);
nand UO_1312 (O_1312,N_9939,N_9958);
and UO_1313 (O_1313,N_9943,N_9914);
and UO_1314 (O_1314,N_9990,N_9950);
nor UO_1315 (O_1315,N_9997,N_9912);
and UO_1316 (O_1316,N_9971,N_9950);
and UO_1317 (O_1317,N_9928,N_9913);
nor UO_1318 (O_1318,N_9952,N_9918);
or UO_1319 (O_1319,N_9967,N_9975);
nand UO_1320 (O_1320,N_9904,N_9912);
nand UO_1321 (O_1321,N_9984,N_9924);
or UO_1322 (O_1322,N_9953,N_9967);
nor UO_1323 (O_1323,N_9926,N_9984);
and UO_1324 (O_1324,N_9996,N_9911);
nor UO_1325 (O_1325,N_9970,N_9950);
or UO_1326 (O_1326,N_9943,N_9995);
nand UO_1327 (O_1327,N_9980,N_9920);
or UO_1328 (O_1328,N_9927,N_9955);
nand UO_1329 (O_1329,N_9954,N_9928);
and UO_1330 (O_1330,N_9934,N_9990);
or UO_1331 (O_1331,N_9986,N_9939);
xnor UO_1332 (O_1332,N_9979,N_9947);
or UO_1333 (O_1333,N_9988,N_9917);
and UO_1334 (O_1334,N_9932,N_9900);
xor UO_1335 (O_1335,N_9965,N_9914);
or UO_1336 (O_1336,N_9935,N_9927);
and UO_1337 (O_1337,N_9950,N_9904);
nor UO_1338 (O_1338,N_9958,N_9997);
xor UO_1339 (O_1339,N_9929,N_9911);
nor UO_1340 (O_1340,N_9901,N_9912);
and UO_1341 (O_1341,N_9920,N_9926);
nand UO_1342 (O_1342,N_9932,N_9952);
and UO_1343 (O_1343,N_9963,N_9936);
xor UO_1344 (O_1344,N_9988,N_9948);
nand UO_1345 (O_1345,N_9985,N_9919);
nor UO_1346 (O_1346,N_9936,N_9940);
or UO_1347 (O_1347,N_9987,N_9997);
nor UO_1348 (O_1348,N_9975,N_9966);
nand UO_1349 (O_1349,N_9936,N_9955);
or UO_1350 (O_1350,N_9910,N_9995);
and UO_1351 (O_1351,N_9998,N_9930);
or UO_1352 (O_1352,N_9992,N_9931);
xor UO_1353 (O_1353,N_9978,N_9907);
or UO_1354 (O_1354,N_9950,N_9919);
or UO_1355 (O_1355,N_9966,N_9933);
nand UO_1356 (O_1356,N_9979,N_9900);
xnor UO_1357 (O_1357,N_9932,N_9924);
nor UO_1358 (O_1358,N_9958,N_9932);
and UO_1359 (O_1359,N_9948,N_9908);
or UO_1360 (O_1360,N_9986,N_9992);
nand UO_1361 (O_1361,N_9932,N_9906);
or UO_1362 (O_1362,N_9915,N_9917);
and UO_1363 (O_1363,N_9912,N_9943);
and UO_1364 (O_1364,N_9953,N_9918);
or UO_1365 (O_1365,N_9936,N_9920);
and UO_1366 (O_1366,N_9925,N_9920);
nand UO_1367 (O_1367,N_9914,N_9960);
xor UO_1368 (O_1368,N_9908,N_9978);
nand UO_1369 (O_1369,N_9994,N_9908);
nor UO_1370 (O_1370,N_9931,N_9988);
nand UO_1371 (O_1371,N_9935,N_9952);
or UO_1372 (O_1372,N_9921,N_9971);
and UO_1373 (O_1373,N_9925,N_9958);
and UO_1374 (O_1374,N_9983,N_9981);
nor UO_1375 (O_1375,N_9922,N_9996);
and UO_1376 (O_1376,N_9996,N_9918);
nand UO_1377 (O_1377,N_9995,N_9969);
or UO_1378 (O_1378,N_9999,N_9902);
nor UO_1379 (O_1379,N_9995,N_9942);
nor UO_1380 (O_1380,N_9904,N_9986);
nand UO_1381 (O_1381,N_9953,N_9936);
and UO_1382 (O_1382,N_9938,N_9941);
nand UO_1383 (O_1383,N_9903,N_9910);
and UO_1384 (O_1384,N_9971,N_9964);
nor UO_1385 (O_1385,N_9994,N_9949);
or UO_1386 (O_1386,N_9988,N_9963);
and UO_1387 (O_1387,N_9917,N_9945);
nor UO_1388 (O_1388,N_9965,N_9987);
nor UO_1389 (O_1389,N_9917,N_9916);
and UO_1390 (O_1390,N_9946,N_9905);
nor UO_1391 (O_1391,N_9967,N_9944);
or UO_1392 (O_1392,N_9989,N_9922);
and UO_1393 (O_1393,N_9906,N_9922);
and UO_1394 (O_1394,N_9922,N_9995);
and UO_1395 (O_1395,N_9952,N_9977);
or UO_1396 (O_1396,N_9925,N_9917);
or UO_1397 (O_1397,N_9979,N_9938);
or UO_1398 (O_1398,N_9976,N_9959);
nand UO_1399 (O_1399,N_9936,N_9904);
and UO_1400 (O_1400,N_9920,N_9997);
nor UO_1401 (O_1401,N_9930,N_9994);
xor UO_1402 (O_1402,N_9979,N_9923);
xnor UO_1403 (O_1403,N_9977,N_9935);
nand UO_1404 (O_1404,N_9998,N_9973);
and UO_1405 (O_1405,N_9982,N_9966);
and UO_1406 (O_1406,N_9995,N_9923);
or UO_1407 (O_1407,N_9953,N_9958);
or UO_1408 (O_1408,N_9912,N_9983);
xnor UO_1409 (O_1409,N_9993,N_9976);
nand UO_1410 (O_1410,N_9990,N_9922);
nand UO_1411 (O_1411,N_9989,N_9986);
nand UO_1412 (O_1412,N_9948,N_9918);
or UO_1413 (O_1413,N_9918,N_9997);
nand UO_1414 (O_1414,N_9978,N_9921);
and UO_1415 (O_1415,N_9934,N_9977);
and UO_1416 (O_1416,N_9928,N_9970);
or UO_1417 (O_1417,N_9997,N_9986);
and UO_1418 (O_1418,N_9959,N_9918);
xnor UO_1419 (O_1419,N_9953,N_9906);
nor UO_1420 (O_1420,N_9989,N_9951);
or UO_1421 (O_1421,N_9949,N_9931);
nand UO_1422 (O_1422,N_9905,N_9995);
nor UO_1423 (O_1423,N_9918,N_9976);
and UO_1424 (O_1424,N_9901,N_9981);
xnor UO_1425 (O_1425,N_9979,N_9937);
or UO_1426 (O_1426,N_9911,N_9938);
nor UO_1427 (O_1427,N_9952,N_9974);
and UO_1428 (O_1428,N_9939,N_9901);
or UO_1429 (O_1429,N_9935,N_9909);
and UO_1430 (O_1430,N_9966,N_9930);
nor UO_1431 (O_1431,N_9973,N_9994);
or UO_1432 (O_1432,N_9939,N_9971);
nor UO_1433 (O_1433,N_9916,N_9925);
xnor UO_1434 (O_1434,N_9980,N_9997);
nand UO_1435 (O_1435,N_9912,N_9993);
or UO_1436 (O_1436,N_9920,N_9937);
nor UO_1437 (O_1437,N_9994,N_9909);
nand UO_1438 (O_1438,N_9906,N_9913);
and UO_1439 (O_1439,N_9992,N_9921);
or UO_1440 (O_1440,N_9973,N_9969);
nor UO_1441 (O_1441,N_9975,N_9904);
nor UO_1442 (O_1442,N_9938,N_9958);
and UO_1443 (O_1443,N_9970,N_9944);
nand UO_1444 (O_1444,N_9914,N_9948);
nand UO_1445 (O_1445,N_9923,N_9958);
nand UO_1446 (O_1446,N_9944,N_9973);
or UO_1447 (O_1447,N_9961,N_9954);
nor UO_1448 (O_1448,N_9957,N_9901);
and UO_1449 (O_1449,N_9963,N_9986);
and UO_1450 (O_1450,N_9930,N_9925);
nor UO_1451 (O_1451,N_9959,N_9914);
and UO_1452 (O_1452,N_9907,N_9912);
nand UO_1453 (O_1453,N_9968,N_9951);
nor UO_1454 (O_1454,N_9916,N_9960);
nand UO_1455 (O_1455,N_9947,N_9995);
nor UO_1456 (O_1456,N_9973,N_9965);
nand UO_1457 (O_1457,N_9925,N_9961);
and UO_1458 (O_1458,N_9930,N_9957);
or UO_1459 (O_1459,N_9972,N_9952);
nor UO_1460 (O_1460,N_9958,N_9989);
or UO_1461 (O_1461,N_9922,N_9903);
nand UO_1462 (O_1462,N_9957,N_9945);
and UO_1463 (O_1463,N_9972,N_9954);
and UO_1464 (O_1464,N_9948,N_9925);
nor UO_1465 (O_1465,N_9945,N_9982);
or UO_1466 (O_1466,N_9980,N_9943);
nand UO_1467 (O_1467,N_9937,N_9953);
and UO_1468 (O_1468,N_9937,N_9965);
nor UO_1469 (O_1469,N_9925,N_9927);
nand UO_1470 (O_1470,N_9936,N_9949);
nand UO_1471 (O_1471,N_9965,N_9924);
nor UO_1472 (O_1472,N_9955,N_9928);
or UO_1473 (O_1473,N_9911,N_9983);
and UO_1474 (O_1474,N_9995,N_9936);
or UO_1475 (O_1475,N_9905,N_9953);
and UO_1476 (O_1476,N_9906,N_9982);
nor UO_1477 (O_1477,N_9900,N_9968);
xnor UO_1478 (O_1478,N_9962,N_9967);
nor UO_1479 (O_1479,N_9997,N_9991);
and UO_1480 (O_1480,N_9907,N_9974);
nand UO_1481 (O_1481,N_9970,N_9956);
and UO_1482 (O_1482,N_9953,N_9925);
nor UO_1483 (O_1483,N_9911,N_9904);
nor UO_1484 (O_1484,N_9950,N_9984);
and UO_1485 (O_1485,N_9914,N_9962);
nor UO_1486 (O_1486,N_9966,N_9987);
xor UO_1487 (O_1487,N_9963,N_9925);
nand UO_1488 (O_1488,N_9959,N_9926);
nor UO_1489 (O_1489,N_9955,N_9965);
nand UO_1490 (O_1490,N_9916,N_9907);
and UO_1491 (O_1491,N_9907,N_9976);
or UO_1492 (O_1492,N_9996,N_9945);
or UO_1493 (O_1493,N_9927,N_9939);
and UO_1494 (O_1494,N_9954,N_9991);
xor UO_1495 (O_1495,N_9955,N_9904);
and UO_1496 (O_1496,N_9991,N_9923);
and UO_1497 (O_1497,N_9978,N_9980);
nand UO_1498 (O_1498,N_9946,N_9966);
or UO_1499 (O_1499,N_9967,N_9941);
endmodule