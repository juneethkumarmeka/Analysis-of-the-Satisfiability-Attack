module basic_500_3000_500_3_levels_1xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nand U0 (N_0,In_21,In_484);
and U1 (N_1,In_96,In_115);
nor U2 (N_2,In_92,In_376);
nor U3 (N_3,In_10,In_150);
or U4 (N_4,In_4,In_226);
and U5 (N_5,In_128,In_318);
or U6 (N_6,In_240,In_109);
nor U7 (N_7,In_310,In_112);
nand U8 (N_8,In_17,In_33);
nand U9 (N_9,In_156,In_476);
nor U10 (N_10,In_397,In_371);
and U11 (N_11,In_111,In_389);
nor U12 (N_12,In_78,In_444);
or U13 (N_13,In_269,In_404);
or U14 (N_14,In_127,In_27);
and U15 (N_15,In_351,In_237);
nor U16 (N_16,In_315,In_171);
and U17 (N_17,In_295,In_222);
nor U18 (N_18,In_352,In_71);
nand U19 (N_19,In_448,In_451);
or U20 (N_20,In_428,In_79);
or U21 (N_21,In_192,In_375);
and U22 (N_22,In_392,In_436);
and U23 (N_23,In_7,In_415);
nor U24 (N_24,In_186,In_427);
nand U25 (N_25,In_348,In_316);
xor U26 (N_26,In_409,In_160);
nor U27 (N_27,In_104,In_234);
nand U28 (N_28,In_132,In_70);
and U29 (N_29,In_162,In_342);
nor U30 (N_30,In_44,In_252);
or U31 (N_31,In_187,In_144);
nor U32 (N_32,In_42,In_473);
or U33 (N_33,In_122,In_102);
nor U34 (N_34,In_277,In_370);
or U35 (N_35,In_307,In_378);
nor U36 (N_36,In_64,In_327);
nand U37 (N_37,In_204,In_218);
or U38 (N_38,In_282,In_168);
nand U39 (N_39,In_394,In_88);
or U40 (N_40,In_76,In_18);
or U41 (N_41,In_485,In_424);
nand U42 (N_42,In_221,In_408);
or U43 (N_43,In_421,In_301);
nor U44 (N_44,In_477,In_199);
nor U45 (N_45,In_442,In_113);
nor U46 (N_46,In_134,In_357);
nor U47 (N_47,In_154,In_490);
and U48 (N_48,In_180,In_114);
nand U49 (N_49,In_95,In_98);
nor U50 (N_50,In_124,In_437);
nor U51 (N_51,In_306,In_77);
nor U52 (N_52,In_243,In_135);
and U53 (N_53,In_280,In_432);
nand U54 (N_54,In_398,In_68);
nor U55 (N_55,In_125,In_82);
nor U56 (N_56,In_416,In_396);
and U57 (N_57,In_184,In_188);
nor U58 (N_58,In_23,In_67);
or U59 (N_59,In_49,In_89);
and U60 (N_60,In_36,In_145);
and U61 (N_61,In_469,In_429);
or U62 (N_62,In_495,In_201);
or U63 (N_63,In_94,In_69);
nor U64 (N_64,In_411,In_28);
nand U65 (N_65,In_385,In_37);
or U66 (N_66,In_219,In_236);
nand U67 (N_67,In_334,In_433);
nand U68 (N_68,In_208,In_337);
nor U69 (N_69,In_32,In_137);
or U70 (N_70,In_272,In_449);
or U71 (N_71,In_443,In_72);
and U72 (N_72,In_123,In_158);
and U73 (N_73,In_462,In_399);
or U74 (N_74,In_209,In_390);
and U75 (N_75,In_11,In_105);
nand U76 (N_76,In_231,In_80);
nor U77 (N_77,In_251,In_74);
and U78 (N_78,In_175,In_141);
nor U79 (N_79,In_482,In_294);
nor U80 (N_80,In_341,In_340);
nor U81 (N_81,In_143,In_212);
nor U82 (N_82,In_110,In_40);
nand U83 (N_83,In_202,In_383);
and U84 (N_84,In_87,In_139);
and U85 (N_85,In_138,In_459);
or U86 (N_86,In_321,In_229);
or U87 (N_87,In_312,In_285);
xor U88 (N_88,In_486,In_483);
or U89 (N_89,In_116,In_60);
xnor U90 (N_90,In_308,In_215);
nand U91 (N_91,In_107,In_176);
nand U92 (N_92,In_230,In_146);
or U93 (N_93,In_197,In_263);
or U94 (N_94,In_470,In_45);
nor U95 (N_95,In_129,In_13);
nor U96 (N_96,In_170,In_90);
nor U97 (N_97,In_386,In_254);
or U98 (N_98,In_338,In_480);
and U99 (N_99,In_468,In_172);
nand U100 (N_100,In_14,In_364);
or U101 (N_101,In_336,In_163);
xnor U102 (N_102,In_190,In_75);
nor U103 (N_103,In_25,In_493);
or U104 (N_104,In_99,In_346);
and U105 (N_105,In_270,In_50);
and U106 (N_106,In_46,In_302);
nor U107 (N_107,In_319,In_475);
or U108 (N_108,In_133,In_457);
or U109 (N_109,In_52,In_216);
nor U110 (N_110,In_178,In_496);
and U111 (N_111,In_401,In_494);
or U112 (N_112,In_273,In_498);
nor U113 (N_113,In_377,In_153);
nor U114 (N_114,In_425,In_29);
nand U115 (N_115,In_55,In_24);
and U116 (N_116,In_242,In_196);
and U117 (N_117,In_9,In_34);
and U118 (N_118,In_136,In_363);
nand U119 (N_119,In_12,In_265);
or U120 (N_120,In_245,In_15);
nor U121 (N_121,In_400,In_366);
or U122 (N_122,In_281,In_164);
or U123 (N_123,In_195,In_63);
and U124 (N_124,In_155,In_350);
and U125 (N_125,In_463,In_335);
and U126 (N_126,In_372,In_381);
or U127 (N_127,In_6,In_26);
nand U128 (N_128,In_311,In_380);
nor U129 (N_129,In_86,In_177);
or U130 (N_130,In_31,In_238);
and U131 (N_131,In_434,In_19);
or U132 (N_132,In_194,In_358);
and U133 (N_133,In_326,In_418);
nand U134 (N_134,In_499,In_174);
nand U135 (N_135,In_354,In_487);
nand U136 (N_136,In_304,In_165);
nor U137 (N_137,In_83,In_417);
and U138 (N_138,In_0,In_287);
nor U139 (N_139,In_183,In_330);
and U140 (N_140,In_467,In_289);
and U141 (N_141,In_262,In_291);
nand U142 (N_142,In_48,In_220);
or U143 (N_143,In_452,In_445);
nor U144 (N_144,In_349,In_423);
nand U145 (N_145,In_198,In_450);
nand U146 (N_146,In_465,In_157);
nand U147 (N_147,In_275,In_402);
and U148 (N_148,In_43,In_223);
or U149 (N_149,In_296,In_455);
or U150 (N_150,In_120,In_331);
nand U151 (N_151,In_447,In_439);
and U152 (N_152,In_393,In_413);
or U153 (N_153,In_461,In_322);
nor U154 (N_154,In_151,In_2);
or U155 (N_155,In_298,In_374);
or U156 (N_156,In_264,In_246);
and U157 (N_157,In_166,In_317);
or U158 (N_158,In_200,In_224);
or U159 (N_159,In_41,In_161);
nand U160 (N_160,In_347,In_206);
nor U161 (N_161,In_203,In_149);
nor U162 (N_162,In_20,In_121);
nand U163 (N_163,In_8,In_305);
nand U164 (N_164,In_456,In_57);
nor U165 (N_165,In_407,In_247);
nor U166 (N_166,In_403,In_148);
or U167 (N_167,In_103,In_359);
nand U168 (N_168,In_292,In_140);
nor U169 (N_169,In_241,In_474);
nor U170 (N_170,In_460,In_369);
or U171 (N_171,In_395,In_131);
nor U172 (N_172,In_259,In_379);
nand U173 (N_173,In_293,In_119);
nor U174 (N_174,In_339,In_384);
and U175 (N_175,In_313,In_446);
and U176 (N_176,In_274,In_492);
nor U177 (N_177,In_333,In_478);
or U178 (N_178,In_300,In_320);
nand U179 (N_179,In_497,In_152);
nor U180 (N_180,In_53,In_325);
nor U181 (N_181,In_343,In_278);
and U182 (N_182,In_235,In_472);
nand U183 (N_183,In_426,In_205);
or U184 (N_184,In_440,In_249);
or U185 (N_185,In_16,In_388);
nor U186 (N_186,In_430,In_435);
and U187 (N_187,In_173,In_51);
nand U188 (N_188,In_458,In_182);
nor U189 (N_189,In_466,In_362);
nor U190 (N_190,In_117,In_367);
and U191 (N_191,In_189,In_248);
and U192 (N_192,In_286,In_232);
nand U193 (N_193,In_169,In_260);
nor U194 (N_194,In_167,In_299);
nor U195 (N_195,In_382,In_39);
or U196 (N_196,In_422,In_332);
nor U197 (N_197,In_453,In_211);
and U198 (N_198,In_279,In_35);
or U199 (N_199,In_214,In_159);
and U200 (N_200,In_360,In_288);
nand U201 (N_201,In_329,In_431);
nand U202 (N_202,In_181,In_207);
and U203 (N_203,In_387,In_276);
nand U204 (N_204,In_66,In_97);
nor U205 (N_205,In_420,In_5);
or U206 (N_206,In_62,In_85);
nor U207 (N_207,In_227,In_344);
and U208 (N_208,In_323,In_479);
and U209 (N_209,In_1,In_59);
nor U210 (N_210,In_65,In_142);
or U211 (N_211,In_283,In_257);
or U212 (N_212,In_22,In_255);
or U213 (N_213,In_253,In_258);
nor U214 (N_214,In_73,In_38);
nand U215 (N_215,In_353,In_324);
and U216 (N_216,In_438,In_250);
nand U217 (N_217,In_3,In_419);
or U218 (N_218,In_213,In_271);
and U219 (N_219,In_108,In_217);
nand U220 (N_220,In_30,In_489);
or U221 (N_221,In_126,In_410);
nor U222 (N_222,In_373,In_365);
or U223 (N_223,In_328,In_488);
nor U224 (N_224,In_54,In_361);
and U225 (N_225,In_355,In_290);
nor U226 (N_226,In_309,In_441);
or U227 (N_227,In_284,In_391);
and U228 (N_228,In_147,In_93);
and U229 (N_229,In_47,In_210);
and U230 (N_230,In_101,In_481);
nand U231 (N_231,In_228,In_58);
nand U232 (N_232,In_406,In_61);
nor U233 (N_233,In_100,In_454);
or U234 (N_234,In_261,In_84);
or U235 (N_235,In_191,In_356);
or U236 (N_236,In_244,In_297);
nand U237 (N_237,In_368,In_268);
or U238 (N_238,In_314,In_405);
or U239 (N_239,In_81,In_193);
or U240 (N_240,In_239,In_225);
nand U241 (N_241,In_303,In_106);
nand U242 (N_242,In_412,In_91);
nand U243 (N_243,In_464,In_118);
nor U244 (N_244,In_256,In_471);
nand U245 (N_245,In_179,In_267);
or U246 (N_246,In_266,In_491);
or U247 (N_247,In_185,In_56);
or U248 (N_248,In_345,In_130);
nand U249 (N_249,In_233,In_414);
nor U250 (N_250,In_426,In_87);
nand U251 (N_251,In_155,In_493);
nor U252 (N_252,In_205,In_451);
and U253 (N_253,In_132,In_385);
or U254 (N_254,In_306,In_303);
nor U255 (N_255,In_438,In_407);
nor U256 (N_256,In_227,In_399);
and U257 (N_257,In_495,In_215);
or U258 (N_258,In_164,In_363);
nor U259 (N_259,In_100,In_1);
nor U260 (N_260,In_457,In_415);
nand U261 (N_261,In_148,In_70);
nand U262 (N_262,In_206,In_87);
nor U263 (N_263,In_288,In_261);
nand U264 (N_264,In_430,In_331);
nand U265 (N_265,In_447,In_311);
nand U266 (N_266,In_150,In_307);
nor U267 (N_267,In_327,In_142);
nor U268 (N_268,In_465,In_103);
and U269 (N_269,In_95,In_450);
nand U270 (N_270,In_204,In_117);
nand U271 (N_271,In_27,In_419);
nand U272 (N_272,In_145,In_415);
nor U273 (N_273,In_119,In_10);
and U274 (N_274,In_28,In_159);
nand U275 (N_275,In_348,In_371);
and U276 (N_276,In_205,In_210);
or U277 (N_277,In_21,In_18);
nor U278 (N_278,In_24,In_247);
or U279 (N_279,In_87,In_41);
and U280 (N_280,In_240,In_285);
nand U281 (N_281,In_252,In_177);
and U282 (N_282,In_491,In_483);
nor U283 (N_283,In_367,In_148);
and U284 (N_284,In_411,In_21);
or U285 (N_285,In_272,In_393);
nor U286 (N_286,In_202,In_339);
nand U287 (N_287,In_267,In_171);
and U288 (N_288,In_427,In_343);
nor U289 (N_289,In_428,In_469);
nand U290 (N_290,In_477,In_207);
nand U291 (N_291,In_258,In_231);
nor U292 (N_292,In_265,In_39);
nor U293 (N_293,In_231,In_305);
nand U294 (N_294,In_481,In_188);
nor U295 (N_295,In_216,In_323);
or U296 (N_296,In_14,In_176);
or U297 (N_297,In_243,In_469);
nor U298 (N_298,In_486,In_295);
nor U299 (N_299,In_237,In_418);
nand U300 (N_300,In_283,In_284);
and U301 (N_301,In_67,In_346);
nor U302 (N_302,In_312,In_194);
and U303 (N_303,In_491,In_200);
and U304 (N_304,In_94,In_100);
and U305 (N_305,In_347,In_331);
or U306 (N_306,In_329,In_217);
nand U307 (N_307,In_436,In_263);
nand U308 (N_308,In_280,In_212);
nor U309 (N_309,In_458,In_301);
nor U310 (N_310,In_100,In_270);
nor U311 (N_311,In_408,In_340);
and U312 (N_312,In_127,In_238);
and U313 (N_313,In_347,In_110);
or U314 (N_314,In_23,In_380);
nor U315 (N_315,In_100,In_71);
and U316 (N_316,In_394,In_85);
nor U317 (N_317,In_328,In_214);
nor U318 (N_318,In_52,In_364);
or U319 (N_319,In_5,In_83);
and U320 (N_320,In_328,In_74);
nor U321 (N_321,In_485,In_366);
and U322 (N_322,In_111,In_476);
or U323 (N_323,In_383,In_376);
nand U324 (N_324,In_177,In_231);
nor U325 (N_325,In_154,In_62);
or U326 (N_326,In_92,In_77);
nor U327 (N_327,In_252,In_426);
and U328 (N_328,In_10,In_445);
nor U329 (N_329,In_55,In_74);
and U330 (N_330,In_28,In_339);
or U331 (N_331,In_245,In_186);
nor U332 (N_332,In_400,In_214);
and U333 (N_333,In_139,In_38);
nor U334 (N_334,In_82,In_14);
nor U335 (N_335,In_237,In_41);
or U336 (N_336,In_204,In_485);
nor U337 (N_337,In_113,In_288);
nor U338 (N_338,In_261,In_140);
or U339 (N_339,In_409,In_202);
nor U340 (N_340,In_137,In_495);
nand U341 (N_341,In_327,In_382);
and U342 (N_342,In_10,In_453);
nor U343 (N_343,In_160,In_463);
or U344 (N_344,In_499,In_134);
nand U345 (N_345,In_350,In_113);
nor U346 (N_346,In_482,In_168);
or U347 (N_347,In_115,In_340);
nor U348 (N_348,In_385,In_396);
or U349 (N_349,In_332,In_474);
nor U350 (N_350,In_183,In_336);
nand U351 (N_351,In_314,In_238);
nand U352 (N_352,In_76,In_363);
and U353 (N_353,In_2,In_38);
or U354 (N_354,In_172,In_200);
nand U355 (N_355,In_485,In_201);
and U356 (N_356,In_174,In_455);
nand U357 (N_357,In_402,In_37);
nand U358 (N_358,In_231,In_105);
and U359 (N_359,In_428,In_230);
or U360 (N_360,In_48,In_288);
nor U361 (N_361,In_59,In_211);
nor U362 (N_362,In_492,In_406);
or U363 (N_363,In_345,In_108);
nor U364 (N_364,In_441,In_115);
or U365 (N_365,In_396,In_44);
nor U366 (N_366,In_417,In_286);
nand U367 (N_367,In_401,In_2);
nor U368 (N_368,In_62,In_319);
nor U369 (N_369,In_28,In_25);
or U370 (N_370,In_360,In_46);
nor U371 (N_371,In_231,In_494);
nor U372 (N_372,In_148,In_358);
xor U373 (N_373,In_19,In_478);
or U374 (N_374,In_114,In_168);
and U375 (N_375,In_455,In_113);
and U376 (N_376,In_338,In_353);
and U377 (N_377,In_439,In_204);
nor U378 (N_378,In_422,In_198);
nand U379 (N_379,In_193,In_332);
and U380 (N_380,In_439,In_404);
and U381 (N_381,In_162,In_254);
and U382 (N_382,In_2,In_261);
or U383 (N_383,In_42,In_429);
nand U384 (N_384,In_285,In_315);
or U385 (N_385,In_346,In_73);
or U386 (N_386,In_301,In_26);
or U387 (N_387,In_426,In_338);
and U388 (N_388,In_193,In_425);
nand U389 (N_389,In_95,In_290);
or U390 (N_390,In_287,In_474);
nand U391 (N_391,In_467,In_278);
and U392 (N_392,In_1,In_163);
and U393 (N_393,In_237,In_75);
nor U394 (N_394,In_414,In_62);
and U395 (N_395,In_479,In_391);
and U396 (N_396,In_14,In_207);
and U397 (N_397,In_484,In_452);
nor U398 (N_398,In_63,In_133);
nand U399 (N_399,In_391,In_303);
and U400 (N_400,In_108,In_202);
nand U401 (N_401,In_130,In_69);
and U402 (N_402,In_335,In_259);
and U403 (N_403,In_123,In_183);
nor U404 (N_404,In_453,In_140);
nor U405 (N_405,In_81,In_177);
nand U406 (N_406,In_107,In_143);
and U407 (N_407,In_44,In_486);
or U408 (N_408,In_370,In_166);
and U409 (N_409,In_466,In_227);
or U410 (N_410,In_179,In_155);
and U411 (N_411,In_154,In_119);
nor U412 (N_412,In_266,In_125);
nor U413 (N_413,In_491,In_394);
nor U414 (N_414,In_86,In_337);
and U415 (N_415,In_429,In_366);
and U416 (N_416,In_288,In_55);
or U417 (N_417,In_335,In_467);
nand U418 (N_418,In_184,In_304);
nand U419 (N_419,In_465,In_458);
and U420 (N_420,In_376,In_307);
or U421 (N_421,In_483,In_239);
and U422 (N_422,In_253,In_35);
and U423 (N_423,In_26,In_2);
and U424 (N_424,In_24,In_489);
and U425 (N_425,In_395,In_33);
or U426 (N_426,In_220,In_158);
or U427 (N_427,In_142,In_127);
nand U428 (N_428,In_266,In_176);
or U429 (N_429,In_358,In_186);
nor U430 (N_430,In_461,In_425);
nand U431 (N_431,In_19,In_273);
and U432 (N_432,In_91,In_245);
or U433 (N_433,In_90,In_384);
and U434 (N_434,In_428,In_496);
nand U435 (N_435,In_253,In_288);
nand U436 (N_436,In_275,In_354);
nor U437 (N_437,In_446,In_172);
or U438 (N_438,In_209,In_461);
nand U439 (N_439,In_334,In_359);
nor U440 (N_440,In_132,In_21);
nor U441 (N_441,In_203,In_463);
and U442 (N_442,In_242,In_373);
nand U443 (N_443,In_57,In_31);
nor U444 (N_444,In_166,In_499);
nor U445 (N_445,In_445,In_350);
nand U446 (N_446,In_481,In_166);
nand U447 (N_447,In_397,In_144);
nor U448 (N_448,In_307,In_275);
and U449 (N_449,In_425,In_334);
nor U450 (N_450,In_222,In_211);
and U451 (N_451,In_5,In_250);
and U452 (N_452,In_390,In_170);
or U453 (N_453,In_98,In_225);
or U454 (N_454,In_252,In_145);
or U455 (N_455,In_351,In_384);
and U456 (N_456,In_62,In_358);
or U457 (N_457,In_404,In_437);
nand U458 (N_458,In_294,In_106);
and U459 (N_459,In_125,In_45);
nor U460 (N_460,In_107,In_251);
nand U461 (N_461,In_172,In_202);
nand U462 (N_462,In_325,In_373);
or U463 (N_463,In_422,In_262);
nand U464 (N_464,In_497,In_388);
or U465 (N_465,In_361,In_294);
and U466 (N_466,In_33,In_428);
or U467 (N_467,In_59,In_330);
or U468 (N_468,In_343,In_447);
nor U469 (N_469,In_400,In_249);
nor U470 (N_470,In_451,In_250);
nor U471 (N_471,In_479,In_225);
nor U472 (N_472,In_246,In_483);
nand U473 (N_473,In_266,In_156);
or U474 (N_474,In_45,In_213);
nand U475 (N_475,In_45,In_414);
or U476 (N_476,In_208,In_435);
nand U477 (N_477,In_79,In_289);
nor U478 (N_478,In_11,In_197);
nor U479 (N_479,In_439,In_448);
or U480 (N_480,In_299,In_247);
nor U481 (N_481,In_219,In_471);
nand U482 (N_482,In_276,In_102);
or U483 (N_483,In_64,In_283);
nor U484 (N_484,In_350,In_136);
or U485 (N_485,In_456,In_231);
or U486 (N_486,In_114,In_22);
and U487 (N_487,In_55,In_79);
nor U488 (N_488,In_118,In_141);
nor U489 (N_489,In_291,In_159);
nor U490 (N_490,In_123,In_420);
or U491 (N_491,In_227,In_131);
nand U492 (N_492,In_176,In_434);
and U493 (N_493,In_320,In_447);
xor U494 (N_494,In_310,In_6);
nand U495 (N_495,In_392,In_334);
or U496 (N_496,In_121,In_357);
and U497 (N_497,In_282,In_55);
and U498 (N_498,In_88,In_23);
nor U499 (N_499,In_220,In_182);
or U500 (N_500,In_172,In_270);
or U501 (N_501,In_181,In_281);
and U502 (N_502,In_349,In_396);
and U503 (N_503,In_113,In_328);
nor U504 (N_504,In_44,In_248);
nor U505 (N_505,In_44,In_463);
or U506 (N_506,In_219,In_268);
nand U507 (N_507,In_166,In_263);
or U508 (N_508,In_127,In_375);
and U509 (N_509,In_166,In_491);
nand U510 (N_510,In_185,In_199);
or U511 (N_511,In_446,In_233);
and U512 (N_512,In_366,In_187);
nor U513 (N_513,In_32,In_239);
nor U514 (N_514,In_5,In_43);
nand U515 (N_515,In_89,In_117);
nand U516 (N_516,In_439,In_36);
and U517 (N_517,In_383,In_419);
and U518 (N_518,In_0,In_270);
and U519 (N_519,In_452,In_228);
nand U520 (N_520,In_436,In_17);
or U521 (N_521,In_25,In_121);
nor U522 (N_522,In_268,In_497);
nand U523 (N_523,In_322,In_447);
nor U524 (N_524,In_361,In_485);
or U525 (N_525,In_73,In_388);
nand U526 (N_526,In_284,In_328);
and U527 (N_527,In_497,In_102);
nor U528 (N_528,In_45,In_354);
and U529 (N_529,In_426,In_310);
or U530 (N_530,In_104,In_345);
or U531 (N_531,In_468,In_477);
nor U532 (N_532,In_72,In_317);
nor U533 (N_533,In_169,In_439);
or U534 (N_534,In_358,In_426);
or U535 (N_535,In_41,In_84);
and U536 (N_536,In_264,In_100);
nand U537 (N_537,In_336,In_421);
and U538 (N_538,In_22,In_373);
and U539 (N_539,In_29,In_175);
and U540 (N_540,In_310,In_432);
or U541 (N_541,In_327,In_220);
or U542 (N_542,In_388,In_120);
nor U543 (N_543,In_211,In_54);
or U544 (N_544,In_152,In_146);
nor U545 (N_545,In_138,In_93);
nor U546 (N_546,In_283,In_101);
nor U547 (N_547,In_27,In_413);
and U548 (N_548,In_405,In_123);
nand U549 (N_549,In_335,In_273);
or U550 (N_550,In_409,In_200);
nand U551 (N_551,In_284,In_288);
nand U552 (N_552,In_97,In_327);
nor U553 (N_553,In_399,In_445);
xor U554 (N_554,In_254,In_18);
nor U555 (N_555,In_485,In_496);
or U556 (N_556,In_16,In_229);
nor U557 (N_557,In_86,In_479);
nand U558 (N_558,In_165,In_294);
and U559 (N_559,In_339,In_26);
nand U560 (N_560,In_348,In_451);
and U561 (N_561,In_347,In_440);
nand U562 (N_562,In_182,In_439);
nor U563 (N_563,In_330,In_84);
nand U564 (N_564,In_488,In_427);
and U565 (N_565,In_48,In_298);
or U566 (N_566,In_263,In_156);
or U567 (N_567,In_476,In_329);
and U568 (N_568,In_198,In_257);
nor U569 (N_569,In_101,In_202);
and U570 (N_570,In_309,In_158);
or U571 (N_571,In_36,In_75);
nand U572 (N_572,In_192,In_13);
and U573 (N_573,In_271,In_225);
or U574 (N_574,In_179,In_58);
or U575 (N_575,In_466,In_376);
and U576 (N_576,In_0,In_159);
nor U577 (N_577,In_456,In_4);
or U578 (N_578,In_385,In_455);
or U579 (N_579,In_378,In_253);
nor U580 (N_580,In_157,In_237);
nor U581 (N_581,In_54,In_34);
nor U582 (N_582,In_333,In_28);
or U583 (N_583,In_135,In_27);
and U584 (N_584,In_100,In_287);
and U585 (N_585,In_243,In_16);
or U586 (N_586,In_56,In_45);
and U587 (N_587,In_207,In_42);
and U588 (N_588,In_327,In_9);
or U589 (N_589,In_253,In_350);
or U590 (N_590,In_429,In_339);
and U591 (N_591,In_22,In_38);
and U592 (N_592,In_241,In_33);
nor U593 (N_593,In_340,In_461);
nor U594 (N_594,In_188,In_457);
nor U595 (N_595,In_233,In_478);
or U596 (N_596,In_51,In_151);
nand U597 (N_597,In_3,In_51);
nand U598 (N_598,In_189,In_81);
and U599 (N_599,In_174,In_82);
nor U600 (N_600,In_381,In_358);
or U601 (N_601,In_387,In_23);
nor U602 (N_602,In_49,In_462);
nor U603 (N_603,In_370,In_453);
and U604 (N_604,In_482,In_241);
nor U605 (N_605,In_229,In_428);
and U606 (N_606,In_156,In_268);
or U607 (N_607,In_452,In_495);
or U608 (N_608,In_94,In_387);
xnor U609 (N_609,In_31,In_364);
nor U610 (N_610,In_419,In_491);
and U611 (N_611,In_207,In_219);
and U612 (N_612,In_127,In_228);
nor U613 (N_613,In_387,In_275);
nand U614 (N_614,In_195,In_374);
nor U615 (N_615,In_35,In_1);
and U616 (N_616,In_368,In_482);
nor U617 (N_617,In_304,In_9);
and U618 (N_618,In_488,In_158);
or U619 (N_619,In_333,In_487);
nand U620 (N_620,In_298,In_138);
and U621 (N_621,In_38,In_417);
nand U622 (N_622,In_109,In_216);
nand U623 (N_623,In_425,In_429);
nand U624 (N_624,In_152,In_142);
nor U625 (N_625,In_376,In_478);
or U626 (N_626,In_72,In_312);
or U627 (N_627,In_12,In_396);
and U628 (N_628,In_271,In_434);
nor U629 (N_629,In_387,In_393);
nor U630 (N_630,In_20,In_43);
nor U631 (N_631,In_242,In_389);
and U632 (N_632,In_322,In_330);
nor U633 (N_633,In_345,In_284);
or U634 (N_634,In_0,In_335);
nor U635 (N_635,In_70,In_401);
or U636 (N_636,In_75,In_9);
or U637 (N_637,In_287,In_244);
xor U638 (N_638,In_212,In_186);
nand U639 (N_639,In_122,In_493);
nor U640 (N_640,In_267,In_78);
and U641 (N_641,In_465,In_301);
and U642 (N_642,In_439,In_77);
nand U643 (N_643,In_419,In_70);
and U644 (N_644,In_95,In_293);
and U645 (N_645,In_117,In_245);
or U646 (N_646,In_9,In_21);
or U647 (N_647,In_198,In_310);
nor U648 (N_648,In_344,In_473);
or U649 (N_649,In_113,In_275);
nand U650 (N_650,In_55,In_180);
and U651 (N_651,In_182,In_273);
nand U652 (N_652,In_360,In_16);
nand U653 (N_653,In_110,In_57);
xor U654 (N_654,In_474,In_164);
nor U655 (N_655,In_313,In_404);
nand U656 (N_656,In_438,In_276);
nand U657 (N_657,In_472,In_490);
or U658 (N_658,In_300,In_310);
nand U659 (N_659,In_121,In_440);
nor U660 (N_660,In_26,In_357);
nor U661 (N_661,In_125,In_185);
and U662 (N_662,In_334,In_294);
and U663 (N_663,In_306,In_388);
nor U664 (N_664,In_21,In_326);
or U665 (N_665,In_244,In_448);
nand U666 (N_666,In_394,In_481);
nand U667 (N_667,In_381,In_91);
and U668 (N_668,In_99,In_410);
nor U669 (N_669,In_138,In_325);
and U670 (N_670,In_235,In_227);
nor U671 (N_671,In_364,In_189);
or U672 (N_672,In_398,In_283);
nand U673 (N_673,In_229,In_98);
and U674 (N_674,In_141,In_158);
nand U675 (N_675,In_485,In_190);
nor U676 (N_676,In_313,In_127);
or U677 (N_677,In_483,In_186);
xor U678 (N_678,In_139,In_239);
and U679 (N_679,In_473,In_82);
nand U680 (N_680,In_53,In_195);
nand U681 (N_681,In_485,In_105);
nor U682 (N_682,In_211,In_147);
and U683 (N_683,In_106,In_435);
nand U684 (N_684,In_436,In_85);
nand U685 (N_685,In_361,In_130);
nand U686 (N_686,In_100,In_88);
nor U687 (N_687,In_411,In_164);
or U688 (N_688,In_408,In_144);
or U689 (N_689,In_203,In_484);
or U690 (N_690,In_112,In_202);
or U691 (N_691,In_453,In_318);
or U692 (N_692,In_183,In_286);
nand U693 (N_693,In_345,In_395);
nand U694 (N_694,In_160,In_189);
or U695 (N_695,In_7,In_180);
or U696 (N_696,In_128,In_419);
or U697 (N_697,In_149,In_369);
or U698 (N_698,In_57,In_203);
and U699 (N_699,In_30,In_343);
or U700 (N_700,In_85,In_270);
nand U701 (N_701,In_304,In_140);
nor U702 (N_702,In_126,In_254);
and U703 (N_703,In_268,In_226);
nor U704 (N_704,In_255,In_421);
and U705 (N_705,In_154,In_57);
nor U706 (N_706,In_289,In_250);
and U707 (N_707,In_119,In_100);
nand U708 (N_708,In_459,In_156);
xor U709 (N_709,In_174,In_485);
or U710 (N_710,In_419,In_92);
nand U711 (N_711,In_89,In_364);
or U712 (N_712,In_411,In_354);
nor U713 (N_713,In_268,In_168);
nand U714 (N_714,In_94,In_420);
and U715 (N_715,In_56,In_474);
nand U716 (N_716,In_464,In_160);
nor U717 (N_717,In_57,In_158);
or U718 (N_718,In_209,In_160);
nor U719 (N_719,In_453,In_81);
nand U720 (N_720,In_290,In_415);
or U721 (N_721,In_120,In_407);
and U722 (N_722,In_220,In_419);
nand U723 (N_723,In_114,In_222);
or U724 (N_724,In_86,In_343);
nand U725 (N_725,In_11,In_31);
nor U726 (N_726,In_154,In_197);
and U727 (N_727,In_402,In_23);
nor U728 (N_728,In_441,In_119);
or U729 (N_729,In_330,In_253);
and U730 (N_730,In_409,In_162);
nor U731 (N_731,In_437,In_168);
nor U732 (N_732,In_61,In_203);
and U733 (N_733,In_58,In_216);
and U734 (N_734,In_413,In_482);
and U735 (N_735,In_197,In_7);
or U736 (N_736,In_50,In_499);
or U737 (N_737,In_455,In_51);
and U738 (N_738,In_78,In_367);
or U739 (N_739,In_68,In_480);
or U740 (N_740,In_193,In_39);
nor U741 (N_741,In_275,In_483);
or U742 (N_742,In_115,In_409);
or U743 (N_743,In_299,In_185);
nand U744 (N_744,In_312,In_149);
nand U745 (N_745,In_191,In_460);
and U746 (N_746,In_4,In_170);
and U747 (N_747,In_456,In_492);
nor U748 (N_748,In_90,In_345);
nor U749 (N_749,In_50,In_183);
nand U750 (N_750,In_177,In_101);
or U751 (N_751,In_130,In_151);
nand U752 (N_752,In_55,In_199);
or U753 (N_753,In_465,In_166);
or U754 (N_754,In_474,In_347);
or U755 (N_755,In_275,In_392);
nand U756 (N_756,In_416,In_323);
and U757 (N_757,In_469,In_495);
or U758 (N_758,In_222,In_371);
and U759 (N_759,In_233,In_382);
or U760 (N_760,In_357,In_170);
nand U761 (N_761,In_368,In_230);
and U762 (N_762,In_116,In_271);
nand U763 (N_763,In_239,In_87);
and U764 (N_764,In_57,In_229);
or U765 (N_765,In_72,In_409);
nor U766 (N_766,In_38,In_333);
nor U767 (N_767,In_83,In_382);
or U768 (N_768,In_232,In_10);
or U769 (N_769,In_7,In_476);
or U770 (N_770,In_27,In_71);
nor U771 (N_771,In_341,In_435);
nand U772 (N_772,In_52,In_386);
and U773 (N_773,In_179,In_169);
and U774 (N_774,In_472,In_282);
nor U775 (N_775,In_284,In_443);
and U776 (N_776,In_394,In_121);
xnor U777 (N_777,In_271,In_370);
nor U778 (N_778,In_382,In_137);
nand U779 (N_779,In_280,In_133);
and U780 (N_780,In_400,In_158);
and U781 (N_781,In_146,In_201);
nor U782 (N_782,In_170,In_449);
and U783 (N_783,In_336,In_23);
or U784 (N_784,In_107,In_248);
nor U785 (N_785,In_249,In_212);
xnor U786 (N_786,In_274,In_358);
and U787 (N_787,In_264,In_272);
and U788 (N_788,In_90,In_368);
and U789 (N_789,In_16,In_444);
nand U790 (N_790,In_50,In_241);
nand U791 (N_791,In_203,In_382);
nand U792 (N_792,In_219,In_159);
or U793 (N_793,In_382,In_230);
and U794 (N_794,In_194,In_140);
nor U795 (N_795,In_472,In_497);
and U796 (N_796,In_162,In_458);
nor U797 (N_797,In_206,In_399);
nand U798 (N_798,In_489,In_271);
nor U799 (N_799,In_144,In_457);
or U800 (N_800,In_100,In_194);
and U801 (N_801,In_85,In_328);
and U802 (N_802,In_162,In_391);
nor U803 (N_803,In_169,In_358);
or U804 (N_804,In_243,In_141);
and U805 (N_805,In_289,In_21);
or U806 (N_806,In_187,In_412);
or U807 (N_807,In_42,In_431);
and U808 (N_808,In_155,In_277);
nor U809 (N_809,In_168,In_337);
and U810 (N_810,In_326,In_127);
or U811 (N_811,In_336,In_76);
nor U812 (N_812,In_319,In_109);
nor U813 (N_813,In_175,In_323);
and U814 (N_814,In_17,In_487);
or U815 (N_815,In_446,In_418);
nor U816 (N_816,In_52,In_349);
nor U817 (N_817,In_223,In_182);
nor U818 (N_818,In_413,In_132);
nand U819 (N_819,In_231,In_420);
nand U820 (N_820,In_406,In_374);
or U821 (N_821,In_209,In_93);
and U822 (N_822,In_440,In_329);
and U823 (N_823,In_297,In_196);
nand U824 (N_824,In_327,In_486);
nand U825 (N_825,In_112,In_232);
and U826 (N_826,In_46,In_222);
nand U827 (N_827,In_152,In_202);
and U828 (N_828,In_2,In_379);
and U829 (N_829,In_189,In_343);
nand U830 (N_830,In_473,In_316);
and U831 (N_831,In_104,In_334);
nor U832 (N_832,In_12,In_415);
and U833 (N_833,In_157,In_490);
nor U834 (N_834,In_31,In_379);
nand U835 (N_835,In_427,In_449);
or U836 (N_836,In_266,In_131);
and U837 (N_837,In_304,In_382);
and U838 (N_838,In_197,In_214);
nand U839 (N_839,In_51,In_311);
and U840 (N_840,In_440,In_310);
and U841 (N_841,In_164,In_130);
or U842 (N_842,In_425,In_101);
nor U843 (N_843,In_98,In_44);
nand U844 (N_844,In_174,In_52);
or U845 (N_845,In_194,In_237);
or U846 (N_846,In_116,In_378);
xnor U847 (N_847,In_83,In_394);
or U848 (N_848,In_484,In_167);
or U849 (N_849,In_389,In_289);
nand U850 (N_850,In_218,In_73);
nor U851 (N_851,In_188,In_80);
nor U852 (N_852,In_41,In_392);
xor U853 (N_853,In_325,In_128);
nand U854 (N_854,In_338,In_416);
nor U855 (N_855,In_247,In_109);
nand U856 (N_856,In_106,In_181);
xnor U857 (N_857,In_183,In_454);
or U858 (N_858,In_162,In_157);
nor U859 (N_859,In_411,In_290);
and U860 (N_860,In_244,In_146);
nand U861 (N_861,In_451,In_382);
nor U862 (N_862,In_57,In_243);
nor U863 (N_863,In_312,In_212);
or U864 (N_864,In_41,In_313);
or U865 (N_865,In_293,In_277);
and U866 (N_866,In_424,In_378);
nor U867 (N_867,In_370,In_371);
nand U868 (N_868,In_465,In_96);
or U869 (N_869,In_431,In_46);
and U870 (N_870,In_259,In_441);
nor U871 (N_871,In_381,In_397);
nor U872 (N_872,In_85,In_268);
nand U873 (N_873,In_193,In_308);
or U874 (N_874,In_254,In_11);
and U875 (N_875,In_337,In_201);
or U876 (N_876,In_448,In_18);
nor U877 (N_877,In_114,In_322);
or U878 (N_878,In_441,In_249);
or U879 (N_879,In_93,In_326);
nor U880 (N_880,In_164,In_40);
and U881 (N_881,In_247,In_438);
or U882 (N_882,In_204,In_115);
and U883 (N_883,In_30,In_307);
and U884 (N_884,In_214,In_47);
nor U885 (N_885,In_30,In_444);
nor U886 (N_886,In_206,In_392);
nand U887 (N_887,In_113,In_463);
nand U888 (N_888,In_59,In_285);
and U889 (N_889,In_205,In_270);
nand U890 (N_890,In_494,In_133);
or U891 (N_891,In_69,In_238);
and U892 (N_892,In_476,In_178);
or U893 (N_893,In_494,In_144);
and U894 (N_894,In_215,In_331);
nor U895 (N_895,In_94,In_158);
or U896 (N_896,In_42,In_482);
and U897 (N_897,In_354,In_173);
or U898 (N_898,In_388,In_298);
or U899 (N_899,In_399,In_137);
or U900 (N_900,In_317,In_439);
nor U901 (N_901,In_293,In_60);
nor U902 (N_902,In_396,In_75);
nand U903 (N_903,In_231,In_57);
or U904 (N_904,In_396,In_26);
nor U905 (N_905,In_109,In_169);
and U906 (N_906,In_207,In_334);
and U907 (N_907,In_32,In_411);
or U908 (N_908,In_68,In_37);
and U909 (N_909,In_157,In_351);
nand U910 (N_910,In_47,In_473);
and U911 (N_911,In_53,In_171);
xor U912 (N_912,In_236,In_54);
and U913 (N_913,In_173,In_322);
nand U914 (N_914,In_67,In_130);
nand U915 (N_915,In_453,In_462);
and U916 (N_916,In_82,In_496);
nor U917 (N_917,In_374,In_349);
or U918 (N_918,In_76,In_136);
nor U919 (N_919,In_22,In_298);
and U920 (N_920,In_75,In_394);
and U921 (N_921,In_0,In_266);
xor U922 (N_922,In_53,In_297);
or U923 (N_923,In_366,In_8);
nor U924 (N_924,In_220,In_280);
nor U925 (N_925,In_494,In_230);
nand U926 (N_926,In_460,In_316);
or U927 (N_927,In_495,In_366);
nand U928 (N_928,In_470,In_443);
nand U929 (N_929,In_479,In_314);
nand U930 (N_930,In_253,In_139);
nand U931 (N_931,In_59,In_134);
nor U932 (N_932,In_65,In_467);
or U933 (N_933,In_21,In_61);
and U934 (N_934,In_77,In_312);
nor U935 (N_935,In_485,In_281);
or U936 (N_936,In_87,In_38);
nor U937 (N_937,In_484,In_206);
nor U938 (N_938,In_77,In_78);
or U939 (N_939,In_248,In_282);
xnor U940 (N_940,In_12,In_111);
or U941 (N_941,In_195,In_201);
nor U942 (N_942,In_216,In_170);
nor U943 (N_943,In_57,In_189);
and U944 (N_944,In_114,In_198);
nand U945 (N_945,In_207,In_432);
and U946 (N_946,In_116,In_39);
or U947 (N_947,In_484,In_360);
and U948 (N_948,In_358,In_219);
nand U949 (N_949,In_294,In_179);
or U950 (N_950,In_50,In_37);
nand U951 (N_951,In_84,In_110);
nor U952 (N_952,In_253,In_468);
and U953 (N_953,In_476,In_250);
or U954 (N_954,In_363,In_427);
nand U955 (N_955,In_329,In_322);
nand U956 (N_956,In_62,In_42);
nor U957 (N_957,In_342,In_144);
and U958 (N_958,In_126,In_496);
and U959 (N_959,In_385,In_162);
and U960 (N_960,In_240,In_185);
nand U961 (N_961,In_447,In_193);
and U962 (N_962,In_418,In_152);
and U963 (N_963,In_91,In_109);
or U964 (N_964,In_82,In_208);
and U965 (N_965,In_118,In_155);
nand U966 (N_966,In_35,In_212);
and U967 (N_967,In_122,In_464);
and U968 (N_968,In_210,In_75);
and U969 (N_969,In_321,In_176);
nor U970 (N_970,In_314,In_155);
and U971 (N_971,In_474,In_387);
and U972 (N_972,In_240,In_448);
and U973 (N_973,In_79,In_479);
and U974 (N_974,In_138,In_492);
or U975 (N_975,In_27,In_310);
nand U976 (N_976,In_306,In_311);
and U977 (N_977,In_299,In_395);
nor U978 (N_978,In_214,In_136);
or U979 (N_979,In_115,In_356);
nor U980 (N_980,In_498,In_230);
nor U981 (N_981,In_122,In_148);
or U982 (N_982,In_281,In_56);
and U983 (N_983,In_489,In_35);
nand U984 (N_984,In_492,In_318);
nor U985 (N_985,In_185,In_2);
or U986 (N_986,In_336,In_27);
or U987 (N_987,In_46,In_451);
nand U988 (N_988,In_24,In_314);
or U989 (N_989,In_97,In_272);
or U990 (N_990,In_276,In_292);
or U991 (N_991,In_499,In_225);
nor U992 (N_992,In_264,In_350);
and U993 (N_993,In_63,In_425);
and U994 (N_994,In_194,In_86);
or U995 (N_995,In_141,In_161);
nor U996 (N_996,In_115,In_466);
or U997 (N_997,In_409,In_18);
nor U998 (N_998,In_295,In_420);
nor U999 (N_999,In_75,In_334);
and U1000 (N_1000,N_917,N_600);
nor U1001 (N_1001,N_10,N_589);
xor U1002 (N_1002,N_410,N_233);
nand U1003 (N_1003,N_773,N_134);
nand U1004 (N_1004,N_873,N_30);
nand U1005 (N_1005,N_473,N_998);
or U1006 (N_1006,N_123,N_674);
nand U1007 (N_1007,N_876,N_165);
nand U1008 (N_1008,N_859,N_567);
nand U1009 (N_1009,N_618,N_796);
nand U1010 (N_1010,N_972,N_70);
or U1011 (N_1011,N_389,N_551);
nand U1012 (N_1012,N_969,N_191);
nor U1013 (N_1013,N_394,N_696);
nor U1014 (N_1014,N_453,N_476);
or U1015 (N_1015,N_336,N_153);
nand U1016 (N_1016,N_43,N_523);
nand U1017 (N_1017,N_264,N_620);
and U1018 (N_1018,N_502,N_26);
or U1019 (N_1019,N_146,N_435);
or U1020 (N_1020,N_727,N_964);
and U1021 (N_1021,N_402,N_803);
and U1022 (N_1022,N_48,N_184);
and U1023 (N_1023,N_662,N_130);
nand U1024 (N_1024,N_2,N_749);
and U1025 (N_1025,N_774,N_456);
nand U1026 (N_1026,N_910,N_614);
and U1027 (N_1027,N_538,N_87);
nor U1028 (N_1028,N_658,N_409);
nor U1029 (N_1029,N_99,N_732);
and U1030 (N_1030,N_4,N_919);
or U1031 (N_1031,N_746,N_572);
nor U1032 (N_1032,N_137,N_817);
nand U1033 (N_1033,N_437,N_826);
nor U1034 (N_1034,N_903,N_425);
or U1035 (N_1035,N_627,N_622);
nor U1036 (N_1036,N_35,N_552);
or U1037 (N_1037,N_503,N_578);
and U1038 (N_1038,N_343,N_815);
and U1039 (N_1039,N_378,N_767);
and U1040 (N_1040,N_734,N_766);
or U1041 (N_1041,N_947,N_654);
or U1042 (N_1042,N_299,N_488);
nand U1043 (N_1043,N_178,N_479);
or U1044 (N_1044,N_305,N_326);
or U1045 (N_1045,N_376,N_112);
or U1046 (N_1046,N_239,N_471);
or U1047 (N_1047,N_21,N_827);
and U1048 (N_1048,N_940,N_457);
or U1049 (N_1049,N_704,N_714);
nor U1050 (N_1050,N_445,N_64);
or U1051 (N_1051,N_121,N_539);
nand U1052 (N_1052,N_267,N_213);
or U1053 (N_1053,N_900,N_562);
nor U1054 (N_1054,N_649,N_939);
nand U1055 (N_1055,N_477,N_609);
or U1056 (N_1056,N_12,N_836);
and U1057 (N_1057,N_591,N_814);
nand U1058 (N_1058,N_624,N_922);
nand U1059 (N_1059,N_985,N_518);
or U1060 (N_1060,N_55,N_177);
or U1061 (N_1061,N_253,N_584);
or U1062 (N_1062,N_133,N_39);
nor U1063 (N_1063,N_269,N_978);
nor U1064 (N_1064,N_856,N_656);
nand U1065 (N_1065,N_263,N_80);
or U1066 (N_1066,N_429,N_695);
or U1067 (N_1067,N_303,N_712);
nand U1068 (N_1068,N_149,N_861);
and U1069 (N_1069,N_744,N_186);
nor U1070 (N_1070,N_327,N_347);
or U1071 (N_1071,N_494,N_970);
nand U1072 (N_1072,N_432,N_158);
or U1073 (N_1073,N_729,N_293);
nor U1074 (N_1074,N_990,N_517);
nand U1075 (N_1075,N_629,N_379);
or U1076 (N_1076,N_190,N_797);
and U1077 (N_1077,N_886,N_474);
xnor U1078 (N_1078,N_434,N_923);
nor U1079 (N_1079,N_314,N_798);
or U1080 (N_1080,N_265,N_759);
nor U1081 (N_1081,N_603,N_845);
or U1082 (N_1082,N_761,N_397);
and U1083 (N_1083,N_325,N_54);
nor U1084 (N_1084,N_849,N_188);
nor U1085 (N_1085,N_199,N_207);
nor U1086 (N_1086,N_300,N_772);
nor U1087 (N_1087,N_937,N_515);
and U1088 (N_1088,N_282,N_8);
nor U1089 (N_1089,N_920,N_735);
nor U1090 (N_1090,N_443,N_291);
or U1091 (N_1091,N_672,N_728);
and U1092 (N_1092,N_667,N_723);
nand U1093 (N_1093,N_167,N_800);
or U1094 (N_1094,N_602,N_463);
nor U1095 (N_1095,N_769,N_963);
nand U1096 (N_1096,N_871,N_257);
or U1097 (N_1097,N_60,N_104);
and U1098 (N_1098,N_850,N_140);
and U1099 (N_1099,N_892,N_740);
nor U1100 (N_1100,N_752,N_840);
or U1101 (N_1101,N_991,N_482);
nand U1102 (N_1102,N_101,N_268);
nor U1103 (N_1103,N_328,N_596);
and U1104 (N_1104,N_863,N_706);
and U1105 (N_1105,N_504,N_292);
nand U1106 (N_1106,N_375,N_933);
nor U1107 (N_1107,N_89,N_32);
or U1108 (N_1108,N_847,N_512);
and U1109 (N_1109,N_610,N_748);
or U1110 (N_1110,N_593,N_957);
and U1111 (N_1111,N_372,N_877);
nor U1112 (N_1112,N_483,N_472);
or U1113 (N_1113,N_717,N_118);
nor U1114 (N_1114,N_392,N_776);
nor U1115 (N_1115,N_787,N_351);
or U1116 (N_1116,N_738,N_408);
or U1117 (N_1117,N_152,N_481);
and U1118 (N_1118,N_485,N_924);
nand U1119 (N_1119,N_681,N_763);
xnor U1120 (N_1120,N_148,N_189);
nand U1121 (N_1121,N_266,N_527);
and U1122 (N_1122,N_66,N_427);
or U1123 (N_1123,N_352,N_242);
nand U1124 (N_1124,N_768,N_451);
or U1125 (N_1125,N_6,N_870);
nand U1126 (N_1126,N_261,N_820);
and U1127 (N_1127,N_374,N_666);
and U1128 (N_1128,N_301,N_321);
or U1129 (N_1129,N_204,N_154);
nand U1130 (N_1130,N_659,N_743);
nand U1131 (N_1131,N_771,N_895);
nor U1132 (N_1132,N_869,N_365);
nor U1133 (N_1133,N_381,N_982);
and U1134 (N_1134,N_499,N_124);
nor U1135 (N_1135,N_284,N_225);
or U1136 (N_1136,N_319,N_819);
nand U1137 (N_1137,N_219,N_887);
nor U1138 (N_1138,N_366,N_673);
nand U1139 (N_1139,N_309,N_271);
nand U1140 (N_1140,N_926,N_984);
nor U1141 (N_1141,N_491,N_329);
or U1142 (N_1142,N_245,N_755);
xor U1143 (N_1143,N_812,N_785);
and U1144 (N_1144,N_931,N_450);
nor U1145 (N_1145,N_916,N_95);
nand U1146 (N_1146,N_573,N_138);
nand U1147 (N_1147,N_805,N_576);
nor U1148 (N_1148,N_139,N_949);
nor U1149 (N_1149,N_332,N_956);
nand U1150 (N_1150,N_193,N_821);
or U1151 (N_1151,N_0,N_493);
nand U1152 (N_1152,N_553,N_313);
or U1153 (N_1153,N_519,N_383);
or U1154 (N_1154,N_357,N_685);
nor U1155 (N_1155,N_75,N_387);
nand U1156 (N_1156,N_49,N_536);
nand U1157 (N_1157,N_902,N_73);
or U1158 (N_1158,N_175,N_825);
or U1159 (N_1159,N_941,N_58);
nor U1160 (N_1160,N_390,N_532);
nand U1161 (N_1161,N_363,N_323);
or U1162 (N_1162,N_641,N_270);
nor U1163 (N_1163,N_929,N_346);
nor U1164 (N_1164,N_534,N_533);
and U1165 (N_1165,N_240,N_643);
and U1166 (N_1166,N_371,N_646);
or U1167 (N_1167,N_569,N_839);
or U1168 (N_1168,N_109,N_571);
and U1169 (N_1169,N_289,N_71);
nor U1170 (N_1170,N_822,N_141);
or U1171 (N_1171,N_625,N_469);
or U1172 (N_1172,N_757,N_230);
nand U1173 (N_1173,N_832,N_331);
nand U1174 (N_1174,N_858,N_637);
and U1175 (N_1175,N_653,N_513);
nand U1176 (N_1176,N_547,N_22);
nand U1177 (N_1177,N_784,N_806);
nor U1178 (N_1178,N_559,N_315);
nor U1179 (N_1179,N_180,N_691);
or U1180 (N_1180,N_975,N_566);
nor U1181 (N_1181,N_281,N_733);
nor U1182 (N_1182,N_831,N_216);
or U1183 (N_1183,N_151,N_893);
nand U1184 (N_1184,N_492,N_74);
nor U1185 (N_1185,N_683,N_795);
nand U1186 (N_1186,N_988,N_63);
nand U1187 (N_1187,N_824,N_241);
and U1188 (N_1188,N_594,N_908);
and U1189 (N_1189,N_879,N_535);
nand U1190 (N_1190,N_354,N_113);
nand U1191 (N_1191,N_516,N_349);
nor U1192 (N_1192,N_385,N_295);
nor U1193 (N_1193,N_514,N_550);
or U1194 (N_1194,N_9,N_753);
or U1195 (N_1195,N_844,N_549);
nor U1196 (N_1196,N_592,N_872);
or U1197 (N_1197,N_632,N_880);
or U1198 (N_1198,N_220,N_361);
nor U1199 (N_1199,N_196,N_913);
nand U1200 (N_1200,N_868,N_855);
nor U1201 (N_1201,N_423,N_545);
or U1202 (N_1202,N_611,N_132);
or U1203 (N_1203,N_278,N_599);
and U1204 (N_1204,N_823,N_799);
nor U1205 (N_1205,N_181,N_454);
and U1206 (N_1206,N_792,N_470);
or U1207 (N_1207,N_501,N_671);
and U1208 (N_1208,N_585,N_317);
and U1209 (N_1209,N_901,N_833);
or U1210 (N_1210,N_126,N_82);
or U1211 (N_1211,N_93,N_809);
nand U1212 (N_1212,N_762,N_966);
nor U1213 (N_1213,N_234,N_403);
or U1214 (N_1214,N_320,N_287);
and U1215 (N_1215,N_83,N_915);
or U1216 (N_1216,N_954,N_159);
nand U1217 (N_1217,N_475,N_422);
nand U1218 (N_1218,N_102,N_262);
nor U1219 (N_1219,N_709,N_987);
nand U1220 (N_1220,N_508,N_680);
and U1221 (N_1221,N_120,N_775);
nor U1222 (N_1222,N_444,N_358);
or U1223 (N_1223,N_693,N_322);
and U1224 (N_1224,N_907,N_384);
or U1225 (N_1225,N_528,N_318);
nor U1226 (N_1226,N_794,N_185);
and U1227 (N_1227,N_143,N_85);
nand U1228 (N_1228,N_202,N_205);
nand U1229 (N_1229,N_952,N_854);
or U1230 (N_1230,N_441,N_192);
nor U1231 (N_1231,N_837,N_50);
or U1232 (N_1232,N_786,N_843);
nor U1233 (N_1233,N_793,N_77);
nand U1234 (N_1234,N_163,N_853);
and U1235 (N_1235,N_285,N_726);
nor U1236 (N_1236,N_811,N_91);
or U1237 (N_1237,N_210,N_235);
nand U1238 (N_1238,N_283,N_986);
nand U1239 (N_1239,N_114,N_248);
nand U1240 (N_1240,N_286,N_490);
and U1241 (N_1241,N_430,N_439);
nand U1242 (N_1242,N_636,N_276);
or U1243 (N_1243,N_623,N_955);
or U1244 (N_1244,N_778,N_851);
or U1245 (N_1245,N_497,N_829);
nand U1246 (N_1246,N_943,N_977);
and U1247 (N_1247,N_14,N_94);
nor U1248 (N_1248,N_580,N_7);
or U1249 (N_1249,N_912,N_976);
and U1250 (N_1250,N_710,N_353);
or U1251 (N_1251,N_781,N_968);
and U1252 (N_1252,N_678,N_330);
and U1253 (N_1253,N_348,N_247);
nor U1254 (N_1254,N_17,N_46);
nor U1255 (N_1255,N_813,N_399);
or U1256 (N_1256,N_628,N_27);
and U1257 (N_1257,N_407,N_335);
nor U1258 (N_1258,N_260,N_586);
or U1259 (N_1259,N_311,N_162);
and U1260 (N_1260,N_57,N_224);
or U1261 (N_1261,N_100,N_345);
or U1262 (N_1262,N_911,N_852);
nor U1263 (N_1263,N_455,N_415);
nor U1264 (N_1264,N_307,N_932);
nor U1265 (N_1265,N_801,N_537);
nand U1266 (N_1266,N_38,N_983);
nand U1267 (N_1267,N_108,N_69);
and U1268 (N_1268,N_925,N_522);
or U1269 (N_1269,N_369,N_431);
nor U1270 (N_1270,N_777,N_828);
or U1271 (N_1271,N_496,N_388);
nand U1272 (N_1272,N_692,N_981);
nand U1273 (N_1273,N_789,N_677);
or U1274 (N_1274,N_486,N_209);
nand U1275 (N_1275,N_464,N_742);
nand U1276 (N_1276,N_360,N_187);
and U1277 (N_1277,N_72,N_557);
nor U1278 (N_1278,N_59,N_197);
nand U1279 (N_1279,N_414,N_560);
or U1280 (N_1280,N_484,N_928);
or U1281 (N_1281,N_842,N_127);
nand U1282 (N_1282,N_297,N_117);
nand U1283 (N_1283,N_90,N_416);
and U1284 (N_1284,N_802,N_555);
and U1285 (N_1285,N_294,N_936);
nor U1286 (N_1286,N_697,N_604);
nand U1287 (N_1287,N_244,N_626);
nand U1288 (N_1288,N_461,N_65);
nand U1289 (N_1289,N_942,N_899);
nor U1290 (N_1290,N_231,N_807);
or U1291 (N_1291,N_129,N_705);
and U1292 (N_1292,N_631,N_834);
or U1293 (N_1293,N_782,N_223);
nand U1294 (N_1294,N_511,N_934);
and U1295 (N_1295,N_174,N_206);
or U1296 (N_1296,N_722,N_810);
nand U1297 (N_1297,N_750,N_841);
and U1298 (N_1298,N_703,N_642);
nor U1299 (N_1299,N_41,N_583);
nor U1300 (N_1300,N_218,N_296);
and U1301 (N_1301,N_340,N_700);
nor U1302 (N_1302,N_846,N_316);
nand U1303 (N_1303,N_563,N_249);
or U1304 (N_1304,N_144,N_42);
nand U1305 (N_1305,N_36,N_421);
and U1306 (N_1306,N_145,N_838);
or U1307 (N_1307,N_707,N_310);
or U1308 (N_1308,N_918,N_607);
nor U1309 (N_1309,N_676,N_721);
and U1310 (N_1310,N_657,N_51);
or U1311 (N_1311,N_951,N_595);
and U1312 (N_1312,N_183,N_756);
and U1313 (N_1313,N_448,N_255);
and U1314 (N_1314,N_478,N_462);
nor U1315 (N_1315,N_170,N_290);
nand U1316 (N_1316,N_546,N_554);
nor U1317 (N_1317,N_783,N_164);
xor U1318 (N_1318,N_312,N_417);
nor U1319 (N_1319,N_24,N_974);
or U1320 (N_1320,N_994,N_867);
or U1321 (N_1321,N_11,N_650);
nand U1322 (N_1322,N_147,N_119);
nor U1323 (N_1323,N_195,N_156);
or U1324 (N_1324,N_716,N_400);
nand U1325 (N_1325,N_79,N_525);
or U1326 (N_1326,N_770,N_914);
or U1327 (N_1327,N_342,N_405);
nand U1328 (N_1328,N_338,N_258);
nand U1329 (N_1329,N_237,N_23);
or U1330 (N_1330,N_608,N_229);
and U1331 (N_1331,N_904,N_274);
nor U1332 (N_1332,N_999,N_699);
and U1333 (N_1333,N_489,N_142);
nand U1334 (N_1334,N_897,N_221);
nand U1335 (N_1335,N_989,N_169);
and U1336 (N_1336,N_160,N_226);
nor U1337 (N_1337,N_406,N_298);
and U1338 (N_1338,N_808,N_745);
or U1339 (N_1339,N_857,N_419);
or U1340 (N_1340,N_304,N_500);
nand U1341 (N_1341,N_339,N_334);
nand U1342 (N_1342,N_447,N_708);
and U1343 (N_1343,N_938,N_370);
or U1344 (N_1344,N_401,N_15);
and U1345 (N_1345,N_395,N_804);
and U1346 (N_1346,N_606,N_651);
nand U1347 (N_1347,N_509,N_272);
and U1348 (N_1348,N_992,N_155);
nand U1349 (N_1349,N_377,N_860);
or U1350 (N_1350,N_212,N_965);
and U1351 (N_1351,N_980,N_115);
and U1352 (N_1352,N_18,N_598);
nand U1353 (N_1353,N_719,N_182);
nand U1354 (N_1354,N_779,N_788);
and U1355 (N_1355,N_574,N_575);
nor U1356 (N_1356,N_944,N_647);
or U1357 (N_1357,N_971,N_862);
and U1358 (N_1358,N_997,N_529);
nand U1359 (N_1359,N_711,N_81);
or U1360 (N_1360,N_105,N_203);
nand U1361 (N_1361,N_921,N_612);
and U1362 (N_1362,N_724,N_173);
nand U1363 (N_1363,N_47,N_53);
and U1364 (N_1364,N_888,N_78);
and U1365 (N_1365,N_33,N_254);
or U1366 (N_1366,N_96,N_541);
or U1367 (N_1367,N_958,N_68);
or U1368 (N_1368,N_945,N_638);
and U1369 (N_1369,N_76,N_864);
and U1370 (N_1370,N_337,N_288);
and U1371 (N_1371,N_498,N_946);
or U1372 (N_1372,N_568,N_67);
and U1373 (N_1373,N_790,N_86);
or U1374 (N_1374,N_758,N_590);
or U1375 (N_1375,N_621,N_106);
nand U1376 (N_1376,N_236,N_521);
and U1377 (N_1377,N_398,N_393);
nand U1378 (N_1378,N_882,N_665);
nor U1379 (N_1379,N_13,N_682);
xor U1380 (N_1380,N_1,N_935);
nor U1381 (N_1381,N_350,N_380);
and U1382 (N_1382,N_420,N_279);
or U1383 (N_1383,N_848,N_601);
or U1384 (N_1384,N_480,N_211);
or U1385 (N_1385,N_356,N_56);
and U1386 (N_1386,N_150,N_29);
nor U1387 (N_1387,N_465,N_780);
nor U1388 (N_1388,N_613,N_259);
nand U1389 (N_1389,N_731,N_20);
nand U1390 (N_1390,N_198,N_215);
nand U1391 (N_1391,N_157,N_252);
nor U1392 (N_1392,N_458,N_232);
or U1393 (N_1393,N_128,N_214);
nor U1394 (N_1394,N_701,N_959);
and U1395 (N_1395,N_644,N_713);
or U1396 (N_1396,N_664,N_40);
or U1397 (N_1397,N_715,N_412);
and U1398 (N_1398,N_564,N_433);
and U1399 (N_1399,N_874,N_449);
nor U1400 (N_1400,N_718,N_565);
nor U1401 (N_1401,N_582,N_865);
or U1402 (N_1402,N_979,N_630);
nand U1403 (N_1403,N_62,N_561);
nand U1404 (N_1404,N_679,N_176);
and U1405 (N_1405,N_588,N_617);
nand U1406 (N_1406,N_885,N_760);
or U1407 (N_1407,N_243,N_250);
xor U1408 (N_1408,N_635,N_16);
or U1409 (N_1409,N_200,N_505);
nor U1410 (N_1410,N_111,N_634);
or U1411 (N_1411,N_684,N_668);
and U1412 (N_1412,N_359,N_131);
and U1413 (N_1413,N_663,N_487);
nand U1414 (N_1414,N_655,N_122);
nor U1415 (N_1415,N_364,N_616);
nor U1416 (N_1416,N_467,N_960);
nand U1417 (N_1417,N_386,N_436);
nor U1418 (N_1418,N_166,N_577);
nand U1419 (N_1419,N_739,N_698);
or U1420 (N_1420,N_905,N_396);
or U1421 (N_1421,N_306,N_308);
nor U1422 (N_1422,N_201,N_570);
and U1423 (N_1423,N_694,N_894);
nand U1424 (N_1424,N_344,N_19);
nor U1425 (N_1425,N_136,N_648);
nand U1426 (N_1426,N_438,N_277);
and U1427 (N_1427,N_222,N_530);
or U1428 (N_1428,N_581,N_5);
or U1429 (N_1429,N_424,N_558);
and U1430 (N_1430,N_878,N_967);
nor U1431 (N_1431,N_442,N_506);
or U1432 (N_1432,N_791,N_228);
and U1433 (N_1433,N_28,N_896);
and U1434 (N_1434,N_661,N_459);
nand U1435 (N_1435,N_891,N_548);
nor U1436 (N_1436,N_103,N_690);
nand U1437 (N_1437,N_741,N_747);
or U1438 (N_1438,N_172,N_702);
or U1439 (N_1439,N_725,N_930);
or U1440 (N_1440,N_256,N_996);
nor U1441 (N_1441,N_520,N_619);
or U1442 (N_1442,N_61,N_835);
or U1443 (N_1443,N_890,N_238);
and U1444 (N_1444,N_413,N_751);
nand U1445 (N_1445,N_906,N_953);
nand U1446 (N_1446,N_973,N_507);
and U1447 (N_1447,N_411,N_107);
nand U1448 (N_1448,N_92,N_689);
nand U1449 (N_1449,N_962,N_217);
or U1450 (N_1450,N_866,N_440);
nand U1451 (N_1451,N_543,N_168);
or U1452 (N_1452,N_452,N_542);
or U1453 (N_1453,N_227,N_526);
or U1454 (N_1454,N_927,N_675);
nor U1455 (N_1455,N_460,N_275);
and U1456 (N_1456,N_639,N_355);
and U1457 (N_1457,N_368,N_730);
or U1458 (N_1458,N_110,N_418);
nand U1459 (N_1459,N_280,N_88);
nand U1460 (N_1460,N_251,N_273);
or U1461 (N_1461,N_125,N_754);
or U1462 (N_1462,N_883,N_830);
nand U1463 (N_1463,N_540,N_446);
nand U1464 (N_1464,N_686,N_597);
and U1465 (N_1465,N_898,N_116);
nor U1466 (N_1466,N_645,N_44);
and U1467 (N_1467,N_171,N_333);
nor U1468 (N_1468,N_993,N_889);
or U1469 (N_1469,N_362,N_652);
and U1470 (N_1470,N_884,N_84);
nand U1471 (N_1471,N_52,N_466);
or U1472 (N_1472,N_816,N_194);
or U1473 (N_1473,N_25,N_909);
and U1474 (N_1474,N_179,N_587);
nor U1475 (N_1475,N_382,N_341);
nor U1476 (N_1476,N_161,N_531);
or U1477 (N_1477,N_524,N_556);
nor U1478 (N_1478,N_948,N_135);
and U1479 (N_1479,N_391,N_605);
and U1480 (N_1480,N_881,N_510);
nand U1481 (N_1481,N_765,N_875);
or U1482 (N_1482,N_31,N_373);
nand U1483 (N_1483,N_302,N_45);
nor U1484 (N_1484,N_961,N_579);
nand U1485 (N_1485,N_818,N_428);
or U1486 (N_1486,N_3,N_995);
nand U1487 (N_1487,N_495,N_736);
and U1488 (N_1488,N_426,N_98);
or U1489 (N_1489,N_468,N_764);
and U1490 (N_1490,N_737,N_37);
and U1491 (N_1491,N_688,N_615);
and U1492 (N_1492,N_950,N_367);
nand U1493 (N_1493,N_640,N_97);
nor U1494 (N_1494,N_687,N_669);
and U1495 (N_1495,N_246,N_670);
and U1496 (N_1496,N_208,N_544);
nand U1497 (N_1497,N_404,N_34);
nor U1498 (N_1498,N_633,N_720);
and U1499 (N_1499,N_324,N_660);
and U1500 (N_1500,N_207,N_655);
nor U1501 (N_1501,N_640,N_642);
nor U1502 (N_1502,N_113,N_24);
nand U1503 (N_1503,N_351,N_950);
nor U1504 (N_1504,N_740,N_103);
nand U1505 (N_1505,N_755,N_247);
and U1506 (N_1506,N_740,N_406);
and U1507 (N_1507,N_834,N_905);
or U1508 (N_1508,N_597,N_48);
or U1509 (N_1509,N_690,N_477);
and U1510 (N_1510,N_265,N_99);
or U1511 (N_1511,N_614,N_700);
nor U1512 (N_1512,N_291,N_717);
or U1513 (N_1513,N_566,N_811);
nor U1514 (N_1514,N_216,N_987);
nor U1515 (N_1515,N_980,N_1);
nor U1516 (N_1516,N_786,N_339);
and U1517 (N_1517,N_927,N_163);
nor U1518 (N_1518,N_760,N_554);
nand U1519 (N_1519,N_965,N_330);
nand U1520 (N_1520,N_920,N_117);
nand U1521 (N_1521,N_560,N_282);
or U1522 (N_1522,N_82,N_264);
nand U1523 (N_1523,N_336,N_43);
and U1524 (N_1524,N_525,N_487);
nor U1525 (N_1525,N_271,N_842);
and U1526 (N_1526,N_329,N_556);
and U1527 (N_1527,N_398,N_327);
nor U1528 (N_1528,N_293,N_665);
nor U1529 (N_1529,N_176,N_403);
nor U1530 (N_1530,N_965,N_853);
nand U1531 (N_1531,N_595,N_164);
nand U1532 (N_1532,N_125,N_421);
nor U1533 (N_1533,N_216,N_756);
and U1534 (N_1534,N_390,N_691);
nand U1535 (N_1535,N_110,N_315);
nor U1536 (N_1536,N_404,N_118);
nand U1537 (N_1537,N_578,N_613);
nor U1538 (N_1538,N_963,N_33);
and U1539 (N_1539,N_860,N_600);
nor U1540 (N_1540,N_789,N_211);
nor U1541 (N_1541,N_841,N_633);
nor U1542 (N_1542,N_653,N_387);
nand U1543 (N_1543,N_809,N_367);
and U1544 (N_1544,N_604,N_107);
or U1545 (N_1545,N_971,N_368);
nor U1546 (N_1546,N_984,N_398);
or U1547 (N_1547,N_398,N_601);
and U1548 (N_1548,N_323,N_264);
nor U1549 (N_1549,N_913,N_695);
or U1550 (N_1550,N_435,N_784);
or U1551 (N_1551,N_927,N_714);
or U1552 (N_1552,N_562,N_138);
or U1553 (N_1553,N_716,N_126);
nand U1554 (N_1554,N_538,N_895);
nand U1555 (N_1555,N_839,N_71);
nand U1556 (N_1556,N_713,N_859);
or U1557 (N_1557,N_779,N_499);
or U1558 (N_1558,N_986,N_166);
nor U1559 (N_1559,N_505,N_51);
or U1560 (N_1560,N_891,N_132);
nand U1561 (N_1561,N_689,N_250);
and U1562 (N_1562,N_6,N_408);
and U1563 (N_1563,N_600,N_425);
and U1564 (N_1564,N_732,N_895);
or U1565 (N_1565,N_265,N_302);
and U1566 (N_1566,N_356,N_475);
and U1567 (N_1567,N_169,N_754);
and U1568 (N_1568,N_359,N_881);
nor U1569 (N_1569,N_958,N_904);
nor U1570 (N_1570,N_151,N_105);
nand U1571 (N_1571,N_156,N_708);
and U1572 (N_1572,N_473,N_246);
and U1573 (N_1573,N_553,N_879);
or U1574 (N_1574,N_179,N_377);
xnor U1575 (N_1575,N_327,N_917);
and U1576 (N_1576,N_199,N_465);
nand U1577 (N_1577,N_968,N_112);
and U1578 (N_1578,N_519,N_872);
nand U1579 (N_1579,N_805,N_539);
nand U1580 (N_1580,N_464,N_903);
or U1581 (N_1581,N_822,N_118);
or U1582 (N_1582,N_29,N_153);
or U1583 (N_1583,N_519,N_617);
nand U1584 (N_1584,N_676,N_868);
nor U1585 (N_1585,N_201,N_494);
nor U1586 (N_1586,N_332,N_108);
nor U1587 (N_1587,N_600,N_782);
or U1588 (N_1588,N_707,N_987);
nor U1589 (N_1589,N_737,N_196);
and U1590 (N_1590,N_469,N_609);
or U1591 (N_1591,N_340,N_894);
and U1592 (N_1592,N_534,N_748);
or U1593 (N_1593,N_420,N_504);
and U1594 (N_1594,N_849,N_334);
nor U1595 (N_1595,N_799,N_230);
nor U1596 (N_1596,N_749,N_368);
or U1597 (N_1597,N_311,N_313);
nand U1598 (N_1598,N_541,N_458);
nor U1599 (N_1599,N_754,N_684);
or U1600 (N_1600,N_90,N_115);
nor U1601 (N_1601,N_93,N_378);
nor U1602 (N_1602,N_994,N_700);
and U1603 (N_1603,N_823,N_659);
and U1604 (N_1604,N_140,N_725);
nor U1605 (N_1605,N_497,N_348);
and U1606 (N_1606,N_31,N_13);
and U1607 (N_1607,N_821,N_81);
nor U1608 (N_1608,N_55,N_817);
and U1609 (N_1609,N_318,N_828);
nor U1610 (N_1610,N_930,N_632);
nand U1611 (N_1611,N_838,N_550);
nor U1612 (N_1612,N_147,N_245);
and U1613 (N_1613,N_891,N_593);
or U1614 (N_1614,N_527,N_864);
and U1615 (N_1615,N_134,N_579);
nand U1616 (N_1616,N_778,N_889);
nand U1617 (N_1617,N_952,N_593);
and U1618 (N_1618,N_447,N_389);
or U1619 (N_1619,N_803,N_905);
nor U1620 (N_1620,N_939,N_886);
nand U1621 (N_1621,N_948,N_921);
or U1622 (N_1622,N_145,N_505);
and U1623 (N_1623,N_258,N_197);
nor U1624 (N_1624,N_436,N_687);
and U1625 (N_1625,N_196,N_275);
and U1626 (N_1626,N_105,N_262);
nor U1627 (N_1627,N_691,N_342);
nand U1628 (N_1628,N_317,N_115);
or U1629 (N_1629,N_978,N_377);
or U1630 (N_1630,N_424,N_954);
nand U1631 (N_1631,N_706,N_264);
nor U1632 (N_1632,N_968,N_208);
xnor U1633 (N_1633,N_537,N_408);
nand U1634 (N_1634,N_947,N_569);
or U1635 (N_1635,N_452,N_200);
nor U1636 (N_1636,N_465,N_934);
nand U1637 (N_1637,N_307,N_1);
or U1638 (N_1638,N_313,N_388);
nand U1639 (N_1639,N_287,N_901);
nand U1640 (N_1640,N_97,N_803);
nor U1641 (N_1641,N_417,N_574);
xnor U1642 (N_1642,N_911,N_904);
or U1643 (N_1643,N_905,N_872);
nand U1644 (N_1644,N_113,N_513);
and U1645 (N_1645,N_783,N_538);
or U1646 (N_1646,N_632,N_60);
nand U1647 (N_1647,N_25,N_552);
nand U1648 (N_1648,N_75,N_213);
or U1649 (N_1649,N_779,N_647);
or U1650 (N_1650,N_947,N_911);
and U1651 (N_1651,N_326,N_795);
xnor U1652 (N_1652,N_730,N_26);
nor U1653 (N_1653,N_857,N_257);
or U1654 (N_1654,N_177,N_627);
or U1655 (N_1655,N_423,N_867);
and U1656 (N_1656,N_845,N_891);
and U1657 (N_1657,N_429,N_257);
or U1658 (N_1658,N_127,N_255);
or U1659 (N_1659,N_858,N_46);
or U1660 (N_1660,N_8,N_13);
and U1661 (N_1661,N_709,N_773);
and U1662 (N_1662,N_245,N_578);
or U1663 (N_1663,N_995,N_752);
and U1664 (N_1664,N_985,N_526);
nand U1665 (N_1665,N_443,N_79);
nor U1666 (N_1666,N_798,N_738);
nor U1667 (N_1667,N_221,N_94);
and U1668 (N_1668,N_961,N_269);
nor U1669 (N_1669,N_935,N_229);
and U1670 (N_1670,N_168,N_575);
nor U1671 (N_1671,N_458,N_388);
nand U1672 (N_1672,N_982,N_515);
or U1673 (N_1673,N_724,N_377);
nor U1674 (N_1674,N_137,N_18);
nand U1675 (N_1675,N_931,N_12);
nor U1676 (N_1676,N_878,N_263);
and U1677 (N_1677,N_995,N_629);
nand U1678 (N_1678,N_52,N_606);
and U1679 (N_1679,N_271,N_748);
and U1680 (N_1680,N_571,N_40);
or U1681 (N_1681,N_828,N_148);
nand U1682 (N_1682,N_573,N_830);
nor U1683 (N_1683,N_833,N_529);
nor U1684 (N_1684,N_574,N_278);
or U1685 (N_1685,N_45,N_392);
nor U1686 (N_1686,N_485,N_522);
and U1687 (N_1687,N_198,N_873);
nand U1688 (N_1688,N_851,N_139);
nand U1689 (N_1689,N_612,N_939);
or U1690 (N_1690,N_449,N_379);
nand U1691 (N_1691,N_642,N_306);
or U1692 (N_1692,N_322,N_332);
or U1693 (N_1693,N_429,N_673);
nor U1694 (N_1694,N_474,N_171);
xor U1695 (N_1695,N_354,N_279);
and U1696 (N_1696,N_71,N_978);
and U1697 (N_1697,N_891,N_259);
nor U1698 (N_1698,N_935,N_554);
nor U1699 (N_1699,N_302,N_183);
nand U1700 (N_1700,N_804,N_129);
nor U1701 (N_1701,N_495,N_297);
nor U1702 (N_1702,N_579,N_567);
nand U1703 (N_1703,N_258,N_161);
nand U1704 (N_1704,N_126,N_318);
nor U1705 (N_1705,N_308,N_687);
nor U1706 (N_1706,N_472,N_727);
and U1707 (N_1707,N_719,N_240);
or U1708 (N_1708,N_990,N_469);
and U1709 (N_1709,N_843,N_60);
and U1710 (N_1710,N_915,N_834);
nand U1711 (N_1711,N_987,N_977);
nor U1712 (N_1712,N_945,N_391);
nand U1713 (N_1713,N_916,N_258);
nand U1714 (N_1714,N_968,N_816);
nand U1715 (N_1715,N_241,N_818);
nor U1716 (N_1716,N_790,N_449);
nand U1717 (N_1717,N_40,N_393);
nand U1718 (N_1718,N_574,N_640);
nand U1719 (N_1719,N_911,N_562);
nand U1720 (N_1720,N_639,N_108);
nand U1721 (N_1721,N_283,N_482);
or U1722 (N_1722,N_946,N_613);
nor U1723 (N_1723,N_899,N_757);
and U1724 (N_1724,N_959,N_260);
and U1725 (N_1725,N_51,N_683);
and U1726 (N_1726,N_273,N_182);
and U1727 (N_1727,N_884,N_983);
nor U1728 (N_1728,N_15,N_29);
xor U1729 (N_1729,N_255,N_923);
and U1730 (N_1730,N_595,N_177);
nor U1731 (N_1731,N_234,N_727);
or U1732 (N_1732,N_779,N_859);
or U1733 (N_1733,N_258,N_208);
nor U1734 (N_1734,N_447,N_557);
xor U1735 (N_1735,N_859,N_726);
or U1736 (N_1736,N_596,N_24);
and U1737 (N_1737,N_741,N_817);
nand U1738 (N_1738,N_735,N_589);
nand U1739 (N_1739,N_617,N_381);
nor U1740 (N_1740,N_167,N_661);
nor U1741 (N_1741,N_602,N_793);
nand U1742 (N_1742,N_526,N_927);
nor U1743 (N_1743,N_554,N_534);
nor U1744 (N_1744,N_396,N_772);
and U1745 (N_1745,N_49,N_330);
nand U1746 (N_1746,N_37,N_710);
and U1747 (N_1747,N_895,N_263);
nor U1748 (N_1748,N_608,N_810);
or U1749 (N_1749,N_754,N_415);
nor U1750 (N_1750,N_837,N_441);
nor U1751 (N_1751,N_153,N_265);
nor U1752 (N_1752,N_505,N_866);
and U1753 (N_1753,N_138,N_731);
nand U1754 (N_1754,N_277,N_848);
and U1755 (N_1755,N_878,N_545);
nor U1756 (N_1756,N_96,N_942);
and U1757 (N_1757,N_369,N_866);
and U1758 (N_1758,N_156,N_716);
nor U1759 (N_1759,N_402,N_174);
or U1760 (N_1760,N_757,N_343);
xnor U1761 (N_1761,N_72,N_388);
nor U1762 (N_1762,N_608,N_642);
nor U1763 (N_1763,N_312,N_191);
or U1764 (N_1764,N_445,N_878);
nor U1765 (N_1765,N_978,N_255);
or U1766 (N_1766,N_86,N_130);
nor U1767 (N_1767,N_516,N_644);
and U1768 (N_1768,N_232,N_304);
nand U1769 (N_1769,N_223,N_482);
or U1770 (N_1770,N_236,N_259);
and U1771 (N_1771,N_276,N_442);
or U1772 (N_1772,N_874,N_155);
nor U1773 (N_1773,N_913,N_319);
nor U1774 (N_1774,N_101,N_15);
nand U1775 (N_1775,N_984,N_484);
and U1776 (N_1776,N_155,N_619);
nor U1777 (N_1777,N_186,N_45);
nor U1778 (N_1778,N_393,N_161);
or U1779 (N_1779,N_272,N_766);
and U1780 (N_1780,N_558,N_265);
nand U1781 (N_1781,N_835,N_446);
nand U1782 (N_1782,N_619,N_742);
nand U1783 (N_1783,N_174,N_903);
and U1784 (N_1784,N_52,N_993);
or U1785 (N_1785,N_635,N_29);
and U1786 (N_1786,N_73,N_360);
and U1787 (N_1787,N_965,N_302);
or U1788 (N_1788,N_781,N_675);
nand U1789 (N_1789,N_210,N_127);
and U1790 (N_1790,N_528,N_411);
nor U1791 (N_1791,N_217,N_450);
nor U1792 (N_1792,N_706,N_617);
or U1793 (N_1793,N_501,N_3);
or U1794 (N_1794,N_330,N_509);
and U1795 (N_1795,N_864,N_450);
or U1796 (N_1796,N_540,N_773);
nor U1797 (N_1797,N_482,N_933);
nor U1798 (N_1798,N_480,N_964);
or U1799 (N_1799,N_776,N_953);
and U1800 (N_1800,N_264,N_246);
nand U1801 (N_1801,N_923,N_164);
nor U1802 (N_1802,N_163,N_653);
and U1803 (N_1803,N_226,N_95);
nand U1804 (N_1804,N_416,N_961);
nand U1805 (N_1805,N_379,N_386);
xnor U1806 (N_1806,N_548,N_673);
and U1807 (N_1807,N_856,N_193);
nor U1808 (N_1808,N_694,N_506);
and U1809 (N_1809,N_777,N_260);
and U1810 (N_1810,N_441,N_591);
xnor U1811 (N_1811,N_331,N_115);
or U1812 (N_1812,N_785,N_130);
nand U1813 (N_1813,N_977,N_524);
and U1814 (N_1814,N_470,N_622);
or U1815 (N_1815,N_281,N_832);
and U1816 (N_1816,N_197,N_948);
or U1817 (N_1817,N_248,N_590);
and U1818 (N_1818,N_898,N_493);
nand U1819 (N_1819,N_159,N_104);
nand U1820 (N_1820,N_819,N_85);
nor U1821 (N_1821,N_140,N_971);
or U1822 (N_1822,N_599,N_402);
or U1823 (N_1823,N_727,N_952);
nor U1824 (N_1824,N_866,N_364);
nand U1825 (N_1825,N_987,N_922);
nor U1826 (N_1826,N_350,N_762);
and U1827 (N_1827,N_743,N_497);
nand U1828 (N_1828,N_129,N_513);
nand U1829 (N_1829,N_846,N_541);
and U1830 (N_1830,N_829,N_584);
nor U1831 (N_1831,N_630,N_943);
nor U1832 (N_1832,N_738,N_992);
nand U1833 (N_1833,N_890,N_989);
nand U1834 (N_1834,N_5,N_334);
nand U1835 (N_1835,N_839,N_89);
and U1836 (N_1836,N_736,N_269);
and U1837 (N_1837,N_452,N_205);
nor U1838 (N_1838,N_69,N_852);
and U1839 (N_1839,N_355,N_392);
or U1840 (N_1840,N_112,N_526);
and U1841 (N_1841,N_487,N_76);
and U1842 (N_1842,N_526,N_712);
or U1843 (N_1843,N_308,N_452);
nor U1844 (N_1844,N_532,N_717);
nand U1845 (N_1845,N_794,N_25);
and U1846 (N_1846,N_409,N_977);
nor U1847 (N_1847,N_236,N_280);
nor U1848 (N_1848,N_974,N_560);
nand U1849 (N_1849,N_353,N_0);
nand U1850 (N_1850,N_285,N_692);
nand U1851 (N_1851,N_850,N_827);
nand U1852 (N_1852,N_806,N_961);
nor U1853 (N_1853,N_178,N_201);
or U1854 (N_1854,N_997,N_293);
nor U1855 (N_1855,N_844,N_982);
nor U1856 (N_1856,N_157,N_839);
nor U1857 (N_1857,N_183,N_181);
nor U1858 (N_1858,N_873,N_515);
nor U1859 (N_1859,N_162,N_502);
and U1860 (N_1860,N_489,N_516);
nor U1861 (N_1861,N_50,N_333);
and U1862 (N_1862,N_639,N_143);
or U1863 (N_1863,N_405,N_248);
nor U1864 (N_1864,N_273,N_104);
and U1865 (N_1865,N_242,N_149);
nor U1866 (N_1866,N_46,N_289);
and U1867 (N_1867,N_688,N_854);
nor U1868 (N_1868,N_917,N_774);
nor U1869 (N_1869,N_223,N_13);
nor U1870 (N_1870,N_676,N_106);
and U1871 (N_1871,N_44,N_277);
nand U1872 (N_1872,N_411,N_479);
nor U1873 (N_1873,N_378,N_99);
or U1874 (N_1874,N_339,N_35);
or U1875 (N_1875,N_76,N_514);
or U1876 (N_1876,N_429,N_804);
nand U1877 (N_1877,N_99,N_375);
or U1878 (N_1878,N_111,N_685);
and U1879 (N_1879,N_754,N_435);
and U1880 (N_1880,N_279,N_582);
nor U1881 (N_1881,N_905,N_228);
nand U1882 (N_1882,N_665,N_356);
and U1883 (N_1883,N_182,N_522);
xnor U1884 (N_1884,N_653,N_44);
nand U1885 (N_1885,N_388,N_487);
nor U1886 (N_1886,N_64,N_757);
nor U1887 (N_1887,N_62,N_977);
nand U1888 (N_1888,N_993,N_931);
and U1889 (N_1889,N_844,N_326);
nor U1890 (N_1890,N_797,N_255);
or U1891 (N_1891,N_510,N_474);
nand U1892 (N_1892,N_155,N_225);
nand U1893 (N_1893,N_703,N_496);
and U1894 (N_1894,N_409,N_695);
and U1895 (N_1895,N_497,N_748);
or U1896 (N_1896,N_380,N_382);
or U1897 (N_1897,N_498,N_68);
nor U1898 (N_1898,N_372,N_970);
nand U1899 (N_1899,N_582,N_661);
nor U1900 (N_1900,N_897,N_830);
and U1901 (N_1901,N_721,N_513);
and U1902 (N_1902,N_817,N_159);
and U1903 (N_1903,N_738,N_531);
and U1904 (N_1904,N_358,N_140);
or U1905 (N_1905,N_398,N_373);
and U1906 (N_1906,N_635,N_986);
and U1907 (N_1907,N_108,N_805);
nand U1908 (N_1908,N_126,N_198);
nand U1909 (N_1909,N_275,N_727);
and U1910 (N_1910,N_468,N_869);
or U1911 (N_1911,N_457,N_298);
nor U1912 (N_1912,N_793,N_369);
nand U1913 (N_1913,N_261,N_230);
nand U1914 (N_1914,N_847,N_544);
xnor U1915 (N_1915,N_601,N_164);
or U1916 (N_1916,N_397,N_687);
and U1917 (N_1917,N_119,N_857);
nor U1918 (N_1918,N_564,N_351);
and U1919 (N_1919,N_222,N_560);
and U1920 (N_1920,N_32,N_853);
or U1921 (N_1921,N_536,N_726);
nand U1922 (N_1922,N_725,N_657);
or U1923 (N_1923,N_719,N_387);
or U1924 (N_1924,N_288,N_526);
nor U1925 (N_1925,N_691,N_733);
or U1926 (N_1926,N_620,N_631);
or U1927 (N_1927,N_17,N_869);
nand U1928 (N_1928,N_48,N_894);
or U1929 (N_1929,N_803,N_567);
or U1930 (N_1930,N_570,N_421);
or U1931 (N_1931,N_726,N_11);
nand U1932 (N_1932,N_423,N_735);
or U1933 (N_1933,N_452,N_847);
or U1934 (N_1934,N_471,N_304);
or U1935 (N_1935,N_433,N_917);
nor U1936 (N_1936,N_935,N_740);
nand U1937 (N_1937,N_348,N_584);
or U1938 (N_1938,N_401,N_684);
or U1939 (N_1939,N_735,N_778);
nand U1940 (N_1940,N_287,N_25);
and U1941 (N_1941,N_330,N_539);
and U1942 (N_1942,N_354,N_562);
nor U1943 (N_1943,N_959,N_673);
or U1944 (N_1944,N_316,N_746);
and U1945 (N_1945,N_613,N_736);
and U1946 (N_1946,N_799,N_380);
or U1947 (N_1947,N_413,N_468);
nor U1948 (N_1948,N_120,N_721);
nor U1949 (N_1949,N_896,N_524);
nor U1950 (N_1950,N_295,N_477);
nand U1951 (N_1951,N_290,N_226);
xor U1952 (N_1952,N_727,N_359);
or U1953 (N_1953,N_349,N_226);
xor U1954 (N_1954,N_199,N_191);
nor U1955 (N_1955,N_393,N_255);
or U1956 (N_1956,N_108,N_391);
nand U1957 (N_1957,N_427,N_488);
and U1958 (N_1958,N_869,N_324);
or U1959 (N_1959,N_944,N_751);
and U1960 (N_1960,N_544,N_942);
nor U1961 (N_1961,N_641,N_724);
or U1962 (N_1962,N_37,N_303);
nand U1963 (N_1963,N_685,N_760);
nor U1964 (N_1964,N_896,N_369);
nand U1965 (N_1965,N_68,N_43);
or U1966 (N_1966,N_776,N_660);
or U1967 (N_1967,N_809,N_628);
and U1968 (N_1968,N_541,N_297);
or U1969 (N_1969,N_510,N_24);
nand U1970 (N_1970,N_85,N_493);
nand U1971 (N_1971,N_326,N_834);
and U1972 (N_1972,N_969,N_398);
nand U1973 (N_1973,N_935,N_202);
or U1974 (N_1974,N_697,N_851);
nand U1975 (N_1975,N_589,N_849);
and U1976 (N_1976,N_121,N_377);
and U1977 (N_1977,N_679,N_414);
nand U1978 (N_1978,N_28,N_789);
or U1979 (N_1979,N_493,N_685);
nor U1980 (N_1980,N_835,N_613);
nor U1981 (N_1981,N_487,N_252);
nand U1982 (N_1982,N_764,N_266);
and U1983 (N_1983,N_162,N_830);
nand U1984 (N_1984,N_48,N_179);
and U1985 (N_1985,N_353,N_519);
and U1986 (N_1986,N_580,N_58);
nor U1987 (N_1987,N_315,N_570);
nor U1988 (N_1988,N_253,N_821);
or U1989 (N_1989,N_655,N_992);
or U1990 (N_1990,N_65,N_574);
and U1991 (N_1991,N_633,N_539);
or U1992 (N_1992,N_296,N_875);
nand U1993 (N_1993,N_300,N_978);
nand U1994 (N_1994,N_369,N_541);
nor U1995 (N_1995,N_799,N_374);
xnor U1996 (N_1996,N_947,N_641);
and U1997 (N_1997,N_95,N_815);
nand U1998 (N_1998,N_981,N_988);
nor U1999 (N_1999,N_873,N_736);
nor U2000 (N_2000,N_1544,N_1000);
and U2001 (N_2001,N_1189,N_1162);
and U2002 (N_2002,N_1071,N_1258);
or U2003 (N_2003,N_1400,N_1718);
nand U2004 (N_2004,N_1920,N_1937);
nor U2005 (N_2005,N_1959,N_1105);
and U2006 (N_2006,N_1781,N_1888);
nand U2007 (N_2007,N_1517,N_1042);
nand U2008 (N_2008,N_1304,N_1091);
or U2009 (N_2009,N_1305,N_1531);
nand U2010 (N_2010,N_1656,N_1238);
nor U2011 (N_2011,N_1955,N_1357);
and U2012 (N_2012,N_1886,N_1722);
nor U2013 (N_2013,N_1856,N_1424);
nor U2014 (N_2014,N_1208,N_1791);
or U2015 (N_2015,N_1599,N_1637);
nand U2016 (N_2016,N_1241,N_1027);
and U2017 (N_2017,N_1472,N_1354);
or U2018 (N_2018,N_1644,N_1288);
nand U2019 (N_2019,N_1402,N_1281);
nor U2020 (N_2020,N_1770,N_1717);
nor U2021 (N_2021,N_1534,N_1651);
nand U2022 (N_2022,N_1983,N_1335);
or U2023 (N_2023,N_1804,N_1261);
nor U2024 (N_2024,N_1487,N_1240);
nor U2025 (N_2025,N_1765,N_1589);
nor U2026 (N_2026,N_1764,N_1643);
nand U2027 (N_2027,N_1380,N_1848);
nor U2028 (N_2028,N_1752,N_1579);
or U2029 (N_2029,N_1786,N_1246);
nand U2030 (N_2030,N_1115,N_1857);
or U2031 (N_2031,N_1009,N_1635);
nand U2032 (N_2032,N_1085,N_1743);
nor U2033 (N_2033,N_1193,N_1634);
and U2034 (N_2034,N_1585,N_1066);
nor U2035 (N_2035,N_1177,N_1662);
and U2036 (N_2036,N_1128,N_1112);
or U2037 (N_2037,N_1974,N_1214);
and U2038 (N_2038,N_1481,N_1120);
nor U2039 (N_2039,N_1389,N_1245);
or U2040 (N_2040,N_1022,N_1188);
nor U2041 (N_2041,N_1501,N_1237);
or U2042 (N_2042,N_1324,N_1202);
nand U2043 (N_2043,N_1165,N_1911);
nor U2044 (N_2044,N_1934,N_1293);
and U2045 (N_2045,N_1545,N_1425);
nand U2046 (N_2046,N_1780,N_1795);
or U2047 (N_2047,N_1853,N_1360);
nand U2048 (N_2048,N_1129,N_1524);
or U2049 (N_2049,N_1055,N_1279);
nor U2050 (N_2050,N_1741,N_1234);
nand U2051 (N_2051,N_1845,N_1280);
or U2052 (N_2052,N_1282,N_1270);
or U2053 (N_2053,N_1842,N_1441);
and U2054 (N_2054,N_1454,N_1126);
or U2055 (N_2055,N_1963,N_1542);
nand U2056 (N_2056,N_1355,N_1701);
and U2057 (N_2057,N_1628,N_1073);
nand U2058 (N_2058,N_1734,N_1285);
nor U2059 (N_2059,N_1026,N_1958);
nor U2060 (N_2060,N_1577,N_1171);
or U2061 (N_2061,N_1563,N_1539);
nor U2062 (N_2062,N_1692,N_1918);
nand U2063 (N_2063,N_1582,N_1051);
or U2064 (N_2064,N_1431,N_1316);
nand U2065 (N_2065,N_1034,N_1823);
and U2066 (N_2066,N_1287,N_1778);
or U2067 (N_2067,N_1190,N_1605);
nand U2068 (N_2068,N_1056,N_1206);
nor U2069 (N_2069,N_1301,N_1302);
or U2070 (N_2070,N_1307,N_1760);
or U2071 (N_2071,N_1383,N_1909);
and U2072 (N_2072,N_1158,N_1254);
nor U2073 (N_2073,N_1331,N_1311);
nand U2074 (N_2074,N_1757,N_1322);
nor U2075 (N_2075,N_1064,N_1233);
and U2076 (N_2076,N_1966,N_1676);
nor U2077 (N_2077,N_1050,N_1871);
or U2078 (N_2078,N_1394,N_1392);
and U2079 (N_2079,N_1679,N_1986);
nand U2080 (N_2080,N_1767,N_1065);
or U2081 (N_2081,N_1609,N_1898);
or U2082 (N_2082,N_1049,N_1434);
nor U2083 (N_2083,N_1385,N_1604);
and U2084 (N_2084,N_1784,N_1365);
and U2085 (N_2085,N_1841,N_1553);
xnor U2086 (N_2086,N_1782,N_1173);
or U2087 (N_2087,N_1862,N_1452);
nor U2088 (N_2088,N_1957,N_1276);
and U2089 (N_2089,N_1366,N_1805);
or U2090 (N_2090,N_1572,N_1426);
or U2091 (N_2091,N_1225,N_1914);
and U2092 (N_2092,N_1011,N_1399);
nand U2093 (N_2093,N_1999,N_1540);
nor U2094 (N_2094,N_1231,N_1555);
and U2095 (N_2095,N_1201,N_1032);
nand U2096 (N_2096,N_1490,N_1445);
or U2097 (N_2097,N_1894,N_1010);
or U2098 (N_2098,N_1950,N_1813);
and U2099 (N_2099,N_1801,N_1720);
or U2100 (N_2100,N_1977,N_1954);
and U2101 (N_2101,N_1507,N_1086);
nand U2102 (N_2102,N_1758,N_1885);
or U2103 (N_2103,N_1825,N_1486);
nor U2104 (N_2104,N_1151,N_1740);
or U2105 (N_2105,N_1672,N_1736);
nor U2106 (N_2106,N_1994,N_1063);
or U2107 (N_2107,N_1807,N_1905);
and U2108 (N_2108,N_1779,N_1873);
or U2109 (N_2109,N_1960,N_1774);
and U2110 (N_2110,N_1913,N_1737);
or U2111 (N_2111,N_1875,N_1495);
or U2112 (N_2112,N_1226,N_1600);
or U2113 (N_2113,N_1012,N_1180);
nor U2114 (N_2114,N_1143,N_1220);
and U2115 (N_2115,N_1378,N_1968);
nor U2116 (N_2116,N_1797,N_1552);
nor U2117 (N_2117,N_1567,N_1127);
or U2118 (N_2118,N_1204,N_1221);
nand U2119 (N_2119,N_1649,N_1297);
and U2120 (N_2120,N_1982,N_1437);
nand U2121 (N_2121,N_1453,N_1154);
or U2122 (N_2122,N_1788,N_1062);
and U2123 (N_2123,N_1705,N_1576);
nor U2124 (N_2124,N_1541,N_1506);
or U2125 (N_2125,N_1447,N_1653);
and U2126 (N_2126,N_1996,N_1723);
nand U2127 (N_2127,N_1989,N_1256);
or U2128 (N_2128,N_1700,N_1038);
nor U2129 (N_2129,N_1732,N_1008);
and U2130 (N_2130,N_1834,N_1559);
nand U2131 (N_2131,N_1090,N_1864);
or U2132 (N_2132,N_1512,N_1754);
and U2133 (N_2133,N_1759,N_1005);
nand U2134 (N_2134,N_1388,N_1586);
and U2135 (N_2135,N_1899,N_1024);
nor U2136 (N_2136,N_1943,N_1728);
nor U2137 (N_2137,N_1810,N_1155);
and U2138 (N_2138,N_1418,N_1761);
nor U2139 (N_2139,N_1537,N_1648);
or U2140 (N_2140,N_1948,N_1466);
or U2141 (N_2141,N_1775,N_1638);
nand U2142 (N_2142,N_1236,N_1688);
and U2143 (N_2143,N_1248,N_1626);
or U2144 (N_2144,N_1997,N_1592);
and U2145 (N_2145,N_1613,N_1346);
nand U2146 (N_2146,N_1928,N_1518);
nand U2147 (N_2147,N_1227,N_1580);
nor U2148 (N_2148,N_1040,N_1255);
or U2149 (N_2149,N_1962,N_1169);
nand U2150 (N_2150,N_1861,N_1944);
nor U2151 (N_2151,N_1423,N_1726);
nand U2152 (N_2152,N_1375,N_1473);
nand U2153 (N_2153,N_1137,N_1854);
or U2154 (N_2154,N_1892,N_1926);
nand U2155 (N_2155,N_1463,N_1902);
nor U2156 (N_2156,N_1891,N_1458);
nor U2157 (N_2157,N_1157,N_1940);
or U2158 (N_2158,N_1361,N_1593);
and U2159 (N_2159,N_1095,N_1596);
nand U2160 (N_2160,N_1059,N_1160);
nand U2161 (N_2161,N_1694,N_1646);
or U2162 (N_2162,N_1876,N_1670);
or U2163 (N_2163,N_1607,N_1205);
nor U2164 (N_2164,N_1578,N_1353);
or U2165 (N_2165,N_1851,N_1074);
nor U2166 (N_2166,N_1315,N_1715);
nand U2167 (N_2167,N_1475,N_1247);
and U2168 (N_2168,N_1152,N_1414);
or U2169 (N_2169,N_1739,N_1884);
and U2170 (N_2170,N_1993,N_1102);
nand U2171 (N_2171,N_1494,N_1422);
or U2172 (N_2172,N_1401,N_1377);
or U2173 (N_2173,N_1069,N_1800);
and U2174 (N_2174,N_1751,N_1624);
nand U2175 (N_2175,N_1719,N_1462);
nand U2176 (N_2176,N_1047,N_1148);
and U2177 (N_2177,N_1440,N_1502);
nor U2178 (N_2178,N_1548,N_1343);
nand U2179 (N_2179,N_1564,N_1748);
nor U2180 (N_2180,N_1043,N_1253);
and U2181 (N_2181,N_1789,N_1749);
or U2182 (N_2182,N_1855,N_1538);
and U2183 (N_2183,N_1114,N_1122);
nor U2184 (N_2184,N_1641,N_1668);
and U2185 (N_2185,N_1199,N_1023);
nor U2186 (N_2186,N_1274,N_1992);
and U2187 (N_2187,N_1953,N_1232);
and U2188 (N_2188,N_1275,N_1265);
or U2189 (N_2189,N_1844,N_1756);
nor U2190 (N_2190,N_1919,N_1883);
nor U2191 (N_2191,N_1669,N_1048);
and U2192 (N_2192,N_1216,N_1893);
nor U2193 (N_2193,N_1250,N_1526);
xor U2194 (N_2194,N_1956,N_1584);
nor U2195 (N_2195,N_1744,N_1570);
or U2196 (N_2196,N_1571,N_1395);
and U2197 (N_2197,N_1470,N_1620);
and U2198 (N_2198,N_1908,N_1619);
or U2199 (N_2199,N_1106,N_1391);
nand U2200 (N_2200,N_1104,N_1773);
or U2201 (N_2201,N_1061,N_1309);
or U2202 (N_2202,N_1182,N_1268);
nor U2203 (N_2203,N_1257,N_1429);
and U2204 (N_2204,N_1725,N_1017);
nor U2205 (N_2205,N_1295,N_1030);
nor U2206 (N_2206,N_1822,N_1769);
or U2207 (N_2207,N_1376,N_1405);
and U2208 (N_2208,N_1738,N_1667);
or U2209 (N_2209,N_1211,N_1410);
or U2210 (N_2210,N_1080,N_1194);
and U2211 (N_2211,N_1528,N_1735);
nand U2212 (N_2212,N_1887,N_1318);
or U2213 (N_2213,N_1820,N_1016);
and U2214 (N_2214,N_1703,N_1614);
or U2215 (N_2215,N_1041,N_1469);
nor U2216 (N_2216,N_1504,N_1547);
or U2217 (N_2217,N_1031,N_1264);
nand U2218 (N_2218,N_1103,N_1792);
or U2219 (N_2219,N_1153,N_1079);
nor U2220 (N_2220,N_1632,N_1092);
or U2221 (N_2221,N_1386,N_1611);
and U2222 (N_2222,N_1149,N_1093);
nor U2223 (N_2223,N_1289,N_1053);
nand U2224 (N_2224,N_1076,N_1729);
nand U2225 (N_2225,N_1590,N_1067);
or U2226 (N_2226,N_1144,N_1186);
or U2227 (N_2227,N_1991,N_1942);
or U2228 (N_2228,N_1438,N_1094);
nor U2229 (N_2229,N_1832,N_1777);
nand U2230 (N_2230,N_1197,N_1793);
or U2231 (N_2231,N_1100,N_1403);
or U2232 (N_2232,N_1852,N_1242);
or U2233 (N_2233,N_1698,N_1896);
nand U2234 (N_2234,N_1436,N_1184);
nand U2235 (N_2235,N_1675,N_1981);
nor U2236 (N_2236,N_1284,N_1099);
nand U2237 (N_2237,N_1606,N_1665);
or U2238 (N_2238,N_1002,N_1058);
nand U2239 (N_2239,N_1818,N_1168);
nand U2240 (N_2240,N_1880,N_1416);
and U2241 (N_2241,N_1147,N_1511);
nor U2242 (N_2242,N_1830,N_1098);
or U2243 (N_2243,N_1762,N_1323);
xnor U2244 (N_2244,N_1573,N_1591);
or U2245 (N_2245,N_1858,N_1872);
or U2246 (N_2246,N_1121,N_1747);
or U2247 (N_2247,N_1616,N_1140);
nor U2248 (N_2248,N_1124,N_1397);
nor U2249 (N_2249,N_1217,N_1686);
nand U2250 (N_2250,N_1835,N_1803);
or U2251 (N_2251,N_1312,N_1923);
nor U2252 (N_2252,N_1681,N_1695);
nand U2253 (N_2253,N_1101,N_1645);
nand U2254 (N_2254,N_1910,N_1785);
or U2255 (N_2255,N_1164,N_1594);
and U2256 (N_2256,N_1671,N_1984);
nor U2257 (N_2257,N_1411,N_1961);
nor U2258 (N_2258,N_1687,N_1156);
nand U2259 (N_2259,N_1136,N_1581);
nand U2260 (N_2260,N_1179,N_1513);
nand U2261 (N_2261,N_1828,N_1198);
nand U2262 (N_2262,N_1721,N_1831);
nand U2263 (N_2263,N_1650,N_1230);
and U2264 (N_2264,N_1111,N_1046);
and U2265 (N_2265,N_1890,N_1271);
or U2266 (N_2266,N_1409,N_1783);
nand U2267 (N_2267,N_1025,N_1569);
and U2268 (N_2268,N_1252,N_1183);
or U2269 (N_2269,N_1975,N_1543);
and U2270 (N_2270,N_1798,N_1146);
or U2271 (N_2271,N_1174,N_1970);
and U2272 (N_2272,N_1678,N_1219);
and U2273 (N_2273,N_1655,N_1618);
and U2274 (N_2274,N_1480,N_1172);
nand U2275 (N_2275,N_1393,N_1460);
nor U2276 (N_2276,N_1863,N_1176);
and U2277 (N_2277,N_1551,N_1461);
nand U2278 (N_2278,N_1224,N_1574);
nor U2279 (N_2279,N_1682,N_1763);
nor U2280 (N_2280,N_1796,N_1249);
nand U2281 (N_2281,N_1556,N_1903);
and U2282 (N_2282,N_1654,N_1433);
or U2283 (N_2283,N_1001,N_1406);
nor U2284 (N_2284,N_1471,N_1658);
or U2285 (N_2285,N_1474,N_1313);
nor U2286 (N_2286,N_1382,N_1768);
and U2287 (N_2287,N_1283,N_1060);
nor U2288 (N_2288,N_1131,N_1195);
and U2289 (N_2289,N_1509,N_1498);
nor U2290 (N_2290,N_1530,N_1491);
nand U2291 (N_2291,N_1941,N_1636);
or U2292 (N_2292,N_1192,N_1118);
and U2293 (N_2293,N_1035,N_1704);
or U2294 (N_2294,N_1499,N_1931);
or U2295 (N_2295,N_1446,N_1371);
and U2296 (N_2296,N_1381,N_1693);
nor U2297 (N_2297,N_1995,N_1263);
or U2298 (N_2298,N_1519,N_1699);
nor U2299 (N_2299,N_1527,N_1266);
nand U2300 (N_2300,N_1652,N_1869);
nand U2301 (N_2301,N_1806,N_1979);
and U2302 (N_2302,N_1623,N_1349);
nor U2303 (N_2303,N_1117,N_1750);
nor U2304 (N_2304,N_1123,N_1477);
and U2305 (N_2305,N_1332,N_1334);
and U2306 (N_2306,N_1013,N_1430);
and U2307 (N_2307,N_1262,N_1326);
and U2308 (N_2308,N_1710,N_1110);
and U2309 (N_2309,N_1344,N_1130);
nand U2310 (N_2310,N_1291,N_1697);
and U2311 (N_2311,N_1847,N_1878);
and U2312 (N_2312,N_1866,N_1412);
nand U2313 (N_2313,N_1338,N_1327);
or U2314 (N_2314,N_1901,N_1533);
nor U2315 (N_2315,N_1210,N_1588);
or U2316 (N_2316,N_1081,N_1610);
nor U2317 (N_2317,N_1178,N_1003);
nor U2318 (N_2318,N_1398,N_1229);
and U2319 (N_2319,N_1286,N_1298);
nand U2320 (N_2320,N_1998,N_1881);
nand U2321 (N_2321,N_1163,N_1451);
or U2322 (N_2322,N_1243,N_1536);
nand U2323 (N_2323,N_1057,N_1496);
nand U2324 (N_2324,N_1575,N_1339);
nor U2325 (N_2325,N_1935,N_1595);
and U2326 (N_2326,N_1340,N_1755);
or U2327 (N_2327,N_1333,N_1990);
nor U2328 (N_2328,N_1390,N_1731);
or U2329 (N_2329,N_1833,N_1921);
and U2330 (N_2330,N_1407,N_1052);
and U2331 (N_2331,N_1364,N_1362);
nor U2332 (N_2332,N_1816,N_1321);
nand U2333 (N_2333,N_1359,N_1971);
or U2334 (N_2334,N_1036,N_1689);
nand U2335 (N_2335,N_1838,N_1415);
and U2336 (N_2336,N_1680,N_1709);
nor U2337 (N_2337,N_1549,N_1419);
nor U2338 (N_2338,N_1325,N_1134);
nor U2339 (N_2339,N_1608,N_1181);
nor U2340 (N_2340,N_1072,N_1683);
and U2341 (N_2341,N_1980,N_1505);
nor U2342 (N_2342,N_1879,N_1037);
or U2343 (N_2343,N_1317,N_1912);
and U2344 (N_2344,N_1617,N_1877);
nor U2345 (N_2345,N_1625,N_1351);
and U2346 (N_2346,N_1379,N_1459);
nor U2347 (N_2347,N_1482,N_1267);
and U2348 (N_2348,N_1196,N_1868);
or U2349 (N_2349,N_1150,N_1347);
and U2350 (N_2350,N_1843,N_1808);
xor U2351 (N_2351,N_1116,N_1622);
and U2352 (N_2352,N_1142,N_1310);
nor U2353 (N_2353,N_1448,N_1292);
nand U2354 (N_2354,N_1520,N_1396);
or U2355 (N_2355,N_1215,N_1139);
and U2356 (N_2356,N_1846,N_1408);
or U2357 (N_2357,N_1684,N_1696);
and U2358 (N_2358,N_1484,N_1087);
nand U2359 (N_2359,N_1952,N_1900);
and U2360 (N_2360,N_1657,N_1239);
nand U2361 (N_2361,N_1358,N_1706);
nand U2362 (N_2362,N_1612,N_1075);
and U2363 (N_2363,N_1916,N_1870);
and U2364 (N_2364,N_1084,N_1691);
nor U2365 (N_2365,N_1456,N_1373);
or U2366 (N_2366,N_1108,N_1907);
nand U2367 (N_2367,N_1077,N_1455);
and U2368 (N_2368,N_1949,N_1175);
nand U2369 (N_2369,N_1521,N_1827);
or U2370 (N_2370,N_1630,N_1020);
or U2371 (N_2371,N_1449,N_1516);
and U2372 (N_2372,N_1787,N_1583);
and U2373 (N_2373,N_1664,N_1203);
or U2374 (N_2374,N_1812,N_1272);
and U2375 (N_2375,N_1068,N_1345);
and U2376 (N_2376,N_1978,N_1021);
xor U2377 (N_2377,N_1303,N_1874);
and U2378 (N_2378,N_1566,N_1413);
nor U2379 (N_2379,N_1702,N_1746);
nor U2380 (N_2380,N_1936,N_1476);
nand U2381 (N_2381,N_1368,N_1922);
or U2382 (N_2382,N_1141,N_1510);
nand U2383 (N_2383,N_1299,N_1132);
or U2384 (N_2384,N_1930,N_1727);
and U2385 (N_2385,N_1337,N_1850);
nand U2386 (N_2386,N_1708,N_1367);
nor U2387 (N_2387,N_1352,N_1170);
nor U2388 (N_2388,N_1925,N_1083);
nand U2389 (N_2389,N_1420,N_1135);
nor U2390 (N_2390,N_1951,N_1976);
nor U2391 (N_2391,N_1404,N_1945);
and U2392 (N_2392,N_1640,N_1985);
nand U2393 (N_2393,N_1044,N_1947);
nand U2394 (N_2394,N_1895,N_1089);
nor U2395 (N_2395,N_1417,N_1492);
and U2396 (N_2396,N_1627,N_1166);
nor U2397 (N_2397,N_1629,N_1222);
nor U2398 (N_2398,N_1223,N_1532);
or U2399 (N_2399,N_1314,N_1826);
and U2400 (N_2400,N_1483,N_1802);
xnor U2401 (N_2401,N_1601,N_1374);
or U2402 (N_2402,N_1320,N_1799);
nand U2403 (N_2403,N_1860,N_1674);
and U2404 (N_2404,N_1113,N_1439);
and U2405 (N_2405,N_1522,N_1435);
or U2406 (N_2406,N_1096,N_1213);
or U2407 (N_2407,N_1815,N_1119);
or U2408 (N_2408,N_1904,N_1933);
or U2409 (N_2409,N_1647,N_1296);
nor U2410 (N_2410,N_1218,N_1467);
or U2411 (N_2411,N_1690,N_1442);
and U2412 (N_2412,N_1514,N_1489);
nand U2413 (N_2413,N_1915,N_1685);
nor U2414 (N_2414,N_1840,N_1939);
or U2415 (N_2415,N_1207,N_1730);
or U2416 (N_2416,N_1809,N_1464);
or U2417 (N_2417,N_1007,N_1714);
nand U2418 (N_2418,N_1712,N_1523);
nor U2419 (N_2419,N_1742,N_1235);
nor U2420 (N_2420,N_1865,N_1427);
nand U2421 (N_2421,N_1018,N_1251);
and U2422 (N_2422,N_1014,N_1209);
or U2423 (N_2423,N_1557,N_1260);
and U2424 (N_2424,N_1228,N_1639);
nor U2425 (N_2425,N_1814,N_1938);
or U2426 (N_2426,N_1319,N_1946);
or U2427 (N_2427,N_1277,N_1713);
nand U2428 (N_2428,N_1485,N_1821);
nand U2429 (N_2429,N_1882,N_1004);
nand U2430 (N_2430,N_1294,N_1964);
nor U2431 (N_2431,N_1724,N_1554);
or U2432 (N_2432,N_1917,N_1350);
or U2433 (N_2433,N_1525,N_1372);
nor U2434 (N_2434,N_1988,N_1273);
nand U2435 (N_2435,N_1631,N_1824);
and U2436 (N_2436,N_1562,N_1039);
and U2437 (N_2437,N_1987,N_1603);
nor U2438 (N_2438,N_1660,N_1300);
or U2439 (N_2439,N_1753,N_1078);
nor U2440 (N_2440,N_1794,N_1082);
nand U2441 (N_2441,N_1811,N_1776);
nand U2442 (N_2442,N_1973,N_1535);
and U2443 (N_2443,N_1488,N_1642);
nor U2444 (N_2444,N_1621,N_1837);
nand U2445 (N_2445,N_1308,N_1771);
or U2446 (N_2446,N_1666,N_1568);
and U2447 (N_2447,N_1829,N_1597);
and U2448 (N_2448,N_1819,N_1924);
or U2449 (N_2449,N_1889,N_1015);
nor U2450 (N_2450,N_1766,N_1212);
nand U2451 (N_2451,N_1045,N_1849);
nor U2452 (N_2452,N_1244,N_1125);
and U2453 (N_2453,N_1306,N_1478);
nor U2454 (N_2454,N_1969,N_1493);
nand U2455 (N_2455,N_1772,N_1508);
and U2456 (N_2456,N_1191,N_1897);
nor U2457 (N_2457,N_1733,N_1259);
nor U2458 (N_2458,N_1341,N_1633);
nand U2459 (N_2459,N_1428,N_1859);
nor U2460 (N_2460,N_1185,N_1457);
nor U2461 (N_2461,N_1529,N_1560);
nor U2462 (N_2462,N_1711,N_1348);
nor U2463 (N_2463,N_1965,N_1546);
nor U2464 (N_2464,N_1932,N_1328);
or U2465 (N_2465,N_1817,N_1330);
nand U2466 (N_2466,N_1278,N_1929);
or U2467 (N_2467,N_1159,N_1479);
nand U2468 (N_2468,N_1587,N_1677);
and U2469 (N_2469,N_1029,N_1387);
nand U2470 (N_2470,N_1867,N_1145);
nor U2471 (N_2471,N_1972,N_1432);
or U2472 (N_2472,N_1615,N_1550);
nor U2473 (N_2473,N_1290,N_1839);
or U2474 (N_2474,N_1269,N_1336);
or U2475 (N_2475,N_1006,N_1836);
and U2476 (N_2476,N_1468,N_1967);
nor U2477 (N_2477,N_1745,N_1503);
or U2478 (N_2478,N_1070,N_1019);
or U2479 (N_2479,N_1187,N_1465);
nor U2480 (N_2480,N_1133,N_1565);
nand U2481 (N_2481,N_1558,N_1500);
nand U2482 (N_2482,N_1161,N_1109);
and U2483 (N_2483,N_1673,N_1329);
nand U2484 (N_2484,N_1054,N_1033);
or U2485 (N_2485,N_1370,N_1028);
and U2486 (N_2486,N_1450,N_1369);
and U2487 (N_2487,N_1384,N_1167);
nand U2488 (N_2488,N_1927,N_1097);
nor U2489 (N_2489,N_1707,N_1515);
nor U2490 (N_2490,N_1598,N_1088);
nand U2491 (N_2491,N_1561,N_1602);
nand U2492 (N_2492,N_1200,N_1138);
nand U2493 (N_2493,N_1661,N_1342);
nor U2494 (N_2494,N_1356,N_1443);
and U2495 (N_2495,N_1421,N_1497);
nor U2496 (N_2496,N_1107,N_1663);
nand U2497 (N_2497,N_1906,N_1716);
and U2498 (N_2498,N_1659,N_1790);
nor U2499 (N_2499,N_1363,N_1444);
and U2500 (N_2500,N_1204,N_1640);
or U2501 (N_2501,N_1205,N_1106);
and U2502 (N_2502,N_1800,N_1878);
or U2503 (N_2503,N_1408,N_1528);
and U2504 (N_2504,N_1679,N_1686);
and U2505 (N_2505,N_1133,N_1833);
nor U2506 (N_2506,N_1759,N_1874);
and U2507 (N_2507,N_1603,N_1936);
nand U2508 (N_2508,N_1908,N_1634);
or U2509 (N_2509,N_1873,N_1143);
and U2510 (N_2510,N_1372,N_1709);
and U2511 (N_2511,N_1971,N_1548);
nor U2512 (N_2512,N_1879,N_1194);
nor U2513 (N_2513,N_1715,N_1022);
nand U2514 (N_2514,N_1836,N_1282);
or U2515 (N_2515,N_1235,N_1666);
nor U2516 (N_2516,N_1542,N_1574);
and U2517 (N_2517,N_1538,N_1350);
nand U2518 (N_2518,N_1912,N_1665);
and U2519 (N_2519,N_1511,N_1123);
nor U2520 (N_2520,N_1654,N_1327);
nor U2521 (N_2521,N_1805,N_1314);
nand U2522 (N_2522,N_1136,N_1232);
and U2523 (N_2523,N_1941,N_1260);
nor U2524 (N_2524,N_1031,N_1314);
nand U2525 (N_2525,N_1389,N_1367);
nand U2526 (N_2526,N_1396,N_1235);
or U2527 (N_2527,N_1570,N_1173);
and U2528 (N_2528,N_1441,N_1120);
and U2529 (N_2529,N_1531,N_1070);
or U2530 (N_2530,N_1615,N_1017);
nand U2531 (N_2531,N_1295,N_1399);
and U2532 (N_2532,N_1096,N_1456);
or U2533 (N_2533,N_1108,N_1361);
nand U2534 (N_2534,N_1674,N_1036);
and U2535 (N_2535,N_1125,N_1479);
nor U2536 (N_2536,N_1000,N_1848);
nand U2537 (N_2537,N_1930,N_1389);
or U2538 (N_2538,N_1921,N_1442);
nand U2539 (N_2539,N_1003,N_1725);
nor U2540 (N_2540,N_1856,N_1650);
nor U2541 (N_2541,N_1624,N_1829);
nand U2542 (N_2542,N_1297,N_1203);
nor U2543 (N_2543,N_1915,N_1421);
and U2544 (N_2544,N_1654,N_1820);
and U2545 (N_2545,N_1745,N_1305);
nand U2546 (N_2546,N_1321,N_1314);
or U2547 (N_2547,N_1355,N_1432);
or U2548 (N_2548,N_1209,N_1845);
nand U2549 (N_2549,N_1232,N_1013);
or U2550 (N_2550,N_1629,N_1922);
and U2551 (N_2551,N_1159,N_1929);
nand U2552 (N_2552,N_1391,N_1545);
nor U2553 (N_2553,N_1980,N_1652);
and U2554 (N_2554,N_1581,N_1907);
or U2555 (N_2555,N_1467,N_1015);
or U2556 (N_2556,N_1399,N_1812);
nor U2557 (N_2557,N_1451,N_1941);
and U2558 (N_2558,N_1664,N_1290);
nand U2559 (N_2559,N_1785,N_1319);
and U2560 (N_2560,N_1830,N_1224);
nor U2561 (N_2561,N_1814,N_1437);
nand U2562 (N_2562,N_1936,N_1239);
nand U2563 (N_2563,N_1376,N_1524);
xnor U2564 (N_2564,N_1797,N_1946);
nor U2565 (N_2565,N_1865,N_1946);
and U2566 (N_2566,N_1928,N_1049);
and U2567 (N_2567,N_1349,N_1040);
nor U2568 (N_2568,N_1274,N_1856);
or U2569 (N_2569,N_1246,N_1009);
and U2570 (N_2570,N_1642,N_1351);
nor U2571 (N_2571,N_1004,N_1831);
xnor U2572 (N_2572,N_1813,N_1626);
nor U2573 (N_2573,N_1561,N_1247);
and U2574 (N_2574,N_1127,N_1625);
or U2575 (N_2575,N_1898,N_1532);
nand U2576 (N_2576,N_1547,N_1402);
or U2577 (N_2577,N_1932,N_1465);
or U2578 (N_2578,N_1882,N_1355);
or U2579 (N_2579,N_1618,N_1793);
nor U2580 (N_2580,N_1041,N_1974);
and U2581 (N_2581,N_1388,N_1175);
nand U2582 (N_2582,N_1428,N_1662);
nor U2583 (N_2583,N_1755,N_1751);
or U2584 (N_2584,N_1069,N_1911);
and U2585 (N_2585,N_1541,N_1333);
nor U2586 (N_2586,N_1502,N_1330);
nor U2587 (N_2587,N_1647,N_1301);
nand U2588 (N_2588,N_1270,N_1514);
or U2589 (N_2589,N_1505,N_1884);
or U2590 (N_2590,N_1145,N_1787);
and U2591 (N_2591,N_1316,N_1100);
nand U2592 (N_2592,N_1647,N_1963);
or U2593 (N_2593,N_1328,N_1882);
and U2594 (N_2594,N_1928,N_1355);
nor U2595 (N_2595,N_1112,N_1730);
nand U2596 (N_2596,N_1564,N_1146);
nor U2597 (N_2597,N_1602,N_1169);
and U2598 (N_2598,N_1450,N_1683);
or U2599 (N_2599,N_1605,N_1438);
nor U2600 (N_2600,N_1555,N_1347);
nor U2601 (N_2601,N_1647,N_1743);
and U2602 (N_2602,N_1719,N_1029);
nor U2603 (N_2603,N_1633,N_1327);
nand U2604 (N_2604,N_1384,N_1773);
or U2605 (N_2605,N_1356,N_1750);
nand U2606 (N_2606,N_1711,N_1746);
or U2607 (N_2607,N_1240,N_1523);
nand U2608 (N_2608,N_1777,N_1025);
nand U2609 (N_2609,N_1739,N_1723);
nand U2610 (N_2610,N_1765,N_1754);
or U2611 (N_2611,N_1321,N_1642);
nor U2612 (N_2612,N_1509,N_1468);
xnor U2613 (N_2613,N_1790,N_1680);
nand U2614 (N_2614,N_1730,N_1637);
and U2615 (N_2615,N_1368,N_1504);
and U2616 (N_2616,N_1706,N_1871);
nand U2617 (N_2617,N_1809,N_1677);
or U2618 (N_2618,N_1691,N_1211);
nand U2619 (N_2619,N_1789,N_1365);
nor U2620 (N_2620,N_1950,N_1045);
and U2621 (N_2621,N_1159,N_1628);
or U2622 (N_2622,N_1352,N_1292);
nand U2623 (N_2623,N_1113,N_1589);
or U2624 (N_2624,N_1393,N_1045);
and U2625 (N_2625,N_1061,N_1710);
and U2626 (N_2626,N_1409,N_1819);
or U2627 (N_2627,N_1101,N_1607);
nand U2628 (N_2628,N_1078,N_1478);
or U2629 (N_2629,N_1895,N_1942);
nand U2630 (N_2630,N_1770,N_1616);
nand U2631 (N_2631,N_1094,N_1218);
nor U2632 (N_2632,N_1938,N_1060);
nor U2633 (N_2633,N_1235,N_1231);
or U2634 (N_2634,N_1592,N_1324);
or U2635 (N_2635,N_1573,N_1211);
nand U2636 (N_2636,N_1200,N_1949);
and U2637 (N_2637,N_1142,N_1602);
nand U2638 (N_2638,N_1686,N_1597);
and U2639 (N_2639,N_1112,N_1737);
nand U2640 (N_2640,N_1070,N_1893);
nand U2641 (N_2641,N_1512,N_1513);
and U2642 (N_2642,N_1213,N_1328);
nor U2643 (N_2643,N_1466,N_1372);
or U2644 (N_2644,N_1778,N_1668);
nand U2645 (N_2645,N_1714,N_1959);
nor U2646 (N_2646,N_1345,N_1600);
or U2647 (N_2647,N_1537,N_1213);
nand U2648 (N_2648,N_1931,N_1872);
nor U2649 (N_2649,N_1016,N_1341);
or U2650 (N_2650,N_1866,N_1515);
or U2651 (N_2651,N_1921,N_1254);
and U2652 (N_2652,N_1687,N_1509);
and U2653 (N_2653,N_1154,N_1407);
and U2654 (N_2654,N_1326,N_1406);
or U2655 (N_2655,N_1048,N_1382);
nor U2656 (N_2656,N_1782,N_1238);
or U2657 (N_2657,N_1097,N_1432);
or U2658 (N_2658,N_1516,N_1261);
and U2659 (N_2659,N_1566,N_1213);
nand U2660 (N_2660,N_1323,N_1542);
nand U2661 (N_2661,N_1000,N_1270);
nor U2662 (N_2662,N_1124,N_1556);
or U2663 (N_2663,N_1808,N_1241);
nand U2664 (N_2664,N_1563,N_1677);
or U2665 (N_2665,N_1397,N_1129);
nand U2666 (N_2666,N_1891,N_1543);
or U2667 (N_2667,N_1200,N_1102);
nand U2668 (N_2668,N_1440,N_1915);
nor U2669 (N_2669,N_1151,N_1539);
or U2670 (N_2670,N_1254,N_1518);
and U2671 (N_2671,N_1803,N_1423);
nor U2672 (N_2672,N_1430,N_1993);
nor U2673 (N_2673,N_1501,N_1729);
and U2674 (N_2674,N_1664,N_1511);
nor U2675 (N_2675,N_1647,N_1763);
or U2676 (N_2676,N_1683,N_1529);
or U2677 (N_2677,N_1575,N_1374);
nand U2678 (N_2678,N_1356,N_1576);
nand U2679 (N_2679,N_1145,N_1186);
nand U2680 (N_2680,N_1136,N_1883);
nand U2681 (N_2681,N_1652,N_1546);
and U2682 (N_2682,N_1724,N_1453);
nand U2683 (N_2683,N_1697,N_1967);
nand U2684 (N_2684,N_1347,N_1106);
nand U2685 (N_2685,N_1679,N_1611);
nand U2686 (N_2686,N_1121,N_1810);
nand U2687 (N_2687,N_1255,N_1870);
nand U2688 (N_2688,N_1884,N_1352);
and U2689 (N_2689,N_1203,N_1146);
nand U2690 (N_2690,N_1117,N_1966);
and U2691 (N_2691,N_1792,N_1539);
nand U2692 (N_2692,N_1583,N_1470);
or U2693 (N_2693,N_1870,N_1593);
nor U2694 (N_2694,N_1446,N_1569);
and U2695 (N_2695,N_1832,N_1906);
or U2696 (N_2696,N_1375,N_1403);
nor U2697 (N_2697,N_1691,N_1742);
nand U2698 (N_2698,N_1869,N_1621);
and U2699 (N_2699,N_1669,N_1900);
or U2700 (N_2700,N_1847,N_1020);
or U2701 (N_2701,N_1864,N_1181);
and U2702 (N_2702,N_1252,N_1045);
or U2703 (N_2703,N_1247,N_1447);
xor U2704 (N_2704,N_1671,N_1206);
or U2705 (N_2705,N_1384,N_1996);
nor U2706 (N_2706,N_1509,N_1612);
and U2707 (N_2707,N_1880,N_1924);
or U2708 (N_2708,N_1119,N_1326);
or U2709 (N_2709,N_1241,N_1019);
nand U2710 (N_2710,N_1979,N_1989);
nand U2711 (N_2711,N_1188,N_1154);
nor U2712 (N_2712,N_1344,N_1935);
nand U2713 (N_2713,N_1200,N_1517);
nor U2714 (N_2714,N_1476,N_1315);
nor U2715 (N_2715,N_1825,N_1008);
and U2716 (N_2716,N_1597,N_1981);
nand U2717 (N_2717,N_1513,N_1987);
nor U2718 (N_2718,N_1380,N_1547);
nand U2719 (N_2719,N_1345,N_1945);
nor U2720 (N_2720,N_1601,N_1074);
nor U2721 (N_2721,N_1133,N_1040);
nand U2722 (N_2722,N_1342,N_1447);
nor U2723 (N_2723,N_1558,N_1806);
nor U2724 (N_2724,N_1933,N_1543);
nor U2725 (N_2725,N_1943,N_1508);
nand U2726 (N_2726,N_1635,N_1479);
and U2727 (N_2727,N_1379,N_1859);
nand U2728 (N_2728,N_1374,N_1126);
nand U2729 (N_2729,N_1273,N_1667);
nand U2730 (N_2730,N_1268,N_1974);
and U2731 (N_2731,N_1321,N_1293);
nor U2732 (N_2732,N_1333,N_1416);
or U2733 (N_2733,N_1941,N_1034);
or U2734 (N_2734,N_1272,N_1308);
nor U2735 (N_2735,N_1598,N_1627);
and U2736 (N_2736,N_1226,N_1738);
nand U2737 (N_2737,N_1008,N_1248);
or U2738 (N_2738,N_1997,N_1879);
nand U2739 (N_2739,N_1708,N_1423);
or U2740 (N_2740,N_1311,N_1679);
and U2741 (N_2741,N_1643,N_1375);
nor U2742 (N_2742,N_1564,N_1167);
nand U2743 (N_2743,N_1186,N_1053);
nor U2744 (N_2744,N_1524,N_1517);
nor U2745 (N_2745,N_1306,N_1377);
nor U2746 (N_2746,N_1157,N_1681);
or U2747 (N_2747,N_1790,N_1259);
or U2748 (N_2748,N_1645,N_1641);
nor U2749 (N_2749,N_1100,N_1719);
nand U2750 (N_2750,N_1093,N_1013);
nand U2751 (N_2751,N_1363,N_1844);
and U2752 (N_2752,N_1983,N_1286);
nor U2753 (N_2753,N_1997,N_1600);
nand U2754 (N_2754,N_1470,N_1545);
or U2755 (N_2755,N_1357,N_1374);
nor U2756 (N_2756,N_1751,N_1547);
nor U2757 (N_2757,N_1989,N_1900);
nor U2758 (N_2758,N_1793,N_1315);
nor U2759 (N_2759,N_1790,N_1577);
and U2760 (N_2760,N_1498,N_1951);
nand U2761 (N_2761,N_1665,N_1945);
or U2762 (N_2762,N_1580,N_1613);
nor U2763 (N_2763,N_1713,N_1654);
or U2764 (N_2764,N_1747,N_1486);
or U2765 (N_2765,N_1017,N_1765);
nand U2766 (N_2766,N_1166,N_1097);
or U2767 (N_2767,N_1191,N_1256);
nor U2768 (N_2768,N_1712,N_1256);
nor U2769 (N_2769,N_1855,N_1500);
or U2770 (N_2770,N_1171,N_1837);
nand U2771 (N_2771,N_1064,N_1442);
and U2772 (N_2772,N_1825,N_1887);
nand U2773 (N_2773,N_1854,N_1647);
nor U2774 (N_2774,N_1248,N_1639);
nor U2775 (N_2775,N_1414,N_1665);
and U2776 (N_2776,N_1641,N_1913);
or U2777 (N_2777,N_1080,N_1562);
nor U2778 (N_2778,N_1009,N_1516);
or U2779 (N_2779,N_1725,N_1274);
nor U2780 (N_2780,N_1383,N_1130);
nor U2781 (N_2781,N_1057,N_1387);
nor U2782 (N_2782,N_1590,N_1630);
or U2783 (N_2783,N_1047,N_1476);
nand U2784 (N_2784,N_1973,N_1518);
nand U2785 (N_2785,N_1467,N_1712);
nand U2786 (N_2786,N_1293,N_1322);
or U2787 (N_2787,N_1838,N_1302);
and U2788 (N_2788,N_1245,N_1186);
nand U2789 (N_2789,N_1776,N_1097);
and U2790 (N_2790,N_1161,N_1110);
or U2791 (N_2791,N_1161,N_1146);
nor U2792 (N_2792,N_1811,N_1597);
and U2793 (N_2793,N_1635,N_1361);
and U2794 (N_2794,N_1228,N_1559);
nor U2795 (N_2795,N_1806,N_1012);
or U2796 (N_2796,N_1550,N_1679);
nand U2797 (N_2797,N_1565,N_1497);
nand U2798 (N_2798,N_1930,N_1781);
and U2799 (N_2799,N_1106,N_1325);
and U2800 (N_2800,N_1924,N_1824);
nor U2801 (N_2801,N_1962,N_1448);
nand U2802 (N_2802,N_1377,N_1098);
nor U2803 (N_2803,N_1671,N_1590);
and U2804 (N_2804,N_1122,N_1507);
and U2805 (N_2805,N_1231,N_1787);
nand U2806 (N_2806,N_1749,N_1061);
or U2807 (N_2807,N_1021,N_1237);
or U2808 (N_2808,N_1265,N_1447);
and U2809 (N_2809,N_1020,N_1077);
nor U2810 (N_2810,N_1750,N_1999);
or U2811 (N_2811,N_1301,N_1095);
or U2812 (N_2812,N_1398,N_1228);
and U2813 (N_2813,N_1304,N_1545);
nand U2814 (N_2814,N_1370,N_1882);
nand U2815 (N_2815,N_1384,N_1233);
nand U2816 (N_2816,N_1771,N_1855);
nor U2817 (N_2817,N_1765,N_1442);
nor U2818 (N_2818,N_1866,N_1605);
and U2819 (N_2819,N_1085,N_1706);
or U2820 (N_2820,N_1371,N_1478);
or U2821 (N_2821,N_1793,N_1451);
and U2822 (N_2822,N_1076,N_1687);
nand U2823 (N_2823,N_1257,N_1095);
xor U2824 (N_2824,N_1276,N_1221);
nand U2825 (N_2825,N_1112,N_1338);
and U2826 (N_2826,N_1905,N_1594);
nand U2827 (N_2827,N_1075,N_1973);
nand U2828 (N_2828,N_1513,N_1622);
and U2829 (N_2829,N_1581,N_1002);
nor U2830 (N_2830,N_1542,N_1230);
nor U2831 (N_2831,N_1492,N_1155);
and U2832 (N_2832,N_1687,N_1079);
and U2833 (N_2833,N_1333,N_1098);
and U2834 (N_2834,N_1127,N_1114);
and U2835 (N_2835,N_1451,N_1450);
or U2836 (N_2836,N_1371,N_1370);
nand U2837 (N_2837,N_1556,N_1301);
nand U2838 (N_2838,N_1699,N_1535);
nor U2839 (N_2839,N_1205,N_1555);
and U2840 (N_2840,N_1850,N_1384);
and U2841 (N_2841,N_1545,N_1983);
and U2842 (N_2842,N_1184,N_1740);
nand U2843 (N_2843,N_1334,N_1394);
nand U2844 (N_2844,N_1799,N_1588);
nand U2845 (N_2845,N_1570,N_1456);
nand U2846 (N_2846,N_1477,N_1836);
nand U2847 (N_2847,N_1814,N_1185);
or U2848 (N_2848,N_1566,N_1726);
nor U2849 (N_2849,N_1321,N_1382);
nor U2850 (N_2850,N_1779,N_1598);
nand U2851 (N_2851,N_1715,N_1918);
nand U2852 (N_2852,N_1048,N_1911);
nand U2853 (N_2853,N_1756,N_1002);
nand U2854 (N_2854,N_1713,N_1970);
nand U2855 (N_2855,N_1579,N_1240);
or U2856 (N_2856,N_1147,N_1647);
nand U2857 (N_2857,N_1382,N_1484);
nand U2858 (N_2858,N_1423,N_1623);
nand U2859 (N_2859,N_1276,N_1715);
nor U2860 (N_2860,N_1178,N_1688);
or U2861 (N_2861,N_1940,N_1669);
and U2862 (N_2862,N_1156,N_1702);
nand U2863 (N_2863,N_1712,N_1277);
or U2864 (N_2864,N_1891,N_1437);
nor U2865 (N_2865,N_1612,N_1744);
nor U2866 (N_2866,N_1711,N_1673);
and U2867 (N_2867,N_1270,N_1988);
and U2868 (N_2868,N_1880,N_1216);
and U2869 (N_2869,N_1341,N_1388);
nand U2870 (N_2870,N_1232,N_1095);
or U2871 (N_2871,N_1580,N_1352);
nor U2872 (N_2872,N_1825,N_1911);
xnor U2873 (N_2873,N_1084,N_1376);
and U2874 (N_2874,N_1952,N_1695);
nor U2875 (N_2875,N_1023,N_1704);
nand U2876 (N_2876,N_1870,N_1881);
nor U2877 (N_2877,N_1019,N_1111);
nor U2878 (N_2878,N_1352,N_1661);
and U2879 (N_2879,N_1865,N_1993);
nor U2880 (N_2880,N_1333,N_1693);
and U2881 (N_2881,N_1095,N_1231);
or U2882 (N_2882,N_1887,N_1157);
nor U2883 (N_2883,N_1976,N_1248);
or U2884 (N_2884,N_1046,N_1134);
and U2885 (N_2885,N_1257,N_1900);
or U2886 (N_2886,N_1755,N_1920);
and U2887 (N_2887,N_1658,N_1773);
and U2888 (N_2888,N_1421,N_1855);
nor U2889 (N_2889,N_1524,N_1923);
nand U2890 (N_2890,N_1240,N_1182);
or U2891 (N_2891,N_1813,N_1047);
and U2892 (N_2892,N_1425,N_1737);
nor U2893 (N_2893,N_1581,N_1855);
nor U2894 (N_2894,N_1668,N_1241);
nor U2895 (N_2895,N_1744,N_1333);
nor U2896 (N_2896,N_1050,N_1069);
or U2897 (N_2897,N_1829,N_1745);
nor U2898 (N_2898,N_1020,N_1386);
nand U2899 (N_2899,N_1877,N_1055);
and U2900 (N_2900,N_1157,N_1367);
or U2901 (N_2901,N_1975,N_1284);
and U2902 (N_2902,N_1167,N_1088);
or U2903 (N_2903,N_1976,N_1209);
nand U2904 (N_2904,N_1733,N_1516);
and U2905 (N_2905,N_1688,N_1964);
nor U2906 (N_2906,N_1017,N_1805);
and U2907 (N_2907,N_1681,N_1864);
nand U2908 (N_2908,N_1918,N_1211);
or U2909 (N_2909,N_1574,N_1955);
nor U2910 (N_2910,N_1043,N_1414);
nand U2911 (N_2911,N_1009,N_1275);
nand U2912 (N_2912,N_1221,N_1636);
or U2913 (N_2913,N_1264,N_1812);
nand U2914 (N_2914,N_1029,N_1232);
and U2915 (N_2915,N_1296,N_1483);
and U2916 (N_2916,N_1990,N_1056);
nor U2917 (N_2917,N_1649,N_1273);
or U2918 (N_2918,N_1858,N_1982);
or U2919 (N_2919,N_1792,N_1467);
nor U2920 (N_2920,N_1758,N_1478);
nor U2921 (N_2921,N_1334,N_1101);
or U2922 (N_2922,N_1856,N_1786);
nor U2923 (N_2923,N_1115,N_1851);
and U2924 (N_2924,N_1140,N_1732);
nor U2925 (N_2925,N_1939,N_1764);
and U2926 (N_2926,N_1321,N_1943);
and U2927 (N_2927,N_1360,N_1855);
xnor U2928 (N_2928,N_1137,N_1077);
or U2929 (N_2929,N_1305,N_1578);
and U2930 (N_2930,N_1998,N_1430);
and U2931 (N_2931,N_1039,N_1364);
and U2932 (N_2932,N_1453,N_1676);
and U2933 (N_2933,N_1818,N_1450);
nor U2934 (N_2934,N_1329,N_1441);
or U2935 (N_2935,N_1449,N_1462);
and U2936 (N_2936,N_1205,N_1633);
and U2937 (N_2937,N_1869,N_1041);
xor U2938 (N_2938,N_1834,N_1571);
or U2939 (N_2939,N_1914,N_1276);
or U2940 (N_2940,N_1547,N_1045);
nand U2941 (N_2941,N_1039,N_1204);
nand U2942 (N_2942,N_1778,N_1960);
or U2943 (N_2943,N_1034,N_1702);
nor U2944 (N_2944,N_1838,N_1091);
nor U2945 (N_2945,N_1171,N_1020);
or U2946 (N_2946,N_1285,N_1133);
and U2947 (N_2947,N_1202,N_1385);
or U2948 (N_2948,N_1761,N_1678);
nand U2949 (N_2949,N_1372,N_1447);
and U2950 (N_2950,N_1034,N_1601);
nand U2951 (N_2951,N_1551,N_1396);
nor U2952 (N_2952,N_1520,N_1287);
and U2953 (N_2953,N_1770,N_1475);
nor U2954 (N_2954,N_1174,N_1193);
nand U2955 (N_2955,N_1444,N_1553);
or U2956 (N_2956,N_1481,N_1451);
nor U2957 (N_2957,N_1925,N_1900);
or U2958 (N_2958,N_1192,N_1057);
and U2959 (N_2959,N_1360,N_1772);
or U2960 (N_2960,N_1603,N_1308);
nand U2961 (N_2961,N_1750,N_1451);
nand U2962 (N_2962,N_1148,N_1761);
or U2963 (N_2963,N_1439,N_1434);
and U2964 (N_2964,N_1971,N_1951);
and U2965 (N_2965,N_1294,N_1438);
nand U2966 (N_2966,N_1942,N_1232);
nor U2967 (N_2967,N_1864,N_1214);
nor U2968 (N_2968,N_1407,N_1743);
and U2969 (N_2969,N_1919,N_1397);
and U2970 (N_2970,N_1831,N_1361);
nand U2971 (N_2971,N_1142,N_1455);
and U2972 (N_2972,N_1993,N_1250);
nand U2973 (N_2973,N_1234,N_1291);
and U2974 (N_2974,N_1147,N_1738);
nand U2975 (N_2975,N_1527,N_1566);
and U2976 (N_2976,N_1949,N_1421);
nor U2977 (N_2977,N_1076,N_1461);
or U2978 (N_2978,N_1334,N_1253);
nor U2979 (N_2979,N_1333,N_1145);
or U2980 (N_2980,N_1574,N_1535);
or U2981 (N_2981,N_1271,N_1998);
xor U2982 (N_2982,N_1619,N_1887);
nand U2983 (N_2983,N_1037,N_1444);
nand U2984 (N_2984,N_1430,N_1005);
and U2985 (N_2985,N_1459,N_1048);
and U2986 (N_2986,N_1860,N_1597);
nand U2987 (N_2987,N_1607,N_1941);
nor U2988 (N_2988,N_1154,N_1527);
nand U2989 (N_2989,N_1104,N_1687);
and U2990 (N_2990,N_1215,N_1084);
and U2991 (N_2991,N_1069,N_1670);
or U2992 (N_2992,N_1735,N_1935);
and U2993 (N_2993,N_1312,N_1801);
and U2994 (N_2994,N_1644,N_1017);
and U2995 (N_2995,N_1974,N_1438);
or U2996 (N_2996,N_1782,N_1529);
nand U2997 (N_2997,N_1085,N_1566);
or U2998 (N_2998,N_1107,N_1362);
nand U2999 (N_2999,N_1832,N_1294);
or UO_0 (O_0,N_2091,N_2433);
or UO_1 (O_1,N_2481,N_2028);
and UO_2 (O_2,N_2453,N_2190);
nor UO_3 (O_3,N_2323,N_2405);
and UO_4 (O_4,N_2548,N_2460);
nand UO_5 (O_5,N_2712,N_2714);
nand UO_6 (O_6,N_2166,N_2600);
nand UO_7 (O_7,N_2719,N_2769);
or UO_8 (O_8,N_2660,N_2207);
xnor UO_9 (O_9,N_2403,N_2140);
nor UO_10 (O_10,N_2715,N_2902);
nand UO_11 (O_11,N_2117,N_2636);
nand UO_12 (O_12,N_2261,N_2567);
nor UO_13 (O_13,N_2517,N_2195);
or UO_14 (O_14,N_2042,N_2374);
or UO_15 (O_15,N_2844,N_2848);
and UO_16 (O_16,N_2574,N_2711);
or UO_17 (O_17,N_2193,N_2988);
nand UO_18 (O_18,N_2057,N_2620);
xor UO_19 (O_19,N_2992,N_2901);
or UO_20 (O_20,N_2577,N_2016);
and UO_21 (O_21,N_2324,N_2299);
nand UO_22 (O_22,N_2488,N_2101);
or UO_23 (O_23,N_2301,N_2784);
or UO_24 (O_24,N_2480,N_2514);
and UO_25 (O_25,N_2742,N_2796);
and UO_26 (O_26,N_2368,N_2381);
nand UO_27 (O_27,N_2777,N_2765);
and UO_28 (O_28,N_2700,N_2322);
or UO_29 (O_29,N_2321,N_2008);
nor UO_30 (O_30,N_2804,N_2229);
nand UO_31 (O_31,N_2734,N_2341);
and UO_32 (O_32,N_2486,N_2098);
nor UO_33 (O_33,N_2694,N_2684);
nor UO_34 (O_34,N_2814,N_2630);
xor UO_35 (O_35,N_2972,N_2967);
and UO_36 (O_36,N_2653,N_2987);
nor UO_37 (O_37,N_2379,N_2958);
nor UO_38 (O_38,N_2546,N_2552);
nand UO_39 (O_39,N_2566,N_2133);
nor UO_40 (O_40,N_2802,N_2451);
and UO_41 (O_41,N_2220,N_2523);
or UO_42 (O_42,N_2065,N_2670);
or UO_43 (O_43,N_2417,N_2276);
nand UO_44 (O_44,N_2162,N_2128);
and UO_45 (O_45,N_2073,N_2390);
nand UO_46 (O_46,N_2497,N_2896);
nand UO_47 (O_47,N_2255,N_2729);
or UO_48 (O_48,N_2833,N_2353);
nand UO_49 (O_49,N_2204,N_2173);
and UO_50 (O_50,N_2538,N_2860);
and UO_51 (O_51,N_2174,N_2828);
and UO_52 (O_52,N_2268,N_2009);
or UO_53 (O_53,N_2392,N_2948);
or UO_54 (O_54,N_2235,N_2373);
nor UO_55 (O_55,N_2909,N_2606);
nor UO_56 (O_56,N_2741,N_2146);
nor UO_57 (O_57,N_2473,N_2103);
nor UO_58 (O_58,N_2085,N_2384);
and UO_59 (O_59,N_2044,N_2647);
or UO_60 (O_60,N_2316,N_2464);
or UO_61 (O_61,N_2233,N_2601);
and UO_62 (O_62,N_2212,N_2527);
nor UO_63 (O_63,N_2865,N_2690);
or UO_64 (O_64,N_2238,N_2617);
or UO_65 (O_65,N_2918,N_2850);
or UO_66 (O_66,N_2342,N_2831);
or UO_67 (O_67,N_2183,N_2021);
and UO_68 (O_68,N_2161,N_2516);
nand UO_69 (O_69,N_2570,N_2315);
or UO_70 (O_70,N_2651,N_2870);
nor UO_71 (O_71,N_2983,N_2130);
nor UO_72 (O_72,N_2770,N_2641);
nor UO_73 (O_73,N_2924,N_2030);
or UO_74 (O_74,N_2885,N_2244);
or UO_75 (O_75,N_2759,N_2032);
xor UO_76 (O_76,N_2350,N_2726);
or UO_77 (O_77,N_2874,N_2683);
or UO_78 (O_78,N_2731,N_2652);
nor UO_79 (O_79,N_2679,N_2087);
nand UO_80 (O_80,N_2922,N_2525);
nor UO_81 (O_81,N_2422,N_2837);
and UO_82 (O_82,N_2014,N_2940);
and UO_83 (O_83,N_2458,N_2171);
or UO_84 (O_84,N_2155,N_2763);
nor UO_85 (O_85,N_2258,N_2702);
xor UO_86 (O_86,N_2084,N_2164);
and UO_87 (O_87,N_2977,N_2083);
nor UO_88 (O_88,N_2176,N_2781);
nand UO_89 (O_89,N_2891,N_2298);
and UO_90 (O_90,N_2476,N_2920);
nor UO_91 (O_91,N_2709,N_2661);
nand UO_92 (O_92,N_2170,N_2724);
or UO_93 (O_93,N_2555,N_2461);
or UO_94 (O_94,N_2160,N_2478);
or UO_95 (O_95,N_2545,N_2657);
nor UO_96 (O_96,N_2397,N_2696);
nand UO_97 (O_97,N_2968,N_2760);
nor UO_98 (O_98,N_2326,N_2036);
or UO_99 (O_99,N_2986,N_2449);
and UO_100 (O_100,N_2109,N_2883);
or UO_101 (O_101,N_2039,N_2903);
nor UO_102 (O_102,N_2937,N_2232);
and UO_103 (O_103,N_2941,N_2629);
or UO_104 (O_104,N_2144,N_2139);
and UO_105 (O_105,N_2296,N_2794);
nand UO_106 (O_106,N_2692,N_2252);
or UO_107 (O_107,N_2845,N_2020);
and UO_108 (O_108,N_2593,N_2248);
nor UO_109 (O_109,N_2380,N_2245);
or UO_110 (O_110,N_2609,N_2088);
or UO_111 (O_111,N_2406,N_2187);
nand UO_112 (O_112,N_2801,N_2100);
nor UO_113 (O_113,N_2001,N_2884);
and UO_114 (O_114,N_2266,N_2366);
and UO_115 (O_115,N_2753,N_2125);
or UO_116 (O_116,N_2633,N_2442);
nor UO_117 (O_117,N_2049,N_2964);
and UO_118 (O_118,N_2465,N_2169);
and UO_119 (O_119,N_2529,N_2826);
or UO_120 (O_120,N_2613,N_2058);
nand UO_121 (O_121,N_2701,N_2662);
nor UO_122 (O_122,N_2762,N_2910);
and UO_123 (O_123,N_2973,N_2107);
or UO_124 (O_124,N_2185,N_2921);
nor UO_125 (O_125,N_2426,N_2857);
and UO_126 (O_126,N_2391,N_2867);
nand UO_127 (O_127,N_2048,N_2257);
nand UO_128 (O_128,N_2912,N_2188);
and UO_129 (O_129,N_2092,N_2498);
or UO_130 (O_130,N_2589,N_2585);
or UO_131 (O_131,N_2289,N_2596);
nor UO_132 (O_132,N_2587,N_2925);
or UO_133 (O_133,N_2303,N_2056);
and UO_134 (O_134,N_2806,N_2787);
nor UO_135 (O_135,N_2886,N_2519);
nand UO_136 (O_136,N_2797,N_2680);
or UO_137 (O_137,N_2678,N_2539);
nor UO_138 (O_138,N_2191,N_2795);
nor UO_139 (O_139,N_2062,N_2310);
and UO_140 (O_140,N_2788,N_2436);
nand UO_141 (O_141,N_2349,N_2732);
or UO_142 (O_142,N_2231,N_2869);
and UO_143 (O_143,N_2111,N_2597);
nor UO_144 (O_144,N_2178,N_2551);
nor UO_145 (O_145,N_2074,N_2950);
and UO_146 (O_146,N_2544,N_2025);
or UO_147 (O_147,N_2468,N_2329);
or UO_148 (O_148,N_2360,N_2510);
or UO_149 (O_149,N_2003,N_2658);
and UO_150 (O_150,N_2496,N_2619);
nand UO_151 (O_151,N_2698,N_2082);
or UO_152 (O_152,N_2829,N_2746);
nand UO_153 (O_153,N_2841,N_2138);
nand UO_154 (O_154,N_2502,N_2864);
and UO_155 (O_155,N_2331,N_2239);
or UO_156 (O_156,N_2512,N_2927);
and UO_157 (O_157,N_2142,N_2495);
and UO_158 (O_158,N_2803,N_2308);
nor UO_159 (O_159,N_2650,N_2509);
or UO_160 (O_160,N_2491,N_2150);
and UO_161 (O_161,N_2106,N_2443);
and UO_162 (O_162,N_2938,N_2751);
nor UO_163 (O_163,N_2881,N_2642);
nor UO_164 (O_164,N_2077,N_2553);
nor UO_165 (O_165,N_2061,N_2962);
or UO_166 (O_166,N_2676,N_2951);
or UO_167 (O_167,N_2500,N_2050);
or UO_168 (O_168,N_2999,N_2236);
or UO_169 (O_169,N_2110,N_2484);
nor UO_170 (O_170,N_2399,N_2995);
and UO_171 (O_171,N_2628,N_2645);
or UO_172 (O_172,N_2595,N_2840);
nor UO_173 (O_173,N_2693,N_2071);
and UO_174 (O_174,N_2915,N_2813);
and UO_175 (O_175,N_2027,N_2718);
and UO_176 (O_176,N_2721,N_2241);
or UO_177 (O_177,N_2492,N_2330);
nand UO_178 (O_178,N_2506,N_2272);
or UO_179 (O_179,N_2401,N_2104);
nor UO_180 (O_180,N_2249,N_2246);
nor UO_181 (O_181,N_2462,N_2580);
nor UO_182 (O_182,N_2681,N_2340);
and UO_183 (O_183,N_2730,N_2383);
or UO_184 (O_184,N_2202,N_2621);
nor UO_185 (O_185,N_2807,N_2618);
and UO_186 (O_186,N_2969,N_2018);
nor UO_187 (O_187,N_2740,N_2563);
or UO_188 (O_188,N_2123,N_2006);
nor UO_189 (O_189,N_2095,N_2966);
or UO_190 (O_190,N_2414,N_2782);
or UO_191 (O_191,N_2254,N_2132);
or UO_192 (O_192,N_2556,N_2875);
nor UO_193 (O_193,N_2389,N_2592);
nand UO_194 (O_194,N_2685,N_2432);
and UO_195 (O_195,N_2371,N_2041);
and UO_196 (O_196,N_2364,N_2842);
or UO_197 (O_197,N_2859,N_2444);
nor UO_198 (O_198,N_2118,N_2262);
nor UO_199 (O_199,N_2518,N_2849);
nor UO_200 (O_200,N_2522,N_2532);
and UO_201 (O_201,N_2916,N_2614);
or UO_202 (O_202,N_2816,N_2682);
or UO_203 (O_203,N_2998,N_2457);
nand UO_204 (O_204,N_2059,N_2243);
nor UO_205 (O_205,N_2993,N_2790);
nand UO_206 (O_206,N_2304,N_2112);
nand UO_207 (O_207,N_2985,N_2791);
nand UO_208 (O_208,N_2005,N_2063);
nor UO_209 (O_209,N_2078,N_2573);
nor UO_210 (O_210,N_2887,N_2505);
nor UO_211 (O_211,N_2817,N_2184);
nand UO_212 (O_212,N_2854,N_2159);
or UO_213 (O_213,N_2452,N_2997);
or UO_214 (O_214,N_2666,N_2309);
and UO_215 (O_215,N_2919,N_2588);
or UO_216 (O_216,N_2477,N_2472);
nor UO_217 (O_217,N_2213,N_2418);
nor UO_218 (O_218,N_2200,N_2705);
or UO_219 (O_219,N_2758,N_2824);
nor UO_220 (O_220,N_2739,N_2012);
or UO_221 (O_221,N_2863,N_2054);
nor UO_222 (O_222,N_2348,N_2428);
nor UO_223 (O_223,N_2914,N_2933);
nand UO_224 (O_224,N_2269,N_2351);
and UO_225 (O_225,N_2369,N_2534);
nor UO_226 (O_226,N_2136,N_2228);
nor UO_227 (O_227,N_2778,N_2953);
or UO_228 (O_228,N_2385,N_2097);
nand UO_229 (O_229,N_2673,N_2386);
nor UO_230 (O_230,N_2093,N_2622);
or UO_231 (O_231,N_2121,N_2314);
or UO_232 (O_232,N_2017,N_2659);
nand UO_233 (O_233,N_2135,N_2485);
or UO_234 (O_234,N_2752,N_2053);
nor UO_235 (O_235,N_2270,N_2627);
nor UO_236 (O_236,N_2010,N_2533);
or UO_237 (O_237,N_2648,N_2507);
nand UO_238 (O_238,N_2143,N_2459);
or UO_239 (O_239,N_2707,N_2668);
or UO_240 (O_240,N_2448,N_2899);
nor UO_241 (O_241,N_2156,N_2148);
nand UO_242 (O_242,N_2735,N_2646);
or UO_243 (O_243,N_2898,N_2590);
and UO_244 (O_244,N_2494,N_2210);
nor UO_245 (O_245,N_2441,N_2602);
nor UO_246 (O_246,N_2780,N_2253);
or UO_247 (O_247,N_2035,N_2764);
or UO_248 (O_248,N_2271,N_2521);
nand UO_249 (O_249,N_2479,N_2812);
or UO_250 (O_250,N_2911,N_2991);
nor UO_251 (O_251,N_2410,N_2305);
and UO_252 (O_252,N_2989,N_2375);
and UO_253 (O_253,N_2163,N_2247);
and UO_254 (O_254,N_2815,N_2810);
or UO_255 (O_255,N_2667,N_2879);
nand UO_256 (O_256,N_2559,N_2530);
nor UO_257 (O_257,N_2749,N_2102);
and UO_258 (O_258,N_2251,N_2435);
nor UO_259 (O_259,N_2105,N_2792);
nand UO_260 (O_260,N_2689,N_2256);
or UO_261 (O_261,N_2728,N_2894);
or UO_262 (O_262,N_2708,N_2930);
nand UO_263 (O_263,N_2339,N_2663);
and UO_264 (O_264,N_2470,N_2540);
nor UO_265 (O_265,N_2821,N_2440);
or UO_266 (O_266,N_2260,N_2004);
nand UO_267 (O_267,N_2293,N_2126);
or UO_268 (O_268,N_2873,N_2240);
nor UO_269 (O_269,N_2358,N_2604);
or UO_270 (O_270,N_2311,N_2026);
or UO_271 (O_271,N_2398,N_2727);
nand UO_272 (O_272,N_2265,N_2334);
or UO_273 (O_273,N_2649,N_2343);
and UO_274 (O_274,N_2736,N_2290);
and UO_275 (O_275,N_2856,N_2766);
nand UO_276 (O_276,N_2750,N_2931);
nor UO_277 (O_277,N_2508,N_2565);
nor UO_278 (O_278,N_2793,N_2755);
nand UO_279 (O_279,N_2294,N_2939);
nor UO_280 (O_280,N_2327,N_2583);
nor UO_281 (O_281,N_2394,N_2949);
and UO_282 (O_282,N_2603,N_2720);
or UO_283 (O_283,N_2474,N_2332);
and UO_284 (O_284,N_2285,N_2560);
nor UO_285 (O_285,N_2800,N_2830);
and UO_286 (O_286,N_2357,N_2838);
or UO_287 (O_287,N_2064,N_2632);
nand UO_288 (O_288,N_2463,N_2851);
and UO_289 (O_289,N_2223,N_2421);
and UO_290 (O_290,N_2129,N_2355);
nor UO_291 (O_291,N_2295,N_2996);
and UO_292 (O_292,N_2328,N_2388);
nand UO_293 (O_293,N_2445,N_2372);
nand UO_294 (O_294,N_2335,N_2945);
nor UO_295 (O_295,N_2674,N_2429);
nor UO_296 (O_296,N_2834,N_2965);
nand UO_297 (O_297,N_2757,N_2697);
nor UO_298 (O_298,N_2225,N_2319);
and UO_299 (O_299,N_2582,N_2482);
nand UO_300 (O_300,N_2929,N_2634);
or UO_301 (O_301,N_2549,N_2716);
nand UO_302 (O_302,N_2536,N_2033);
and UO_303 (O_303,N_2317,N_2007);
nand UO_304 (O_304,N_2513,N_2124);
nand UO_305 (O_305,N_2354,N_2172);
nand UO_306 (O_306,N_2362,N_2827);
nand UO_307 (O_307,N_2768,N_2230);
nand UO_308 (O_308,N_2571,N_2378);
nand UO_309 (O_309,N_2141,N_2704);
nor UO_310 (O_310,N_2843,N_2242);
or UO_311 (O_311,N_2165,N_2099);
nand UO_312 (O_312,N_2043,N_2655);
or UO_313 (O_313,N_2877,N_2511);
nand UO_314 (O_314,N_2263,N_2320);
nand UO_315 (O_315,N_2640,N_2744);
nor UO_316 (O_316,N_2923,N_2120);
nand UO_317 (O_317,N_2932,N_2297);
nand UO_318 (O_318,N_2687,N_2888);
nand UO_319 (O_319,N_2423,N_2656);
and UO_320 (O_320,N_2313,N_2713);
or UO_321 (O_321,N_2671,N_2917);
nor UO_322 (O_322,N_2221,N_2905);
or UO_323 (O_323,N_2205,N_2818);
or UO_324 (O_324,N_2974,N_2970);
and UO_325 (O_325,N_2631,N_2267);
and UO_326 (O_326,N_2038,N_2675);
nor UO_327 (O_327,N_2638,N_2963);
or UO_328 (O_328,N_2688,N_2819);
or UO_329 (O_329,N_2281,N_2738);
and UO_330 (O_330,N_2504,N_2822);
nand UO_331 (O_331,N_2094,N_2643);
nand UO_332 (O_332,N_2454,N_2575);
and UO_333 (O_333,N_2637,N_2345);
nor UO_334 (O_334,N_2586,N_2893);
and UO_335 (O_335,N_2081,N_2572);
nor UO_336 (O_336,N_2218,N_2537);
and UO_337 (O_337,N_2367,N_2475);
or UO_338 (O_338,N_2743,N_2665);
or UO_339 (O_339,N_2890,N_2944);
or UO_340 (O_340,N_2934,N_2209);
and UO_341 (O_341,N_2558,N_2811);
nand UO_342 (O_342,N_2168,N_2203);
or UO_343 (O_343,N_2325,N_2359);
or UO_344 (O_344,N_2022,N_2175);
nand UO_345 (O_345,N_2733,N_2113);
xnor UO_346 (O_346,N_2913,N_2946);
and UO_347 (O_347,N_2347,N_2832);
nand UO_348 (O_348,N_2906,N_2576);
and UO_349 (O_349,N_2723,N_2562);
nor UO_350 (O_350,N_2561,N_2564);
nor UO_351 (O_351,N_2250,N_2706);
and UO_352 (O_352,N_2072,N_2608);
nand UO_353 (O_353,N_2579,N_2157);
nand UO_354 (O_354,N_2352,N_2227);
or UO_355 (O_355,N_2089,N_2234);
and UO_356 (O_356,N_2908,N_2023);
nor UO_357 (O_357,N_2192,N_2745);
or UO_358 (O_358,N_2356,N_2975);
or UO_359 (O_359,N_2447,N_2490);
xnor UO_360 (O_360,N_2434,N_2365);
or UO_361 (O_361,N_2956,N_2080);
and UO_362 (O_362,N_2060,N_2935);
or UO_363 (O_363,N_2224,N_2264);
nand UO_364 (O_364,N_2412,N_2942);
nand UO_365 (O_365,N_2499,N_2288);
nor UO_366 (O_366,N_2425,N_2882);
and UO_367 (O_367,N_2798,N_2695);
nor UO_368 (O_368,N_2710,N_2131);
and UO_369 (O_369,N_2154,N_2015);
nor UO_370 (O_370,N_2377,N_2981);
and UO_371 (O_371,N_2382,N_2431);
xnor UO_372 (O_372,N_2404,N_2407);
or UO_373 (O_373,N_2194,N_2591);
and UO_374 (O_374,N_2501,N_2976);
and UO_375 (O_375,N_2990,N_2569);
or UO_376 (O_376,N_2846,N_2526);
nand UO_377 (O_377,N_2892,N_2411);
and UO_378 (O_378,N_2855,N_2134);
nor UO_379 (O_379,N_2167,N_2889);
and UO_380 (O_380,N_2427,N_2610);
nor UO_381 (O_381,N_2029,N_2754);
nand UO_382 (O_382,N_2936,N_2413);
nor UO_383 (O_383,N_2153,N_2489);
nand UO_384 (O_384,N_2158,N_2907);
and UO_385 (O_385,N_2274,N_2273);
nand UO_386 (O_386,N_2108,N_2438);
nor UO_387 (O_387,N_2147,N_2926);
nand UO_388 (O_388,N_2858,N_2615);
or UO_389 (O_389,N_2598,N_2137);
and UO_390 (O_390,N_2419,N_2612);
or UO_391 (O_391,N_2420,N_2809);
or UO_392 (O_392,N_2145,N_2280);
nand UO_393 (O_393,N_2467,N_2761);
or UO_394 (O_394,N_2402,N_2363);
and UO_395 (O_395,N_2943,N_2114);
nor UO_396 (O_396,N_2069,N_2198);
and UO_397 (O_397,N_2971,N_2408);
or UO_398 (O_398,N_2395,N_2226);
and UO_399 (O_399,N_2469,N_2528);
or UO_400 (O_400,N_2122,N_2952);
or UO_401 (O_401,N_2779,N_2493);
nor UO_402 (O_402,N_2186,N_2664);
or UO_403 (O_403,N_2196,N_2346);
nand UO_404 (O_404,N_2487,N_2836);
nand UO_405 (O_405,N_2748,N_2872);
and UO_406 (O_406,N_2557,N_2978);
nand UO_407 (O_407,N_2955,N_2283);
nor UO_408 (O_408,N_2237,N_2287);
or UO_409 (O_409,N_2086,N_2051);
nor UO_410 (O_410,N_2878,N_2333);
nand UO_411 (O_411,N_2079,N_2214);
nand UO_412 (O_412,N_2222,N_2835);
and UO_413 (O_413,N_2045,N_2119);
nand UO_414 (O_414,N_2635,N_2437);
or UO_415 (O_415,N_2279,N_2786);
or UO_416 (O_416,N_2075,N_2286);
and UO_417 (O_417,N_2982,N_2773);
and UO_418 (O_418,N_2772,N_2669);
or UO_419 (O_419,N_2868,N_2483);
nand UO_420 (O_420,N_2455,N_2789);
and UO_421 (O_421,N_2361,N_2013);
and UO_422 (O_422,N_2424,N_2199);
nand UO_423 (O_423,N_2980,N_2880);
nor UO_424 (O_424,N_2284,N_2578);
nand UO_425 (O_425,N_2775,N_2639);
nor UO_426 (O_426,N_2520,N_2776);
or UO_427 (O_427,N_2605,N_2626);
or UO_428 (O_428,N_2904,N_2531);
nand UO_429 (O_429,N_2961,N_2219);
nand UO_430 (O_430,N_2542,N_2002);
nor UO_431 (O_431,N_2396,N_2034);
or UO_432 (O_432,N_2182,N_2066);
and UO_433 (O_433,N_2439,N_2307);
and UO_434 (O_434,N_2376,N_2616);
or UO_435 (O_435,N_2691,N_2699);
and UO_436 (O_436,N_2550,N_2217);
xor UO_437 (O_437,N_2031,N_2337);
or UO_438 (O_438,N_2278,N_2852);
or UO_439 (O_439,N_2861,N_2292);
and UO_440 (O_440,N_2466,N_2046);
nor UO_441 (O_441,N_2686,N_2876);
nand UO_442 (O_442,N_2040,N_2954);
or UO_443 (O_443,N_2047,N_2300);
nor UO_444 (O_444,N_2847,N_2839);
nor UO_445 (O_445,N_2070,N_2211);
nand UO_446 (O_446,N_2197,N_2947);
nor UO_447 (O_447,N_2076,N_2400);
or UO_448 (O_448,N_2672,N_2524);
nor UO_449 (O_449,N_2959,N_2344);
nand UO_450 (O_450,N_2180,N_2599);
nand UO_451 (O_451,N_2011,N_2928);
nand UO_452 (O_452,N_2446,N_2654);
nand UO_453 (O_453,N_2277,N_2216);
nor UO_454 (O_454,N_2096,N_2052);
or UO_455 (O_455,N_2866,N_2393);
nor UO_456 (O_456,N_2725,N_2338);
and UO_457 (O_457,N_2805,N_2703);
and UO_458 (O_458,N_2960,N_2623);
nand UO_459 (O_459,N_2215,N_2152);
nand UO_460 (O_460,N_2611,N_2024);
nor UO_461 (O_461,N_2541,N_2090);
and UO_462 (O_462,N_2282,N_2181);
nor UO_463 (O_463,N_2037,N_2717);
and UO_464 (O_464,N_2825,N_2994);
nor UO_465 (O_465,N_2554,N_2430);
nand UO_466 (O_466,N_2318,N_2607);
or UO_467 (O_467,N_2547,N_2116);
or UO_468 (O_468,N_2450,N_2456);
and UO_469 (O_469,N_2000,N_2206);
or UO_470 (O_470,N_2055,N_2275);
nand UO_471 (O_471,N_2900,N_2068);
nor UO_472 (O_472,N_2179,N_2149);
nor UO_473 (O_473,N_2515,N_2737);
or UO_474 (O_474,N_2808,N_2862);
or UO_475 (O_475,N_2336,N_2783);
nand UO_476 (O_476,N_2471,N_2259);
nor UO_477 (O_477,N_2625,N_2584);
and UO_478 (O_478,N_2177,N_2535);
and UO_479 (O_479,N_2416,N_2415);
nor UO_480 (O_480,N_2151,N_2771);
nand UO_481 (O_481,N_2302,N_2581);
or UO_482 (O_482,N_2785,N_2624);
nand UO_483 (O_483,N_2543,N_2897);
nor UO_484 (O_484,N_2189,N_2208);
and UO_485 (O_485,N_2677,N_2747);
nand UO_486 (O_486,N_2823,N_2409);
nor UO_487 (O_487,N_2127,N_2767);
or UO_488 (O_488,N_2984,N_2774);
nor UO_489 (O_489,N_2853,N_2067);
xnor UO_490 (O_490,N_2799,N_2370);
and UO_491 (O_491,N_2979,N_2312);
nand UO_492 (O_492,N_2957,N_2387);
or UO_493 (O_493,N_2871,N_2306);
nor UO_494 (O_494,N_2820,N_2019);
nor UO_495 (O_495,N_2644,N_2895);
or UO_496 (O_496,N_2503,N_2291);
and UO_497 (O_497,N_2722,N_2568);
or UO_498 (O_498,N_2756,N_2115);
and UO_499 (O_499,N_2594,N_2201);
endmodule