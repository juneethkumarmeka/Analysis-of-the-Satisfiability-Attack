module basic_1500_15000_2000_3_levels_10xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10002,N_10003,N_10004,N_10005,N_10006,N_10008,N_10010,N_10011,N_10013,N_10014,N_10015,N_10017,N_10018,N_10019,N_10020,N_10021,N_10023,N_10024,N_10025,N_10026,N_10027,N_10030,N_10031,N_10032,N_10033,N_10035,N_10036,N_10038,N_10039,N_10040,N_10041,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10053,N_10055,N_10057,N_10060,N_10061,N_10063,N_10064,N_10065,N_10066,N_10067,N_10069,N_10070,N_10071,N_10072,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10081,N_10083,N_10084,N_10085,N_10086,N_10088,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10115,N_10116,N_10117,N_10118,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10150,N_10152,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10171,N_10172,N_10175,N_10176,N_10179,N_10180,N_10181,N_10182,N_10183,N_10185,N_10186,N_10187,N_10188,N_10189,N_10193,N_10195,N_10196,N_10197,N_10198,N_10200,N_10201,N_10203,N_10204,N_10205,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10214,N_10216,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10238,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10249,N_10250,N_10251,N_10252,N_10253,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10319,N_10320,N_10321,N_10323,N_10325,N_10326,N_10327,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10354,N_10355,N_10357,N_10358,N_10359,N_10361,N_10362,N_10364,N_10365,N_10368,N_10369,N_10372,N_10373,N_10374,N_10376,N_10377,N_10378,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10393,N_10394,N_10395,N_10396,N_10397,N_10399,N_10401,N_10403,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10419,N_10420,N_10422,N_10423,N_10424,N_10425,N_10426,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10454,N_10455,N_10456,N_10457,N_10458,N_10460,N_10461,N_10462,N_10463,N_10464,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10473,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10484,N_10485,N_10486,N_10488,N_10489,N_10490,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10510,N_10511,N_10512,N_10513,N_10514,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10532,N_10533,N_10534,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10543,N_10544,N_10545,N_10547,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10564,N_10565,N_10567,N_10568,N_10569,N_10570,N_10571,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10581,N_10583,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10593,N_10594,N_10595,N_10596,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10629,N_10630,N_10631,N_10632,N_10634,N_10635,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10652,N_10653,N_10655,N_10656,N_10657,N_10658,N_10659,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10681,N_10682,N_10685,N_10686,N_10688,N_10690,N_10692,N_10693,N_10694,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10715,N_10717,N_10718,N_10719,N_10721,N_10723,N_10724,N_10725,N_10727,N_10728,N_10729,N_10730,N_10731,N_10733,N_10735,N_10736,N_10739,N_10740,N_10743,N_10744,N_10745,N_10747,N_10748,N_10749,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10759,N_10762,N_10763,N_10764,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10776,N_10777,N_10778,N_10779,N_10780,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10806,N_10807,N_10808,N_10809,N_10811,N_10812,N_10813,N_10814,N_10816,N_10818,N_10819,N_10820,N_10821,N_10823,N_10824,N_10825,N_10826,N_10828,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10873,N_10874,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10884,N_10885,N_10887,N_10889,N_10890,N_10891,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10908,N_10909,N_10911,N_10912,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10924,N_10925,N_10926,N_10928,N_10929,N_10931,N_10932,N_10933,N_10934,N_10936,N_10937,N_10938,N_10939,N_10941,N_10942,N_10943,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11003,N_11004,N_11005,N_11006,N_11007,N_11009,N_11010,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11024,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11034,N_11035,N_11036,N_11037,N_11038,N_11042,N_11043,N_11044,N_11045,N_11046,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11062,N_11063,N_11064,N_11065,N_11067,N_11068,N_11070,N_11071,N_11072,N_11074,N_11075,N_11078,N_11079,N_11082,N_11084,N_11085,N_11087,N_11088,N_11089,N_11091,N_11092,N_11093,N_11094,N_11097,N_11098,N_11099,N_11100,N_11102,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11113,N_11114,N_11116,N_11117,N_11118,N_11119,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11128,N_11129,N_11131,N_11133,N_11134,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11143,N_11144,N_11147,N_11148,N_11151,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11164,N_11165,N_11166,N_11168,N_11170,N_11171,N_11173,N_11174,N_11175,N_11176,N_11177,N_11179,N_11180,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11189,N_11190,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11252,N_11253,N_11254,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11270,N_11271,N_11273,N_11275,N_11276,N_11277,N_11281,N_11283,N_11284,N_11285,N_11286,N_11287,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11301,N_11302,N_11303,N_11305,N_11306,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11324,N_11325,N_11326,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11348,N_11350,N_11353,N_11354,N_11355,N_11356,N_11358,N_11359,N_11362,N_11363,N_11365,N_11366,N_11368,N_11369,N_11370,N_11371,N_11373,N_11374,N_11376,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11389,N_11391,N_11392,N_11393,N_11396,N_11397,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11416,N_11417,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11438,N_11439,N_11441,N_11442,N_11443,N_11445,N_11446,N_11447,N_11448,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11476,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11511,N_11512,N_11513,N_11514,N_11516,N_11517,N_11518,N_11519,N_11522,N_11523,N_11524,N_11527,N_11529,N_11530,N_11531,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11540,N_11541,N_11542,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11555,N_11557,N_11558,N_11559,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11569,N_11570,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11605,N_11606,N_11608,N_11609,N_11610,N_11611,N_11613,N_11614,N_11615,N_11616,N_11617,N_11619,N_11620,N_11621,N_11622,N_11623,N_11626,N_11627,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11636,N_11637,N_11638,N_11640,N_11641,N_11642,N_11643,N_11646,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11668,N_11669,N_11670,N_11672,N_11673,N_11675,N_11676,N_11677,N_11678,N_11679,N_11681,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11696,N_11697,N_11698,N_11700,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11717,N_11718,N_11719,N_11720,N_11721,N_11723,N_11725,N_11726,N_11728,N_11729,N_11730,N_11731,N_11732,N_11734,N_11736,N_11737,N_11738,N_11740,N_11741,N_11742,N_11743,N_11745,N_11746,N_11747,N_11749,N_11750,N_11752,N_11753,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11765,N_11766,N_11767,N_11768,N_11770,N_11772,N_11773,N_11774,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11794,N_11795,N_11796,N_11797,N_11798,N_11800,N_11801,N_11802,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11816,N_11817,N_11818,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11829,N_11830,N_11831,N_11832,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11844,N_11845,N_11846,N_11847,N_11848,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11878,N_11879,N_11880,N_11881,N_11882,N_11885,N_11886,N_11887,N_11888,N_11889,N_11894,N_11895,N_11896,N_11897,N_11899,N_11900,N_11901,N_11902,N_11903,N_11905,N_11906,N_11907,N_11908,N_11909,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11929,N_11930,N_11933,N_11934,N_11935,N_11936,N_11937,N_11940,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11952,N_11953,N_11954,N_11955,N_11958,N_11959,N_11961,N_11962,N_11963,N_11965,N_11966,N_11967,N_11970,N_11971,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11982,N_11983,N_11984,N_11985,N_11987,N_11988,N_11989,N_11990,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12001,N_12002,N_12003,N_12004,N_12005,N_12007,N_12008,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12019,N_12020,N_12021,N_12022,N_12024,N_12025,N_12026,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12045,N_12046,N_12047,N_12049,N_12050,N_12051,N_12052,N_12054,N_12056,N_12057,N_12058,N_12060,N_12061,N_12063,N_12064,N_12065,N_12066,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12078,N_12079,N_12080,N_12081,N_12082,N_12084,N_12085,N_12086,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12104,N_12105,N_12106,N_12107,N_12109,N_12111,N_12112,N_12113,N_12114,N_12115,N_12117,N_12119,N_12120,N_12122,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12132,N_12133,N_12134,N_12136,N_12138,N_12141,N_12142,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12179,N_12181,N_12182,N_12185,N_12186,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12201,N_12203,N_12204,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12227,N_12228,N_12229,N_12232,N_12233,N_12234,N_12235,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12244,N_12245,N_12246,N_12248,N_12249,N_12251,N_12252,N_12254,N_12255,N_12256,N_12258,N_12259,N_12260,N_12261,N_12263,N_12264,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12287,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12306,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12361,N_12362,N_12363,N_12365,N_12366,N_12367,N_12368,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12377,N_12378,N_12381,N_12383,N_12384,N_12385,N_12387,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12413,N_12415,N_12416,N_12417,N_12419,N_12420,N_12421,N_12422,N_12424,N_12425,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12457,N_12458,N_12460,N_12462,N_12464,N_12465,N_12466,N_12467,N_12468,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12486,N_12488,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12500,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12553,N_12554,N_12557,N_12559,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12580,N_12581,N_12582,N_12583,N_12584,N_12586,N_12587,N_12588,N_12590,N_12591,N_12592,N_12594,N_12595,N_12596,N_12597,N_12598,N_12600,N_12601,N_12602,N_12604,N_12605,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12624,N_12625,N_12626,N_12627,N_12628,N_12630,N_12631,N_12633,N_12634,N_12635,N_12637,N_12638,N_12640,N_12641,N_12642,N_12643,N_12645,N_12648,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12658,N_12660,N_12661,N_12663,N_12664,N_12665,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12684,N_12685,N_12689,N_12690,N_12691,N_12692,N_12694,N_12695,N_12698,N_12700,N_12701,N_12702,N_12703,N_12706,N_12708,N_12709,N_12710,N_12711,N_12713,N_12714,N_12715,N_12717,N_12720,N_12721,N_12723,N_12724,N_12725,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12746,N_12747,N_12748,N_12750,N_12751,N_12752,N_12754,N_12755,N_12756,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12766,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12779,N_12780,N_12781,N_12783,N_12784,N_12785,N_12786,N_12787,N_12789,N_12792,N_12794,N_12796,N_12797,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12809,N_12810,N_12812,N_12814,N_12817,N_12818,N_12819,N_12820,N_12822,N_12823,N_12824,N_12825,N_12826,N_12828,N_12829,N_12830,N_12831,N_12832,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12862,N_12863,N_12864,N_12866,N_12867,N_12868,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12897,N_12898,N_12899,N_12901,N_12902,N_12905,N_12906,N_12908,N_12909,N_12911,N_12913,N_12915,N_12916,N_12918,N_12919,N_12921,N_12923,N_12924,N_12925,N_12926,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12980,N_12981,N_12982,N_12983,N_12984,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12996,N_12998,N_12999,N_13000,N_13001,N_13002,N_13004,N_13005,N_13006,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13021,N_13022,N_13025,N_13026,N_13027,N_13029,N_13030,N_13031,N_13033,N_13034,N_13035,N_13036,N_13037,N_13039,N_13040,N_13041,N_13043,N_13045,N_13046,N_13047,N_13048,N_13049,N_13051,N_13052,N_13053,N_13056,N_13057,N_13058,N_13059,N_13060,N_13062,N_13063,N_13064,N_13065,N_13066,N_13068,N_13069,N_13070,N_13071,N_13073,N_13074,N_13076,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13085,N_13086,N_13087,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13099,N_13100,N_13101,N_13103,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13125,N_13126,N_13128,N_13130,N_13131,N_13132,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13144,N_13145,N_13146,N_13147,N_13149,N_13150,N_13151,N_13152,N_13154,N_13155,N_13156,N_13157,N_13158,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13169,N_13171,N_13172,N_13174,N_13176,N_13177,N_13178,N_13179,N_13180,N_13182,N_13183,N_13185,N_13186,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13204,N_13205,N_13206,N_13208,N_13210,N_13211,N_13212,N_13215,N_13216,N_13217,N_13220,N_13221,N_13223,N_13224,N_13225,N_13226,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13238,N_13239,N_13241,N_13242,N_13243,N_13244,N_13245,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13264,N_13265,N_13266,N_13267,N_13269,N_13270,N_13271,N_13272,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13283,N_13284,N_13285,N_13286,N_13287,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13312,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13323,N_13325,N_13326,N_13327,N_13328,N_13331,N_13332,N_13333,N_13334,N_13336,N_13337,N_13338,N_13339,N_13342,N_13343,N_13344,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13375,N_13376,N_13377,N_13378,N_13379,N_13381,N_13382,N_13384,N_13385,N_13387,N_13388,N_13389,N_13390,N_13392,N_13393,N_13394,N_13396,N_13397,N_13398,N_13399,N_13400,N_13402,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13411,N_13412,N_13413,N_13414,N_13417,N_13419,N_13420,N_13421,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13433,N_13434,N_13435,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13452,N_13454,N_13455,N_13457,N_13460,N_13463,N_13464,N_13466,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13503,N_13504,N_13505,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13534,N_13535,N_13536,N_13537,N_13538,N_13542,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13561,N_13563,N_13564,N_13566,N_13567,N_13569,N_13570,N_13571,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13604,N_13606,N_13609,N_13611,N_13612,N_13613,N_13615,N_13616,N_13617,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13638,N_13639,N_13640,N_13641,N_13643,N_13646,N_13647,N_13648,N_13649,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13663,N_13665,N_13666,N_13667,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13689,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13699,N_13700,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13710,N_13711,N_13712,N_13713,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13736,N_13737,N_13739,N_13740,N_13743,N_13744,N_13745,N_13747,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13827,N_13828,N_13829,N_13830,N_13831,N_13833,N_13835,N_13836,N_13837,N_13838,N_13839,N_13841,N_13843,N_13844,N_13846,N_13847,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13867,N_13868,N_13869,N_13870,N_13871,N_13873,N_13874,N_13875,N_13877,N_13879,N_13880,N_13881,N_13882,N_13883,N_13885,N_13887,N_13888,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13901,N_13902,N_13903,N_13904,N_13906,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13919,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13931,N_13932,N_13934,N_13935,N_13936,N_13938,N_13939,N_13943,N_13944,N_13947,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13959,N_13960,N_13961,N_13962,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13971,N_13974,N_13975,N_13976,N_13977,N_13978,N_13980,N_13981,N_13983,N_13984,N_13986,N_13987,N_13988,N_13989,N_13990,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14003,N_14004,N_14005,N_14010,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14022,N_14024,N_14026,N_14027,N_14028,N_14029,N_14030,N_14032,N_14033,N_14034,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14046,N_14047,N_14049,N_14051,N_14052,N_14053,N_14054,N_14056,N_14057,N_14058,N_14059,N_14060,N_14062,N_14065,N_14066,N_14067,N_14068,N_14070,N_14072,N_14073,N_14074,N_14076,N_14077,N_14079,N_14081,N_14083,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14103,N_14104,N_14107,N_14108,N_14109,N_14110,N_14112,N_14113,N_14114,N_14115,N_14117,N_14118,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14146,N_14147,N_14148,N_14149,N_14150,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14160,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14182,N_14183,N_14184,N_14186,N_14187,N_14190,N_14191,N_14192,N_14194,N_14195,N_14197,N_14198,N_14199,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14209,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14218,N_14219,N_14221,N_14222,N_14223,N_14224,N_14227,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14247,N_14248,N_14250,N_14251,N_14252,N_14253,N_14255,N_14256,N_14257,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14271,N_14272,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14294,N_14295,N_14297,N_14298,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14319,N_14320,N_14321,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14335,N_14336,N_14337,N_14339,N_14341,N_14343,N_14344,N_14345,N_14347,N_14348,N_14349,N_14351,N_14352,N_14354,N_14355,N_14356,N_14357,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14371,N_14374,N_14375,N_14376,N_14378,N_14379,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14388,N_14389,N_14390,N_14391,N_14392,N_14395,N_14396,N_14398,N_14403,N_14404,N_14405,N_14406,N_14408,N_14414,N_14417,N_14418,N_14419,N_14420,N_14421,N_14423,N_14424,N_14425,N_14426,N_14427,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14441,N_14442,N_14443,N_14444,N_14446,N_14448,N_14449,N_14450,N_14451,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14478,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14489,N_14492,N_14494,N_14495,N_14496,N_14497,N_14500,N_14501,N_14502,N_14503,N_14504,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14514,N_14515,N_14516,N_14517,N_14518,N_14520,N_14522,N_14523,N_14524,N_14525,N_14526,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14546,N_14547,N_14548,N_14550,N_14553,N_14554,N_14555,N_14557,N_14560,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14569,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14581,N_14582,N_14584,N_14585,N_14586,N_14587,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14597,N_14598,N_14599,N_14600,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14610,N_14611,N_14612,N_14613,N_14615,N_14616,N_14617,N_14618,N_14619,N_14621,N_14622,N_14623,N_14624,N_14626,N_14628,N_14629,N_14631,N_14632,N_14633,N_14634,N_14635,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14644,N_14646,N_14647,N_14649,N_14650,N_14651,N_14652,N_14653,N_14656,N_14657,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14674,N_14675,N_14676,N_14678,N_14679,N_14682,N_14683,N_14684,N_14685,N_14686,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14700,N_14701,N_14703,N_14705,N_14706,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14715,N_14716,N_14717,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14727,N_14728,N_14730,N_14731,N_14732,N_14733,N_14735,N_14736,N_14737,N_14740,N_14741,N_14742,N_14743,N_14745,N_14746,N_14747,N_14749,N_14750,N_14751,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14765,N_14766,N_14767,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14791,N_14793,N_14794,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14814,N_14815,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14825,N_14826,N_14827,N_14828,N_14831,N_14832,N_14833,N_14835,N_14836,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14850,N_14851,N_14852,N_14855,N_14856,N_14857,N_14860,N_14861,N_14862,N_14863,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14876,N_14879,N_14880,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14891,N_14892,N_14893,N_14894,N_14895,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14913,N_14914,N_14915,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14924,N_14925,N_14926,N_14927,N_14928,N_14930,N_14931,N_14932,N_14933,N_14934,N_14936,N_14937,N_14938,N_14940,N_14942,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14994,N_14995,N_14996,N_14999;
nor U0 (N_0,In_301,In_312);
or U1 (N_1,In_1368,In_378);
xor U2 (N_2,In_1325,In_1477);
nand U3 (N_3,In_950,In_1085);
xor U4 (N_4,In_201,In_894);
or U5 (N_5,In_387,In_124);
nand U6 (N_6,In_725,In_715);
nor U7 (N_7,In_1250,In_1416);
nor U8 (N_8,In_411,In_15);
nor U9 (N_9,In_795,In_654);
nor U10 (N_10,In_41,In_1392);
nand U11 (N_11,In_473,In_1);
nor U12 (N_12,In_1478,In_838);
or U13 (N_13,In_860,In_911);
xor U14 (N_14,In_1297,In_1256);
nand U15 (N_15,In_585,In_937);
nand U16 (N_16,In_204,In_8);
nor U17 (N_17,In_1048,In_1291);
xnor U18 (N_18,In_766,In_568);
and U19 (N_19,In_804,In_452);
nand U20 (N_20,In_606,In_44);
xnor U21 (N_21,In_1424,In_1058);
or U22 (N_22,In_1492,In_683);
xnor U23 (N_23,In_589,In_70);
xor U24 (N_24,In_1307,In_418);
nand U25 (N_25,In_861,In_135);
xor U26 (N_26,In_601,In_668);
nor U27 (N_27,In_495,In_408);
xnor U28 (N_28,In_644,In_1480);
nand U29 (N_29,In_233,In_770);
or U30 (N_30,In_366,In_1181);
and U31 (N_31,In_256,In_599);
or U32 (N_32,In_363,In_690);
nand U33 (N_33,In_496,In_1482);
nand U34 (N_34,In_1022,In_40);
nand U35 (N_35,In_323,In_518);
or U36 (N_36,In_1269,In_882);
xor U37 (N_37,In_430,In_271);
nand U38 (N_38,In_346,In_531);
and U39 (N_39,In_1199,In_1225);
nor U40 (N_40,In_564,In_1407);
xor U41 (N_41,In_1105,In_587);
or U42 (N_42,In_805,In_611);
xor U43 (N_43,In_629,In_358);
xnor U44 (N_44,In_1244,In_855);
or U45 (N_45,In_429,In_602);
nand U46 (N_46,In_1342,In_143);
or U47 (N_47,In_272,In_171);
and U48 (N_48,In_1361,In_862);
or U49 (N_49,In_491,In_685);
nor U50 (N_50,In_153,In_1292);
and U51 (N_51,In_845,In_537);
and U52 (N_52,In_1205,In_1403);
or U53 (N_53,In_431,In_1345);
xor U54 (N_54,In_994,In_1108);
nand U55 (N_55,In_1163,In_873);
nand U56 (N_56,In_1087,In_1193);
nand U57 (N_57,In_836,In_1444);
xnor U58 (N_58,In_438,In_1024);
nor U59 (N_59,In_130,In_659);
xnor U60 (N_60,In_933,In_0);
nand U61 (N_61,In_675,In_1071);
or U62 (N_62,In_425,In_54);
or U63 (N_63,In_243,In_317);
and U64 (N_64,In_95,In_1235);
and U65 (N_65,In_1341,In_1204);
nor U66 (N_66,In_575,In_907);
and U67 (N_67,In_1122,In_405);
xor U68 (N_68,In_539,In_931);
and U69 (N_69,In_1270,In_981);
xnor U70 (N_70,In_901,In_1401);
and U71 (N_71,In_940,In_370);
nand U72 (N_72,In_1386,In_511);
or U73 (N_73,In_517,In_1165);
and U74 (N_74,In_225,In_1317);
or U75 (N_75,In_79,In_109);
xnor U76 (N_76,In_580,In_864);
xor U77 (N_77,In_923,In_414);
nand U78 (N_78,In_749,In_549);
nand U79 (N_79,In_485,In_1430);
or U80 (N_80,In_906,In_817);
and U81 (N_81,In_276,In_247);
and U82 (N_82,In_979,In_1343);
xnor U83 (N_83,In_1406,In_434);
nor U84 (N_84,In_141,In_157);
nand U85 (N_85,In_277,In_784);
nand U86 (N_86,In_635,In_971);
xnor U87 (N_87,In_1035,In_1174);
or U88 (N_88,In_710,In_532);
xnor U89 (N_89,In_1428,In_1083);
nand U90 (N_90,In_780,In_691);
xor U91 (N_91,In_454,In_605);
nand U92 (N_92,In_581,In_1383);
or U93 (N_93,In_577,In_1027);
xor U94 (N_94,In_23,In_169);
or U95 (N_95,In_1064,In_188);
or U96 (N_96,In_791,In_748);
xor U97 (N_97,In_946,In_392);
xnor U98 (N_98,In_724,In_953);
and U99 (N_99,In_1337,In_758);
nor U100 (N_100,In_1151,In_910);
or U101 (N_101,In_1272,In_1121);
nor U102 (N_102,In_85,In_379);
nor U103 (N_103,In_355,In_240);
and U104 (N_104,In_959,In_353);
and U105 (N_105,In_754,In_1218);
xnor U106 (N_106,In_1037,In_324);
nand U107 (N_107,In_622,In_973);
nor U108 (N_108,In_961,In_643);
nor U109 (N_109,In_50,In_853);
or U110 (N_110,In_1190,In_1426);
and U111 (N_111,In_995,In_1240);
nand U112 (N_112,In_936,In_819);
nor U113 (N_113,In_42,In_1373);
or U114 (N_114,In_1398,In_990);
nand U115 (N_115,In_273,In_949);
nor U116 (N_116,In_1491,In_789);
and U117 (N_117,In_929,In_627);
or U118 (N_118,In_71,In_1143);
nand U119 (N_119,In_206,In_1023);
and U120 (N_120,In_499,In_1200);
or U121 (N_121,In_311,In_787);
or U122 (N_122,In_35,In_829);
and U123 (N_123,In_1068,In_958);
nand U124 (N_124,In_648,In_1470);
nor U125 (N_125,In_1391,In_360);
nor U126 (N_126,In_1147,In_1276);
nand U127 (N_127,In_94,In_132);
or U128 (N_128,In_470,In_249);
nor U129 (N_129,In_1034,In_1113);
nor U130 (N_130,In_802,In_1496);
nand U131 (N_131,In_129,In_1212);
xnor U132 (N_132,In_1326,In_1446);
and U133 (N_133,In_964,In_1054);
and U134 (N_134,In_730,In_1006);
and U135 (N_135,In_679,In_560);
nor U136 (N_136,In_352,In_55);
and U137 (N_137,In_615,In_872);
nand U138 (N_138,In_123,In_297);
or U139 (N_139,In_11,In_737);
and U140 (N_140,In_614,In_1473);
nand U141 (N_141,In_1031,In_835);
and U142 (N_142,In_242,In_1155);
and U143 (N_143,In_1374,In_992);
nand U144 (N_144,In_680,In_6);
and U145 (N_145,In_1384,In_788);
nand U146 (N_146,In_306,In_1241);
nor U147 (N_147,In_404,In_180);
and U148 (N_148,In_515,In_925);
or U149 (N_149,In_672,In_451);
and U150 (N_150,In_1211,In_179);
xnor U151 (N_151,In_351,In_800);
and U152 (N_152,In_1456,In_1298);
and U153 (N_153,In_843,In_856);
nor U154 (N_154,In_650,In_919);
or U155 (N_155,In_419,In_86);
nand U156 (N_156,In_76,In_1397);
xor U157 (N_157,In_701,In_117);
nor U158 (N_158,In_818,In_290);
or U159 (N_159,In_883,In_479);
xor U160 (N_160,In_367,In_1172);
and U161 (N_161,In_497,In_167);
nor U162 (N_162,In_729,In_87);
and U163 (N_163,In_91,In_384);
and U164 (N_164,In_1041,In_337);
or U165 (N_165,In_93,In_1295);
nor U166 (N_166,In_1260,In_420);
nand U167 (N_167,In_455,In_1176);
nor U168 (N_168,In_1045,In_1251);
and U169 (N_169,In_228,In_52);
xor U170 (N_170,In_716,In_1277);
xor U171 (N_171,In_33,In_956);
xnor U172 (N_172,In_1339,In_1351);
nand U173 (N_173,In_695,In_1310);
nand U174 (N_174,In_274,In_174);
xor U175 (N_175,In_380,In_612);
and U176 (N_176,In_1100,In_1187);
and U177 (N_177,In_707,In_877);
xnor U178 (N_178,In_904,In_1372);
nor U179 (N_179,In_1033,In_1153);
nand U180 (N_180,In_1171,In_583);
xor U181 (N_181,In_1154,In_1452);
and U182 (N_182,In_376,In_483);
nor U183 (N_183,In_1168,In_199);
xor U184 (N_184,In_579,In_968);
nand U185 (N_185,In_742,In_196);
nand U186 (N_186,In_390,In_1380);
xor U187 (N_187,In_756,In_874);
and U188 (N_188,In_53,In_723);
and U189 (N_189,In_1110,In_726);
nor U190 (N_190,In_1040,In_1135);
or U191 (N_191,In_28,In_1405);
xnor U192 (N_192,In_345,In_1381);
and U193 (N_193,In_281,In_745);
xnor U194 (N_194,In_183,In_636);
and U195 (N_195,In_69,In_56);
or U196 (N_196,In_238,In_667);
xnor U197 (N_197,In_1166,In_1050);
xor U198 (N_198,In_712,In_542);
and U199 (N_199,In_484,In_458);
nor U200 (N_200,In_439,In_676);
xnor U201 (N_201,In_572,In_1081);
nor U202 (N_202,In_1278,In_762);
and U203 (N_203,In_1042,In_996);
xnor U204 (N_204,In_757,In_212);
nor U205 (N_205,In_251,In_170);
xor U206 (N_206,In_61,In_565);
and U207 (N_207,In_1059,In_626);
nand U208 (N_208,In_653,In_806);
nor U209 (N_209,In_475,In_1436);
and U210 (N_210,In_464,In_932);
and U211 (N_211,In_507,In_21);
and U212 (N_212,In_768,In_796);
nor U213 (N_213,In_1078,In_467);
and U214 (N_214,In_1495,In_1335);
xor U215 (N_215,In_1371,In_1215);
nor U216 (N_216,In_781,In_3);
nand U217 (N_217,In_808,In_498);
or U218 (N_218,In_12,In_1002);
or U219 (N_219,In_226,In_381);
and U220 (N_220,In_1088,In_1097);
xor U221 (N_221,In_1161,In_785);
or U222 (N_222,In_423,In_852);
and U223 (N_223,In_661,In_538);
nand U224 (N_224,In_330,In_1464);
or U225 (N_225,In_239,In_1318);
or U226 (N_226,In_1125,In_375);
and U227 (N_227,In_164,In_377);
nand U228 (N_228,In_908,In_1104);
or U229 (N_229,In_651,In_190);
nor U230 (N_230,In_930,In_283);
or U231 (N_231,In_1420,In_698);
nand U232 (N_232,In_1055,In_590);
xnor U233 (N_233,In_1453,In_435);
nor U234 (N_234,In_669,In_39);
nand U235 (N_235,In_1152,In_1167);
xnor U236 (N_236,In_826,In_104);
or U237 (N_237,In_89,In_368);
nor U238 (N_238,In_417,In_1228);
nand U239 (N_239,In_871,In_177);
or U240 (N_240,In_1312,In_1399);
xor U241 (N_241,In_986,In_192);
xnor U242 (N_242,In_825,In_131);
and U243 (N_243,In_105,In_1356);
xnor U244 (N_244,In_1237,In_771);
nand U245 (N_245,In_1017,In_286);
and U246 (N_246,In_1474,In_1112);
nor U247 (N_247,In_948,In_461);
nand U248 (N_248,In_533,In_628);
xor U249 (N_249,In_1299,In_1001);
nand U250 (N_250,In_786,In_1304);
and U251 (N_251,In_149,In_915);
and U252 (N_252,In_254,In_1029);
nor U253 (N_253,In_284,In_342);
xnor U254 (N_254,In_714,In_513);
xnor U255 (N_255,In_547,In_975);
nor U256 (N_256,In_255,In_999);
xor U257 (N_257,In_176,In_1283);
xnor U258 (N_258,In_219,In_588);
or U259 (N_259,In_1447,In_1425);
or U260 (N_260,In_1130,In_673);
xnor U261 (N_261,In_450,In_943);
xor U262 (N_262,In_1289,In_1092);
and U263 (N_263,In_744,In_407);
xor U264 (N_264,In_1046,In_101);
nor U265 (N_265,In_529,In_1210);
and U266 (N_266,In_584,In_751);
or U267 (N_267,In_445,In_998);
or U268 (N_268,In_993,In_798);
nor U269 (N_269,In_58,In_300);
and U270 (N_270,In_942,In_116);
or U271 (N_271,In_1202,In_294);
xor U272 (N_272,In_389,In_316);
and U273 (N_273,In_245,In_1208);
or U274 (N_274,In_369,In_1094);
and U275 (N_275,In_630,In_1493);
xor U276 (N_276,In_236,In_893);
nor U277 (N_277,In_250,In_598);
nand U278 (N_278,In_159,In_1093);
nand U279 (N_279,In_1049,In_66);
or U280 (N_280,In_1460,In_98);
nor U281 (N_281,In_618,In_684);
xor U282 (N_282,In_1475,In_1305);
nor U283 (N_283,In_974,In_733);
nor U284 (N_284,In_1259,In_1004);
xnor U285 (N_285,In_1221,In_112);
nand U286 (N_286,In_1109,In_115);
or U287 (N_287,In_1432,In_1330);
nand U288 (N_288,In_508,In_540);
or U289 (N_289,In_81,In_374);
xnor U290 (N_290,In_734,In_1141);
nand U291 (N_291,In_1149,In_952);
xnor U292 (N_292,In_1129,In_332);
and U293 (N_293,In_821,In_444);
or U294 (N_294,In_1077,In_700);
xnor U295 (N_295,In_147,In_1349);
nand U296 (N_296,In_1288,In_761);
or U297 (N_297,In_99,In_7);
nor U298 (N_298,In_74,In_570);
or U299 (N_299,In_260,In_1003);
nor U300 (N_300,In_456,In_1451);
or U301 (N_301,In_708,In_1411);
xor U302 (N_302,In_945,In_970);
and U303 (N_303,In_664,In_361);
and U304 (N_304,In_1179,In_72);
nand U305 (N_305,In_448,In_519);
or U306 (N_306,In_82,In_1198);
nor U307 (N_307,In_1137,In_1025);
nand U308 (N_308,In_501,In_402);
xnor U309 (N_309,In_65,In_645);
xnor U310 (N_310,In_400,In_1316);
and U311 (N_311,In_1309,In_834);
nor U312 (N_312,In_4,In_1255);
xnor U313 (N_313,In_962,In_1306);
or U314 (N_314,In_111,In_526);
nand U315 (N_315,In_1136,In_866);
and U316 (N_316,In_898,In_678);
xnor U317 (N_317,In_759,In_727);
xnor U318 (N_318,In_1146,In_1095);
xor U319 (N_319,In_1178,In_857);
xor U320 (N_320,In_899,In_1115);
xnor U321 (N_321,In_1102,In_1346);
nand U322 (N_322,In_299,In_298);
xnor U323 (N_323,In_84,In_134);
xor U324 (N_324,In_574,In_1497);
xnor U325 (N_325,In_399,In_1131);
nand U326 (N_326,In_1385,In_1323);
nand U327 (N_327,In_75,In_1026);
or U328 (N_328,In_1072,In_1489);
xnor U329 (N_329,In_1281,In_1140);
xor U330 (N_330,In_902,In_118);
nor U331 (N_331,In_1375,In_334);
nor U332 (N_332,In_24,In_362);
nor U333 (N_333,In_1160,In_1329);
or U334 (N_334,In_935,In_34);
and U335 (N_335,In_1051,In_220);
and U336 (N_336,In_32,In_1123);
xor U337 (N_337,In_763,In_1030);
or U338 (N_338,In_282,In_980);
xnor U339 (N_339,In_1360,In_1261);
xor U340 (N_340,In_310,In_987);
xnor U341 (N_341,In_903,In_476);
and U342 (N_342,In_868,In_248);
nand U343 (N_343,In_582,In_2);
nand U344 (N_344,In_382,In_1457);
or U345 (N_345,In_1127,In_1472);
or U346 (N_346,In_1286,In_349);
and U347 (N_347,In_280,In_1271);
nand U348 (N_348,In_1454,In_918);
xor U349 (N_349,In_1038,In_815);
and U350 (N_350,In_343,In_891);
and U351 (N_351,In_63,In_1359);
nor U352 (N_352,In_632,In_1364);
or U353 (N_353,In_1435,In_1173);
or U354 (N_354,In_1099,In_851);
nand U355 (N_355,In_230,In_421);
and U356 (N_356,In_215,In_1175);
and U357 (N_357,In_29,In_128);
or U358 (N_358,In_794,In_793);
and U359 (N_359,In_988,In_554);
nor U360 (N_360,In_1427,In_1379);
or U361 (N_361,In_1128,In_881);
or U362 (N_362,In_1015,In_1053);
xor U363 (N_363,In_1438,In_594);
nor U364 (N_364,In_774,In_728);
nand U365 (N_365,In_1084,In_1018);
and U366 (N_366,In_198,In_1485);
xnor U367 (N_367,In_1431,In_173);
xnor U368 (N_368,In_184,In_223);
or U369 (N_369,In_5,In_45);
nor U370 (N_370,In_321,In_150);
xor U371 (N_371,In_658,In_704);
nor U372 (N_372,In_1465,In_500);
xnor U373 (N_373,In_711,In_963);
xnor U374 (N_374,In_1043,In_846);
nand U375 (N_375,In_217,In_889);
xor U376 (N_376,In_489,In_603);
nor U377 (N_377,In_820,In_760);
nand U378 (N_378,In_152,In_1180);
or U379 (N_379,In_333,In_1409);
and U380 (N_380,In_1363,In_912);
or U381 (N_381,In_315,In_709);
and U382 (N_382,In_1086,In_463);
or U383 (N_383,In_985,In_764);
nand U384 (N_384,In_638,In_205);
nor U385 (N_385,In_9,In_849);
nand U386 (N_386,In_263,In_1219);
xor U387 (N_387,In_1367,In_1182);
nor U388 (N_388,In_457,In_465);
and U389 (N_389,In_279,In_858);
and U390 (N_390,In_488,In_469);
and U391 (N_391,In_520,In_722);
nand U392 (N_392,In_1194,In_859);
nand U393 (N_393,In_341,In_1134);
xor U394 (N_394,In_307,In_1148);
nand U395 (N_395,In_832,In_1120);
and U396 (N_396,In_1340,In_1468);
nand U397 (N_397,In_401,In_1209);
nor U398 (N_398,In_625,In_790);
nand U399 (N_399,In_516,In_113);
and U400 (N_400,In_126,In_1213);
nor U401 (N_401,In_1124,In_552);
or U402 (N_402,In_304,In_1333);
nor U403 (N_403,In_1448,In_1303);
nand U404 (N_404,In_1378,In_1234);
nand U405 (N_405,In_1423,In_897);
xnor U406 (N_406,In_222,In_831);
and U407 (N_407,In_427,In_266);
xor U408 (N_408,In_100,In_140);
nor U409 (N_409,In_267,In_211);
nor U410 (N_410,In_151,In_524);
xnor U411 (N_411,In_553,In_1471);
or U412 (N_412,In_717,In_1126);
nor U413 (N_413,In_663,In_446);
and U414 (N_414,In_978,In_291);
xnor U415 (N_415,In_792,In_1206);
and U416 (N_416,In_319,In_133);
and U417 (N_417,In_593,In_1469);
nor U418 (N_418,In_1061,In_80);
nor U419 (N_419,In_302,In_1188);
nor U420 (N_420,In_189,In_36);
nand U421 (N_421,In_1005,In_1264);
nor U422 (N_422,In_1311,In_1020);
nor U423 (N_423,In_285,In_1036);
nor U424 (N_424,In_314,In_1296);
or U425 (N_425,In_1239,In_848);
nor U426 (N_426,In_1192,In_178);
xnor U427 (N_427,In_1197,In_1201);
nand U428 (N_428,In_595,In_1463);
xor U429 (N_429,In_803,In_747);
nor U430 (N_430,In_325,In_1066);
and U431 (N_431,In_928,In_536);
nor U432 (N_432,In_563,In_666);
nand U433 (N_433,In_1459,In_305);
or U434 (N_434,In_824,In_976);
nand U435 (N_435,In_1191,In_1358);
and U436 (N_436,In_822,In_1315);
and U437 (N_437,In_735,In_1439);
and U438 (N_438,In_809,In_1189);
or U439 (N_439,In_966,In_534);
xnor U440 (N_440,In_1394,In_840);
nor U441 (N_441,In_165,In_197);
xor U442 (N_442,In_1273,In_827);
xnor U443 (N_443,In_481,In_895);
xor U444 (N_444,In_77,In_559);
nor U445 (N_445,In_320,In_1322);
nor U446 (N_446,In_1057,In_288);
nor U447 (N_447,In_557,In_916);
nand U448 (N_448,In_121,In_1009);
nor U449 (N_449,In_1417,In_1467);
or U450 (N_450,In_37,In_295);
and U451 (N_451,In_138,In_416);
xor U452 (N_452,In_1461,In_810);
or U453 (N_453,In_1275,In_1252);
nand U454 (N_454,In_409,In_1107);
nor U455 (N_455,In_1410,In_797);
xor U456 (N_456,In_1257,In_403);
xor U457 (N_457,In_1314,In_550);
or U458 (N_458,In_913,In_813);
xor U459 (N_459,In_494,In_106);
nor U460 (N_460,In_1158,In_275);
or U461 (N_461,In_879,In_551);
xnor U462 (N_462,In_246,In_652);
nor U463 (N_463,In_122,In_778);
xor U464 (N_464,In_1357,In_693);
xor U465 (N_465,In_478,In_1065);
and U466 (N_466,In_433,In_505);
or U467 (N_467,In_202,In_686);
and U468 (N_468,In_1203,In_1119);
nand U469 (N_469,In_1159,In_1111);
and U470 (N_470,In_359,In_646);
nor U471 (N_471,In_329,In_103);
and U472 (N_472,In_460,In_1014);
or U473 (N_473,In_1230,In_472);
nor U474 (N_474,In_1321,In_1393);
nand U475 (N_475,In_1195,In_136);
nand U476 (N_476,In_1254,In_17);
xnor U477 (N_477,In_234,In_1488);
and U478 (N_478,In_617,In_703);
and U479 (N_479,In_657,In_1243);
nand U480 (N_480,In_767,In_527);
xor U481 (N_481,In_1056,In_1076);
or U482 (N_482,In_750,In_200);
nor U483 (N_483,In_1369,In_847);
and U484 (N_484,In_772,In_186);
and U485 (N_485,In_1449,In_471);
or U486 (N_486,In_156,In_1332);
nand U487 (N_487,In_268,In_57);
xor U488 (N_488,In_1074,In_1418);
nor U489 (N_489,In_807,In_509);
nand U490 (N_490,In_410,In_208);
and U491 (N_491,In_493,In_90);
nor U492 (N_492,In_142,In_1060);
nand U493 (N_493,In_694,In_1481);
nor U494 (N_494,In_1348,In_1070);
and U495 (N_495,In_944,In_428);
or U496 (N_496,In_47,In_398);
xor U497 (N_497,In_487,In_437);
xor U498 (N_498,In_1067,In_1222);
nor U499 (N_499,In_623,In_114);
or U500 (N_500,In_193,In_639);
nor U501 (N_501,In_1039,In_1287);
nor U502 (N_502,In_779,In_642);
and U503 (N_503,In_842,In_1390);
nand U504 (N_504,In_187,In_1382);
or U505 (N_505,In_1344,In_1415);
nor U506 (N_506,In_548,In_1262);
nand U507 (N_507,In_261,In_878);
nand U508 (N_508,In_965,In_145);
or U509 (N_509,In_955,In_231);
nor U510 (N_510,In_327,In_718);
nand U511 (N_511,In_1242,In_22);
xor U512 (N_512,In_609,In_396);
or U513 (N_513,In_811,In_1091);
nor U514 (N_514,In_732,In_608);
or U515 (N_515,In_1362,In_922);
xnor U516 (N_516,In_637,In_139);
nand U517 (N_517,In_96,In_350);
or U518 (N_518,In_674,In_168);
and U519 (N_519,In_1101,In_969);
or U520 (N_520,In_477,In_1139);
and U521 (N_521,In_385,In_1479);
nor U522 (N_522,In_506,In_1293);
and U523 (N_523,In_466,In_699);
and U524 (N_524,In_869,In_681);
and U525 (N_525,In_702,In_1214);
or U526 (N_526,In_960,In_383);
nand U527 (N_527,In_364,In_586);
nand U528 (N_528,In_18,In_107);
and U529 (N_529,In_677,In_616);
nand U530 (N_530,In_1236,In_293);
xnor U531 (N_531,In_1082,In_1353);
nand U532 (N_532,In_556,In_1336);
nor U533 (N_533,In_492,In_1466);
or U534 (N_534,In_982,In_1280);
xnor U535 (N_535,In_365,In_649);
and U536 (N_536,In_14,In_921);
and U537 (N_537,In_1462,In_633);
xor U538 (N_538,In_814,In_696);
and U539 (N_539,In_1080,In_1079);
and U540 (N_540,In_182,In_530);
nand U541 (N_541,In_670,In_917);
nor U542 (N_542,In_989,In_442);
xor U543 (N_543,In_522,In_504);
nor U544 (N_544,In_865,In_1156);
nand U545 (N_545,In_1494,In_1249);
nand U546 (N_546,In_1258,In_1185);
and U547 (N_547,In_947,In_1389);
or U548 (N_548,In_591,In_1402);
xor U549 (N_549,In_1458,In_1116);
and U550 (N_550,In_783,In_296);
nor U551 (N_551,In_573,In_1090);
nor U552 (N_552,In_1370,In_213);
or U553 (N_553,In_896,In_957);
or U554 (N_554,In_490,In_1350);
nor U555 (N_555,In_83,In_289);
nand U556 (N_556,In_340,In_393);
xor U557 (N_557,In_543,In_1443);
and U558 (N_558,In_1063,In_503);
xnor U559 (N_559,In_292,In_373);
xnor U560 (N_560,In_731,In_1177);
nand U561 (N_561,In_839,In_597);
and U562 (N_562,In_1441,In_713);
xnor U563 (N_563,In_1376,In_799);
or U564 (N_564,In_755,In_338);
or U565 (N_565,In_596,In_119);
xnor U566 (N_566,In_765,In_1266);
or U567 (N_567,In_1487,In_59);
xor U568 (N_568,In_544,In_1217);
and U569 (N_569,In_474,In_102);
and U570 (N_570,In_191,In_1233);
or U571 (N_571,In_1013,In_1331);
nand U572 (N_572,In_227,In_900);
and U573 (N_573,In_655,In_1223);
nand U574 (N_574,In_528,In_541);
or U575 (N_575,In_1396,In_78);
or U576 (N_576,In_1455,In_347);
nand U577 (N_577,In_163,In_1499);
nand U578 (N_578,In_1434,In_844);
xnor U579 (N_579,In_1000,In_412);
or U580 (N_580,In_1245,In_318);
nor U581 (N_581,In_833,In_909);
xnor U582 (N_582,In_278,In_110);
and U583 (N_583,In_620,In_120);
or U584 (N_584,In_326,In_1142);
nor U585 (N_585,In_158,In_837);
and U586 (N_586,In_535,In_743);
nor U587 (N_587,In_1227,In_951);
or U588 (N_588,In_569,In_613);
nor U589 (N_589,In_441,In_1265);
xor U590 (N_590,In_348,In_344);
and U591 (N_591,In_1282,In_870);
and U592 (N_592,In_60,In_1334);
nor U593 (N_593,In_48,In_769);
nor U594 (N_594,In_706,In_746);
and U595 (N_595,In_413,In_1395);
nor U596 (N_596,In_604,In_1162);
nand U597 (N_597,In_920,In_1008);
nand U598 (N_598,In_462,In_752);
nor U599 (N_599,In_841,In_938);
nand U600 (N_600,In_887,In_812);
xnor U601 (N_601,In_1138,In_308);
xnor U602 (N_602,In_449,In_546);
nand U603 (N_603,In_776,In_252);
nor U604 (N_604,In_67,In_660);
and U605 (N_605,In_19,In_1267);
xnor U606 (N_606,In_357,In_941);
and U607 (N_607,In_1073,In_10);
nor U608 (N_608,In_1414,In_13);
or U609 (N_609,In_1355,In_1352);
nand U610 (N_610,In_127,In_830);
and U611 (N_611,In_194,In_1184);
xor U612 (N_612,In_38,In_313);
xnor U613 (N_613,In_972,In_1186);
nor U614 (N_614,In_1231,In_502);
nand U615 (N_615,In_607,In_692);
xor U616 (N_616,In_303,In_1377);
and U617 (N_617,In_521,In_1387);
xnor U618 (N_618,In_426,In_828);
xnor U619 (N_619,In_97,In_1490);
and U620 (N_620,In_641,In_927);
xnor U621 (N_621,In_1338,In_1096);
nor U622 (N_622,In_394,In_1300);
and U623 (N_623,In_482,In_875);
or U624 (N_624,In_892,In_224);
xor U625 (N_625,In_432,In_905);
xor U626 (N_626,In_459,In_354);
and U627 (N_627,In_185,In_1232);
nand U628 (N_628,In_926,In_740);
nand U629 (N_629,In_671,In_241);
and U630 (N_630,In_73,In_1413);
or U631 (N_631,In_30,In_801);
nor U632 (N_632,In_823,In_154);
or U633 (N_633,In_372,In_1170);
or U634 (N_634,In_391,In_1089);
nand U635 (N_635,In_1263,In_1238);
nor U636 (N_636,In_92,In_1145);
or U637 (N_637,In_997,In_1285);
nand U638 (N_638,In_777,In_339);
and U639 (N_639,In_523,In_697);
nor U640 (N_640,In_736,In_214);
nand U641 (N_641,In_1226,In_967);
xor U642 (N_642,In_244,In_1450);
nand U643 (N_643,In_257,In_656);
xnor U644 (N_644,In_1075,In_578);
nand U645 (N_645,In_328,In_146);
or U646 (N_646,In_610,In_1019);
nor U647 (N_647,In_1486,In_1319);
xnor U648 (N_648,In_600,In_880);
nand U649 (N_649,In_914,In_1308);
nor U650 (N_650,In_934,In_687);
nand U651 (N_651,In_125,In_619);
and U652 (N_652,In_1445,In_356);
nor U653 (N_653,In_924,In_43);
nor U654 (N_654,In_51,In_1442);
xor U655 (N_655,In_46,In_1247);
xor U656 (N_656,In_773,In_662);
nor U657 (N_657,In_1028,In_443);
xor U658 (N_658,In_1484,In_221);
or U659 (N_659,In_1274,In_689);
nand U660 (N_660,In_1229,In_1302);
xor U661 (N_661,In_525,In_1021);
and U662 (N_662,In_144,In_1117);
nand U663 (N_663,In_705,In_265);
or U664 (N_664,In_1164,In_984);
or U665 (N_665,In_1347,In_1012);
and U666 (N_666,In_49,In_1047);
and U667 (N_667,In_453,In_1132);
and U668 (N_668,In_1169,In_567);
or U669 (N_669,In_309,In_1157);
nand U670 (N_670,In_721,In_566);
and U671 (N_671,In_210,In_983);
nor U672 (N_672,In_371,In_1429);
xor U673 (N_673,In_1421,In_1400);
or U674 (N_674,In_939,In_1483);
xnor U675 (N_675,In_287,In_335);
nand U676 (N_676,In_1412,In_1150);
nor U677 (N_677,In_1103,In_886);
xor U678 (N_678,In_1433,In_161);
and U679 (N_679,In_181,In_331);
or U680 (N_680,In_336,In_1422);
and U681 (N_681,In_720,In_422);
or U682 (N_682,In_1440,In_1114);
nand U683 (N_683,In_397,In_561);
nand U684 (N_684,In_867,In_424);
nor U685 (N_685,In_253,In_1290);
or U686 (N_686,In_1196,In_1224);
and U687 (N_687,In_108,In_440);
or U688 (N_688,In_218,In_1437);
nor U689 (N_689,In_1419,In_386);
nand U690 (N_690,In_624,In_634);
or U691 (N_691,In_175,In_62);
or U692 (N_692,In_1301,In_1354);
and U693 (N_693,In_562,In_155);
and U694 (N_694,In_665,In_216);
nand U695 (N_695,In_1010,In_406);
or U696 (N_696,In_1016,In_1007);
nand U697 (N_697,In_688,In_447);
or U698 (N_698,In_162,In_719);
or U699 (N_699,In_160,In_207);
nor U700 (N_700,In_1498,In_388);
xnor U701 (N_701,In_1365,In_977);
nor U702 (N_702,In_850,In_1098);
nor U703 (N_703,In_1144,In_1246);
and U704 (N_704,In_739,In_1404);
or U705 (N_705,In_1044,In_264);
nor U706 (N_706,In_1284,In_514);
or U707 (N_707,In_753,In_395);
nor U708 (N_708,In_1313,In_558);
nor U709 (N_709,In_64,In_20);
and U710 (N_710,In_1279,In_782);
or U711 (N_711,In_26,In_88);
xnor U712 (N_712,In_631,In_1327);
xor U713 (N_713,In_237,In_1408);
or U714 (N_714,In_738,In_885);
xor U715 (N_715,In_1052,In_621);
and U716 (N_716,In_415,In_1207);
or U717 (N_717,In_1366,In_1328);
and U718 (N_718,In_25,In_510);
nand U719 (N_719,In_172,In_1248);
nand U720 (N_720,In_258,In_1118);
nor U721 (N_721,In_232,In_1320);
or U722 (N_722,In_31,In_1069);
nor U723 (N_723,In_1324,In_1253);
xnor U724 (N_724,In_148,In_571);
xnor U725 (N_725,In_863,In_1476);
nand U726 (N_726,In_486,In_954);
nand U727 (N_727,In_991,In_1220);
xor U728 (N_728,In_876,In_884);
or U729 (N_729,In_1133,In_68);
xnor U730 (N_730,In_209,In_16);
and U731 (N_731,In_27,In_229);
and U732 (N_732,In_555,In_322);
nor U733 (N_733,In_1216,In_235);
xor U734 (N_734,In_1062,In_203);
nor U735 (N_735,In_259,In_166);
nand U736 (N_736,In_480,In_775);
nor U737 (N_737,In_1011,In_137);
or U738 (N_738,In_545,In_890);
or U739 (N_739,In_1183,In_262);
nand U740 (N_740,In_436,In_592);
nand U741 (N_741,In_647,In_576);
nor U742 (N_742,In_1294,In_741);
or U743 (N_743,In_1106,In_1268);
nand U744 (N_744,In_640,In_682);
and U745 (N_745,In_269,In_270);
nand U746 (N_746,In_512,In_1032);
xor U747 (N_747,In_1388,In_468);
nand U748 (N_748,In_888,In_195);
nor U749 (N_749,In_816,In_854);
or U750 (N_750,In_376,In_1218);
xnor U751 (N_751,In_1007,In_1408);
nor U752 (N_752,In_1462,In_291);
xor U753 (N_753,In_923,In_1167);
xnor U754 (N_754,In_1086,In_496);
nor U755 (N_755,In_1382,In_1243);
or U756 (N_756,In_652,In_1284);
xor U757 (N_757,In_1279,In_582);
or U758 (N_758,In_1335,In_382);
or U759 (N_759,In_464,In_1185);
xor U760 (N_760,In_1297,In_869);
or U761 (N_761,In_1445,In_157);
or U762 (N_762,In_405,In_779);
nand U763 (N_763,In_1310,In_812);
xor U764 (N_764,In_227,In_257);
xnor U765 (N_765,In_873,In_1178);
and U766 (N_766,In_361,In_1186);
nand U767 (N_767,In_1382,In_621);
nor U768 (N_768,In_1439,In_1290);
and U769 (N_769,In_256,In_1146);
xnor U770 (N_770,In_1452,In_294);
xor U771 (N_771,In_1164,In_280);
or U772 (N_772,In_691,In_318);
xor U773 (N_773,In_755,In_561);
xnor U774 (N_774,In_1407,In_1130);
nand U775 (N_775,In_883,In_902);
and U776 (N_776,In_1010,In_878);
nor U777 (N_777,In_1308,In_1478);
xor U778 (N_778,In_591,In_157);
and U779 (N_779,In_28,In_794);
and U780 (N_780,In_1099,In_1471);
nor U781 (N_781,In_277,In_73);
xor U782 (N_782,In_787,In_849);
or U783 (N_783,In_800,In_50);
xor U784 (N_784,In_217,In_1476);
or U785 (N_785,In_686,In_1405);
xor U786 (N_786,In_1167,In_783);
xnor U787 (N_787,In_639,In_765);
or U788 (N_788,In_848,In_472);
xor U789 (N_789,In_968,In_9);
nand U790 (N_790,In_832,In_440);
xor U791 (N_791,In_765,In_440);
or U792 (N_792,In_1065,In_1493);
nor U793 (N_793,In_531,In_300);
nand U794 (N_794,In_1055,In_293);
and U795 (N_795,In_793,In_371);
or U796 (N_796,In_1221,In_920);
or U797 (N_797,In_1187,In_738);
and U798 (N_798,In_90,In_1220);
xnor U799 (N_799,In_1055,In_816);
nand U800 (N_800,In_1204,In_872);
and U801 (N_801,In_1285,In_1277);
xor U802 (N_802,In_1215,In_914);
or U803 (N_803,In_645,In_1123);
and U804 (N_804,In_1419,In_336);
and U805 (N_805,In_1274,In_667);
or U806 (N_806,In_988,In_1183);
nand U807 (N_807,In_813,In_735);
or U808 (N_808,In_1236,In_618);
or U809 (N_809,In_1421,In_128);
nor U810 (N_810,In_22,In_1326);
nor U811 (N_811,In_585,In_1428);
or U812 (N_812,In_91,In_405);
xnor U813 (N_813,In_1276,In_755);
nand U814 (N_814,In_113,In_1264);
and U815 (N_815,In_382,In_1237);
and U816 (N_816,In_744,In_427);
xnor U817 (N_817,In_1245,In_660);
nor U818 (N_818,In_1118,In_1044);
nor U819 (N_819,In_1484,In_835);
and U820 (N_820,In_1496,In_1091);
nor U821 (N_821,In_1406,In_521);
nand U822 (N_822,In_1129,In_1110);
or U823 (N_823,In_1017,In_568);
xor U824 (N_824,In_1186,In_1456);
nand U825 (N_825,In_785,In_686);
nor U826 (N_826,In_870,In_671);
or U827 (N_827,In_1149,In_1257);
nand U828 (N_828,In_1427,In_531);
xnor U829 (N_829,In_343,In_1441);
nor U830 (N_830,In_765,In_1089);
nor U831 (N_831,In_494,In_1426);
and U832 (N_832,In_399,In_947);
xor U833 (N_833,In_1159,In_114);
nor U834 (N_834,In_200,In_302);
nand U835 (N_835,In_72,In_560);
xor U836 (N_836,In_50,In_1250);
xor U837 (N_837,In_620,In_1138);
nand U838 (N_838,In_402,In_1075);
and U839 (N_839,In_1067,In_1338);
nand U840 (N_840,In_1134,In_735);
and U841 (N_841,In_164,In_180);
nor U842 (N_842,In_417,In_943);
or U843 (N_843,In_1116,In_136);
nor U844 (N_844,In_902,In_1106);
and U845 (N_845,In_482,In_180);
nand U846 (N_846,In_1279,In_1257);
nand U847 (N_847,In_167,In_854);
or U848 (N_848,In_1458,In_604);
nand U849 (N_849,In_87,In_1060);
nor U850 (N_850,In_731,In_977);
nand U851 (N_851,In_383,In_1300);
nor U852 (N_852,In_948,In_90);
nor U853 (N_853,In_355,In_484);
xnor U854 (N_854,In_1187,In_1005);
and U855 (N_855,In_1338,In_1371);
or U856 (N_856,In_1202,In_1426);
nor U857 (N_857,In_715,In_1164);
or U858 (N_858,In_924,In_1056);
and U859 (N_859,In_560,In_326);
and U860 (N_860,In_1101,In_1068);
xor U861 (N_861,In_919,In_886);
nor U862 (N_862,In_898,In_624);
nand U863 (N_863,In_1173,In_1067);
nor U864 (N_864,In_275,In_397);
and U865 (N_865,In_738,In_146);
and U866 (N_866,In_527,In_45);
or U867 (N_867,In_545,In_1048);
or U868 (N_868,In_402,In_1192);
nand U869 (N_869,In_715,In_769);
nand U870 (N_870,In_1031,In_527);
or U871 (N_871,In_442,In_133);
and U872 (N_872,In_1277,In_588);
and U873 (N_873,In_445,In_43);
nand U874 (N_874,In_290,In_1231);
xor U875 (N_875,In_1371,In_341);
nand U876 (N_876,In_623,In_1466);
nand U877 (N_877,In_1296,In_382);
nor U878 (N_878,In_684,In_1391);
nand U879 (N_879,In_191,In_1065);
or U880 (N_880,In_1413,In_324);
or U881 (N_881,In_503,In_459);
nor U882 (N_882,In_1246,In_1103);
nand U883 (N_883,In_27,In_320);
nand U884 (N_884,In_400,In_310);
or U885 (N_885,In_83,In_508);
nor U886 (N_886,In_1269,In_52);
or U887 (N_887,In_470,In_1074);
or U888 (N_888,In_394,In_191);
or U889 (N_889,In_1442,In_34);
xnor U890 (N_890,In_208,In_583);
nand U891 (N_891,In_200,In_1392);
nor U892 (N_892,In_101,In_899);
nand U893 (N_893,In_1489,In_26);
xnor U894 (N_894,In_1345,In_1002);
nor U895 (N_895,In_671,In_539);
or U896 (N_896,In_403,In_55);
and U897 (N_897,In_545,In_208);
or U898 (N_898,In_543,In_536);
or U899 (N_899,In_803,In_273);
nor U900 (N_900,In_609,In_1121);
or U901 (N_901,In_306,In_148);
nand U902 (N_902,In_892,In_839);
nand U903 (N_903,In_1184,In_716);
xor U904 (N_904,In_1492,In_1089);
nor U905 (N_905,In_479,In_0);
or U906 (N_906,In_118,In_1163);
xor U907 (N_907,In_209,In_251);
and U908 (N_908,In_1241,In_1004);
xnor U909 (N_909,In_1189,In_409);
nor U910 (N_910,In_733,In_451);
nor U911 (N_911,In_1068,In_200);
nand U912 (N_912,In_1379,In_376);
nor U913 (N_913,In_1246,In_652);
nor U914 (N_914,In_1209,In_1352);
xnor U915 (N_915,In_234,In_561);
and U916 (N_916,In_8,In_611);
nor U917 (N_917,In_567,In_937);
nand U918 (N_918,In_496,In_394);
nor U919 (N_919,In_1436,In_1339);
nand U920 (N_920,In_561,In_892);
xor U921 (N_921,In_668,In_351);
nor U922 (N_922,In_974,In_637);
xor U923 (N_923,In_1027,In_1339);
nand U924 (N_924,In_982,In_381);
xnor U925 (N_925,In_804,In_728);
nand U926 (N_926,In_1004,In_852);
xnor U927 (N_927,In_415,In_257);
xor U928 (N_928,In_555,In_1305);
nand U929 (N_929,In_932,In_1075);
and U930 (N_930,In_1253,In_372);
xor U931 (N_931,In_1388,In_847);
or U932 (N_932,In_830,In_780);
nand U933 (N_933,In_1420,In_428);
or U934 (N_934,In_352,In_568);
xor U935 (N_935,In_1464,In_1287);
nand U936 (N_936,In_318,In_948);
nand U937 (N_937,In_790,In_950);
nor U938 (N_938,In_748,In_716);
nand U939 (N_939,In_668,In_950);
or U940 (N_940,In_1148,In_1244);
or U941 (N_941,In_600,In_386);
and U942 (N_942,In_652,In_1008);
and U943 (N_943,In_1328,In_1056);
nor U944 (N_944,In_972,In_805);
and U945 (N_945,In_1279,In_992);
and U946 (N_946,In_737,In_964);
nand U947 (N_947,In_1347,In_1256);
xor U948 (N_948,In_1365,In_1007);
and U949 (N_949,In_520,In_647);
or U950 (N_950,In_516,In_1118);
nand U951 (N_951,In_664,In_625);
xor U952 (N_952,In_178,In_52);
or U953 (N_953,In_941,In_675);
nand U954 (N_954,In_1205,In_434);
or U955 (N_955,In_1147,In_470);
or U956 (N_956,In_112,In_1477);
nand U957 (N_957,In_231,In_1055);
nand U958 (N_958,In_360,In_1295);
xnor U959 (N_959,In_942,In_519);
nor U960 (N_960,In_351,In_498);
xnor U961 (N_961,In_527,In_915);
nand U962 (N_962,In_621,In_1233);
or U963 (N_963,In_855,In_1478);
and U964 (N_964,In_800,In_482);
nand U965 (N_965,In_1093,In_269);
and U966 (N_966,In_1006,In_1146);
nor U967 (N_967,In_219,In_1460);
nor U968 (N_968,In_1130,In_420);
nor U969 (N_969,In_670,In_1375);
nand U970 (N_970,In_199,In_558);
xnor U971 (N_971,In_1267,In_914);
or U972 (N_972,In_125,In_784);
nand U973 (N_973,In_793,In_1119);
and U974 (N_974,In_885,In_143);
nor U975 (N_975,In_387,In_597);
nor U976 (N_976,In_752,In_1050);
or U977 (N_977,In_1046,In_300);
xnor U978 (N_978,In_1227,In_791);
or U979 (N_979,In_1240,In_1394);
or U980 (N_980,In_850,In_111);
xnor U981 (N_981,In_1239,In_942);
and U982 (N_982,In_1016,In_449);
xnor U983 (N_983,In_815,In_1355);
or U984 (N_984,In_851,In_1200);
or U985 (N_985,In_1114,In_544);
nand U986 (N_986,In_522,In_85);
nand U987 (N_987,In_838,In_1487);
xnor U988 (N_988,In_489,In_1269);
xor U989 (N_989,In_1132,In_634);
nand U990 (N_990,In_1255,In_1283);
nor U991 (N_991,In_631,In_1490);
xnor U992 (N_992,In_472,In_997);
xor U993 (N_993,In_633,In_575);
or U994 (N_994,In_1089,In_50);
and U995 (N_995,In_961,In_1319);
or U996 (N_996,In_558,In_1298);
or U997 (N_997,In_1156,In_522);
nor U998 (N_998,In_717,In_833);
nor U999 (N_999,In_264,In_1401);
and U1000 (N_1000,In_1355,In_375);
nand U1001 (N_1001,In_273,In_310);
or U1002 (N_1002,In_1319,In_1374);
nand U1003 (N_1003,In_21,In_101);
or U1004 (N_1004,In_1147,In_301);
nand U1005 (N_1005,In_880,In_1124);
xor U1006 (N_1006,In_787,In_1311);
nor U1007 (N_1007,In_999,In_300);
or U1008 (N_1008,In_962,In_335);
or U1009 (N_1009,In_743,In_1036);
nor U1010 (N_1010,In_124,In_762);
and U1011 (N_1011,In_378,In_223);
nor U1012 (N_1012,In_980,In_722);
nor U1013 (N_1013,In_859,In_1207);
xnor U1014 (N_1014,In_1285,In_1405);
or U1015 (N_1015,In_160,In_1163);
nand U1016 (N_1016,In_87,In_818);
xnor U1017 (N_1017,In_1146,In_1295);
and U1018 (N_1018,In_1089,In_853);
nand U1019 (N_1019,In_462,In_1464);
or U1020 (N_1020,In_137,In_1466);
and U1021 (N_1021,In_776,In_1242);
or U1022 (N_1022,In_764,In_8);
and U1023 (N_1023,In_1478,In_959);
nor U1024 (N_1024,In_231,In_961);
or U1025 (N_1025,In_638,In_1412);
xnor U1026 (N_1026,In_1191,In_1193);
and U1027 (N_1027,In_791,In_853);
nor U1028 (N_1028,In_1256,In_441);
nor U1029 (N_1029,In_668,In_518);
xnor U1030 (N_1030,In_650,In_667);
nand U1031 (N_1031,In_374,In_120);
xnor U1032 (N_1032,In_483,In_1145);
and U1033 (N_1033,In_135,In_305);
nand U1034 (N_1034,In_1023,In_607);
nand U1035 (N_1035,In_1341,In_756);
nand U1036 (N_1036,In_155,In_737);
or U1037 (N_1037,In_585,In_1152);
and U1038 (N_1038,In_1224,In_1198);
or U1039 (N_1039,In_1305,In_154);
nand U1040 (N_1040,In_853,In_1152);
xor U1041 (N_1041,In_541,In_796);
or U1042 (N_1042,In_1069,In_1144);
nand U1043 (N_1043,In_502,In_548);
nand U1044 (N_1044,In_1250,In_1283);
xor U1045 (N_1045,In_649,In_550);
and U1046 (N_1046,In_68,In_612);
xnor U1047 (N_1047,In_1050,In_818);
xor U1048 (N_1048,In_828,In_343);
nand U1049 (N_1049,In_1455,In_515);
or U1050 (N_1050,In_630,In_752);
nor U1051 (N_1051,In_1061,In_718);
xnor U1052 (N_1052,In_532,In_683);
or U1053 (N_1053,In_790,In_412);
nor U1054 (N_1054,In_413,In_97);
or U1055 (N_1055,In_1278,In_1425);
and U1056 (N_1056,In_818,In_467);
nor U1057 (N_1057,In_1193,In_666);
xor U1058 (N_1058,In_926,In_902);
and U1059 (N_1059,In_1397,In_590);
nand U1060 (N_1060,In_917,In_383);
and U1061 (N_1061,In_926,In_1122);
xnor U1062 (N_1062,In_1044,In_566);
nor U1063 (N_1063,In_776,In_1246);
nand U1064 (N_1064,In_133,In_1004);
and U1065 (N_1065,In_650,In_327);
xnor U1066 (N_1066,In_1163,In_1244);
and U1067 (N_1067,In_1427,In_1436);
or U1068 (N_1068,In_151,In_250);
nor U1069 (N_1069,In_1037,In_774);
nor U1070 (N_1070,In_1399,In_880);
nand U1071 (N_1071,In_1436,In_1291);
nand U1072 (N_1072,In_166,In_727);
nor U1073 (N_1073,In_662,In_77);
or U1074 (N_1074,In_1338,In_450);
nand U1075 (N_1075,In_135,In_359);
nand U1076 (N_1076,In_655,In_168);
nor U1077 (N_1077,In_1364,In_1433);
nand U1078 (N_1078,In_1325,In_63);
and U1079 (N_1079,In_620,In_1405);
nor U1080 (N_1080,In_1460,In_1285);
or U1081 (N_1081,In_1176,In_1351);
or U1082 (N_1082,In_1151,In_1460);
nand U1083 (N_1083,In_284,In_885);
nand U1084 (N_1084,In_342,In_1122);
xor U1085 (N_1085,In_289,In_67);
nor U1086 (N_1086,In_1057,In_1132);
nor U1087 (N_1087,In_523,In_541);
or U1088 (N_1088,In_785,In_351);
nand U1089 (N_1089,In_134,In_1042);
and U1090 (N_1090,In_951,In_1334);
nor U1091 (N_1091,In_894,In_11);
nor U1092 (N_1092,In_967,In_261);
nor U1093 (N_1093,In_769,In_427);
xor U1094 (N_1094,In_974,In_670);
nand U1095 (N_1095,In_939,In_382);
xor U1096 (N_1096,In_181,In_512);
and U1097 (N_1097,In_297,In_1139);
nand U1098 (N_1098,In_888,In_817);
xor U1099 (N_1099,In_1182,In_1221);
or U1100 (N_1100,In_150,In_25);
and U1101 (N_1101,In_1022,In_267);
nor U1102 (N_1102,In_503,In_227);
or U1103 (N_1103,In_571,In_27);
xnor U1104 (N_1104,In_975,In_530);
xnor U1105 (N_1105,In_1435,In_746);
nor U1106 (N_1106,In_1468,In_606);
nor U1107 (N_1107,In_513,In_0);
and U1108 (N_1108,In_339,In_1457);
nand U1109 (N_1109,In_1179,In_675);
or U1110 (N_1110,In_736,In_1338);
xor U1111 (N_1111,In_1095,In_321);
xor U1112 (N_1112,In_852,In_1217);
nand U1113 (N_1113,In_93,In_344);
or U1114 (N_1114,In_573,In_950);
nand U1115 (N_1115,In_879,In_1065);
and U1116 (N_1116,In_975,In_1465);
xnor U1117 (N_1117,In_1181,In_216);
or U1118 (N_1118,In_1017,In_1179);
xor U1119 (N_1119,In_1110,In_863);
xnor U1120 (N_1120,In_337,In_1089);
nand U1121 (N_1121,In_661,In_1157);
or U1122 (N_1122,In_783,In_1161);
xor U1123 (N_1123,In_237,In_112);
and U1124 (N_1124,In_1200,In_690);
nor U1125 (N_1125,In_994,In_1127);
and U1126 (N_1126,In_290,In_203);
nor U1127 (N_1127,In_37,In_211);
or U1128 (N_1128,In_402,In_1324);
xor U1129 (N_1129,In_1159,In_180);
or U1130 (N_1130,In_246,In_218);
or U1131 (N_1131,In_111,In_623);
nand U1132 (N_1132,In_183,In_649);
nor U1133 (N_1133,In_1112,In_989);
nand U1134 (N_1134,In_71,In_1268);
nor U1135 (N_1135,In_457,In_173);
or U1136 (N_1136,In_484,In_1455);
and U1137 (N_1137,In_190,In_71);
or U1138 (N_1138,In_941,In_413);
and U1139 (N_1139,In_1304,In_715);
nor U1140 (N_1140,In_192,In_1244);
nor U1141 (N_1141,In_1469,In_667);
nand U1142 (N_1142,In_1141,In_983);
and U1143 (N_1143,In_1326,In_130);
nor U1144 (N_1144,In_1003,In_1234);
and U1145 (N_1145,In_85,In_679);
nand U1146 (N_1146,In_1009,In_1243);
xor U1147 (N_1147,In_1394,In_592);
nor U1148 (N_1148,In_296,In_683);
or U1149 (N_1149,In_691,In_811);
or U1150 (N_1150,In_465,In_759);
nand U1151 (N_1151,In_1319,In_29);
or U1152 (N_1152,In_738,In_676);
and U1153 (N_1153,In_1371,In_853);
nand U1154 (N_1154,In_1367,In_1172);
and U1155 (N_1155,In_1301,In_378);
nor U1156 (N_1156,In_824,In_743);
or U1157 (N_1157,In_195,In_1115);
nand U1158 (N_1158,In_1488,In_564);
and U1159 (N_1159,In_336,In_785);
nor U1160 (N_1160,In_1144,In_543);
xnor U1161 (N_1161,In_1098,In_295);
and U1162 (N_1162,In_1118,In_178);
xnor U1163 (N_1163,In_1244,In_1414);
or U1164 (N_1164,In_785,In_1158);
nor U1165 (N_1165,In_1001,In_123);
or U1166 (N_1166,In_207,In_1382);
nor U1167 (N_1167,In_273,In_1463);
xor U1168 (N_1168,In_845,In_1077);
nor U1169 (N_1169,In_1150,In_1006);
or U1170 (N_1170,In_375,In_782);
nand U1171 (N_1171,In_780,In_1235);
nand U1172 (N_1172,In_828,In_988);
xor U1173 (N_1173,In_903,In_1164);
xor U1174 (N_1174,In_1237,In_1090);
nor U1175 (N_1175,In_1037,In_706);
nor U1176 (N_1176,In_1281,In_629);
or U1177 (N_1177,In_307,In_469);
nand U1178 (N_1178,In_263,In_60);
xor U1179 (N_1179,In_531,In_369);
xor U1180 (N_1180,In_1318,In_15);
and U1181 (N_1181,In_494,In_2);
and U1182 (N_1182,In_872,In_1007);
or U1183 (N_1183,In_1130,In_899);
and U1184 (N_1184,In_1164,In_436);
or U1185 (N_1185,In_1439,In_998);
nor U1186 (N_1186,In_25,In_341);
nor U1187 (N_1187,In_131,In_928);
nor U1188 (N_1188,In_1118,In_314);
or U1189 (N_1189,In_1387,In_1020);
and U1190 (N_1190,In_1371,In_929);
nor U1191 (N_1191,In_779,In_1403);
nand U1192 (N_1192,In_707,In_1299);
nand U1193 (N_1193,In_287,In_394);
or U1194 (N_1194,In_789,In_231);
xnor U1195 (N_1195,In_427,In_355);
xor U1196 (N_1196,In_1170,In_569);
xor U1197 (N_1197,In_402,In_1305);
and U1198 (N_1198,In_166,In_198);
xnor U1199 (N_1199,In_756,In_417);
or U1200 (N_1200,In_1048,In_160);
nand U1201 (N_1201,In_675,In_1077);
nand U1202 (N_1202,In_1390,In_881);
nand U1203 (N_1203,In_199,In_549);
nor U1204 (N_1204,In_1290,In_209);
nand U1205 (N_1205,In_1316,In_1031);
or U1206 (N_1206,In_1100,In_246);
or U1207 (N_1207,In_559,In_821);
nor U1208 (N_1208,In_89,In_988);
or U1209 (N_1209,In_160,In_118);
or U1210 (N_1210,In_362,In_899);
and U1211 (N_1211,In_486,In_610);
or U1212 (N_1212,In_370,In_4);
and U1213 (N_1213,In_136,In_1216);
nand U1214 (N_1214,In_373,In_370);
nor U1215 (N_1215,In_883,In_1417);
or U1216 (N_1216,In_578,In_125);
and U1217 (N_1217,In_1314,In_1409);
or U1218 (N_1218,In_362,In_1395);
xnor U1219 (N_1219,In_239,In_200);
and U1220 (N_1220,In_792,In_1090);
nor U1221 (N_1221,In_331,In_123);
nor U1222 (N_1222,In_805,In_1375);
or U1223 (N_1223,In_851,In_946);
xor U1224 (N_1224,In_1428,In_365);
nor U1225 (N_1225,In_496,In_883);
xnor U1226 (N_1226,In_269,In_1373);
and U1227 (N_1227,In_716,In_1189);
nor U1228 (N_1228,In_632,In_502);
nand U1229 (N_1229,In_514,In_1073);
nand U1230 (N_1230,In_1020,In_165);
nand U1231 (N_1231,In_165,In_1478);
xor U1232 (N_1232,In_313,In_400);
xor U1233 (N_1233,In_244,In_116);
xor U1234 (N_1234,In_1070,In_1471);
or U1235 (N_1235,In_487,In_690);
xnor U1236 (N_1236,In_1477,In_919);
nand U1237 (N_1237,In_327,In_1288);
or U1238 (N_1238,In_464,In_1165);
nor U1239 (N_1239,In_368,In_139);
nor U1240 (N_1240,In_517,In_476);
xor U1241 (N_1241,In_1416,In_248);
xnor U1242 (N_1242,In_664,In_1290);
nand U1243 (N_1243,In_936,In_1470);
nand U1244 (N_1244,In_1279,In_1422);
or U1245 (N_1245,In_905,In_482);
nand U1246 (N_1246,In_1210,In_1002);
and U1247 (N_1247,In_1205,In_53);
nand U1248 (N_1248,In_608,In_896);
nand U1249 (N_1249,In_791,In_1499);
xor U1250 (N_1250,In_969,In_1002);
xor U1251 (N_1251,In_1388,In_818);
xnor U1252 (N_1252,In_1159,In_868);
xnor U1253 (N_1253,In_687,In_36);
nor U1254 (N_1254,In_945,In_682);
or U1255 (N_1255,In_59,In_1489);
nand U1256 (N_1256,In_409,In_348);
and U1257 (N_1257,In_923,In_942);
or U1258 (N_1258,In_290,In_906);
nand U1259 (N_1259,In_1230,In_1064);
nand U1260 (N_1260,In_742,In_400);
nand U1261 (N_1261,In_777,In_1242);
and U1262 (N_1262,In_291,In_570);
and U1263 (N_1263,In_801,In_682);
or U1264 (N_1264,In_98,In_444);
nand U1265 (N_1265,In_1295,In_447);
and U1266 (N_1266,In_88,In_1416);
xor U1267 (N_1267,In_1306,In_776);
xor U1268 (N_1268,In_13,In_1034);
nand U1269 (N_1269,In_56,In_748);
or U1270 (N_1270,In_112,In_734);
nand U1271 (N_1271,In_1044,In_1017);
or U1272 (N_1272,In_505,In_793);
xnor U1273 (N_1273,In_1404,In_921);
and U1274 (N_1274,In_685,In_81);
and U1275 (N_1275,In_122,In_503);
nand U1276 (N_1276,In_347,In_560);
or U1277 (N_1277,In_271,In_967);
nand U1278 (N_1278,In_49,In_820);
nand U1279 (N_1279,In_650,In_798);
and U1280 (N_1280,In_538,In_61);
or U1281 (N_1281,In_1170,In_415);
or U1282 (N_1282,In_708,In_1111);
nand U1283 (N_1283,In_1341,In_683);
xnor U1284 (N_1284,In_1039,In_1087);
and U1285 (N_1285,In_1498,In_777);
nor U1286 (N_1286,In_722,In_1067);
or U1287 (N_1287,In_300,In_1372);
nor U1288 (N_1288,In_269,In_1396);
nand U1289 (N_1289,In_1042,In_591);
or U1290 (N_1290,In_92,In_280);
or U1291 (N_1291,In_514,In_1369);
xor U1292 (N_1292,In_257,In_1455);
nor U1293 (N_1293,In_855,In_1286);
and U1294 (N_1294,In_889,In_810);
or U1295 (N_1295,In_235,In_512);
nor U1296 (N_1296,In_1360,In_212);
nand U1297 (N_1297,In_471,In_1141);
nand U1298 (N_1298,In_430,In_437);
nand U1299 (N_1299,In_671,In_922);
nor U1300 (N_1300,In_1114,In_42);
or U1301 (N_1301,In_974,In_1140);
xor U1302 (N_1302,In_812,In_1309);
xnor U1303 (N_1303,In_898,In_198);
nand U1304 (N_1304,In_12,In_26);
nor U1305 (N_1305,In_15,In_527);
nand U1306 (N_1306,In_626,In_59);
or U1307 (N_1307,In_1428,In_1437);
nor U1308 (N_1308,In_840,In_1134);
and U1309 (N_1309,In_418,In_1065);
or U1310 (N_1310,In_694,In_548);
nand U1311 (N_1311,In_874,In_138);
nor U1312 (N_1312,In_623,In_951);
nand U1313 (N_1313,In_554,In_617);
nand U1314 (N_1314,In_882,In_1441);
nor U1315 (N_1315,In_755,In_426);
xnor U1316 (N_1316,In_694,In_771);
and U1317 (N_1317,In_1111,In_863);
and U1318 (N_1318,In_1299,In_62);
xnor U1319 (N_1319,In_1283,In_1038);
or U1320 (N_1320,In_791,In_1336);
xnor U1321 (N_1321,In_308,In_998);
or U1322 (N_1322,In_865,In_622);
nand U1323 (N_1323,In_200,In_1119);
xnor U1324 (N_1324,In_648,In_48);
nor U1325 (N_1325,In_1258,In_496);
nand U1326 (N_1326,In_673,In_333);
xor U1327 (N_1327,In_849,In_72);
xnor U1328 (N_1328,In_338,In_478);
nor U1329 (N_1329,In_685,In_175);
nor U1330 (N_1330,In_766,In_478);
nor U1331 (N_1331,In_811,In_341);
or U1332 (N_1332,In_168,In_1050);
or U1333 (N_1333,In_205,In_1459);
nor U1334 (N_1334,In_1015,In_741);
or U1335 (N_1335,In_841,In_775);
xnor U1336 (N_1336,In_147,In_542);
or U1337 (N_1337,In_1408,In_410);
nand U1338 (N_1338,In_523,In_837);
nand U1339 (N_1339,In_575,In_877);
nand U1340 (N_1340,In_1434,In_1061);
nand U1341 (N_1341,In_1428,In_1251);
nand U1342 (N_1342,In_664,In_1339);
nor U1343 (N_1343,In_613,In_44);
and U1344 (N_1344,In_1458,In_554);
nor U1345 (N_1345,In_669,In_1070);
xnor U1346 (N_1346,In_1185,In_703);
xnor U1347 (N_1347,In_961,In_914);
nor U1348 (N_1348,In_1374,In_1014);
nor U1349 (N_1349,In_58,In_944);
nor U1350 (N_1350,In_629,In_1438);
nor U1351 (N_1351,In_1467,In_843);
nand U1352 (N_1352,In_1005,In_112);
nor U1353 (N_1353,In_1039,In_948);
nand U1354 (N_1354,In_935,In_262);
xor U1355 (N_1355,In_439,In_18);
or U1356 (N_1356,In_1459,In_133);
nor U1357 (N_1357,In_428,In_355);
nand U1358 (N_1358,In_1081,In_946);
nor U1359 (N_1359,In_401,In_599);
nor U1360 (N_1360,In_984,In_417);
xor U1361 (N_1361,In_1429,In_1074);
xor U1362 (N_1362,In_59,In_752);
or U1363 (N_1363,In_1191,In_589);
and U1364 (N_1364,In_1187,In_938);
nand U1365 (N_1365,In_196,In_1049);
or U1366 (N_1366,In_727,In_213);
nand U1367 (N_1367,In_552,In_1395);
nand U1368 (N_1368,In_226,In_1304);
nand U1369 (N_1369,In_851,In_710);
and U1370 (N_1370,In_842,In_1294);
or U1371 (N_1371,In_299,In_1083);
nor U1372 (N_1372,In_592,In_562);
or U1373 (N_1373,In_506,In_213);
xnor U1374 (N_1374,In_116,In_1444);
xor U1375 (N_1375,In_1284,In_1138);
xor U1376 (N_1376,In_621,In_99);
or U1377 (N_1377,In_574,In_1444);
and U1378 (N_1378,In_141,In_778);
or U1379 (N_1379,In_170,In_407);
nand U1380 (N_1380,In_954,In_366);
and U1381 (N_1381,In_646,In_682);
xnor U1382 (N_1382,In_214,In_476);
nand U1383 (N_1383,In_1105,In_856);
xor U1384 (N_1384,In_979,In_9);
nand U1385 (N_1385,In_985,In_604);
xor U1386 (N_1386,In_24,In_637);
xnor U1387 (N_1387,In_814,In_95);
nor U1388 (N_1388,In_1008,In_365);
or U1389 (N_1389,In_10,In_347);
nor U1390 (N_1390,In_154,In_454);
and U1391 (N_1391,In_1326,In_1005);
nand U1392 (N_1392,In_1370,In_1358);
nor U1393 (N_1393,In_705,In_1086);
nand U1394 (N_1394,In_1168,In_423);
nand U1395 (N_1395,In_32,In_576);
or U1396 (N_1396,In_1482,In_162);
and U1397 (N_1397,In_1247,In_324);
and U1398 (N_1398,In_952,In_110);
nor U1399 (N_1399,In_700,In_1197);
nor U1400 (N_1400,In_1494,In_442);
nand U1401 (N_1401,In_1149,In_989);
xnor U1402 (N_1402,In_1083,In_467);
xor U1403 (N_1403,In_921,In_761);
or U1404 (N_1404,In_1148,In_840);
or U1405 (N_1405,In_741,In_1236);
nand U1406 (N_1406,In_35,In_938);
and U1407 (N_1407,In_106,In_1081);
or U1408 (N_1408,In_381,In_797);
xnor U1409 (N_1409,In_1400,In_1228);
and U1410 (N_1410,In_775,In_698);
xor U1411 (N_1411,In_594,In_739);
and U1412 (N_1412,In_752,In_1124);
nor U1413 (N_1413,In_1359,In_788);
nand U1414 (N_1414,In_58,In_957);
and U1415 (N_1415,In_667,In_1312);
nor U1416 (N_1416,In_121,In_575);
or U1417 (N_1417,In_1399,In_288);
or U1418 (N_1418,In_1050,In_48);
xor U1419 (N_1419,In_858,In_963);
nand U1420 (N_1420,In_274,In_195);
and U1421 (N_1421,In_275,In_777);
and U1422 (N_1422,In_1166,In_846);
nor U1423 (N_1423,In_699,In_645);
nor U1424 (N_1424,In_1099,In_1008);
xor U1425 (N_1425,In_609,In_358);
nand U1426 (N_1426,In_346,In_1320);
nor U1427 (N_1427,In_1368,In_717);
or U1428 (N_1428,In_293,In_24);
nand U1429 (N_1429,In_1278,In_1246);
and U1430 (N_1430,In_1139,In_66);
xnor U1431 (N_1431,In_998,In_460);
xnor U1432 (N_1432,In_710,In_812);
and U1433 (N_1433,In_1168,In_1396);
nand U1434 (N_1434,In_1262,In_743);
and U1435 (N_1435,In_127,In_1058);
nor U1436 (N_1436,In_115,In_129);
or U1437 (N_1437,In_892,In_301);
nand U1438 (N_1438,In_385,In_805);
nor U1439 (N_1439,In_712,In_1102);
or U1440 (N_1440,In_889,In_543);
and U1441 (N_1441,In_317,In_526);
xnor U1442 (N_1442,In_136,In_367);
xor U1443 (N_1443,In_494,In_853);
nand U1444 (N_1444,In_224,In_488);
or U1445 (N_1445,In_1432,In_29);
and U1446 (N_1446,In_1204,In_1065);
nor U1447 (N_1447,In_1064,In_58);
xnor U1448 (N_1448,In_692,In_107);
nor U1449 (N_1449,In_1011,In_671);
nand U1450 (N_1450,In_1347,In_118);
or U1451 (N_1451,In_1491,In_1146);
or U1452 (N_1452,In_534,In_877);
and U1453 (N_1453,In_1306,In_1333);
and U1454 (N_1454,In_1342,In_1018);
xnor U1455 (N_1455,In_213,In_551);
and U1456 (N_1456,In_156,In_58);
nand U1457 (N_1457,In_789,In_1234);
and U1458 (N_1458,In_970,In_908);
nand U1459 (N_1459,In_1202,In_1325);
nor U1460 (N_1460,In_717,In_1300);
nor U1461 (N_1461,In_794,In_1251);
and U1462 (N_1462,In_1050,In_1144);
and U1463 (N_1463,In_944,In_1377);
xor U1464 (N_1464,In_885,In_538);
nand U1465 (N_1465,In_980,In_492);
and U1466 (N_1466,In_908,In_852);
xor U1467 (N_1467,In_1353,In_1085);
nand U1468 (N_1468,In_921,In_535);
nand U1469 (N_1469,In_1209,In_926);
and U1470 (N_1470,In_574,In_253);
nand U1471 (N_1471,In_1413,In_745);
or U1472 (N_1472,In_986,In_352);
xor U1473 (N_1473,In_51,In_778);
nor U1474 (N_1474,In_1455,In_1035);
xor U1475 (N_1475,In_449,In_1325);
nor U1476 (N_1476,In_812,In_1394);
xnor U1477 (N_1477,In_762,In_479);
or U1478 (N_1478,In_836,In_338);
xor U1479 (N_1479,In_99,In_1202);
nand U1480 (N_1480,In_980,In_630);
xor U1481 (N_1481,In_921,In_287);
and U1482 (N_1482,In_993,In_13);
xor U1483 (N_1483,In_268,In_388);
or U1484 (N_1484,In_1440,In_1088);
and U1485 (N_1485,In_169,In_695);
and U1486 (N_1486,In_1369,In_563);
xnor U1487 (N_1487,In_207,In_138);
xor U1488 (N_1488,In_1158,In_924);
or U1489 (N_1489,In_1479,In_854);
and U1490 (N_1490,In_424,In_1018);
nand U1491 (N_1491,In_931,In_189);
nor U1492 (N_1492,In_168,In_173);
nand U1493 (N_1493,In_1141,In_129);
nand U1494 (N_1494,In_798,In_1499);
and U1495 (N_1495,In_55,In_962);
xor U1496 (N_1496,In_1085,In_405);
and U1497 (N_1497,In_26,In_611);
or U1498 (N_1498,In_1275,In_1284);
nor U1499 (N_1499,In_1049,In_343);
nand U1500 (N_1500,In_519,In_539);
or U1501 (N_1501,In_1273,In_1306);
or U1502 (N_1502,In_590,In_1484);
and U1503 (N_1503,In_234,In_1111);
nor U1504 (N_1504,In_1385,In_1016);
xor U1505 (N_1505,In_849,In_280);
or U1506 (N_1506,In_959,In_1106);
xnor U1507 (N_1507,In_254,In_1350);
or U1508 (N_1508,In_205,In_1000);
nor U1509 (N_1509,In_952,In_1288);
xor U1510 (N_1510,In_532,In_870);
nand U1511 (N_1511,In_1301,In_258);
nand U1512 (N_1512,In_664,In_549);
xor U1513 (N_1513,In_765,In_643);
nor U1514 (N_1514,In_1365,In_521);
nor U1515 (N_1515,In_785,In_757);
nand U1516 (N_1516,In_1269,In_160);
nand U1517 (N_1517,In_274,In_1027);
or U1518 (N_1518,In_790,In_767);
and U1519 (N_1519,In_1144,In_1499);
xnor U1520 (N_1520,In_1099,In_1259);
nor U1521 (N_1521,In_232,In_351);
or U1522 (N_1522,In_1281,In_175);
nor U1523 (N_1523,In_51,In_1260);
or U1524 (N_1524,In_269,In_413);
xnor U1525 (N_1525,In_69,In_732);
and U1526 (N_1526,In_1437,In_851);
xnor U1527 (N_1527,In_656,In_200);
nor U1528 (N_1528,In_394,In_1483);
nor U1529 (N_1529,In_1184,In_1253);
xnor U1530 (N_1530,In_208,In_637);
nor U1531 (N_1531,In_1191,In_1170);
nand U1532 (N_1532,In_937,In_1427);
nor U1533 (N_1533,In_35,In_1467);
xor U1534 (N_1534,In_679,In_1011);
nor U1535 (N_1535,In_1302,In_56);
or U1536 (N_1536,In_1270,In_663);
and U1537 (N_1537,In_479,In_736);
nand U1538 (N_1538,In_369,In_1099);
xor U1539 (N_1539,In_354,In_1092);
and U1540 (N_1540,In_315,In_1264);
and U1541 (N_1541,In_313,In_951);
nand U1542 (N_1542,In_208,In_515);
or U1543 (N_1543,In_34,In_1171);
and U1544 (N_1544,In_896,In_636);
nand U1545 (N_1545,In_393,In_92);
and U1546 (N_1546,In_788,In_1076);
or U1547 (N_1547,In_1449,In_345);
nand U1548 (N_1548,In_1079,In_364);
nor U1549 (N_1549,In_180,In_12);
and U1550 (N_1550,In_1293,In_426);
or U1551 (N_1551,In_199,In_747);
nor U1552 (N_1552,In_909,In_76);
and U1553 (N_1553,In_251,In_959);
or U1554 (N_1554,In_426,In_949);
nor U1555 (N_1555,In_550,In_889);
nor U1556 (N_1556,In_1191,In_1077);
nor U1557 (N_1557,In_1439,In_1230);
or U1558 (N_1558,In_785,In_1368);
and U1559 (N_1559,In_114,In_778);
nor U1560 (N_1560,In_150,In_1115);
and U1561 (N_1561,In_564,In_515);
xnor U1562 (N_1562,In_204,In_1246);
or U1563 (N_1563,In_232,In_1409);
nand U1564 (N_1564,In_807,In_211);
xnor U1565 (N_1565,In_166,In_536);
and U1566 (N_1566,In_852,In_1331);
nor U1567 (N_1567,In_1067,In_690);
or U1568 (N_1568,In_313,In_229);
nand U1569 (N_1569,In_542,In_1225);
xor U1570 (N_1570,In_907,In_1339);
or U1571 (N_1571,In_398,In_1467);
nor U1572 (N_1572,In_1011,In_702);
nand U1573 (N_1573,In_1358,In_205);
and U1574 (N_1574,In_239,In_50);
nand U1575 (N_1575,In_863,In_127);
nand U1576 (N_1576,In_1333,In_1002);
nand U1577 (N_1577,In_444,In_1113);
or U1578 (N_1578,In_1137,In_902);
nand U1579 (N_1579,In_498,In_68);
and U1580 (N_1580,In_1414,In_949);
xor U1581 (N_1581,In_1233,In_1075);
nand U1582 (N_1582,In_334,In_644);
or U1583 (N_1583,In_30,In_912);
nand U1584 (N_1584,In_825,In_143);
and U1585 (N_1585,In_957,In_786);
and U1586 (N_1586,In_1229,In_597);
nand U1587 (N_1587,In_1228,In_702);
nand U1588 (N_1588,In_523,In_778);
nand U1589 (N_1589,In_1320,In_64);
xnor U1590 (N_1590,In_1285,In_549);
nand U1591 (N_1591,In_1092,In_833);
or U1592 (N_1592,In_1307,In_728);
or U1593 (N_1593,In_513,In_1300);
xor U1594 (N_1594,In_93,In_504);
nor U1595 (N_1595,In_807,In_771);
nor U1596 (N_1596,In_812,In_390);
and U1597 (N_1597,In_1065,In_1449);
xor U1598 (N_1598,In_841,In_673);
nand U1599 (N_1599,In_404,In_1060);
xor U1600 (N_1600,In_1015,In_73);
xor U1601 (N_1601,In_1128,In_383);
or U1602 (N_1602,In_943,In_609);
nor U1603 (N_1603,In_107,In_1083);
or U1604 (N_1604,In_523,In_588);
and U1605 (N_1605,In_1293,In_220);
nand U1606 (N_1606,In_632,In_216);
or U1607 (N_1607,In_517,In_701);
or U1608 (N_1608,In_471,In_1010);
nor U1609 (N_1609,In_1387,In_918);
nand U1610 (N_1610,In_65,In_1411);
nor U1611 (N_1611,In_925,In_732);
and U1612 (N_1612,In_94,In_714);
or U1613 (N_1613,In_1464,In_177);
or U1614 (N_1614,In_847,In_848);
and U1615 (N_1615,In_1134,In_805);
nor U1616 (N_1616,In_580,In_735);
or U1617 (N_1617,In_581,In_977);
xor U1618 (N_1618,In_885,In_26);
and U1619 (N_1619,In_1447,In_1268);
nor U1620 (N_1620,In_647,In_819);
xor U1621 (N_1621,In_1157,In_1375);
nand U1622 (N_1622,In_1249,In_542);
nand U1623 (N_1623,In_878,In_1085);
nor U1624 (N_1624,In_916,In_134);
xnor U1625 (N_1625,In_41,In_1497);
nand U1626 (N_1626,In_195,In_1071);
xnor U1627 (N_1627,In_1227,In_401);
nor U1628 (N_1628,In_46,In_699);
xor U1629 (N_1629,In_856,In_254);
nand U1630 (N_1630,In_113,In_803);
or U1631 (N_1631,In_697,In_366);
nand U1632 (N_1632,In_148,In_8);
nand U1633 (N_1633,In_1491,In_864);
xnor U1634 (N_1634,In_104,In_1298);
or U1635 (N_1635,In_1192,In_445);
and U1636 (N_1636,In_1185,In_1004);
xnor U1637 (N_1637,In_244,In_1007);
or U1638 (N_1638,In_434,In_937);
nand U1639 (N_1639,In_184,In_432);
nand U1640 (N_1640,In_1305,In_278);
and U1641 (N_1641,In_1063,In_1033);
xor U1642 (N_1642,In_1457,In_1393);
and U1643 (N_1643,In_1480,In_1117);
and U1644 (N_1644,In_954,In_616);
and U1645 (N_1645,In_865,In_572);
nand U1646 (N_1646,In_768,In_556);
nor U1647 (N_1647,In_1144,In_65);
or U1648 (N_1648,In_547,In_433);
xnor U1649 (N_1649,In_793,In_581);
and U1650 (N_1650,In_969,In_192);
and U1651 (N_1651,In_306,In_1289);
and U1652 (N_1652,In_1245,In_401);
xnor U1653 (N_1653,In_1299,In_597);
nor U1654 (N_1654,In_715,In_1408);
nand U1655 (N_1655,In_7,In_707);
and U1656 (N_1656,In_949,In_1235);
xor U1657 (N_1657,In_1061,In_1171);
nand U1658 (N_1658,In_936,In_145);
xnor U1659 (N_1659,In_900,In_467);
xor U1660 (N_1660,In_981,In_531);
nand U1661 (N_1661,In_712,In_481);
nand U1662 (N_1662,In_1387,In_1353);
nor U1663 (N_1663,In_4,In_1287);
and U1664 (N_1664,In_263,In_1283);
or U1665 (N_1665,In_1466,In_44);
or U1666 (N_1666,In_877,In_819);
or U1667 (N_1667,In_1432,In_568);
xor U1668 (N_1668,In_674,In_319);
or U1669 (N_1669,In_1045,In_698);
xor U1670 (N_1670,In_1360,In_49);
xor U1671 (N_1671,In_808,In_660);
and U1672 (N_1672,In_1271,In_1275);
and U1673 (N_1673,In_1458,In_1188);
and U1674 (N_1674,In_1275,In_1266);
or U1675 (N_1675,In_1120,In_1290);
or U1676 (N_1676,In_770,In_1305);
nand U1677 (N_1677,In_760,In_631);
or U1678 (N_1678,In_687,In_28);
nand U1679 (N_1679,In_507,In_79);
and U1680 (N_1680,In_399,In_737);
or U1681 (N_1681,In_629,In_238);
xnor U1682 (N_1682,In_402,In_708);
nand U1683 (N_1683,In_884,In_165);
nand U1684 (N_1684,In_100,In_1091);
nand U1685 (N_1685,In_512,In_1026);
xnor U1686 (N_1686,In_338,In_1195);
xor U1687 (N_1687,In_845,In_757);
nand U1688 (N_1688,In_298,In_609);
and U1689 (N_1689,In_1400,In_1372);
nor U1690 (N_1690,In_595,In_349);
or U1691 (N_1691,In_1378,In_562);
nand U1692 (N_1692,In_945,In_1327);
xor U1693 (N_1693,In_468,In_65);
nand U1694 (N_1694,In_1275,In_1436);
nand U1695 (N_1695,In_696,In_406);
and U1696 (N_1696,In_1123,In_1402);
and U1697 (N_1697,In_1443,In_466);
nor U1698 (N_1698,In_1003,In_783);
or U1699 (N_1699,In_1332,In_944);
and U1700 (N_1700,In_1156,In_1336);
xor U1701 (N_1701,In_1021,In_789);
nand U1702 (N_1702,In_832,In_256);
nand U1703 (N_1703,In_342,In_1054);
or U1704 (N_1704,In_156,In_669);
nand U1705 (N_1705,In_1163,In_557);
or U1706 (N_1706,In_1184,In_563);
or U1707 (N_1707,In_567,In_942);
xor U1708 (N_1708,In_865,In_795);
nor U1709 (N_1709,In_1228,In_1107);
or U1710 (N_1710,In_774,In_151);
nand U1711 (N_1711,In_26,In_531);
nor U1712 (N_1712,In_1417,In_442);
xnor U1713 (N_1713,In_998,In_1145);
nor U1714 (N_1714,In_841,In_190);
nor U1715 (N_1715,In_789,In_1051);
xnor U1716 (N_1716,In_1264,In_1150);
nor U1717 (N_1717,In_41,In_850);
nor U1718 (N_1718,In_388,In_178);
and U1719 (N_1719,In_735,In_710);
xnor U1720 (N_1720,In_133,In_466);
or U1721 (N_1721,In_626,In_589);
or U1722 (N_1722,In_1104,In_1085);
nor U1723 (N_1723,In_119,In_1359);
nor U1724 (N_1724,In_476,In_202);
and U1725 (N_1725,In_529,In_851);
and U1726 (N_1726,In_1252,In_753);
nand U1727 (N_1727,In_1192,In_485);
xnor U1728 (N_1728,In_296,In_1358);
nor U1729 (N_1729,In_787,In_1143);
and U1730 (N_1730,In_812,In_1240);
nor U1731 (N_1731,In_99,In_283);
and U1732 (N_1732,In_421,In_829);
or U1733 (N_1733,In_1133,In_1450);
nand U1734 (N_1734,In_584,In_1034);
xor U1735 (N_1735,In_542,In_1078);
xnor U1736 (N_1736,In_383,In_1092);
xnor U1737 (N_1737,In_767,In_879);
xnor U1738 (N_1738,In_991,In_424);
nand U1739 (N_1739,In_1221,In_1219);
nor U1740 (N_1740,In_501,In_639);
nor U1741 (N_1741,In_647,In_277);
or U1742 (N_1742,In_528,In_413);
or U1743 (N_1743,In_850,In_559);
nor U1744 (N_1744,In_12,In_1441);
nor U1745 (N_1745,In_633,In_460);
xor U1746 (N_1746,In_1128,In_1493);
or U1747 (N_1747,In_1448,In_881);
xnor U1748 (N_1748,In_952,In_1419);
nand U1749 (N_1749,In_385,In_790);
and U1750 (N_1750,In_563,In_330);
nor U1751 (N_1751,In_609,In_1066);
nor U1752 (N_1752,In_1274,In_204);
or U1753 (N_1753,In_648,In_185);
and U1754 (N_1754,In_61,In_1311);
xor U1755 (N_1755,In_1344,In_552);
nor U1756 (N_1756,In_224,In_799);
nand U1757 (N_1757,In_929,In_282);
or U1758 (N_1758,In_771,In_1188);
nand U1759 (N_1759,In_1303,In_1134);
nand U1760 (N_1760,In_290,In_611);
nor U1761 (N_1761,In_259,In_925);
xor U1762 (N_1762,In_109,In_120);
xor U1763 (N_1763,In_1322,In_916);
xor U1764 (N_1764,In_1496,In_1214);
or U1765 (N_1765,In_1014,In_11);
nor U1766 (N_1766,In_1366,In_121);
nand U1767 (N_1767,In_6,In_1463);
nor U1768 (N_1768,In_999,In_208);
and U1769 (N_1769,In_732,In_300);
nor U1770 (N_1770,In_1451,In_1008);
nor U1771 (N_1771,In_613,In_779);
and U1772 (N_1772,In_1364,In_1223);
nor U1773 (N_1773,In_3,In_1088);
or U1774 (N_1774,In_142,In_623);
nor U1775 (N_1775,In_757,In_423);
and U1776 (N_1776,In_1160,In_165);
xnor U1777 (N_1777,In_842,In_843);
xnor U1778 (N_1778,In_634,In_604);
xor U1779 (N_1779,In_1438,In_92);
or U1780 (N_1780,In_1256,In_284);
or U1781 (N_1781,In_702,In_1199);
xor U1782 (N_1782,In_312,In_133);
nand U1783 (N_1783,In_891,In_487);
nor U1784 (N_1784,In_730,In_556);
nor U1785 (N_1785,In_868,In_1447);
xnor U1786 (N_1786,In_868,In_283);
xor U1787 (N_1787,In_1316,In_129);
or U1788 (N_1788,In_627,In_633);
and U1789 (N_1789,In_1188,In_1245);
and U1790 (N_1790,In_919,In_154);
or U1791 (N_1791,In_369,In_927);
xnor U1792 (N_1792,In_1443,In_836);
xor U1793 (N_1793,In_730,In_73);
or U1794 (N_1794,In_609,In_684);
nor U1795 (N_1795,In_260,In_650);
xnor U1796 (N_1796,In_519,In_735);
and U1797 (N_1797,In_445,In_101);
and U1798 (N_1798,In_702,In_83);
and U1799 (N_1799,In_132,In_714);
nand U1800 (N_1800,In_178,In_248);
and U1801 (N_1801,In_1172,In_174);
nor U1802 (N_1802,In_519,In_483);
nand U1803 (N_1803,In_647,In_207);
or U1804 (N_1804,In_1389,In_344);
nand U1805 (N_1805,In_791,In_960);
nand U1806 (N_1806,In_864,In_1403);
or U1807 (N_1807,In_574,In_698);
nand U1808 (N_1808,In_326,In_1101);
nor U1809 (N_1809,In_816,In_1460);
or U1810 (N_1810,In_698,In_1131);
or U1811 (N_1811,In_289,In_806);
xnor U1812 (N_1812,In_1366,In_881);
nor U1813 (N_1813,In_787,In_39);
nand U1814 (N_1814,In_69,In_1388);
and U1815 (N_1815,In_1075,In_999);
and U1816 (N_1816,In_803,In_78);
or U1817 (N_1817,In_491,In_1259);
xor U1818 (N_1818,In_362,In_1250);
nand U1819 (N_1819,In_466,In_1459);
or U1820 (N_1820,In_414,In_1446);
nor U1821 (N_1821,In_102,In_765);
xor U1822 (N_1822,In_533,In_1248);
or U1823 (N_1823,In_929,In_99);
nand U1824 (N_1824,In_700,In_515);
xor U1825 (N_1825,In_1393,In_954);
and U1826 (N_1826,In_165,In_682);
xor U1827 (N_1827,In_1315,In_1284);
nor U1828 (N_1828,In_1180,In_1302);
nand U1829 (N_1829,In_968,In_1164);
and U1830 (N_1830,In_392,In_51);
nor U1831 (N_1831,In_230,In_359);
and U1832 (N_1832,In_839,In_311);
nand U1833 (N_1833,In_1493,In_1250);
xor U1834 (N_1834,In_596,In_953);
xor U1835 (N_1835,In_910,In_487);
nand U1836 (N_1836,In_5,In_588);
and U1837 (N_1837,In_64,In_1264);
or U1838 (N_1838,In_1200,In_272);
and U1839 (N_1839,In_163,In_1081);
or U1840 (N_1840,In_384,In_764);
or U1841 (N_1841,In_96,In_1262);
nand U1842 (N_1842,In_387,In_346);
nor U1843 (N_1843,In_1280,In_129);
and U1844 (N_1844,In_832,In_123);
and U1845 (N_1845,In_1485,In_999);
xor U1846 (N_1846,In_1132,In_616);
nor U1847 (N_1847,In_1496,In_783);
nand U1848 (N_1848,In_480,In_824);
nor U1849 (N_1849,In_553,In_707);
or U1850 (N_1850,In_272,In_1299);
xnor U1851 (N_1851,In_968,In_269);
or U1852 (N_1852,In_748,In_273);
nor U1853 (N_1853,In_1017,In_157);
xnor U1854 (N_1854,In_131,In_1436);
and U1855 (N_1855,In_681,In_1208);
nor U1856 (N_1856,In_577,In_1421);
xor U1857 (N_1857,In_1155,In_254);
nand U1858 (N_1858,In_1348,In_391);
xor U1859 (N_1859,In_786,In_202);
nand U1860 (N_1860,In_262,In_727);
nor U1861 (N_1861,In_631,In_570);
nor U1862 (N_1862,In_615,In_1294);
nand U1863 (N_1863,In_964,In_1336);
nor U1864 (N_1864,In_987,In_1274);
nand U1865 (N_1865,In_1109,In_1007);
nor U1866 (N_1866,In_875,In_209);
nand U1867 (N_1867,In_10,In_1276);
nand U1868 (N_1868,In_1040,In_20);
nand U1869 (N_1869,In_1458,In_706);
and U1870 (N_1870,In_198,In_605);
or U1871 (N_1871,In_269,In_1002);
and U1872 (N_1872,In_468,In_152);
xor U1873 (N_1873,In_1127,In_785);
xnor U1874 (N_1874,In_842,In_1420);
and U1875 (N_1875,In_430,In_296);
nor U1876 (N_1876,In_172,In_286);
xnor U1877 (N_1877,In_209,In_927);
and U1878 (N_1878,In_1211,In_937);
nor U1879 (N_1879,In_1041,In_1121);
or U1880 (N_1880,In_700,In_47);
nor U1881 (N_1881,In_1060,In_102);
or U1882 (N_1882,In_85,In_95);
and U1883 (N_1883,In_916,In_1461);
and U1884 (N_1884,In_614,In_388);
xnor U1885 (N_1885,In_871,In_1485);
or U1886 (N_1886,In_1000,In_699);
nor U1887 (N_1887,In_236,In_108);
or U1888 (N_1888,In_661,In_600);
and U1889 (N_1889,In_439,In_1166);
nand U1890 (N_1890,In_101,In_695);
nor U1891 (N_1891,In_1441,In_210);
and U1892 (N_1892,In_800,In_1179);
nor U1893 (N_1893,In_1422,In_332);
nand U1894 (N_1894,In_959,In_1320);
xor U1895 (N_1895,In_196,In_174);
nand U1896 (N_1896,In_241,In_728);
xor U1897 (N_1897,In_542,In_804);
xor U1898 (N_1898,In_167,In_1392);
or U1899 (N_1899,In_1076,In_293);
and U1900 (N_1900,In_347,In_1250);
nor U1901 (N_1901,In_28,In_596);
xnor U1902 (N_1902,In_975,In_95);
nor U1903 (N_1903,In_641,In_1014);
and U1904 (N_1904,In_1127,In_711);
and U1905 (N_1905,In_678,In_806);
nand U1906 (N_1906,In_252,In_657);
and U1907 (N_1907,In_1381,In_306);
xor U1908 (N_1908,In_1305,In_1095);
nor U1909 (N_1909,In_471,In_1366);
and U1910 (N_1910,In_190,In_322);
nand U1911 (N_1911,In_660,In_838);
nor U1912 (N_1912,In_528,In_634);
nand U1913 (N_1913,In_1493,In_807);
and U1914 (N_1914,In_564,In_888);
and U1915 (N_1915,In_281,In_1288);
or U1916 (N_1916,In_298,In_237);
xnor U1917 (N_1917,In_1488,In_1070);
nand U1918 (N_1918,In_683,In_1416);
or U1919 (N_1919,In_119,In_1183);
nor U1920 (N_1920,In_1385,In_1338);
and U1921 (N_1921,In_988,In_1047);
or U1922 (N_1922,In_753,In_7);
or U1923 (N_1923,In_292,In_166);
or U1924 (N_1924,In_613,In_550);
or U1925 (N_1925,In_975,In_1322);
nor U1926 (N_1926,In_1052,In_293);
or U1927 (N_1927,In_1292,In_21);
nor U1928 (N_1928,In_875,In_436);
nor U1929 (N_1929,In_860,In_875);
nor U1930 (N_1930,In_307,In_432);
and U1931 (N_1931,In_1155,In_1015);
nor U1932 (N_1932,In_18,In_182);
and U1933 (N_1933,In_227,In_1102);
xor U1934 (N_1934,In_296,In_649);
and U1935 (N_1935,In_934,In_1035);
nor U1936 (N_1936,In_578,In_489);
or U1937 (N_1937,In_279,In_15);
nand U1938 (N_1938,In_968,In_551);
nand U1939 (N_1939,In_1253,In_126);
nand U1940 (N_1940,In_237,In_57);
nand U1941 (N_1941,In_719,In_341);
xor U1942 (N_1942,In_1063,In_1249);
xor U1943 (N_1943,In_891,In_1445);
and U1944 (N_1944,In_893,In_1055);
or U1945 (N_1945,In_1064,In_451);
xor U1946 (N_1946,In_166,In_1092);
nand U1947 (N_1947,In_590,In_1335);
and U1948 (N_1948,In_395,In_1107);
nand U1949 (N_1949,In_372,In_1180);
nand U1950 (N_1950,In_1266,In_295);
and U1951 (N_1951,In_777,In_36);
nor U1952 (N_1952,In_646,In_797);
and U1953 (N_1953,In_1406,In_89);
nor U1954 (N_1954,In_86,In_277);
or U1955 (N_1955,In_1077,In_136);
nand U1956 (N_1956,In_466,In_928);
nand U1957 (N_1957,In_1141,In_841);
and U1958 (N_1958,In_55,In_779);
or U1959 (N_1959,In_77,In_704);
and U1960 (N_1960,In_203,In_313);
or U1961 (N_1961,In_617,In_219);
or U1962 (N_1962,In_1301,In_1071);
and U1963 (N_1963,In_289,In_1157);
and U1964 (N_1964,In_518,In_546);
xor U1965 (N_1965,In_357,In_740);
nor U1966 (N_1966,In_1323,In_1278);
nand U1967 (N_1967,In_1111,In_1477);
and U1968 (N_1968,In_730,In_307);
xnor U1969 (N_1969,In_1369,In_353);
and U1970 (N_1970,In_1468,In_1261);
nor U1971 (N_1971,In_1292,In_1428);
nand U1972 (N_1972,In_1466,In_758);
nand U1973 (N_1973,In_1311,In_1389);
nor U1974 (N_1974,In_1182,In_608);
or U1975 (N_1975,In_1192,In_694);
xnor U1976 (N_1976,In_1161,In_549);
and U1977 (N_1977,In_113,In_1184);
and U1978 (N_1978,In_1462,In_927);
nor U1979 (N_1979,In_902,In_324);
nor U1980 (N_1980,In_1466,In_33);
xnor U1981 (N_1981,In_44,In_208);
nand U1982 (N_1982,In_1306,In_1111);
xor U1983 (N_1983,In_1109,In_1281);
nor U1984 (N_1984,In_1028,In_1130);
xor U1985 (N_1985,In_1391,In_81);
xnor U1986 (N_1986,In_966,In_488);
and U1987 (N_1987,In_1233,In_1299);
xor U1988 (N_1988,In_1084,In_545);
and U1989 (N_1989,In_1297,In_1262);
nand U1990 (N_1990,In_1009,In_275);
xor U1991 (N_1991,In_830,In_647);
nor U1992 (N_1992,In_382,In_177);
or U1993 (N_1993,In_74,In_725);
nor U1994 (N_1994,In_603,In_1105);
nand U1995 (N_1995,In_1467,In_1280);
nand U1996 (N_1996,In_277,In_106);
or U1997 (N_1997,In_747,In_824);
and U1998 (N_1998,In_653,In_1282);
nor U1999 (N_1999,In_249,In_316);
nand U2000 (N_2000,In_52,In_796);
nor U2001 (N_2001,In_659,In_842);
or U2002 (N_2002,In_1067,In_670);
xor U2003 (N_2003,In_1397,In_176);
nor U2004 (N_2004,In_715,In_628);
nor U2005 (N_2005,In_50,In_312);
xnor U2006 (N_2006,In_1191,In_781);
or U2007 (N_2007,In_48,In_546);
and U2008 (N_2008,In_1406,In_600);
nand U2009 (N_2009,In_1499,In_261);
nand U2010 (N_2010,In_287,In_520);
nand U2011 (N_2011,In_1326,In_409);
nand U2012 (N_2012,In_602,In_1026);
or U2013 (N_2013,In_210,In_1001);
nor U2014 (N_2014,In_384,In_359);
and U2015 (N_2015,In_1143,In_111);
and U2016 (N_2016,In_637,In_64);
nor U2017 (N_2017,In_1186,In_1159);
or U2018 (N_2018,In_326,In_790);
nand U2019 (N_2019,In_289,In_1472);
nor U2020 (N_2020,In_1030,In_159);
nor U2021 (N_2021,In_1338,In_1025);
or U2022 (N_2022,In_1035,In_1461);
or U2023 (N_2023,In_1360,In_899);
and U2024 (N_2024,In_1115,In_1111);
nor U2025 (N_2025,In_1132,In_1364);
xnor U2026 (N_2026,In_835,In_389);
xor U2027 (N_2027,In_16,In_108);
or U2028 (N_2028,In_180,In_1448);
nand U2029 (N_2029,In_1474,In_1175);
xnor U2030 (N_2030,In_916,In_152);
and U2031 (N_2031,In_1252,In_1148);
xnor U2032 (N_2032,In_612,In_1444);
or U2033 (N_2033,In_240,In_38);
xnor U2034 (N_2034,In_1202,In_1127);
nand U2035 (N_2035,In_539,In_790);
xnor U2036 (N_2036,In_1256,In_762);
and U2037 (N_2037,In_1252,In_841);
or U2038 (N_2038,In_1223,In_422);
and U2039 (N_2039,In_894,In_1154);
and U2040 (N_2040,In_733,In_391);
nand U2041 (N_2041,In_69,In_1462);
nor U2042 (N_2042,In_678,In_689);
and U2043 (N_2043,In_528,In_1020);
nand U2044 (N_2044,In_257,In_1007);
xnor U2045 (N_2045,In_305,In_1205);
nor U2046 (N_2046,In_1026,In_1412);
nand U2047 (N_2047,In_1241,In_379);
or U2048 (N_2048,In_1019,In_1284);
and U2049 (N_2049,In_820,In_338);
nand U2050 (N_2050,In_716,In_1486);
xor U2051 (N_2051,In_1263,In_561);
nor U2052 (N_2052,In_1122,In_172);
or U2053 (N_2053,In_556,In_963);
nor U2054 (N_2054,In_428,In_868);
and U2055 (N_2055,In_830,In_583);
nand U2056 (N_2056,In_689,In_764);
nor U2057 (N_2057,In_1356,In_1417);
or U2058 (N_2058,In_1212,In_58);
nand U2059 (N_2059,In_1467,In_1069);
or U2060 (N_2060,In_1027,In_906);
nor U2061 (N_2061,In_1491,In_46);
or U2062 (N_2062,In_908,In_914);
and U2063 (N_2063,In_1291,In_738);
nand U2064 (N_2064,In_479,In_1483);
nor U2065 (N_2065,In_1468,In_217);
nor U2066 (N_2066,In_1312,In_166);
or U2067 (N_2067,In_132,In_1095);
nand U2068 (N_2068,In_1356,In_188);
xor U2069 (N_2069,In_759,In_686);
xor U2070 (N_2070,In_48,In_74);
nor U2071 (N_2071,In_521,In_1209);
or U2072 (N_2072,In_836,In_1218);
or U2073 (N_2073,In_768,In_1078);
nand U2074 (N_2074,In_348,In_991);
xnor U2075 (N_2075,In_951,In_1326);
nor U2076 (N_2076,In_820,In_473);
or U2077 (N_2077,In_563,In_1173);
or U2078 (N_2078,In_311,In_1174);
or U2079 (N_2079,In_982,In_1109);
xnor U2080 (N_2080,In_129,In_767);
xor U2081 (N_2081,In_1329,In_1385);
or U2082 (N_2082,In_1158,In_805);
nor U2083 (N_2083,In_1296,In_972);
or U2084 (N_2084,In_1446,In_534);
nor U2085 (N_2085,In_469,In_1005);
and U2086 (N_2086,In_543,In_704);
nand U2087 (N_2087,In_724,In_1401);
nor U2088 (N_2088,In_377,In_0);
nor U2089 (N_2089,In_1119,In_638);
and U2090 (N_2090,In_482,In_399);
xnor U2091 (N_2091,In_726,In_554);
nor U2092 (N_2092,In_1258,In_367);
nand U2093 (N_2093,In_474,In_1324);
nand U2094 (N_2094,In_1082,In_1313);
nor U2095 (N_2095,In_503,In_631);
nor U2096 (N_2096,In_1060,In_809);
or U2097 (N_2097,In_1124,In_951);
xnor U2098 (N_2098,In_923,In_674);
nand U2099 (N_2099,In_260,In_141);
and U2100 (N_2100,In_202,In_103);
and U2101 (N_2101,In_312,In_1228);
xnor U2102 (N_2102,In_1072,In_1264);
nor U2103 (N_2103,In_288,In_243);
xnor U2104 (N_2104,In_82,In_1019);
nor U2105 (N_2105,In_1135,In_569);
nor U2106 (N_2106,In_366,In_1227);
and U2107 (N_2107,In_465,In_325);
nand U2108 (N_2108,In_1294,In_758);
and U2109 (N_2109,In_280,In_974);
nor U2110 (N_2110,In_479,In_1460);
xor U2111 (N_2111,In_202,In_1324);
or U2112 (N_2112,In_1118,In_313);
and U2113 (N_2113,In_1233,In_823);
nand U2114 (N_2114,In_108,In_254);
and U2115 (N_2115,In_1147,In_1314);
or U2116 (N_2116,In_101,In_370);
or U2117 (N_2117,In_395,In_1267);
and U2118 (N_2118,In_1141,In_126);
nand U2119 (N_2119,In_136,In_379);
and U2120 (N_2120,In_148,In_917);
nor U2121 (N_2121,In_1121,In_235);
xor U2122 (N_2122,In_911,In_640);
or U2123 (N_2123,In_240,In_990);
xor U2124 (N_2124,In_522,In_1149);
or U2125 (N_2125,In_942,In_868);
nand U2126 (N_2126,In_1364,In_1242);
and U2127 (N_2127,In_924,In_1210);
or U2128 (N_2128,In_688,In_539);
nand U2129 (N_2129,In_918,In_7);
nand U2130 (N_2130,In_1085,In_1207);
nor U2131 (N_2131,In_708,In_938);
and U2132 (N_2132,In_606,In_1082);
and U2133 (N_2133,In_1460,In_565);
nor U2134 (N_2134,In_895,In_729);
nor U2135 (N_2135,In_681,In_1360);
or U2136 (N_2136,In_993,In_401);
or U2137 (N_2137,In_116,In_1038);
xnor U2138 (N_2138,In_915,In_1076);
and U2139 (N_2139,In_661,In_68);
and U2140 (N_2140,In_383,In_1421);
and U2141 (N_2141,In_1452,In_236);
and U2142 (N_2142,In_740,In_819);
and U2143 (N_2143,In_183,In_1143);
nor U2144 (N_2144,In_626,In_509);
or U2145 (N_2145,In_898,In_958);
nor U2146 (N_2146,In_430,In_502);
nand U2147 (N_2147,In_829,In_462);
or U2148 (N_2148,In_1263,In_706);
nor U2149 (N_2149,In_451,In_629);
and U2150 (N_2150,In_1479,In_72);
nor U2151 (N_2151,In_572,In_807);
nor U2152 (N_2152,In_1008,In_51);
or U2153 (N_2153,In_1415,In_893);
nand U2154 (N_2154,In_973,In_57);
or U2155 (N_2155,In_1470,In_1033);
nor U2156 (N_2156,In_667,In_329);
nand U2157 (N_2157,In_18,In_239);
nand U2158 (N_2158,In_811,In_872);
or U2159 (N_2159,In_465,In_417);
nand U2160 (N_2160,In_677,In_458);
or U2161 (N_2161,In_1002,In_57);
and U2162 (N_2162,In_991,In_205);
and U2163 (N_2163,In_1021,In_175);
and U2164 (N_2164,In_551,In_1414);
nand U2165 (N_2165,In_702,In_1095);
or U2166 (N_2166,In_768,In_601);
nor U2167 (N_2167,In_753,In_10);
nor U2168 (N_2168,In_432,In_914);
or U2169 (N_2169,In_287,In_1065);
or U2170 (N_2170,In_765,In_207);
nand U2171 (N_2171,In_1236,In_27);
nor U2172 (N_2172,In_1491,In_1338);
xnor U2173 (N_2173,In_960,In_155);
or U2174 (N_2174,In_1165,In_613);
nor U2175 (N_2175,In_1256,In_1065);
xor U2176 (N_2176,In_396,In_1270);
or U2177 (N_2177,In_1351,In_1420);
nor U2178 (N_2178,In_127,In_912);
and U2179 (N_2179,In_559,In_1037);
xnor U2180 (N_2180,In_275,In_662);
xnor U2181 (N_2181,In_165,In_473);
nand U2182 (N_2182,In_174,In_167);
nand U2183 (N_2183,In_355,In_410);
or U2184 (N_2184,In_590,In_206);
nand U2185 (N_2185,In_1104,In_1238);
nand U2186 (N_2186,In_100,In_754);
and U2187 (N_2187,In_502,In_1302);
or U2188 (N_2188,In_1251,In_111);
or U2189 (N_2189,In_941,In_220);
nor U2190 (N_2190,In_836,In_1174);
nor U2191 (N_2191,In_1381,In_628);
xnor U2192 (N_2192,In_18,In_1403);
nand U2193 (N_2193,In_694,In_652);
and U2194 (N_2194,In_496,In_432);
or U2195 (N_2195,In_275,In_478);
and U2196 (N_2196,In_345,In_838);
xor U2197 (N_2197,In_365,In_1055);
xor U2198 (N_2198,In_177,In_915);
nor U2199 (N_2199,In_1263,In_77);
nor U2200 (N_2200,In_561,In_489);
or U2201 (N_2201,In_1376,In_562);
nor U2202 (N_2202,In_518,In_644);
xnor U2203 (N_2203,In_974,In_73);
or U2204 (N_2204,In_1159,In_178);
and U2205 (N_2205,In_370,In_41);
nand U2206 (N_2206,In_1456,In_620);
and U2207 (N_2207,In_832,In_306);
and U2208 (N_2208,In_256,In_1456);
nand U2209 (N_2209,In_164,In_906);
nand U2210 (N_2210,In_971,In_415);
nand U2211 (N_2211,In_1132,In_1134);
nor U2212 (N_2212,In_206,In_184);
xnor U2213 (N_2213,In_1422,In_1169);
or U2214 (N_2214,In_560,In_195);
and U2215 (N_2215,In_1290,In_931);
and U2216 (N_2216,In_728,In_527);
nor U2217 (N_2217,In_429,In_804);
nor U2218 (N_2218,In_626,In_937);
and U2219 (N_2219,In_699,In_1174);
or U2220 (N_2220,In_16,In_728);
nand U2221 (N_2221,In_688,In_133);
nand U2222 (N_2222,In_208,In_31);
nand U2223 (N_2223,In_31,In_1468);
nor U2224 (N_2224,In_178,In_24);
xor U2225 (N_2225,In_1096,In_49);
and U2226 (N_2226,In_565,In_890);
and U2227 (N_2227,In_271,In_1280);
and U2228 (N_2228,In_1210,In_313);
or U2229 (N_2229,In_802,In_402);
or U2230 (N_2230,In_1291,In_1410);
nor U2231 (N_2231,In_1235,In_826);
and U2232 (N_2232,In_1123,In_598);
nor U2233 (N_2233,In_735,In_220);
xor U2234 (N_2234,In_1447,In_152);
nor U2235 (N_2235,In_1131,In_534);
nor U2236 (N_2236,In_1225,In_269);
or U2237 (N_2237,In_220,In_655);
or U2238 (N_2238,In_206,In_380);
nand U2239 (N_2239,In_287,In_1295);
or U2240 (N_2240,In_981,In_523);
nor U2241 (N_2241,In_1146,In_229);
xor U2242 (N_2242,In_648,In_1216);
nand U2243 (N_2243,In_397,In_315);
xor U2244 (N_2244,In_201,In_607);
nor U2245 (N_2245,In_544,In_1027);
nand U2246 (N_2246,In_1287,In_1134);
and U2247 (N_2247,In_1051,In_1267);
and U2248 (N_2248,In_248,In_1211);
or U2249 (N_2249,In_1280,In_337);
xor U2250 (N_2250,In_1022,In_888);
and U2251 (N_2251,In_572,In_1454);
or U2252 (N_2252,In_1347,In_546);
xnor U2253 (N_2253,In_1261,In_616);
nand U2254 (N_2254,In_1054,In_340);
xor U2255 (N_2255,In_114,In_330);
or U2256 (N_2256,In_175,In_904);
nor U2257 (N_2257,In_406,In_754);
nor U2258 (N_2258,In_1057,In_683);
xor U2259 (N_2259,In_1078,In_277);
nand U2260 (N_2260,In_992,In_912);
xor U2261 (N_2261,In_1192,In_635);
or U2262 (N_2262,In_478,In_1249);
nand U2263 (N_2263,In_213,In_4);
xor U2264 (N_2264,In_1364,In_485);
nand U2265 (N_2265,In_1168,In_865);
xor U2266 (N_2266,In_1203,In_622);
and U2267 (N_2267,In_710,In_350);
and U2268 (N_2268,In_1190,In_491);
nor U2269 (N_2269,In_1214,In_1468);
and U2270 (N_2270,In_765,In_189);
and U2271 (N_2271,In_206,In_68);
xor U2272 (N_2272,In_908,In_435);
or U2273 (N_2273,In_424,In_673);
or U2274 (N_2274,In_999,In_483);
nor U2275 (N_2275,In_42,In_656);
nor U2276 (N_2276,In_948,In_612);
nor U2277 (N_2277,In_1481,In_401);
nand U2278 (N_2278,In_184,In_980);
and U2279 (N_2279,In_1115,In_1280);
and U2280 (N_2280,In_1244,In_1239);
xor U2281 (N_2281,In_1314,In_90);
xnor U2282 (N_2282,In_1151,In_627);
or U2283 (N_2283,In_889,In_421);
and U2284 (N_2284,In_388,In_218);
and U2285 (N_2285,In_925,In_22);
nor U2286 (N_2286,In_223,In_671);
xor U2287 (N_2287,In_148,In_475);
xnor U2288 (N_2288,In_26,In_889);
nor U2289 (N_2289,In_97,In_1411);
nand U2290 (N_2290,In_1251,In_445);
nor U2291 (N_2291,In_165,In_900);
or U2292 (N_2292,In_209,In_1487);
nor U2293 (N_2293,In_777,In_319);
nand U2294 (N_2294,In_732,In_178);
or U2295 (N_2295,In_1239,In_626);
nor U2296 (N_2296,In_775,In_916);
xnor U2297 (N_2297,In_94,In_573);
or U2298 (N_2298,In_1419,In_781);
and U2299 (N_2299,In_517,In_1136);
and U2300 (N_2300,In_1300,In_971);
xnor U2301 (N_2301,In_141,In_1422);
and U2302 (N_2302,In_1302,In_1381);
nor U2303 (N_2303,In_500,In_491);
or U2304 (N_2304,In_1160,In_710);
and U2305 (N_2305,In_628,In_957);
nor U2306 (N_2306,In_785,In_197);
xor U2307 (N_2307,In_680,In_337);
or U2308 (N_2308,In_133,In_126);
and U2309 (N_2309,In_1365,In_659);
nor U2310 (N_2310,In_319,In_1495);
nand U2311 (N_2311,In_385,In_197);
nand U2312 (N_2312,In_1349,In_807);
or U2313 (N_2313,In_1038,In_163);
or U2314 (N_2314,In_1081,In_616);
or U2315 (N_2315,In_625,In_971);
xnor U2316 (N_2316,In_402,In_767);
or U2317 (N_2317,In_122,In_898);
nand U2318 (N_2318,In_304,In_1237);
xor U2319 (N_2319,In_311,In_1465);
nor U2320 (N_2320,In_74,In_1159);
and U2321 (N_2321,In_913,In_91);
xor U2322 (N_2322,In_294,In_598);
xnor U2323 (N_2323,In_1063,In_1262);
nand U2324 (N_2324,In_1121,In_698);
or U2325 (N_2325,In_76,In_687);
or U2326 (N_2326,In_1408,In_655);
nand U2327 (N_2327,In_695,In_83);
or U2328 (N_2328,In_629,In_1021);
nor U2329 (N_2329,In_972,In_286);
nor U2330 (N_2330,In_744,In_1453);
or U2331 (N_2331,In_782,In_657);
xor U2332 (N_2332,In_511,In_1153);
xnor U2333 (N_2333,In_207,In_10);
or U2334 (N_2334,In_1101,In_1179);
xor U2335 (N_2335,In_361,In_173);
nor U2336 (N_2336,In_1275,In_826);
and U2337 (N_2337,In_607,In_444);
nor U2338 (N_2338,In_96,In_736);
xnor U2339 (N_2339,In_277,In_469);
nand U2340 (N_2340,In_741,In_1438);
nor U2341 (N_2341,In_156,In_795);
nand U2342 (N_2342,In_136,In_1138);
nor U2343 (N_2343,In_1393,In_459);
nand U2344 (N_2344,In_1309,In_337);
nor U2345 (N_2345,In_1471,In_1189);
nor U2346 (N_2346,In_1374,In_707);
nor U2347 (N_2347,In_888,In_918);
nand U2348 (N_2348,In_727,In_967);
xnor U2349 (N_2349,In_1077,In_1296);
xnor U2350 (N_2350,In_1374,In_1414);
nor U2351 (N_2351,In_1019,In_1265);
nor U2352 (N_2352,In_1353,In_543);
nand U2353 (N_2353,In_1284,In_306);
or U2354 (N_2354,In_667,In_1255);
and U2355 (N_2355,In_224,In_116);
xnor U2356 (N_2356,In_156,In_559);
or U2357 (N_2357,In_6,In_1255);
and U2358 (N_2358,In_1208,In_912);
nand U2359 (N_2359,In_323,In_953);
and U2360 (N_2360,In_1089,In_103);
xor U2361 (N_2361,In_379,In_128);
or U2362 (N_2362,In_118,In_46);
xor U2363 (N_2363,In_248,In_827);
nand U2364 (N_2364,In_46,In_910);
xor U2365 (N_2365,In_140,In_751);
nand U2366 (N_2366,In_611,In_1040);
nor U2367 (N_2367,In_1331,In_1180);
nand U2368 (N_2368,In_1283,In_144);
xor U2369 (N_2369,In_1494,In_1124);
or U2370 (N_2370,In_915,In_1047);
nand U2371 (N_2371,In_852,In_97);
nand U2372 (N_2372,In_827,In_271);
and U2373 (N_2373,In_981,In_959);
and U2374 (N_2374,In_101,In_572);
xor U2375 (N_2375,In_215,In_1407);
or U2376 (N_2376,In_1091,In_332);
nand U2377 (N_2377,In_1092,In_1156);
or U2378 (N_2378,In_456,In_63);
xor U2379 (N_2379,In_217,In_442);
and U2380 (N_2380,In_846,In_79);
and U2381 (N_2381,In_382,In_1281);
nor U2382 (N_2382,In_154,In_1434);
nand U2383 (N_2383,In_1214,In_1296);
or U2384 (N_2384,In_1117,In_1249);
nor U2385 (N_2385,In_1167,In_1424);
xor U2386 (N_2386,In_447,In_902);
or U2387 (N_2387,In_56,In_72);
and U2388 (N_2388,In_1417,In_1252);
nand U2389 (N_2389,In_1404,In_444);
or U2390 (N_2390,In_666,In_398);
and U2391 (N_2391,In_939,In_474);
xor U2392 (N_2392,In_161,In_387);
nand U2393 (N_2393,In_1436,In_937);
xnor U2394 (N_2394,In_1399,In_1003);
xor U2395 (N_2395,In_1192,In_906);
or U2396 (N_2396,In_850,In_1458);
nor U2397 (N_2397,In_77,In_872);
nor U2398 (N_2398,In_1482,In_1247);
nor U2399 (N_2399,In_669,In_405);
and U2400 (N_2400,In_1498,In_1438);
xor U2401 (N_2401,In_663,In_923);
and U2402 (N_2402,In_674,In_1406);
xnor U2403 (N_2403,In_192,In_1027);
nand U2404 (N_2404,In_503,In_1215);
or U2405 (N_2405,In_251,In_534);
nor U2406 (N_2406,In_56,In_293);
nor U2407 (N_2407,In_270,In_435);
nand U2408 (N_2408,In_228,In_652);
or U2409 (N_2409,In_1457,In_283);
nand U2410 (N_2410,In_340,In_1245);
nor U2411 (N_2411,In_266,In_1380);
xnor U2412 (N_2412,In_1149,In_1346);
nand U2413 (N_2413,In_122,In_1146);
or U2414 (N_2414,In_281,In_117);
xor U2415 (N_2415,In_49,In_1150);
or U2416 (N_2416,In_141,In_1366);
xor U2417 (N_2417,In_1013,In_521);
nor U2418 (N_2418,In_1492,In_209);
xor U2419 (N_2419,In_1302,In_568);
nand U2420 (N_2420,In_1236,In_894);
xor U2421 (N_2421,In_1266,In_492);
and U2422 (N_2422,In_1082,In_377);
nand U2423 (N_2423,In_1184,In_746);
nand U2424 (N_2424,In_1034,In_1174);
nand U2425 (N_2425,In_69,In_1238);
xnor U2426 (N_2426,In_317,In_1315);
and U2427 (N_2427,In_1260,In_458);
nor U2428 (N_2428,In_490,In_167);
xnor U2429 (N_2429,In_286,In_1055);
and U2430 (N_2430,In_160,In_92);
xor U2431 (N_2431,In_632,In_553);
nand U2432 (N_2432,In_174,In_806);
or U2433 (N_2433,In_681,In_789);
and U2434 (N_2434,In_931,In_798);
xnor U2435 (N_2435,In_213,In_614);
nor U2436 (N_2436,In_619,In_498);
nor U2437 (N_2437,In_1201,In_1006);
nand U2438 (N_2438,In_867,In_392);
or U2439 (N_2439,In_1207,In_616);
nor U2440 (N_2440,In_701,In_709);
nor U2441 (N_2441,In_374,In_141);
or U2442 (N_2442,In_1070,In_1406);
nor U2443 (N_2443,In_742,In_1407);
xor U2444 (N_2444,In_498,In_985);
nor U2445 (N_2445,In_897,In_246);
xor U2446 (N_2446,In_562,In_1197);
nor U2447 (N_2447,In_1485,In_1099);
nor U2448 (N_2448,In_592,In_1307);
nor U2449 (N_2449,In_859,In_1176);
xnor U2450 (N_2450,In_732,In_1276);
and U2451 (N_2451,In_1064,In_321);
nand U2452 (N_2452,In_476,In_454);
or U2453 (N_2453,In_1464,In_606);
and U2454 (N_2454,In_645,In_320);
or U2455 (N_2455,In_27,In_1402);
and U2456 (N_2456,In_214,In_718);
or U2457 (N_2457,In_853,In_258);
nand U2458 (N_2458,In_867,In_821);
or U2459 (N_2459,In_1175,In_1062);
nor U2460 (N_2460,In_845,In_494);
xor U2461 (N_2461,In_248,In_1447);
nand U2462 (N_2462,In_506,In_841);
nand U2463 (N_2463,In_1383,In_630);
and U2464 (N_2464,In_654,In_368);
nand U2465 (N_2465,In_762,In_670);
and U2466 (N_2466,In_282,In_1040);
nor U2467 (N_2467,In_707,In_1280);
xnor U2468 (N_2468,In_798,In_1301);
nand U2469 (N_2469,In_29,In_412);
xnor U2470 (N_2470,In_755,In_287);
or U2471 (N_2471,In_1225,In_772);
nand U2472 (N_2472,In_840,In_383);
nand U2473 (N_2473,In_971,In_1056);
nand U2474 (N_2474,In_872,In_881);
nor U2475 (N_2475,In_263,In_1175);
or U2476 (N_2476,In_902,In_1224);
xor U2477 (N_2477,In_1415,In_418);
or U2478 (N_2478,In_1303,In_1367);
xor U2479 (N_2479,In_1060,In_577);
and U2480 (N_2480,In_1171,In_132);
and U2481 (N_2481,In_1077,In_537);
and U2482 (N_2482,In_61,In_122);
or U2483 (N_2483,In_8,In_777);
and U2484 (N_2484,In_1317,In_532);
xnor U2485 (N_2485,In_127,In_1066);
xor U2486 (N_2486,In_1371,In_233);
or U2487 (N_2487,In_801,In_845);
or U2488 (N_2488,In_688,In_1196);
or U2489 (N_2489,In_700,In_1194);
and U2490 (N_2490,In_744,In_102);
and U2491 (N_2491,In_945,In_1273);
nand U2492 (N_2492,In_648,In_361);
and U2493 (N_2493,In_1055,In_1427);
nor U2494 (N_2494,In_731,In_682);
nor U2495 (N_2495,In_1273,In_756);
xor U2496 (N_2496,In_319,In_504);
xor U2497 (N_2497,In_401,In_621);
xor U2498 (N_2498,In_130,In_715);
or U2499 (N_2499,In_1222,In_502);
or U2500 (N_2500,In_1184,In_847);
or U2501 (N_2501,In_1385,In_1331);
or U2502 (N_2502,In_557,In_1189);
xnor U2503 (N_2503,In_537,In_735);
or U2504 (N_2504,In_1052,In_50);
xor U2505 (N_2505,In_19,In_812);
or U2506 (N_2506,In_1153,In_774);
and U2507 (N_2507,In_828,In_347);
nor U2508 (N_2508,In_1452,In_477);
nand U2509 (N_2509,In_533,In_1106);
nand U2510 (N_2510,In_167,In_608);
xnor U2511 (N_2511,In_1251,In_1);
and U2512 (N_2512,In_280,In_362);
nor U2513 (N_2513,In_695,In_554);
xnor U2514 (N_2514,In_997,In_914);
or U2515 (N_2515,In_1466,In_992);
xnor U2516 (N_2516,In_79,In_235);
and U2517 (N_2517,In_204,In_214);
nor U2518 (N_2518,In_760,In_1042);
nor U2519 (N_2519,In_12,In_889);
nor U2520 (N_2520,In_161,In_1041);
nand U2521 (N_2521,In_200,In_1085);
nand U2522 (N_2522,In_253,In_1477);
and U2523 (N_2523,In_1358,In_1463);
or U2524 (N_2524,In_1037,In_1071);
and U2525 (N_2525,In_687,In_1102);
and U2526 (N_2526,In_1347,In_9);
or U2527 (N_2527,In_500,In_392);
xor U2528 (N_2528,In_1193,In_1004);
nor U2529 (N_2529,In_806,In_784);
xnor U2530 (N_2530,In_471,In_402);
and U2531 (N_2531,In_1086,In_738);
and U2532 (N_2532,In_604,In_1185);
and U2533 (N_2533,In_979,In_1076);
or U2534 (N_2534,In_290,In_1044);
or U2535 (N_2535,In_367,In_453);
and U2536 (N_2536,In_389,In_65);
and U2537 (N_2537,In_584,In_333);
and U2538 (N_2538,In_1448,In_226);
nand U2539 (N_2539,In_1227,In_965);
or U2540 (N_2540,In_569,In_87);
nand U2541 (N_2541,In_819,In_524);
xnor U2542 (N_2542,In_768,In_132);
and U2543 (N_2543,In_1059,In_1178);
xor U2544 (N_2544,In_281,In_1278);
and U2545 (N_2545,In_825,In_521);
or U2546 (N_2546,In_1353,In_317);
and U2547 (N_2547,In_881,In_1341);
nand U2548 (N_2548,In_1421,In_727);
nor U2549 (N_2549,In_302,In_512);
nand U2550 (N_2550,In_646,In_531);
nor U2551 (N_2551,In_894,In_53);
or U2552 (N_2552,In_827,In_1459);
and U2553 (N_2553,In_538,In_876);
and U2554 (N_2554,In_989,In_1340);
xnor U2555 (N_2555,In_1166,In_1248);
nor U2556 (N_2556,In_779,In_700);
or U2557 (N_2557,In_381,In_327);
xor U2558 (N_2558,In_1494,In_573);
xor U2559 (N_2559,In_735,In_843);
xor U2560 (N_2560,In_442,In_1110);
or U2561 (N_2561,In_512,In_1488);
nor U2562 (N_2562,In_1000,In_295);
nor U2563 (N_2563,In_777,In_269);
nor U2564 (N_2564,In_552,In_1195);
nor U2565 (N_2565,In_813,In_132);
xor U2566 (N_2566,In_486,In_749);
nand U2567 (N_2567,In_689,In_1145);
or U2568 (N_2568,In_324,In_1281);
or U2569 (N_2569,In_530,In_50);
nand U2570 (N_2570,In_904,In_1344);
nor U2571 (N_2571,In_813,In_736);
xnor U2572 (N_2572,In_1397,In_1319);
nor U2573 (N_2573,In_189,In_169);
or U2574 (N_2574,In_1178,In_1025);
xor U2575 (N_2575,In_380,In_217);
nand U2576 (N_2576,In_312,In_556);
or U2577 (N_2577,In_1122,In_417);
nand U2578 (N_2578,In_858,In_875);
nor U2579 (N_2579,In_1285,In_459);
and U2580 (N_2580,In_1422,In_1448);
and U2581 (N_2581,In_911,In_238);
and U2582 (N_2582,In_416,In_372);
and U2583 (N_2583,In_1498,In_621);
nor U2584 (N_2584,In_879,In_583);
nor U2585 (N_2585,In_721,In_310);
nor U2586 (N_2586,In_1392,In_625);
nor U2587 (N_2587,In_1047,In_1150);
and U2588 (N_2588,In_546,In_1364);
xnor U2589 (N_2589,In_76,In_751);
nand U2590 (N_2590,In_403,In_466);
or U2591 (N_2591,In_1429,In_577);
or U2592 (N_2592,In_357,In_1265);
xor U2593 (N_2593,In_32,In_1181);
xor U2594 (N_2594,In_17,In_1287);
nand U2595 (N_2595,In_1066,In_26);
and U2596 (N_2596,In_1295,In_1465);
nand U2597 (N_2597,In_941,In_422);
and U2598 (N_2598,In_1478,In_693);
xor U2599 (N_2599,In_1320,In_697);
nor U2600 (N_2600,In_507,In_993);
nand U2601 (N_2601,In_204,In_624);
or U2602 (N_2602,In_1180,In_1308);
or U2603 (N_2603,In_214,In_675);
nand U2604 (N_2604,In_116,In_1432);
nand U2605 (N_2605,In_515,In_1393);
nor U2606 (N_2606,In_1489,In_1194);
nand U2607 (N_2607,In_742,In_615);
or U2608 (N_2608,In_986,In_294);
and U2609 (N_2609,In_240,In_568);
or U2610 (N_2610,In_579,In_889);
nand U2611 (N_2611,In_236,In_1075);
nand U2612 (N_2612,In_930,In_384);
nor U2613 (N_2613,In_828,In_941);
nand U2614 (N_2614,In_308,In_543);
nand U2615 (N_2615,In_1467,In_124);
or U2616 (N_2616,In_779,In_1258);
nand U2617 (N_2617,In_462,In_1465);
xnor U2618 (N_2618,In_247,In_523);
nor U2619 (N_2619,In_265,In_782);
xnor U2620 (N_2620,In_1123,In_266);
or U2621 (N_2621,In_770,In_310);
and U2622 (N_2622,In_129,In_1446);
nor U2623 (N_2623,In_947,In_340);
and U2624 (N_2624,In_1384,In_1309);
nor U2625 (N_2625,In_68,In_939);
nand U2626 (N_2626,In_1366,In_1405);
nand U2627 (N_2627,In_666,In_701);
xor U2628 (N_2628,In_838,In_54);
nand U2629 (N_2629,In_1291,In_113);
and U2630 (N_2630,In_456,In_844);
nor U2631 (N_2631,In_1141,In_529);
nand U2632 (N_2632,In_1029,In_624);
nand U2633 (N_2633,In_778,In_188);
or U2634 (N_2634,In_911,In_681);
and U2635 (N_2635,In_10,In_561);
nor U2636 (N_2636,In_596,In_714);
and U2637 (N_2637,In_1472,In_450);
nand U2638 (N_2638,In_1244,In_964);
nor U2639 (N_2639,In_926,In_692);
or U2640 (N_2640,In_1466,In_1195);
or U2641 (N_2641,In_251,In_1223);
nand U2642 (N_2642,In_834,In_123);
xor U2643 (N_2643,In_80,In_842);
and U2644 (N_2644,In_352,In_130);
nor U2645 (N_2645,In_985,In_179);
nand U2646 (N_2646,In_557,In_342);
or U2647 (N_2647,In_1148,In_1216);
nor U2648 (N_2648,In_369,In_638);
nor U2649 (N_2649,In_116,In_459);
nand U2650 (N_2650,In_1356,In_975);
nor U2651 (N_2651,In_752,In_1193);
nor U2652 (N_2652,In_304,In_309);
nor U2653 (N_2653,In_708,In_839);
nor U2654 (N_2654,In_485,In_1084);
nor U2655 (N_2655,In_367,In_12);
xnor U2656 (N_2656,In_1438,In_792);
nor U2657 (N_2657,In_1468,In_1325);
nand U2658 (N_2658,In_378,In_487);
nor U2659 (N_2659,In_724,In_950);
nand U2660 (N_2660,In_1490,In_999);
xor U2661 (N_2661,In_966,In_1223);
nor U2662 (N_2662,In_1003,In_912);
and U2663 (N_2663,In_1389,In_574);
and U2664 (N_2664,In_94,In_645);
and U2665 (N_2665,In_264,In_378);
xor U2666 (N_2666,In_1167,In_113);
nor U2667 (N_2667,In_308,In_913);
nand U2668 (N_2668,In_469,In_55);
or U2669 (N_2669,In_1347,In_717);
nand U2670 (N_2670,In_1163,In_339);
xor U2671 (N_2671,In_1025,In_51);
nand U2672 (N_2672,In_616,In_602);
nand U2673 (N_2673,In_608,In_1202);
nand U2674 (N_2674,In_23,In_813);
nor U2675 (N_2675,In_39,In_479);
or U2676 (N_2676,In_1062,In_926);
and U2677 (N_2677,In_196,In_1020);
or U2678 (N_2678,In_74,In_958);
nor U2679 (N_2679,In_939,In_543);
or U2680 (N_2680,In_254,In_780);
and U2681 (N_2681,In_751,In_203);
nand U2682 (N_2682,In_96,In_566);
or U2683 (N_2683,In_440,In_96);
or U2684 (N_2684,In_298,In_594);
or U2685 (N_2685,In_1149,In_218);
xor U2686 (N_2686,In_1109,In_849);
nor U2687 (N_2687,In_740,In_148);
or U2688 (N_2688,In_520,In_1317);
nor U2689 (N_2689,In_737,In_463);
and U2690 (N_2690,In_1413,In_880);
xnor U2691 (N_2691,In_1066,In_1073);
nand U2692 (N_2692,In_1474,In_150);
xor U2693 (N_2693,In_1426,In_522);
and U2694 (N_2694,In_1168,In_238);
nand U2695 (N_2695,In_458,In_1317);
and U2696 (N_2696,In_831,In_770);
nand U2697 (N_2697,In_83,In_1459);
xor U2698 (N_2698,In_69,In_365);
nand U2699 (N_2699,In_1421,In_908);
nand U2700 (N_2700,In_361,In_564);
or U2701 (N_2701,In_997,In_393);
nor U2702 (N_2702,In_635,In_1027);
xor U2703 (N_2703,In_167,In_248);
nand U2704 (N_2704,In_637,In_1354);
or U2705 (N_2705,In_258,In_779);
nand U2706 (N_2706,In_696,In_1355);
nand U2707 (N_2707,In_886,In_1402);
and U2708 (N_2708,In_1204,In_1160);
nor U2709 (N_2709,In_177,In_290);
nand U2710 (N_2710,In_1135,In_525);
xnor U2711 (N_2711,In_1355,In_593);
nand U2712 (N_2712,In_72,In_153);
nor U2713 (N_2713,In_94,In_795);
and U2714 (N_2714,In_1278,In_550);
or U2715 (N_2715,In_491,In_478);
xnor U2716 (N_2716,In_1370,In_356);
or U2717 (N_2717,In_693,In_740);
and U2718 (N_2718,In_360,In_383);
and U2719 (N_2719,In_430,In_1208);
nor U2720 (N_2720,In_752,In_972);
xnor U2721 (N_2721,In_186,In_352);
nand U2722 (N_2722,In_17,In_572);
and U2723 (N_2723,In_1473,In_689);
and U2724 (N_2724,In_1357,In_1238);
or U2725 (N_2725,In_197,In_1256);
or U2726 (N_2726,In_211,In_1410);
xnor U2727 (N_2727,In_388,In_404);
or U2728 (N_2728,In_94,In_262);
nor U2729 (N_2729,In_1033,In_410);
xor U2730 (N_2730,In_486,In_1089);
and U2731 (N_2731,In_1415,In_983);
or U2732 (N_2732,In_647,In_1106);
or U2733 (N_2733,In_1151,In_637);
xnor U2734 (N_2734,In_1483,In_1310);
xor U2735 (N_2735,In_109,In_1293);
and U2736 (N_2736,In_378,In_317);
nor U2737 (N_2737,In_75,In_524);
xor U2738 (N_2738,In_282,In_96);
and U2739 (N_2739,In_146,In_1298);
xor U2740 (N_2740,In_88,In_1225);
or U2741 (N_2741,In_580,In_550);
nand U2742 (N_2742,In_258,In_755);
and U2743 (N_2743,In_220,In_538);
nor U2744 (N_2744,In_187,In_1422);
nand U2745 (N_2745,In_88,In_177);
nand U2746 (N_2746,In_700,In_806);
or U2747 (N_2747,In_1357,In_9);
xor U2748 (N_2748,In_1370,In_1319);
nand U2749 (N_2749,In_669,In_826);
nand U2750 (N_2750,In_1453,In_363);
or U2751 (N_2751,In_1222,In_90);
and U2752 (N_2752,In_381,In_1354);
or U2753 (N_2753,In_674,In_26);
nand U2754 (N_2754,In_1357,In_319);
nor U2755 (N_2755,In_536,In_189);
nor U2756 (N_2756,In_455,In_976);
nor U2757 (N_2757,In_1421,In_418);
nor U2758 (N_2758,In_126,In_301);
nor U2759 (N_2759,In_469,In_47);
nor U2760 (N_2760,In_699,In_223);
nor U2761 (N_2761,In_843,In_603);
nor U2762 (N_2762,In_1002,In_1477);
nand U2763 (N_2763,In_1067,In_640);
nand U2764 (N_2764,In_658,In_959);
nor U2765 (N_2765,In_410,In_1370);
or U2766 (N_2766,In_1263,In_1129);
nor U2767 (N_2767,In_1477,In_802);
or U2768 (N_2768,In_919,In_194);
nand U2769 (N_2769,In_86,In_218);
or U2770 (N_2770,In_1225,In_173);
or U2771 (N_2771,In_877,In_1015);
nor U2772 (N_2772,In_1442,In_461);
xnor U2773 (N_2773,In_1465,In_695);
nand U2774 (N_2774,In_982,In_442);
nand U2775 (N_2775,In_220,In_21);
xnor U2776 (N_2776,In_532,In_1100);
and U2777 (N_2777,In_1455,In_236);
xor U2778 (N_2778,In_1368,In_350);
nor U2779 (N_2779,In_653,In_155);
xnor U2780 (N_2780,In_1055,In_1380);
and U2781 (N_2781,In_747,In_361);
and U2782 (N_2782,In_1286,In_1341);
xor U2783 (N_2783,In_295,In_630);
xnor U2784 (N_2784,In_1004,In_1382);
xor U2785 (N_2785,In_907,In_911);
xnor U2786 (N_2786,In_1099,In_257);
nor U2787 (N_2787,In_192,In_1277);
and U2788 (N_2788,In_1278,In_900);
nor U2789 (N_2789,In_565,In_362);
nor U2790 (N_2790,In_1464,In_971);
and U2791 (N_2791,In_904,In_1492);
or U2792 (N_2792,In_925,In_937);
xor U2793 (N_2793,In_562,In_282);
nor U2794 (N_2794,In_1044,In_490);
nor U2795 (N_2795,In_185,In_1159);
or U2796 (N_2796,In_64,In_374);
nand U2797 (N_2797,In_937,In_166);
and U2798 (N_2798,In_278,In_953);
nand U2799 (N_2799,In_1178,In_869);
nor U2800 (N_2800,In_334,In_1127);
nor U2801 (N_2801,In_255,In_104);
xnor U2802 (N_2802,In_184,In_1270);
or U2803 (N_2803,In_760,In_691);
or U2804 (N_2804,In_529,In_126);
and U2805 (N_2805,In_964,In_827);
and U2806 (N_2806,In_700,In_531);
nor U2807 (N_2807,In_6,In_940);
nor U2808 (N_2808,In_1121,In_1384);
xor U2809 (N_2809,In_1472,In_624);
xnor U2810 (N_2810,In_423,In_148);
and U2811 (N_2811,In_832,In_316);
or U2812 (N_2812,In_1477,In_71);
nor U2813 (N_2813,In_1217,In_891);
nand U2814 (N_2814,In_1075,In_1436);
nor U2815 (N_2815,In_1298,In_69);
and U2816 (N_2816,In_1397,In_164);
xor U2817 (N_2817,In_886,In_705);
nor U2818 (N_2818,In_1113,In_23);
nor U2819 (N_2819,In_191,In_489);
nand U2820 (N_2820,In_327,In_1458);
or U2821 (N_2821,In_515,In_290);
nor U2822 (N_2822,In_549,In_522);
nor U2823 (N_2823,In_221,In_1494);
and U2824 (N_2824,In_796,In_1105);
nor U2825 (N_2825,In_618,In_939);
xnor U2826 (N_2826,In_1130,In_1251);
or U2827 (N_2827,In_962,In_1259);
nor U2828 (N_2828,In_1448,In_1155);
or U2829 (N_2829,In_519,In_53);
or U2830 (N_2830,In_630,In_362);
nor U2831 (N_2831,In_964,In_694);
nor U2832 (N_2832,In_895,In_704);
xnor U2833 (N_2833,In_1133,In_290);
xor U2834 (N_2834,In_496,In_125);
xor U2835 (N_2835,In_866,In_1164);
nor U2836 (N_2836,In_802,In_717);
or U2837 (N_2837,In_260,In_1280);
xnor U2838 (N_2838,In_1438,In_1129);
nand U2839 (N_2839,In_558,In_352);
nand U2840 (N_2840,In_81,In_420);
nor U2841 (N_2841,In_967,In_1425);
and U2842 (N_2842,In_306,In_1174);
nor U2843 (N_2843,In_556,In_682);
nor U2844 (N_2844,In_345,In_1016);
nand U2845 (N_2845,In_1070,In_439);
or U2846 (N_2846,In_414,In_44);
nand U2847 (N_2847,In_1040,In_1213);
xnor U2848 (N_2848,In_992,In_701);
xor U2849 (N_2849,In_1243,In_1462);
and U2850 (N_2850,In_1374,In_868);
and U2851 (N_2851,In_707,In_291);
xor U2852 (N_2852,In_1463,In_1313);
and U2853 (N_2853,In_712,In_573);
and U2854 (N_2854,In_1299,In_739);
nor U2855 (N_2855,In_833,In_547);
or U2856 (N_2856,In_642,In_399);
nor U2857 (N_2857,In_1473,In_943);
nand U2858 (N_2858,In_950,In_1286);
nor U2859 (N_2859,In_1253,In_619);
xor U2860 (N_2860,In_1363,In_434);
nor U2861 (N_2861,In_322,In_117);
xnor U2862 (N_2862,In_1484,In_814);
xnor U2863 (N_2863,In_1416,In_952);
and U2864 (N_2864,In_426,In_771);
xnor U2865 (N_2865,In_836,In_1302);
xnor U2866 (N_2866,In_235,In_768);
nor U2867 (N_2867,In_1058,In_423);
and U2868 (N_2868,In_322,In_227);
xnor U2869 (N_2869,In_66,In_1061);
nand U2870 (N_2870,In_1084,In_620);
or U2871 (N_2871,In_655,In_1124);
nand U2872 (N_2872,In_690,In_1322);
xnor U2873 (N_2873,In_1350,In_161);
nand U2874 (N_2874,In_306,In_1319);
and U2875 (N_2875,In_662,In_43);
nor U2876 (N_2876,In_570,In_491);
nor U2877 (N_2877,In_35,In_542);
xor U2878 (N_2878,In_253,In_808);
or U2879 (N_2879,In_92,In_864);
xnor U2880 (N_2880,In_1381,In_48);
nand U2881 (N_2881,In_939,In_344);
and U2882 (N_2882,In_1136,In_811);
xor U2883 (N_2883,In_1483,In_475);
and U2884 (N_2884,In_749,In_1311);
xor U2885 (N_2885,In_951,In_269);
or U2886 (N_2886,In_216,In_273);
or U2887 (N_2887,In_519,In_768);
xor U2888 (N_2888,In_1451,In_371);
nor U2889 (N_2889,In_1314,In_107);
or U2890 (N_2890,In_603,In_670);
and U2891 (N_2891,In_1111,In_216);
or U2892 (N_2892,In_1419,In_956);
nand U2893 (N_2893,In_276,In_1449);
nand U2894 (N_2894,In_1215,In_849);
or U2895 (N_2895,In_757,In_395);
nand U2896 (N_2896,In_218,In_1490);
nand U2897 (N_2897,In_332,In_959);
or U2898 (N_2898,In_1277,In_629);
nor U2899 (N_2899,In_891,In_1446);
or U2900 (N_2900,In_1027,In_887);
or U2901 (N_2901,In_125,In_176);
nor U2902 (N_2902,In_1105,In_642);
and U2903 (N_2903,In_394,In_224);
nand U2904 (N_2904,In_532,In_604);
or U2905 (N_2905,In_884,In_1333);
nor U2906 (N_2906,In_134,In_1435);
nand U2907 (N_2907,In_1499,In_1284);
or U2908 (N_2908,In_142,In_851);
nor U2909 (N_2909,In_866,In_10);
or U2910 (N_2910,In_756,In_1071);
nand U2911 (N_2911,In_1391,In_179);
or U2912 (N_2912,In_192,In_894);
nor U2913 (N_2913,In_1059,In_1438);
xor U2914 (N_2914,In_824,In_933);
xnor U2915 (N_2915,In_122,In_645);
nand U2916 (N_2916,In_688,In_169);
nand U2917 (N_2917,In_662,In_8);
or U2918 (N_2918,In_471,In_848);
nor U2919 (N_2919,In_77,In_1095);
nand U2920 (N_2920,In_821,In_530);
xor U2921 (N_2921,In_1004,In_1167);
and U2922 (N_2922,In_1332,In_1461);
xor U2923 (N_2923,In_1208,In_1020);
and U2924 (N_2924,In_81,In_1173);
and U2925 (N_2925,In_333,In_278);
xnor U2926 (N_2926,In_321,In_1459);
and U2927 (N_2927,In_194,In_353);
xor U2928 (N_2928,In_1248,In_913);
nand U2929 (N_2929,In_357,In_231);
nor U2930 (N_2930,In_298,In_1455);
and U2931 (N_2931,In_1002,In_950);
nand U2932 (N_2932,In_837,In_1380);
and U2933 (N_2933,In_1186,In_55);
nor U2934 (N_2934,In_1499,In_193);
and U2935 (N_2935,In_1288,In_1221);
nand U2936 (N_2936,In_626,In_136);
and U2937 (N_2937,In_1372,In_888);
xor U2938 (N_2938,In_1495,In_793);
or U2939 (N_2939,In_1282,In_824);
nor U2940 (N_2940,In_719,In_50);
nand U2941 (N_2941,In_1466,In_486);
or U2942 (N_2942,In_768,In_49);
xor U2943 (N_2943,In_991,In_631);
or U2944 (N_2944,In_606,In_1432);
nor U2945 (N_2945,In_319,In_936);
nor U2946 (N_2946,In_171,In_1030);
or U2947 (N_2947,In_410,In_89);
xnor U2948 (N_2948,In_1361,In_278);
xnor U2949 (N_2949,In_727,In_144);
or U2950 (N_2950,In_673,In_1401);
nor U2951 (N_2951,In_263,In_1023);
nor U2952 (N_2952,In_1037,In_1214);
nand U2953 (N_2953,In_583,In_1024);
nand U2954 (N_2954,In_730,In_659);
nor U2955 (N_2955,In_972,In_1474);
xor U2956 (N_2956,In_1118,In_706);
and U2957 (N_2957,In_27,In_958);
or U2958 (N_2958,In_1112,In_513);
or U2959 (N_2959,In_1081,In_1156);
or U2960 (N_2960,In_315,In_737);
and U2961 (N_2961,In_1224,In_736);
or U2962 (N_2962,In_1329,In_736);
or U2963 (N_2963,In_924,In_416);
and U2964 (N_2964,In_1372,In_262);
and U2965 (N_2965,In_100,In_605);
and U2966 (N_2966,In_1434,In_262);
and U2967 (N_2967,In_1417,In_1461);
and U2968 (N_2968,In_1236,In_714);
nand U2969 (N_2969,In_1024,In_1268);
and U2970 (N_2970,In_1216,In_69);
or U2971 (N_2971,In_702,In_27);
nor U2972 (N_2972,In_1242,In_1174);
nor U2973 (N_2973,In_951,In_1108);
nor U2974 (N_2974,In_931,In_178);
nor U2975 (N_2975,In_33,In_1153);
xor U2976 (N_2976,In_350,In_479);
or U2977 (N_2977,In_79,In_602);
xnor U2978 (N_2978,In_24,In_346);
nand U2979 (N_2979,In_1400,In_1091);
nor U2980 (N_2980,In_604,In_508);
xor U2981 (N_2981,In_888,In_1166);
or U2982 (N_2982,In_817,In_1059);
or U2983 (N_2983,In_1457,In_984);
xor U2984 (N_2984,In_158,In_1283);
and U2985 (N_2985,In_484,In_877);
nand U2986 (N_2986,In_774,In_129);
nand U2987 (N_2987,In_705,In_168);
xnor U2988 (N_2988,In_105,In_16);
nand U2989 (N_2989,In_1109,In_676);
xor U2990 (N_2990,In_955,In_132);
nor U2991 (N_2991,In_475,In_404);
and U2992 (N_2992,In_56,In_724);
nor U2993 (N_2993,In_1265,In_3);
or U2994 (N_2994,In_580,In_999);
nand U2995 (N_2995,In_564,In_1497);
nor U2996 (N_2996,In_199,In_293);
xnor U2997 (N_2997,In_1284,In_826);
or U2998 (N_2998,In_740,In_784);
and U2999 (N_2999,In_1407,In_248);
nand U3000 (N_3000,In_846,In_1295);
and U3001 (N_3001,In_1113,In_1242);
nor U3002 (N_3002,In_1134,In_1373);
nand U3003 (N_3003,In_1334,In_1214);
xor U3004 (N_3004,In_812,In_993);
or U3005 (N_3005,In_261,In_832);
nand U3006 (N_3006,In_490,In_1093);
or U3007 (N_3007,In_232,In_205);
and U3008 (N_3008,In_1010,In_0);
nand U3009 (N_3009,In_1308,In_667);
nor U3010 (N_3010,In_830,In_300);
nor U3011 (N_3011,In_112,In_84);
nor U3012 (N_3012,In_186,In_890);
and U3013 (N_3013,In_624,In_38);
nand U3014 (N_3014,In_844,In_1167);
or U3015 (N_3015,In_1152,In_159);
xor U3016 (N_3016,In_1117,In_192);
or U3017 (N_3017,In_1407,In_1255);
nor U3018 (N_3018,In_1211,In_1036);
or U3019 (N_3019,In_908,In_424);
or U3020 (N_3020,In_702,In_577);
and U3021 (N_3021,In_339,In_286);
or U3022 (N_3022,In_716,In_106);
nand U3023 (N_3023,In_762,In_636);
xnor U3024 (N_3024,In_705,In_945);
or U3025 (N_3025,In_532,In_1187);
and U3026 (N_3026,In_1073,In_12);
and U3027 (N_3027,In_1453,In_365);
or U3028 (N_3028,In_230,In_351);
or U3029 (N_3029,In_198,In_1177);
or U3030 (N_3030,In_151,In_834);
nand U3031 (N_3031,In_828,In_1417);
nor U3032 (N_3032,In_802,In_1069);
or U3033 (N_3033,In_867,In_957);
or U3034 (N_3034,In_202,In_1381);
or U3035 (N_3035,In_270,In_1158);
and U3036 (N_3036,In_1422,In_356);
xnor U3037 (N_3037,In_1086,In_575);
and U3038 (N_3038,In_538,In_108);
and U3039 (N_3039,In_677,In_1369);
nand U3040 (N_3040,In_1151,In_368);
and U3041 (N_3041,In_810,In_1318);
nand U3042 (N_3042,In_1112,In_93);
nor U3043 (N_3043,In_394,In_321);
xnor U3044 (N_3044,In_149,In_520);
xor U3045 (N_3045,In_513,In_455);
or U3046 (N_3046,In_402,In_1116);
and U3047 (N_3047,In_429,In_773);
nor U3048 (N_3048,In_724,In_343);
nor U3049 (N_3049,In_1475,In_1318);
nand U3050 (N_3050,In_1155,In_635);
and U3051 (N_3051,In_1460,In_0);
xor U3052 (N_3052,In_1072,In_389);
or U3053 (N_3053,In_588,In_872);
nor U3054 (N_3054,In_178,In_1314);
xnor U3055 (N_3055,In_977,In_1202);
nor U3056 (N_3056,In_946,In_776);
or U3057 (N_3057,In_479,In_450);
nor U3058 (N_3058,In_464,In_674);
nand U3059 (N_3059,In_756,In_1445);
nand U3060 (N_3060,In_1137,In_911);
xor U3061 (N_3061,In_589,In_736);
xor U3062 (N_3062,In_91,In_1299);
nor U3063 (N_3063,In_1089,In_140);
or U3064 (N_3064,In_712,In_471);
nand U3065 (N_3065,In_92,In_1383);
nand U3066 (N_3066,In_1134,In_320);
nor U3067 (N_3067,In_81,In_928);
nand U3068 (N_3068,In_175,In_1084);
or U3069 (N_3069,In_726,In_1088);
or U3070 (N_3070,In_1476,In_1125);
or U3071 (N_3071,In_413,In_1332);
and U3072 (N_3072,In_1066,In_1356);
xnor U3073 (N_3073,In_996,In_432);
nand U3074 (N_3074,In_874,In_804);
nor U3075 (N_3075,In_773,In_1426);
nor U3076 (N_3076,In_133,In_241);
or U3077 (N_3077,In_897,In_1491);
or U3078 (N_3078,In_1109,In_48);
and U3079 (N_3079,In_584,In_1435);
or U3080 (N_3080,In_22,In_1243);
and U3081 (N_3081,In_428,In_545);
nor U3082 (N_3082,In_648,In_794);
nor U3083 (N_3083,In_73,In_796);
and U3084 (N_3084,In_425,In_645);
and U3085 (N_3085,In_58,In_234);
or U3086 (N_3086,In_259,In_1473);
and U3087 (N_3087,In_355,In_457);
nor U3088 (N_3088,In_1432,In_99);
xnor U3089 (N_3089,In_1421,In_142);
and U3090 (N_3090,In_1049,In_1224);
xor U3091 (N_3091,In_1087,In_501);
nor U3092 (N_3092,In_1383,In_1407);
and U3093 (N_3093,In_1414,In_14);
xnor U3094 (N_3094,In_417,In_555);
and U3095 (N_3095,In_384,In_281);
and U3096 (N_3096,In_1081,In_1159);
nor U3097 (N_3097,In_924,In_548);
and U3098 (N_3098,In_375,In_1336);
nand U3099 (N_3099,In_1454,In_1368);
and U3100 (N_3100,In_624,In_766);
nor U3101 (N_3101,In_1245,In_20);
and U3102 (N_3102,In_546,In_543);
and U3103 (N_3103,In_1092,In_530);
or U3104 (N_3104,In_1225,In_1146);
or U3105 (N_3105,In_864,In_348);
or U3106 (N_3106,In_1071,In_837);
and U3107 (N_3107,In_14,In_322);
nand U3108 (N_3108,In_1341,In_73);
nand U3109 (N_3109,In_597,In_1050);
nor U3110 (N_3110,In_569,In_952);
nand U3111 (N_3111,In_40,In_188);
nor U3112 (N_3112,In_1346,In_967);
xnor U3113 (N_3113,In_216,In_1314);
nand U3114 (N_3114,In_180,In_728);
nand U3115 (N_3115,In_364,In_1176);
xnor U3116 (N_3116,In_1371,In_1381);
nand U3117 (N_3117,In_105,In_1160);
xor U3118 (N_3118,In_721,In_70);
nor U3119 (N_3119,In_750,In_636);
nand U3120 (N_3120,In_875,In_842);
nor U3121 (N_3121,In_1190,In_1147);
xor U3122 (N_3122,In_828,In_1220);
nor U3123 (N_3123,In_181,In_300);
or U3124 (N_3124,In_1077,In_1195);
nand U3125 (N_3125,In_352,In_1114);
xnor U3126 (N_3126,In_496,In_874);
xnor U3127 (N_3127,In_684,In_1151);
xnor U3128 (N_3128,In_738,In_215);
and U3129 (N_3129,In_1279,In_1107);
and U3130 (N_3130,In_612,In_951);
and U3131 (N_3131,In_1054,In_1301);
nand U3132 (N_3132,In_1155,In_114);
nand U3133 (N_3133,In_624,In_1356);
or U3134 (N_3134,In_1314,In_766);
xnor U3135 (N_3135,In_85,In_693);
nor U3136 (N_3136,In_385,In_1462);
xor U3137 (N_3137,In_1067,In_11);
or U3138 (N_3138,In_440,In_126);
and U3139 (N_3139,In_864,In_1461);
and U3140 (N_3140,In_757,In_723);
nor U3141 (N_3141,In_53,In_222);
xnor U3142 (N_3142,In_1415,In_761);
or U3143 (N_3143,In_1148,In_1245);
and U3144 (N_3144,In_1129,In_1077);
and U3145 (N_3145,In_183,In_1286);
and U3146 (N_3146,In_1358,In_1395);
or U3147 (N_3147,In_1111,In_167);
xor U3148 (N_3148,In_1263,In_459);
nor U3149 (N_3149,In_1344,In_489);
and U3150 (N_3150,In_79,In_1253);
or U3151 (N_3151,In_118,In_16);
nand U3152 (N_3152,In_746,In_1414);
nand U3153 (N_3153,In_21,In_1404);
and U3154 (N_3154,In_69,In_186);
or U3155 (N_3155,In_228,In_559);
nor U3156 (N_3156,In_156,In_770);
xor U3157 (N_3157,In_1360,In_1312);
and U3158 (N_3158,In_1103,In_811);
nor U3159 (N_3159,In_1195,In_1481);
xnor U3160 (N_3160,In_1133,In_1401);
nor U3161 (N_3161,In_1405,In_65);
nor U3162 (N_3162,In_525,In_1209);
nor U3163 (N_3163,In_670,In_90);
or U3164 (N_3164,In_609,In_1148);
nand U3165 (N_3165,In_1449,In_594);
or U3166 (N_3166,In_1417,In_305);
or U3167 (N_3167,In_38,In_1104);
nand U3168 (N_3168,In_140,In_1166);
or U3169 (N_3169,In_336,In_1389);
or U3170 (N_3170,In_1221,In_1397);
nor U3171 (N_3171,In_206,In_245);
nand U3172 (N_3172,In_951,In_1060);
nand U3173 (N_3173,In_1337,In_643);
and U3174 (N_3174,In_1061,In_1203);
or U3175 (N_3175,In_425,In_595);
nor U3176 (N_3176,In_775,In_1066);
nand U3177 (N_3177,In_784,In_300);
xnor U3178 (N_3178,In_1040,In_285);
nor U3179 (N_3179,In_706,In_667);
or U3180 (N_3180,In_212,In_572);
nor U3181 (N_3181,In_461,In_1222);
or U3182 (N_3182,In_860,In_1211);
nand U3183 (N_3183,In_572,In_1054);
and U3184 (N_3184,In_719,In_364);
xor U3185 (N_3185,In_981,In_769);
or U3186 (N_3186,In_1292,In_658);
xnor U3187 (N_3187,In_1311,In_788);
xor U3188 (N_3188,In_1244,In_1472);
nor U3189 (N_3189,In_449,In_707);
and U3190 (N_3190,In_936,In_652);
nor U3191 (N_3191,In_514,In_994);
xnor U3192 (N_3192,In_1100,In_1482);
nand U3193 (N_3193,In_1312,In_66);
nor U3194 (N_3194,In_1122,In_1106);
nand U3195 (N_3195,In_552,In_888);
nand U3196 (N_3196,In_1429,In_1431);
nand U3197 (N_3197,In_1226,In_469);
and U3198 (N_3198,In_1160,In_609);
or U3199 (N_3199,In_1259,In_257);
xor U3200 (N_3200,In_390,In_243);
and U3201 (N_3201,In_1096,In_1256);
xor U3202 (N_3202,In_963,In_349);
nor U3203 (N_3203,In_167,In_251);
xor U3204 (N_3204,In_707,In_752);
and U3205 (N_3205,In_184,In_1347);
or U3206 (N_3206,In_691,In_1341);
nand U3207 (N_3207,In_18,In_911);
and U3208 (N_3208,In_1272,In_448);
and U3209 (N_3209,In_573,In_497);
nor U3210 (N_3210,In_487,In_1331);
and U3211 (N_3211,In_1053,In_365);
and U3212 (N_3212,In_1337,In_610);
nor U3213 (N_3213,In_238,In_135);
xor U3214 (N_3214,In_443,In_942);
and U3215 (N_3215,In_43,In_1254);
or U3216 (N_3216,In_1174,In_599);
or U3217 (N_3217,In_631,In_645);
nand U3218 (N_3218,In_68,In_1063);
nand U3219 (N_3219,In_138,In_192);
or U3220 (N_3220,In_1232,In_1053);
or U3221 (N_3221,In_786,In_159);
nand U3222 (N_3222,In_1026,In_593);
nor U3223 (N_3223,In_502,In_481);
xnor U3224 (N_3224,In_1253,In_305);
or U3225 (N_3225,In_664,In_706);
and U3226 (N_3226,In_1021,In_244);
nand U3227 (N_3227,In_648,In_157);
nand U3228 (N_3228,In_1086,In_1489);
or U3229 (N_3229,In_1302,In_1442);
nand U3230 (N_3230,In_1001,In_55);
and U3231 (N_3231,In_251,In_831);
nor U3232 (N_3232,In_453,In_863);
xnor U3233 (N_3233,In_933,In_105);
or U3234 (N_3234,In_1185,In_616);
or U3235 (N_3235,In_577,In_488);
xor U3236 (N_3236,In_1445,In_1107);
and U3237 (N_3237,In_1344,In_319);
xnor U3238 (N_3238,In_1481,In_143);
nand U3239 (N_3239,In_591,In_147);
or U3240 (N_3240,In_441,In_1311);
xor U3241 (N_3241,In_1192,In_861);
nand U3242 (N_3242,In_553,In_1179);
xor U3243 (N_3243,In_1112,In_467);
or U3244 (N_3244,In_1094,In_1125);
xnor U3245 (N_3245,In_711,In_838);
and U3246 (N_3246,In_849,In_156);
and U3247 (N_3247,In_53,In_544);
or U3248 (N_3248,In_645,In_1372);
xnor U3249 (N_3249,In_517,In_245);
xor U3250 (N_3250,In_1429,In_1384);
and U3251 (N_3251,In_904,In_803);
xnor U3252 (N_3252,In_1468,In_1274);
or U3253 (N_3253,In_1042,In_593);
nor U3254 (N_3254,In_758,In_702);
nand U3255 (N_3255,In_1185,In_982);
nor U3256 (N_3256,In_752,In_796);
or U3257 (N_3257,In_137,In_634);
nor U3258 (N_3258,In_125,In_214);
or U3259 (N_3259,In_38,In_9);
and U3260 (N_3260,In_1024,In_12);
or U3261 (N_3261,In_670,In_523);
nand U3262 (N_3262,In_545,In_1060);
or U3263 (N_3263,In_324,In_119);
nor U3264 (N_3264,In_973,In_327);
xnor U3265 (N_3265,In_696,In_1289);
or U3266 (N_3266,In_1440,In_1040);
xor U3267 (N_3267,In_854,In_917);
and U3268 (N_3268,In_789,In_239);
nor U3269 (N_3269,In_1199,In_588);
xnor U3270 (N_3270,In_520,In_1208);
or U3271 (N_3271,In_1460,In_5);
nand U3272 (N_3272,In_1291,In_575);
nand U3273 (N_3273,In_692,In_745);
or U3274 (N_3274,In_790,In_818);
nand U3275 (N_3275,In_994,In_141);
xnor U3276 (N_3276,In_878,In_843);
nand U3277 (N_3277,In_1388,In_1096);
xor U3278 (N_3278,In_229,In_327);
or U3279 (N_3279,In_888,In_180);
or U3280 (N_3280,In_615,In_61);
nand U3281 (N_3281,In_1168,In_279);
and U3282 (N_3282,In_418,In_1105);
nand U3283 (N_3283,In_506,In_449);
nor U3284 (N_3284,In_244,In_373);
xor U3285 (N_3285,In_1396,In_1467);
or U3286 (N_3286,In_860,In_797);
nand U3287 (N_3287,In_787,In_980);
or U3288 (N_3288,In_1453,In_340);
or U3289 (N_3289,In_366,In_367);
or U3290 (N_3290,In_1488,In_906);
nand U3291 (N_3291,In_1385,In_917);
and U3292 (N_3292,In_184,In_710);
nand U3293 (N_3293,In_987,In_1229);
nor U3294 (N_3294,In_77,In_113);
nor U3295 (N_3295,In_315,In_1031);
xnor U3296 (N_3296,In_1043,In_356);
nor U3297 (N_3297,In_837,In_506);
xor U3298 (N_3298,In_868,In_1371);
or U3299 (N_3299,In_919,In_744);
or U3300 (N_3300,In_432,In_266);
and U3301 (N_3301,In_994,In_645);
xor U3302 (N_3302,In_55,In_802);
nor U3303 (N_3303,In_657,In_586);
nand U3304 (N_3304,In_104,In_1491);
or U3305 (N_3305,In_118,In_927);
or U3306 (N_3306,In_831,In_1457);
or U3307 (N_3307,In_1486,In_1002);
or U3308 (N_3308,In_618,In_178);
or U3309 (N_3309,In_955,In_414);
nand U3310 (N_3310,In_423,In_1304);
nand U3311 (N_3311,In_763,In_775);
nand U3312 (N_3312,In_43,In_379);
nand U3313 (N_3313,In_1323,In_512);
nand U3314 (N_3314,In_921,In_813);
or U3315 (N_3315,In_87,In_957);
nand U3316 (N_3316,In_1410,In_1192);
xnor U3317 (N_3317,In_208,In_69);
and U3318 (N_3318,In_683,In_1408);
nand U3319 (N_3319,In_1063,In_444);
nor U3320 (N_3320,In_47,In_1223);
or U3321 (N_3321,In_1334,In_285);
or U3322 (N_3322,In_1491,In_1492);
nor U3323 (N_3323,In_1006,In_453);
xnor U3324 (N_3324,In_1380,In_999);
or U3325 (N_3325,In_24,In_902);
or U3326 (N_3326,In_1,In_823);
nand U3327 (N_3327,In_1229,In_1101);
or U3328 (N_3328,In_999,In_1098);
nor U3329 (N_3329,In_81,In_563);
xor U3330 (N_3330,In_1334,In_1375);
and U3331 (N_3331,In_1046,In_947);
and U3332 (N_3332,In_895,In_213);
nor U3333 (N_3333,In_16,In_581);
nor U3334 (N_3334,In_81,In_239);
nor U3335 (N_3335,In_1192,In_1317);
xor U3336 (N_3336,In_976,In_1052);
nor U3337 (N_3337,In_568,In_1085);
nand U3338 (N_3338,In_864,In_811);
and U3339 (N_3339,In_318,In_576);
nand U3340 (N_3340,In_758,In_454);
and U3341 (N_3341,In_92,In_7);
xnor U3342 (N_3342,In_719,In_5);
and U3343 (N_3343,In_1262,In_480);
nand U3344 (N_3344,In_886,In_1264);
nor U3345 (N_3345,In_861,In_985);
or U3346 (N_3346,In_198,In_801);
and U3347 (N_3347,In_831,In_1045);
or U3348 (N_3348,In_599,In_752);
or U3349 (N_3349,In_423,In_412);
or U3350 (N_3350,In_994,In_1297);
xnor U3351 (N_3351,In_427,In_952);
nor U3352 (N_3352,In_90,In_818);
nor U3353 (N_3353,In_1452,In_49);
xnor U3354 (N_3354,In_82,In_1320);
and U3355 (N_3355,In_1493,In_692);
nand U3356 (N_3356,In_1381,In_788);
nor U3357 (N_3357,In_93,In_519);
or U3358 (N_3358,In_1192,In_259);
nor U3359 (N_3359,In_895,In_436);
and U3360 (N_3360,In_866,In_435);
nor U3361 (N_3361,In_1278,In_1184);
xor U3362 (N_3362,In_124,In_590);
nand U3363 (N_3363,In_1208,In_636);
xor U3364 (N_3364,In_474,In_312);
xnor U3365 (N_3365,In_84,In_1495);
or U3366 (N_3366,In_860,In_32);
nor U3367 (N_3367,In_412,In_267);
nor U3368 (N_3368,In_1125,In_680);
and U3369 (N_3369,In_1225,In_1198);
and U3370 (N_3370,In_1296,In_1408);
nand U3371 (N_3371,In_870,In_6);
and U3372 (N_3372,In_245,In_680);
or U3373 (N_3373,In_558,In_1037);
or U3374 (N_3374,In_79,In_994);
xnor U3375 (N_3375,In_237,In_1487);
xnor U3376 (N_3376,In_885,In_60);
nand U3377 (N_3377,In_880,In_146);
xor U3378 (N_3378,In_79,In_1151);
or U3379 (N_3379,In_884,In_657);
xnor U3380 (N_3380,In_20,In_930);
xor U3381 (N_3381,In_627,In_339);
nand U3382 (N_3382,In_113,In_478);
or U3383 (N_3383,In_667,In_450);
or U3384 (N_3384,In_1008,In_37);
nand U3385 (N_3385,In_106,In_1299);
xnor U3386 (N_3386,In_967,In_142);
xnor U3387 (N_3387,In_60,In_695);
nand U3388 (N_3388,In_620,In_1467);
and U3389 (N_3389,In_1391,In_54);
xor U3390 (N_3390,In_837,In_154);
and U3391 (N_3391,In_619,In_185);
nand U3392 (N_3392,In_1252,In_1288);
nor U3393 (N_3393,In_570,In_774);
nor U3394 (N_3394,In_352,In_1081);
xor U3395 (N_3395,In_72,In_390);
xor U3396 (N_3396,In_1306,In_689);
nand U3397 (N_3397,In_1298,In_424);
and U3398 (N_3398,In_194,In_129);
nor U3399 (N_3399,In_202,In_1392);
nand U3400 (N_3400,In_175,In_1183);
and U3401 (N_3401,In_1060,In_281);
or U3402 (N_3402,In_1494,In_754);
and U3403 (N_3403,In_270,In_364);
nand U3404 (N_3404,In_1400,In_351);
nand U3405 (N_3405,In_1426,In_1038);
xnor U3406 (N_3406,In_666,In_530);
or U3407 (N_3407,In_463,In_230);
nor U3408 (N_3408,In_761,In_22);
or U3409 (N_3409,In_110,In_1166);
nand U3410 (N_3410,In_990,In_1339);
and U3411 (N_3411,In_620,In_222);
xnor U3412 (N_3412,In_1495,In_194);
nor U3413 (N_3413,In_536,In_1227);
nand U3414 (N_3414,In_734,In_299);
xor U3415 (N_3415,In_1104,In_928);
and U3416 (N_3416,In_1204,In_617);
nand U3417 (N_3417,In_65,In_125);
nand U3418 (N_3418,In_477,In_639);
and U3419 (N_3419,In_88,In_723);
xnor U3420 (N_3420,In_1232,In_733);
nor U3421 (N_3421,In_1037,In_1108);
and U3422 (N_3422,In_1352,In_1206);
and U3423 (N_3423,In_319,In_474);
or U3424 (N_3424,In_303,In_1236);
nand U3425 (N_3425,In_1214,In_1088);
or U3426 (N_3426,In_883,In_10);
and U3427 (N_3427,In_1083,In_1463);
nor U3428 (N_3428,In_110,In_973);
xnor U3429 (N_3429,In_765,In_1499);
xor U3430 (N_3430,In_79,In_301);
nor U3431 (N_3431,In_774,In_720);
nand U3432 (N_3432,In_119,In_674);
or U3433 (N_3433,In_74,In_1295);
nand U3434 (N_3434,In_1035,In_655);
xor U3435 (N_3435,In_1035,In_679);
and U3436 (N_3436,In_1307,In_1434);
and U3437 (N_3437,In_344,In_927);
xnor U3438 (N_3438,In_605,In_1179);
or U3439 (N_3439,In_1078,In_1046);
and U3440 (N_3440,In_777,In_135);
or U3441 (N_3441,In_1346,In_205);
xnor U3442 (N_3442,In_460,In_699);
or U3443 (N_3443,In_671,In_1230);
or U3444 (N_3444,In_1244,In_10);
nand U3445 (N_3445,In_647,In_701);
nor U3446 (N_3446,In_55,In_1452);
xnor U3447 (N_3447,In_1254,In_76);
nand U3448 (N_3448,In_567,In_333);
nor U3449 (N_3449,In_1104,In_304);
xor U3450 (N_3450,In_515,In_500);
and U3451 (N_3451,In_757,In_1176);
nor U3452 (N_3452,In_1385,In_351);
or U3453 (N_3453,In_293,In_569);
nor U3454 (N_3454,In_268,In_1291);
and U3455 (N_3455,In_1328,In_1166);
xnor U3456 (N_3456,In_474,In_1359);
nand U3457 (N_3457,In_1221,In_535);
nor U3458 (N_3458,In_646,In_168);
and U3459 (N_3459,In_805,In_378);
nand U3460 (N_3460,In_379,In_1287);
nor U3461 (N_3461,In_1186,In_558);
or U3462 (N_3462,In_62,In_1183);
xor U3463 (N_3463,In_1428,In_711);
and U3464 (N_3464,In_1490,In_1196);
or U3465 (N_3465,In_170,In_1403);
xor U3466 (N_3466,In_1445,In_1039);
or U3467 (N_3467,In_210,In_668);
xor U3468 (N_3468,In_511,In_278);
nor U3469 (N_3469,In_1070,In_433);
nor U3470 (N_3470,In_795,In_535);
nor U3471 (N_3471,In_1271,In_983);
nand U3472 (N_3472,In_655,In_616);
nor U3473 (N_3473,In_469,In_1223);
nand U3474 (N_3474,In_21,In_1314);
nand U3475 (N_3475,In_561,In_1069);
or U3476 (N_3476,In_226,In_364);
or U3477 (N_3477,In_1089,In_634);
or U3478 (N_3478,In_42,In_1271);
xor U3479 (N_3479,In_933,In_1261);
nand U3480 (N_3480,In_1471,In_496);
nand U3481 (N_3481,In_1257,In_842);
and U3482 (N_3482,In_1071,In_839);
and U3483 (N_3483,In_520,In_702);
nor U3484 (N_3484,In_893,In_1249);
or U3485 (N_3485,In_1413,In_416);
and U3486 (N_3486,In_1357,In_545);
and U3487 (N_3487,In_954,In_210);
xor U3488 (N_3488,In_122,In_795);
nand U3489 (N_3489,In_156,In_1492);
nand U3490 (N_3490,In_828,In_143);
nor U3491 (N_3491,In_906,In_11);
nor U3492 (N_3492,In_393,In_1085);
or U3493 (N_3493,In_1226,In_35);
nand U3494 (N_3494,In_1400,In_1135);
nand U3495 (N_3495,In_152,In_690);
xnor U3496 (N_3496,In_700,In_258);
nor U3497 (N_3497,In_1185,In_160);
or U3498 (N_3498,In_145,In_720);
nand U3499 (N_3499,In_1459,In_482);
or U3500 (N_3500,In_1382,In_736);
nor U3501 (N_3501,In_954,In_1272);
and U3502 (N_3502,In_1031,In_1406);
nor U3503 (N_3503,In_404,In_19);
xnor U3504 (N_3504,In_960,In_557);
xor U3505 (N_3505,In_74,In_966);
nand U3506 (N_3506,In_1442,In_1369);
and U3507 (N_3507,In_350,In_888);
nand U3508 (N_3508,In_416,In_1365);
and U3509 (N_3509,In_1470,In_101);
nor U3510 (N_3510,In_655,In_1498);
xor U3511 (N_3511,In_593,In_616);
nand U3512 (N_3512,In_25,In_182);
and U3513 (N_3513,In_99,In_789);
or U3514 (N_3514,In_110,In_127);
or U3515 (N_3515,In_595,In_1175);
nand U3516 (N_3516,In_1288,In_286);
and U3517 (N_3517,In_1308,In_121);
and U3518 (N_3518,In_1310,In_667);
nor U3519 (N_3519,In_1071,In_1056);
or U3520 (N_3520,In_6,In_171);
or U3521 (N_3521,In_1149,In_280);
nor U3522 (N_3522,In_60,In_867);
and U3523 (N_3523,In_663,In_1182);
xor U3524 (N_3524,In_990,In_1207);
nor U3525 (N_3525,In_770,In_253);
nand U3526 (N_3526,In_64,In_690);
nor U3527 (N_3527,In_246,In_1193);
nor U3528 (N_3528,In_960,In_1219);
nand U3529 (N_3529,In_850,In_624);
or U3530 (N_3530,In_1177,In_1260);
and U3531 (N_3531,In_1201,In_1092);
or U3532 (N_3532,In_713,In_1413);
xor U3533 (N_3533,In_752,In_862);
or U3534 (N_3534,In_484,In_624);
and U3535 (N_3535,In_1257,In_1441);
nor U3536 (N_3536,In_335,In_423);
and U3537 (N_3537,In_71,In_953);
or U3538 (N_3538,In_1321,In_788);
nand U3539 (N_3539,In_927,In_841);
or U3540 (N_3540,In_199,In_1222);
nand U3541 (N_3541,In_1262,In_1033);
xor U3542 (N_3542,In_1081,In_954);
xnor U3543 (N_3543,In_860,In_1430);
nor U3544 (N_3544,In_955,In_1199);
xnor U3545 (N_3545,In_1149,In_1021);
or U3546 (N_3546,In_444,In_295);
nor U3547 (N_3547,In_1051,In_1141);
or U3548 (N_3548,In_1332,In_1071);
or U3549 (N_3549,In_495,In_908);
or U3550 (N_3550,In_336,In_578);
xnor U3551 (N_3551,In_263,In_1062);
nor U3552 (N_3552,In_356,In_963);
nand U3553 (N_3553,In_1111,In_545);
or U3554 (N_3554,In_1366,In_1037);
and U3555 (N_3555,In_1377,In_463);
xor U3556 (N_3556,In_590,In_865);
or U3557 (N_3557,In_1323,In_604);
and U3558 (N_3558,In_944,In_1044);
nor U3559 (N_3559,In_1375,In_459);
or U3560 (N_3560,In_249,In_1233);
nand U3561 (N_3561,In_1252,In_176);
or U3562 (N_3562,In_1095,In_746);
nor U3563 (N_3563,In_397,In_1309);
or U3564 (N_3564,In_211,In_95);
or U3565 (N_3565,In_891,In_1320);
and U3566 (N_3566,In_448,In_1140);
nand U3567 (N_3567,In_156,In_1319);
nand U3568 (N_3568,In_1254,In_665);
nand U3569 (N_3569,In_640,In_93);
or U3570 (N_3570,In_329,In_482);
and U3571 (N_3571,In_935,In_327);
and U3572 (N_3572,In_431,In_140);
and U3573 (N_3573,In_644,In_1274);
and U3574 (N_3574,In_124,In_1489);
or U3575 (N_3575,In_111,In_525);
and U3576 (N_3576,In_752,In_302);
nand U3577 (N_3577,In_1297,In_1366);
nand U3578 (N_3578,In_129,In_87);
nor U3579 (N_3579,In_976,In_422);
nor U3580 (N_3580,In_801,In_745);
and U3581 (N_3581,In_164,In_1367);
and U3582 (N_3582,In_786,In_679);
nand U3583 (N_3583,In_909,In_1428);
nor U3584 (N_3584,In_736,In_1416);
or U3585 (N_3585,In_582,In_938);
and U3586 (N_3586,In_1198,In_289);
or U3587 (N_3587,In_11,In_14);
xor U3588 (N_3588,In_895,In_1009);
or U3589 (N_3589,In_939,In_1363);
or U3590 (N_3590,In_119,In_1020);
xor U3591 (N_3591,In_408,In_77);
xor U3592 (N_3592,In_633,In_467);
nand U3593 (N_3593,In_847,In_1407);
xor U3594 (N_3594,In_1384,In_1207);
xor U3595 (N_3595,In_826,In_847);
nor U3596 (N_3596,In_1338,In_956);
nand U3597 (N_3597,In_1435,In_1131);
xnor U3598 (N_3598,In_830,In_335);
nand U3599 (N_3599,In_386,In_554);
xor U3600 (N_3600,In_618,In_205);
xnor U3601 (N_3601,In_198,In_136);
xor U3602 (N_3602,In_69,In_1465);
nand U3603 (N_3603,In_814,In_264);
and U3604 (N_3604,In_752,In_136);
and U3605 (N_3605,In_1057,In_456);
nor U3606 (N_3606,In_1033,In_161);
or U3607 (N_3607,In_1381,In_16);
or U3608 (N_3608,In_555,In_542);
nor U3609 (N_3609,In_415,In_46);
xnor U3610 (N_3610,In_608,In_573);
or U3611 (N_3611,In_375,In_99);
and U3612 (N_3612,In_360,In_1432);
or U3613 (N_3613,In_1253,In_845);
and U3614 (N_3614,In_58,In_690);
nand U3615 (N_3615,In_140,In_97);
xnor U3616 (N_3616,In_1136,In_397);
or U3617 (N_3617,In_62,In_756);
and U3618 (N_3618,In_182,In_461);
nand U3619 (N_3619,In_699,In_915);
or U3620 (N_3620,In_1416,In_1257);
xnor U3621 (N_3621,In_605,In_1325);
or U3622 (N_3622,In_1193,In_146);
nor U3623 (N_3623,In_365,In_313);
and U3624 (N_3624,In_1059,In_203);
nor U3625 (N_3625,In_1476,In_1025);
and U3626 (N_3626,In_770,In_1316);
nor U3627 (N_3627,In_890,In_1022);
nand U3628 (N_3628,In_168,In_1186);
nor U3629 (N_3629,In_52,In_341);
xnor U3630 (N_3630,In_612,In_278);
nor U3631 (N_3631,In_925,In_844);
or U3632 (N_3632,In_800,In_1488);
nor U3633 (N_3633,In_999,In_570);
nand U3634 (N_3634,In_74,In_1443);
nor U3635 (N_3635,In_588,In_770);
xnor U3636 (N_3636,In_1183,In_800);
and U3637 (N_3637,In_148,In_1162);
or U3638 (N_3638,In_201,In_355);
or U3639 (N_3639,In_167,In_568);
and U3640 (N_3640,In_1271,In_436);
or U3641 (N_3641,In_989,In_832);
nand U3642 (N_3642,In_278,In_380);
and U3643 (N_3643,In_286,In_589);
nand U3644 (N_3644,In_1480,In_242);
nor U3645 (N_3645,In_62,In_1200);
or U3646 (N_3646,In_734,In_383);
xnor U3647 (N_3647,In_1441,In_217);
nor U3648 (N_3648,In_92,In_595);
or U3649 (N_3649,In_765,In_466);
nand U3650 (N_3650,In_712,In_959);
nand U3651 (N_3651,In_822,In_925);
nor U3652 (N_3652,In_1053,In_1400);
nand U3653 (N_3653,In_99,In_759);
nor U3654 (N_3654,In_123,In_1169);
xor U3655 (N_3655,In_1345,In_1346);
nor U3656 (N_3656,In_542,In_534);
nor U3657 (N_3657,In_1391,In_1084);
xor U3658 (N_3658,In_53,In_151);
xor U3659 (N_3659,In_783,In_79);
nand U3660 (N_3660,In_687,In_1380);
and U3661 (N_3661,In_1462,In_512);
or U3662 (N_3662,In_251,In_770);
and U3663 (N_3663,In_106,In_376);
and U3664 (N_3664,In_1478,In_730);
and U3665 (N_3665,In_237,In_606);
xor U3666 (N_3666,In_840,In_1413);
nor U3667 (N_3667,In_800,In_451);
or U3668 (N_3668,In_986,In_685);
nor U3669 (N_3669,In_943,In_1253);
nand U3670 (N_3670,In_1342,In_902);
and U3671 (N_3671,In_737,In_336);
or U3672 (N_3672,In_245,In_753);
xnor U3673 (N_3673,In_1200,In_562);
xnor U3674 (N_3674,In_663,In_1453);
and U3675 (N_3675,In_882,In_420);
nand U3676 (N_3676,In_53,In_1022);
nor U3677 (N_3677,In_457,In_1013);
nor U3678 (N_3678,In_1473,In_222);
and U3679 (N_3679,In_1225,In_390);
xor U3680 (N_3680,In_85,In_561);
xor U3681 (N_3681,In_761,In_212);
nor U3682 (N_3682,In_735,In_538);
and U3683 (N_3683,In_558,In_142);
or U3684 (N_3684,In_907,In_1019);
xor U3685 (N_3685,In_1491,In_367);
xnor U3686 (N_3686,In_789,In_1433);
and U3687 (N_3687,In_157,In_690);
or U3688 (N_3688,In_1452,In_1226);
nor U3689 (N_3689,In_1252,In_669);
or U3690 (N_3690,In_1125,In_2);
or U3691 (N_3691,In_946,In_768);
nand U3692 (N_3692,In_263,In_1124);
xor U3693 (N_3693,In_1284,In_759);
nand U3694 (N_3694,In_393,In_150);
xnor U3695 (N_3695,In_1415,In_1311);
or U3696 (N_3696,In_574,In_530);
and U3697 (N_3697,In_326,In_894);
and U3698 (N_3698,In_935,In_1066);
or U3699 (N_3699,In_3,In_1226);
nand U3700 (N_3700,In_503,In_26);
or U3701 (N_3701,In_1038,In_39);
xor U3702 (N_3702,In_1241,In_285);
and U3703 (N_3703,In_1316,In_398);
nand U3704 (N_3704,In_785,In_499);
xnor U3705 (N_3705,In_1189,In_1409);
nor U3706 (N_3706,In_168,In_1340);
nand U3707 (N_3707,In_1449,In_684);
or U3708 (N_3708,In_1278,In_972);
nand U3709 (N_3709,In_813,In_1428);
nand U3710 (N_3710,In_65,In_295);
xor U3711 (N_3711,In_709,In_963);
nor U3712 (N_3712,In_890,In_837);
xnor U3713 (N_3713,In_581,In_504);
or U3714 (N_3714,In_16,In_748);
nand U3715 (N_3715,In_401,In_351);
nand U3716 (N_3716,In_98,In_1286);
nand U3717 (N_3717,In_1417,In_1022);
and U3718 (N_3718,In_106,In_819);
nor U3719 (N_3719,In_693,In_1492);
and U3720 (N_3720,In_1482,In_986);
and U3721 (N_3721,In_936,In_800);
and U3722 (N_3722,In_489,In_1444);
xnor U3723 (N_3723,In_1306,In_1275);
or U3724 (N_3724,In_543,In_1249);
and U3725 (N_3725,In_883,In_550);
xnor U3726 (N_3726,In_1494,In_1439);
nor U3727 (N_3727,In_1445,In_1013);
nor U3728 (N_3728,In_1368,In_732);
nand U3729 (N_3729,In_93,In_460);
xnor U3730 (N_3730,In_1145,In_1462);
nand U3731 (N_3731,In_663,In_1446);
nand U3732 (N_3732,In_1297,In_1334);
nor U3733 (N_3733,In_152,In_319);
nor U3734 (N_3734,In_611,In_394);
xnor U3735 (N_3735,In_294,In_571);
xnor U3736 (N_3736,In_1092,In_214);
nor U3737 (N_3737,In_1002,In_94);
xor U3738 (N_3738,In_1168,In_1138);
or U3739 (N_3739,In_1114,In_589);
xnor U3740 (N_3740,In_7,In_421);
or U3741 (N_3741,In_246,In_201);
and U3742 (N_3742,In_896,In_227);
xnor U3743 (N_3743,In_1408,In_844);
xnor U3744 (N_3744,In_1492,In_926);
nor U3745 (N_3745,In_398,In_918);
xor U3746 (N_3746,In_299,In_650);
and U3747 (N_3747,In_1117,In_1495);
and U3748 (N_3748,In_959,In_979);
or U3749 (N_3749,In_1350,In_1482);
and U3750 (N_3750,In_547,In_554);
nand U3751 (N_3751,In_110,In_838);
or U3752 (N_3752,In_1302,In_155);
and U3753 (N_3753,In_1489,In_217);
nor U3754 (N_3754,In_341,In_787);
or U3755 (N_3755,In_1097,In_511);
and U3756 (N_3756,In_757,In_388);
or U3757 (N_3757,In_1076,In_1344);
xnor U3758 (N_3758,In_1423,In_617);
nand U3759 (N_3759,In_318,In_1349);
and U3760 (N_3760,In_708,In_1089);
and U3761 (N_3761,In_855,In_167);
xnor U3762 (N_3762,In_194,In_460);
nand U3763 (N_3763,In_1435,In_743);
nor U3764 (N_3764,In_1099,In_115);
nor U3765 (N_3765,In_1005,In_1335);
nor U3766 (N_3766,In_1260,In_809);
nand U3767 (N_3767,In_528,In_609);
or U3768 (N_3768,In_1220,In_46);
xnor U3769 (N_3769,In_380,In_856);
or U3770 (N_3770,In_1047,In_810);
nor U3771 (N_3771,In_733,In_1293);
nor U3772 (N_3772,In_1354,In_1196);
and U3773 (N_3773,In_1198,In_1177);
xnor U3774 (N_3774,In_1450,In_7);
nor U3775 (N_3775,In_323,In_996);
nand U3776 (N_3776,In_510,In_800);
nand U3777 (N_3777,In_691,In_927);
nand U3778 (N_3778,In_1222,In_1435);
xnor U3779 (N_3779,In_1051,In_317);
or U3780 (N_3780,In_1350,In_985);
xnor U3781 (N_3781,In_1278,In_1103);
nor U3782 (N_3782,In_908,In_655);
nor U3783 (N_3783,In_213,In_871);
and U3784 (N_3784,In_198,In_1073);
xor U3785 (N_3785,In_442,In_1047);
and U3786 (N_3786,In_291,In_370);
xor U3787 (N_3787,In_1391,In_1433);
nor U3788 (N_3788,In_1467,In_785);
nor U3789 (N_3789,In_292,In_1366);
or U3790 (N_3790,In_811,In_285);
and U3791 (N_3791,In_919,In_992);
xor U3792 (N_3792,In_124,In_574);
or U3793 (N_3793,In_1408,In_1328);
or U3794 (N_3794,In_1200,In_4);
nor U3795 (N_3795,In_1410,In_266);
nand U3796 (N_3796,In_994,In_889);
xnor U3797 (N_3797,In_1076,In_472);
nor U3798 (N_3798,In_627,In_44);
nor U3799 (N_3799,In_395,In_293);
or U3800 (N_3800,In_114,In_597);
xnor U3801 (N_3801,In_303,In_518);
nand U3802 (N_3802,In_1135,In_784);
or U3803 (N_3803,In_1485,In_1270);
and U3804 (N_3804,In_1091,In_292);
nand U3805 (N_3805,In_20,In_863);
xnor U3806 (N_3806,In_460,In_1227);
and U3807 (N_3807,In_1071,In_1016);
or U3808 (N_3808,In_796,In_272);
xor U3809 (N_3809,In_1451,In_1032);
and U3810 (N_3810,In_1391,In_160);
and U3811 (N_3811,In_1355,In_241);
nand U3812 (N_3812,In_305,In_499);
xor U3813 (N_3813,In_1120,In_272);
or U3814 (N_3814,In_751,In_723);
nor U3815 (N_3815,In_374,In_586);
and U3816 (N_3816,In_1103,In_1430);
nand U3817 (N_3817,In_905,In_1488);
xnor U3818 (N_3818,In_415,In_1239);
nand U3819 (N_3819,In_589,In_1468);
nor U3820 (N_3820,In_571,In_416);
nand U3821 (N_3821,In_281,In_599);
or U3822 (N_3822,In_1490,In_285);
nand U3823 (N_3823,In_51,In_721);
or U3824 (N_3824,In_1209,In_1395);
or U3825 (N_3825,In_1206,In_32);
xnor U3826 (N_3826,In_395,In_961);
and U3827 (N_3827,In_1224,In_161);
nand U3828 (N_3828,In_550,In_815);
or U3829 (N_3829,In_470,In_388);
xnor U3830 (N_3830,In_1002,In_0);
nand U3831 (N_3831,In_377,In_1213);
xor U3832 (N_3832,In_386,In_244);
and U3833 (N_3833,In_316,In_1187);
nor U3834 (N_3834,In_51,In_1391);
or U3835 (N_3835,In_568,In_1278);
xor U3836 (N_3836,In_49,In_788);
or U3837 (N_3837,In_445,In_883);
xor U3838 (N_3838,In_570,In_406);
xor U3839 (N_3839,In_401,In_1238);
nand U3840 (N_3840,In_1462,In_311);
xnor U3841 (N_3841,In_496,In_1072);
or U3842 (N_3842,In_540,In_1161);
nor U3843 (N_3843,In_1039,In_939);
nand U3844 (N_3844,In_81,In_1327);
xnor U3845 (N_3845,In_245,In_275);
and U3846 (N_3846,In_334,In_755);
and U3847 (N_3847,In_915,In_406);
nor U3848 (N_3848,In_338,In_562);
xor U3849 (N_3849,In_1096,In_1102);
xnor U3850 (N_3850,In_173,In_1104);
nand U3851 (N_3851,In_1063,In_1472);
xor U3852 (N_3852,In_734,In_1387);
nor U3853 (N_3853,In_895,In_1346);
nor U3854 (N_3854,In_79,In_564);
xnor U3855 (N_3855,In_676,In_72);
xor U3856 (N_3856,In_558,In_1239);
xnor U3857 (N_3857,In_1384,In_830);
nor U3858 (N_3858,In_1441,In_534);
xor U3859 (N_3859,In_617,In_255);
nor U3860 (N_3860,In_443,In_438);
and U3861 (N_3861,In_1096,In_1055);
and U3862 (N_3862,In_589,In_629);
nand U3863 (N_3863,In_520,In_307);
and U3864 (N_3864,In_1436,In_157);
xor U3865 (N_3865,In_715,In_213);
or U3866 (N_3866,In_365,In_8);
or U3867 (N_3867,In_1462,In_1263);
and U3868 (N_3868,In_929,In_1325);
or U3869 (N_3869,In_1160,In_184);
or U3870 (N_3870,In_1287,In_692);
xor U3871 (N_3871,In_688,In_1116);
xor U3872 (N_3872,In_756,In_65);
nor U3873 (N_3873,In_1036,In_65);
and U3874 (N_3874,In_773,In_374);
nand U3875 (N_3875,In_74,In_1479);
xnor U3876 (N_3876,In_1011,In_1413);
nand U3877 (N_3877,In_1357,In_530);
or U3878 (N_3878,In_690,In_1262);
xor U3879 (N_3879,In_391,In_1375);
nor U3880 (N_3880,In_1387,In_75);
nand U3881 (N_3881,In_389,In_431);
nor U3882 (N_3882,In_1343,In_981);
nand U3883 (N_3883,In_1398,In_836);
nand U3884 (N_3884,In_1246,In_1271);
xnor U3885 (N_3885,In_194,In_224);
and U3886 (N_3886,In_663,In_1036);
xor U3887 (N_3887,In_382,In_1389);
or U3888 (N_3888,In_237,In_1141);
or U3889 (N_3889,In_516,In_535);
xor U3890 (N_3890,In_184,In_246);
xnor U3891 (N_3891,In_569,In_434);
and U3892 (N_3892,In_373,In_1467);
or U3893 (N_3893,In_345,In_330);
xnor U3894 (N_3894,In_1051,In_275);
and U3895 (N_3895,In_445,In_1475);
and U3896 (N_3896,In_1240,In_1347);
xnor U3897 (N_3897,In_775,In_658);
nand U3898 (N_3898,In_474,In_545);
nor U3899 (N_3899,In_174,In_1286);
nand U3900 (N_3900,In_774,In_559);
or U3901 (N_3901,In_233,In_1070);
nand U3902 (N_3902,In_1060,In_258);
and U3903 (N_3903,In_441,In_627);
or U3904 (N_3904,In_1301,In_1041);
nor U3905 (N_3905,In_287,In_616);
nor U3906 (N_3906,In_1281,In_946);
or U3907 (N_3907,In_1454,In_77);
nor U3908 (N_3908,In_153,In_1491);
xor U3909 (N_3909,In_363,In_370);
or U3910 (N_3910,In_89,In_1083);
nand U3911 (N_3911,In_504,In_1352);
nand U3912 (N_3912,In_909,In_1177);
nor U3913 (N_3913,In_908,In_941);
xnor U3914 (N_3914,In_87,In_898);
nor U3915 (N_3915,In_722,In_1396);
and U3916 (N_3916,In_648,In_421);
and U3917 (N_3917,In_525,In_997);
nand U3918 (N_3918,In_294,In_277);
nand U3919 (N_3919,In_67,In_1112);
and U3920 (N_3920,In_144,In_1298);
nand U3921 (N_3921,In_1334,In_592);
or U3922 (N_3922,In_564,In_510);
and U3923 (N_3923,In_346,In_949);
nand U3924 (N_3924,In_58,In_292);
or U3925 (N_3925,In_1258,In_821);
or U3926 (N_3926,In_234,In_1053);
xnor U3927 (N_3927,In_1131,In_913);
or U3928 (N_3928,In_75,In_244);
nor U3929 (N_3929,In_7,In_900);
or U3930 (N_3930,In_896,In_1327);
nor U3931 (N_3931,In_140,In_398);
and U3932 (N_3932,In_1376,In_1447);
xor U3933 (N_3933,In_116,In_631);
nand U3934 (N_3934,In_859,In_784);
xor U3935 (N_3935,In_71,In_891);
or U3936 (N_3936,In_70,In_1288);
or U3937 (N_3937,In_1369,In_60);
xor U3938 (N_3938,In_636,In_1133);
and U3939 (N_3939,In_1069,In_131);
nor U3940 (N_3940,In_82,In_240);
nand U3941 (N_3941,In_975,In_853);
xnor U3942 (N_3942,In_1382,In_347);
or U3943 (N_3943,In_1497,In_1363);
nor U3944 (N_3944,In_1487,In_133);
xnor U3945 (N_3945,In_196,In_761);
xor U3946 (N_3946,In_51,In_972);
and U3947 (N_3947,In_834,In_634);
nor U3948 (N_3948,In_572,In_955);
nand U3949 (N_3949,In_46,In_778);
nor U3950 (N_3950,In_215,In_271);
or U3951 (N_3951,In_187,In_488);
and U3952 (N_3952,In_322,In_508);
xor U3953 (N_3953,In_283,In_1147);
and U3954 (N_3954,In_1104,In_818);
nor U3955 (N_3955,In_407,In_526);
nor U3956 (N_3956,In_203,In_1110);
and U3957 (N_3957,In_1043,In_143);
xnor U3958 (N_3958,In_394,In_97);
and U3959 (N_3959,In_694,In_912);
xnor U3960 (N_3960,In_1445,In_413);
nor U3961 (N_3961,In_1006,In_709);
or U3962 (N_3962,In_108,In_1323);
and U3963 (N_3963,In_1480,In_903);
xor U3964 (N_3964,In_1430,In_404);
nor U3965 (N_3965,In_60,In_1025);
or U3966 (N_3966,In_1472,In_749);
nor U3967 (N_3967,In_322,In_514);
and U3968 (N_3968,In_1358,In_1340);
nand U3969 (N_3969,In_220,In_722);
or U3970 (N_3970,In_1247,In_1454);
or U3971 (N_3971,In_834,In_1137);
or U3972 (N_3972,In_224,In_871);
or U3973 (N_3973,In_1205,In_1335);
xor U3974 (N_3974,In_559,In_419);
or U3975 (N_3975,In_22,In_305);
or U3976 (N_3976,In_708,In_92);
nand U3977 (N_3977,In_1124,In_1015);
or U3978 (N_3978,In_1310,In_994);
nor U3979 (N_3979,In_436,In_991);
or U3980 (N_3980,In_877,In_933);
nand U3981 (N_3981,In_817,In_932);
nand U3982 (N_3982,In_974,In_257);
nand U3983 (N_3983,In_579,In_674);
and U3984 (N_3984,In_711,In_439);
nand U3985 (N_3985,In_1309,In_770);
and U3986 (N_3986,In_1052,In_127);
nand U3987 (N_3987,In_84,In_325);
and U3988 (N_3988,In_1396,In_520);
xor U3989 (N_3989,In_1337,In_501);
and U3990 (N_3990,In_808,In_323);
and U3991 (N_3991,In_1125,In_484);
nand U3992 (N_3992,In_369,In_445);
and U3993 (N_3993,In_821,In_967);
and U3994 (N_3994,In_1292,In_1438);
or U3995 (N_3995,In_1082,In_1266);
nor U3996 (N_3996,In_1444,In_1498);
and U3997 (N_3997,In_195,In_1486);
xnor U3998 (N_3998,In_142,In_1273);
and U3999 (N_3999,In_535,In_1467);
or U4000 (N_4000,In_519,In_344);
nor U4001 (N_4001,In_1365,In_914);
xor U4002 (N_4002,In_249,In_329);
or U4003 (N_4003,In_1347,In_231);
nand U4004 (N_4004,In_403,In_910);
nor U4005 (N_4005,In_1217,In_284);
nand U4006 (N_4006,In_205,In_59);
nand U4007 (N_4007,In_1325,In_1178);
nand U4008 (N_4008,In_347,In_1074);
nand U4009 (N_4009,In_728,In_869);
nor U4010 (N_4010,In_1392,In_413);
xnor U4011 (N_4011,In_653,In_827);
or U4012 (N_4012,In_518,In_976);
or U4013 (N_4013,In_648,In_85);
and U4014 (N_4014,In_1088,In_1482);
or U4015 (N_4015,In_261,In_1484);
xor U4016 (N_4016,In_1374,In_269);
nor U4017 (N_4017,In_187,In_1057);
nor U4018 (N_4018,In_319,In_735);
nand U4019 (N_4019,In_666,In_702);
xnor U4020 (N_4020,In_759,In_1035);
and U4021 (N_4021,In_770,In_884);
or U4022 (N_4022,In_134,In_949);
xnor U4023 (N_4023,In_587,In_636);
nand U4024 (N_4024,In_632,In_1119);
nor U4025 (N_4025,In_1432,In_591);
xnor U4026 (N_4026,In_217,In_823);
or U4027 (N_4027,In_1278,In_211);
nand U4028 (N_4028,In_634,In_393);
nand U4029 (N_4029,In_657,In_1081);
or U4030 (N_4030,In_1362,In_251);
or U4031 (N_4031,In_782,In_313);
and U4032 (N_4032,In_182,In_1484);
nor U4033 (N_4033,In_1420,In_795);
and U4034 (N_4034,In_1463,In_842);
and U4035 (N_4035,In_431,In_56);
and U4036 (N_4036,In_517,In_734);
and U4037 (N_4037,In_132,In_1182);
nor U4038 (N_4038,In_1034,In_602);
nand U4039 (N_4039,In_652,In_1381);
nor U4040 (N_4040,In_788,In_130);
xnor U4041 (N_4041,In_1307,In_519);
xnor U4042 (N_4042,In_1127,In_844);
xnor U4043 (N_4043,In_1358,In_1266);
nand U4044 (N_4044,In_556,In_936);
nand U4045 (N_4045,In_782,In_558);
nand U4046 (N_4046,In_1243,In_31);
nand U4047 (N_4047,In_328,In_187);
nor U4048 (N_4048,In_127,In_757);
xnor U4049 (N_4049,In_45,In_850);
nand U4050 (N_4050,In_540,In_767);
xor U4051 (N_4051,In_1471,In_1186);
nand U4052 (N_4052,In_59,In_165);
and U4053 (N_4053,In_553,In_349);
and U4054 (N_4054,In_1091,In_1181);
or U4055 (N_4055,In_1355,In_730);
xor U4056 (N_4056,In_1423,In_91);
nand U4057 (N_4057,In_1251,In_202);
nand U4058 (N_4058,In_643,In_1496);
or U4059 (N_4059,In_1183,In_769);
nor U4060 (N_4060,In_636,In_1338);
or U4061 (N_4061,In_1316,In_1307);
nor U4062 (N_4062,In_1142,In_1102);
and U4063 (N_4063,In_1266,In_307);
nor U4064 (N_4064,In_669,In_57);
or U4065 (N_4065,In_70,In_208);
and U4066 (N_4066,In_687,In_786);
xor U4067 (N_4067,In_987,In_1051);
or U4068 (N_4068,In_1244,In_1264);
or U4069 (N_4069,In_404,In_68);
or U4070 (N_4070,In_392,In_93);
or U4071 (N_4071,In_282,In_1132);
nand U4072 (N_4072,In_979,In_93);
or U4073 (N_4073,In_1302,In_525);
xor U4074 (N_4074,In_363,In_1324);
nor U4075 (N_4075,In_1481,In_151);
nand U4076 (N_4076,In_502,In_1241);
nand U4077 (N_4077,In_1038,In_978);
and U4078 (N_4078,In_877,In_320);
and U4079 (N_4079,In_606,In_88);
and U4080 (N_4080,In_869,In_667);
xnor U4081 (N_4081,In_701,In_1447);
nor U4082 (N_4082,In_590,In_736);
xnor U4083 (N_4083,In_869,In_355);
and U4084 (N_4084,In_655,In_719);
nand U4085 (N_4085,In_765,In_1343);
and U4086 (N_4086,In_1351,In_990);
or U4087 (N_4087,In_202,In_561);
and U4088 (N_4088,In_1488,In_338);
and U4089 (N_4089,In_653,In_1176);
nor U4090 (N_4090,In_1385,In_943);
or U4091 (N_4091,In_188,In_899);
and U4092 (N_4092,In_1437,In_1100);
nand U4093 (N_4093,In_360,In_815);
or U4094 (N_4094,In_350,In_1289);
xor U4095 (N_4095,In_482,In_1380);
nand U4096 (N_4096,In_193,In_1252);
nand U4097 (N_4097,In_1451,In_1279);
nor U4098 (N_4098,In_1419,In_352);
nor U4099 (N_4099,In_430,In_1229);
nand U4100 (N_4100,In_20,In_1318);
nand U4101 (N_4101,In_1368,In_503);
and U4102 (N_4102,In_569,In_1299);
nor U4103 (N_4103,In_1460,In_883);
nor U4104 (N_4104,In_113,In_1185);
nor U4105 (N_4105,In_1221,In_523);
nand U4106 (N_4106,In_1003,In_1304);
nor U4107 (N_4107,In_665,In_1246);
and U4108 (N_4108,In_413,In_443);
or U4109 (N_4109,In_326,In_1190);
and U4110 (N_4110,In_929,In_1011);
nor U4111 (N_4111,In_453,In_552);
nand U4112 (N_4112,In_802,In_171);
and U4113 (N_4113,In_878,In_116);
xnor U4114 (N_4114,In_507,In_1161);
xor U4115 (N_4115,In_1472,In_1036);
nand U4116 (N_4116,In_1306,In_1196);
nor U4117 (N_4117,In_1310,In_1039);
xnor U4118 (N_4118,In_1141,In_340);
or U4119 (N_4119,In_271,In_314);
and U4120 (N_4120,In_47,In_1137);
or U4121 (N_4121,In_683,In_34);
or U4122 (N_4122,In_482,In_473);
xor U4123 (N_4123,In_1037,In_112);
xnor U4124 (N_4124,In_469,In_765);
nor U4125 (N_4125,In_558,In_769);
nand U4126 (N_4126,In_1322,In_1049);
xnor U4127 (N_4127,In_1425,In_504);
xor U4128 (N_4128,In_1101,In_1005);
and U4129 (N_4129,In_81,In_128);
and U4130 (N_4130,In_1161,In_1265);
or U4131 (N_4131,In_620,In_568);
or U4132 (N_4132,In_149,In_90);
nor U4133 (N_4133,In_263,In_1471);
nand U4134 (N_4134,In_657,In_1469);
nand U4135 (N_4135,In_190,In_392);
xor U4136 (N_4136,In_578,In_73);
xnor U4137 (N_4137,In_678,In_398);
nor U4138 (N_4138,In_31,In_1175);
nor U4139 (N_4139,In_1356,In_119);
and U4140 (N_4140,In_447,In_129);
nor U4141 (N_4141,In_46,In_1162);
nor U4142 (N_4142,In_505,In_261);
and U4143 (N_4143,In_106,In_1247);
or U4144 (N_4144,In_683,In_1288);
or U4145 (N_4145,In_627,In_101);
nor U4146 (N_4146,In_785,In_1358);
or U4147 (N_4147,In_129,In_1246);
and U4148 (N_4148,In_739,In_28);
nand U4149 (N_4149,In_900,In_104);
or U4150 (N_4150,In_669,In_20);
xnor U4151 (N_4151,In_1295,In_311);
xnor U4152 (N_4152,In_1434,In_715);
nor U4153 (N_4153,In_1288,In_1074);
or U4154 (N_4154,In_735,In_1211);
nand U4155 (N_4155,In_740,In_1260);
or U4156 (N_4156,In_298,In_765);
or U4157 (N_4157,In_193,In_1173);
xor U4158 (N_4158,In_1126,In_470);
nor U4159 (N_4159,In_1027,In_1486);
or U4160 (N_4160,In_1113,In_419);
or U4161 (N_4161,In_535,In_689);
nand U4162 (N_4162,In_279,In_254);
or U4163 (N_4163,In_1294,In_401);
or U4164 (N_4164,In_1390,In_133);
nand U4165 (N_4165,In_447,In_363);
or U4166 (N_4166,In_883,In_1314);
and U4167 (N_4167,In_48,In_584);
nand U4168 (N_4168,In_847,In_116);
xor U4169 (N_4169,In_197,In_1439);
xor U4170 (N_4170,In_1103,In_65);
nand U4171 (N_4171,In_356,In_1134);
nand U4172 (N_4172,In_556,In_59);
or U4173 (N_4173,In_240,In_684);
nand U4174 (N_4174,In_1097,In_1382);
nand U4175 (N_4175,In_325,In_1023);
nor U4176 (N_4176,In_1153,In_286);
nor U4177 (N_4177,In_1306,In_1151);
nor U4178 (N_4178,In_341,In_881);
nand U4179 (N_4179,In_312,In_878);
nand U4180 (N_4180,In_1341,In_1328);
xor U4181 (N_4181,In_1074,In_425);
xnor U4182 (N_4182,In_1293,In_636);
nand U4183 (N_4183,In_190,In_1333);
and U4184 (N_4184,In_281,In_1239);
xnor U4185 (N_4185,In_1027,In_99);
and U4186 (N_4186,In_771,In_878);
xor U4187 (N_4187,In_219,In_1162);
xnor U4188 (N_4188,In_580,In_1134);
or U4189 (N_4189,In_1313,In_912);
xnor U4190 (N_4190,In_517,In_319);
nand U4191 (N_4191,In_23,In_732);
nand U4192 (N_4192,In_1263,In_373);
xor U4193 (N_4193,In_854,In_1263);
or U4194 (N_4194,In_415,In_802);
nor U4195 (N_4195,In_1264,In_1121);
or U4196 (N_4196,In_98,In_404);
and U4197 (N_4197,In_746,In_1364);
nor U4198 (N_4198,In_864,In_687);
nand U4199 (N_4199,In_490,In_757);
xor U4200 (N_4200,In_1106,In_1279);
xor U4201 (N_4201,In_1128,In_884);
nor U4202 (N_4202,In_825,In_151);
and U4203 (N_4203,In_1442,In_1412);
or U4204 (N_4204,In_1208,In_239);
or U4205 (N_4205,In_1146,In_203);
and U4206 (N_4206,In_941,In_191);
xor U4207 (N_4207,In_1282,In_205);
and U4208 (N_4208,In_543,In_759);
nor U4209 (N_4209,In_625,In_765);
nor U4210 (N_4210,In_602,In_390);
xnor U4211 (N_4211,In_158,In_549);
or U4212 (N_4212,In_1450,In_1367);
nand U4213 (N_4213,In_698,In_405);
nor U4214 (N_4214,In_253,In_482);
and U4215 (N_4215,In_1370,In_535);
nor U4216 (N_4216,In_1234,In_703);
xor U4217 (N_4217,In_832,In_1164);
xor U4218 (N_4218,In_910,In_744);
or U4219 (N_4219,In_391,In_785);
and U4220 (N_4220,In_383,In_1133);
nor U4221 (N_4221,In_485,In_1056);
or U4222 (N_4222,In_855,In_314);
nand U4223 (N_4223,In_1479,In_1294);
or U4224 (N_4224,In_715,In_807);
xnor U4225 (N_4225,In_1084,In_863);
nor U4226 (N_4226,In_236,In_461);
nor U4227 (N_4227,In_698,In_885);
and U4228 (N_4228,In_1026,In_1266);
or U4229 (N_4229,In_1434,In_475);
nor U4230 (N_4230,In_1232,In_369);
nand U4231 (N_4231,In_503,In_699);
nand U4232 (N_4232,In_443,In_1420);
nor U4233 (N_4233,In_719,In_1130);
or U4234 (N_4234,In_418,In_92);
or U4235 (N_4235,In_1338,In_175);
nor U4236 (N_4236,In_81,In_934);
and U4237 (N_4237,In_778,In_1388);
or U4238 (N_4238,In_1058,In_132);
xnor U4239 (N_4239,In_882,In_1267);
nand U4240 (N_4240,In_1490,In_1200);
nand U4241 (N_4241,In_1265,In_1134);
nor U4242 (N_4242,In_1458,In_1159);
xnor U4243 (N_4243,In_1477,In_1109);
xor U4244 (N_4244,In_1254,In_860);
nor U4245 (N_4245,In_1209,In_111);
xnor U4246 (N_4246,In_580,In_710);
and U4247 (N_4247,In_231,In_1138);
nor U4248 (N_4248,In_846,In_173);
or U4249 (N_4249,In_415,In_847);
and U4250 (N_4250,In_54,In_559);
nor U4251 (N_4251,In_1368,In_1280);
nand U4252 (N_4252,In_89,In_1060);
or U4253 (N_4253,In_1417,In_484);
nor U4254 (N_4254,In_1014,In_1369);
and U4255 (N_4255,In_1400,In_812);
and U4256 (N_4256,In_313,In_779);
or U4257 (N_4257,In_282,In_1411);
xnor U4258 (N_4258,In_431,In_1041);
and U4259 (N_4259,In_1443,In_182);
nor U4260 (N_4260,In_767,In_388);
or U4261 (N_4261,In_20,In_965);
nand U4262 (N_4262,In_435,In_467);
or U4263 (N_4263,In_452,In_1182);
and U4264 (N_4264,In_1047,In_677);
nor U4265 (N_4265,In_1321,In_12);
xor U4266 (N_4266,In_637,In_1385);
nor U4267 (N_4267,In_1204,In_934);
nand U4268 (N_4268,In_269,In_1449);
xor U4269 (N_4269,In_574,In_593);
or U4270 (N_4270,In_112,In_1343);
xor U4271 (N_4271,In_786,In_273);
xnor U4272 (N_4272,In_933,In_283);
or U4273 (N_4273,In_402,In_1434);
nor U4274 (N_4274,In_854,In_418);
nand U4275 (N_4275,In_1271,In_367);
nor U4276 (N_4276,In_717,In_36);
and U4277 (N_4277,In_734,In_381);
nor U4278 (N_4278,In_368,In_562);
and U4279 (N_4279,In_1308,In_635);
or U4280 (N_4280,In_800,In_310);
nor U4281 (N_4281,In_876,In_624);
and U4282 (N_4282,In_800,In_291);
nand U4283 (N_4283,In_25,In_23);
and U4284 (N_4284,In_864,In_972);
nor U4285 (N_4285,In_1406,In_1047);
or U4286 (N_4286,In_92,In_55);
xor U4287 (N_4287,In_1421,In_624);
nand U4288 (N_4288,In_504,In_828);
or U4289 (N_4289,In_1409,In_459);
and U4290 (N_4290,In_1221,In_417);
xnor U4291 (N_4291,In_194,In_610);
and U4292 (N_4292,In_253,In_1457);
xor U4293 (N_4293,In_491,In_880);
xnor U4294 (N_4294,In_1494,In_1147);
xnor U4295 (N_4295,In_719,In_1344);
nand U4296 (N_4296,In_232,In_654);
and U4297 (N_4297,In_675,In_1060);
xor U4298 (N_4298,In_231,In_1018);
or U4299 (N_4299,In_451,In_446);
and U4300 (N_4300,In_809,In_995);
and U4301 (N_4301,In_382,In_1204);
and U4302 (N_4302,In_785,In_983);
and U4303 (N_4303,In_1146,In_183);
or U4304 (N_4304,In_1127,In_1453);
nand U4305 (N_4305,In_1404,In_907);
xnor U4306 (N_4306,In_1212,In_1082);
nor U4307 (N_4307,In_462,In_346);
xor U4308 (N_4308,In_970,In_564);
nor U4309 (N_4309,In_1215,In_140);
or U4310 (N_4310,In_963,In_163);
and U4311 (N_4311,In_817,In_61);
nor U4312 (N_4312,In_857,In_656);
nand U4313 (N_4313,In_1141,In_705);
nor U4314 (N_4314,In_293,In_1429);
nor U4315 (N_4315,In_218,In_1284);
or U4316 (N_4316,In_1028,In_574);
nor U4317 (N_4317,In_527,In_410);
nor U4318 (N_4318,In_292,In_530);
xor U4319 (N_4319,In_710,In_345);
xor U4320 (N_4320,In_445,In_1136);
nand U4321 (N_4321,In_630,In_1087);
xnor U4322 (N_4322,In_623,In_902);
nand U4323 (N_4323,In_1002,In_1006);
xor U4324 (N_4324,In_307,In_900);
nand U4325 (N_4325,In_1254,In_609);
xnor U4326 (N_4326,In_1252,In_1395);
and U4327 (N_4327,In_697,In_19);
and U4328 (N_4328,In_270,In_751);
xor U4329 (N_4329,In_270,In_1282);
and U4330 (N_4330,In_1414,In_1311);
nor U4331 (N_4331,In_77,In_776);
or U4332 (N_4332,In_1029,In_746);
xnor U4333 (N_4333,In_864,In_328);
xor U4334 (N_4334,In_62,In_1382);
or U4335 (N_4335,In_1430,In_1088);
xnor U4336 (N_4336,In_1080,In_787);
and U4337 (N_4337,In_463,In_1369);
and U4338 (N_4338,In_1273,In_327);
xnor U4339 (N_4339,In_455,In_721);
nand U4340 (N_4340,In_72,In_1390);
and U4341 (N_4341,In_235,In_267);
and U4342 (N_4342,In_1336,In_712);
nand U4343 (N_4343,In_819,In_817);
xor U4344 (N_4344,In_1373,In_670);
nor U4345 (N_4345,In_6,In_1141);
nand U4346 (N_4346,In_1065,In_1486);
nand U4347 (N_4347,In_128,In_807);
nand U4348 (N_4348,In_91,In_342);
xor U4349 (N_4349,In_612,In_1179);
or U4350 (N_4350,In_469,In_339);
nor U4351 (N_4351,In_1358,In_918);
and U4352 (N_4352,In_767,In_800);
nand U4353 (N_4353,In_1115,In_523);
nand U4354 (N_4354,In_1333,In_465);
nor U4355 (N_4355,In_259,In_719);
nand U4356 (N_4356,In_663,In_1039);
nand U4357 (N_4357,In_333,In_479);
and U4358 (N_4358,In_1162,In_930);
xor U4359 (N_4359,In_295,In_558);
xor U4360 (N_4360,In_1088,In_408);
xor U4361 (N_4361,In_451,In_622);
or U4362 (N_4362,In_1093,In_1250);
and U4363 (N_4363,In_776,In_579);
and U4364 (N_4364,In_102,In_1195);
nand U4365 (N_4365,In_828,In_363);
or U4366 (N_4366,In_498,In_913);
nand U4367 (N_4367,In_888,In_1474);
and U4368 (N_4368,In_372,In_1276);
and U4369 (N_4369,In_37,In_1338);
nor U4370 (N_4370,In_958,In_703);
nor U4371 (N_4371,In_232,In_217);
and U4372 (N_4372,In_773,In_515);
or U4373 (N_4373,In_447,In_1344);
and U4374 (N_4374,In_1476,In_1074);
xor U4375 (N_4375,In_33,In_586);
and U4376 (N_4376,In_3,In_730);
nand U4377 (N_4377,In_1296,In_422);
or U4378 (N_4378,In_232,In_435);
xnor U4379 (N_4379,In_405,In_249);
or U4380 (N_4380,In_2,In_273);
or U4381 (N_4381,In_473,In_723);
nor U4382 (N_4382,In_1057,In_1330);
xor U4383 (N_4383,In_980,In_1096);
xor U4384 (N_4384,In_1148,In_65);
nand U4385 (N_4385,In_1363,In_70);
or U4386 (N_4386,In_1375,In_490);
and U4387 (N_4387,In_986,In_1061);
xor U4388 (N_4388,In_316,In_201);
and U4389 (N_4389,In_1478,In_375);
nor U4390 (N_4390,In_323,In_862);
and U4391 (N_4391,In_1030,In_137);
or U4392 (N_4392,In_1042,In_68);
and U4393 (N_4393,In_1231,In_182);
and U4394 (N_4394,In_576,In_546);
nand U4395 (N_4395,In_656,In_395);
nand U4396 (N_4396,In_1358,In_997);
nor U4397 (N_4397,In_104,In_1444);
xnor U4398 (N_4398,In_714,In_484);
nor U4399 (N_4399,In_1191,In_1171);
nand U4400 (N_4400,In_53,In_1399);
nand U4401 (N_4401,In_840,In_906);
or U4402 (N_4402,In_1059,In_1328);
nor U4403 (N_4403,In_169,In_418);
nand U4404 (N_4404,In_983,In_701);
nand U4405 (N_4405,In_311,In_529);
and U4406 (N_4406,In_1490,In_602);
nand U4407 (N_4407,In_815,In_1158);
nand U4408 (N_4408,In_103,In_1094);
xnor U4409 (N_4409,In_1348,In_649);
xnor U4410 (N_4410,In_950,In_618);
or U4411 (N_4411,In_850,In_435);
nor U4412 (N_4412,In_1479,In_793);
and U4413 (N_4413,In_695,In_1141);
xor U4414 (N_4414,In_736,In_468);
and U4415 (N_4415,In_1193,In_619);
xor U4416 (N_4416,In_1262,In_1489);
nand U4417 (N_4417,In_709,In_468);
or U4418 (N_4418,In_444,In_1020);
nand U4419 (N_4419,In_646,In_821);
xor U4420 (N_4420,In_661,In_974);
nor U4421 (N_4421,In_1489,In_1183);
or U4422 (N_4422,In_1097,In_999);
and U4423 (N_4423,In_1374,In_617);
and U4424 (N_4424,In_156,In_1426);
nor U4425 (N_4425,In_926,In_123);
xor U4426 (N_4426,In_202,In_330);
nor U4427 (N_4427,In_291,In_401);
nor U4428 (N_4428,In_369,In_1264);
and U4429 (N_4429,In_682,In_12);
or U4430 (N_4430,In_995,In_1359);
nand U4431 (N_4431,In_1044,In_844);
xnor U4432 (N_4432,In_145,In_593);
and U4433 (N_4433,In_1268,In_144);
nand U4434 (N_4434,In_883,In_811);
xor U4435 (N_4435,In_266,In_990);
and U4436 (N_4436,In_1164,In_1278);
nand U4437 (N_4437,In_477,In_1190);
xor U4438 (N_4438,In_1407,In_190);
xnor U4439 (N_4439,In_232,In_811);
or U4440 (N_4440,In_1032,In_1059);
and U4441 (N_4441,In_459,In_82);
nand U4442 (N_4442,In_311,In_301);
or U4443 (N_4443,In_1165,In_167);
nor U4444 (N_4444,In_1072,In_383);
and U4445 (N_4445,In_547,In_784);
and U4446 (N_4446,In_1431,In_1105);
or U4447 (N_4447,In_1498,In_518);
nor U4448 (N_4448,In_479,In_187);
and U4449 (N_4449,In_537,In_309);
xor U4450 (N_4450,In_1225,In_959);
xor U4451 (N_4451,In_1492,In_49);
nand U4452 (N_4452,In_169,In_798);
nand U4453 (N_4453,In_1303,In_569);
xor U4454 (N_4454,In_1174,In_767);
nand U4455 (N_4455,In_284,In_402);
and U4456 (N_4456,In_174,In_1341);
and U4457 (N_4457,In_981,In_845);
and U4458 (N_4458,In_542,In_1010);
and U4459 (N_4459,In_1407,In_1422);
nand U4460 (N_4460,In_1401,In_193);
or U4461 (N_4461,In_257,In_1103);
and U4462 (N_4462,In_1100,In_391);
nand U4463 (N_4463,In_1489,In_1324);
and U4464 (N_4464,In_80,In_421);
xor U4465 (N_4465,In_698,In_72);
nand U4466 (N_4466,In_661,In_167);
xor U4467 (N_4467,In_447,In_951);
nor U4468 (N_4468,In_59,In_193);
nor U4469 (N_4469,In_350,In_629);
or U4470 (N_4470,In_1353,In_11);
xor U4471 (N_4471,In_282,In_130);
nor U4472 (N_4472,In_744,In_667);
or U4473 (N_4473,In_893,In_1377);
xnor U4474 (N_4474,In_723,In_479);
nand U4475 (N_4475,In_491,In_482);
or U4476 (N_4476,In_108,In_817);
or U4477 (N_4477,In_723,In_1191);
xnor U4478 (N_4478,In_104,In_715);
nand U4479 (N_4479,In_107,In_534);
or U4480 (N_4480,In_546,In_1461);
xnor U4481 (N_4481,In_176,In_788);
or U4482 (N_4482,In_66,In_200);
or U4483 (N_4483,In_16,In_127);
nor U4484 (N_4484,In_866,In_204);
and U4485 (N_4485,In_825,In_159);
and U4486 (N_4486,In_996,In_264);
and U4487 (N_4487,In_1236,In_1116);
or U4488 (N_4488,In_1345,In_67);
or U4489 (N_4489,In_546,In_397);
nand U4490 (N_4490,In_63,In_877);
nor U4491 (N_4491,In_355,In_513);
nor U4492 (N_4492,In_1320,In_473);
xor U4493 (N_4493,In_100,In_1035);
xnor U4494 (N_4494,In_1494,In_1381);
nand U4495 (N_4495,In_471,In_387);
nand U4496 (N_4496,In_1119,In_402);
or U4497 (N_4497,In_757,In_1427);
and U4498 (N_4498,In_792,In_1172);
or U4499 (N_4499,In_1306,In_621);
or U4500 (N_4500,In_1136,In_401);
nand U4501 (N_4501,In_197,In_1273);
nand U4502 (N_4502,In_1328,In_1000);
xor U4503 (N_4503,In_39,In_782);
xor U4504 (N_4504,In_286,In_597);
nand U4505 (N_4505,In_141,In_1142);
nor U4506 (N_4506,In_1006,In_1295);
nor U4507 (N_4507,In_448,In_1250);
and U4508 (N_4508,In_989,In_708);
nand U4509 (N_4509,In_1114,In_1220);
and U4510 (N_4510,In_120,In_1482);
nor U4511 (N_4511,In_528,In_43);
or U4512 (N_4512,In_1095,In_1303);
xnor U4513 (N_4513,In_1132,In_888);
nor U4514 (N_4514,In_842,In_386);
xor U4515 (N_4515,In_633,In_473);
xor U4516 (N_4516,In_942,In_218);
xor U4517 (N_4517,In_936,In_465);
xor U4518 (N_4518,In_1364,In_1156);
nor U4519 (N_4519,In_1228,In_282);
nor U4520 (N_4520,In_1053,In_605);
and U4521 (N_4521,In_277,In_863);
and U4522 (N_4522,In_69,In_572);
nand U4523 (N_4523,In_49,In_1457);
nand U4524 (N_4524,In_414,In_1389);
nand U4525 (N_4525,In_1029,In_924);
and U4526 (N_4526,In_136,In_1219);
xor U4527 (N_4527,In_583,In_12);
xnor U4528 (N_4528,In_1040,In_184);
and U4529 (N_4529,In_1068,In_884);
and U4530 (N_4530,In_412,In_723);
nand U4531 (N_4531,In_1313,In_96);
or U4532 (N_4532,In_963,In_1323);
nand U4533 (N_4533,In_166,In_539);
nor U4534 (N_4534,In_864,In_347);
xnor U4535 (N_4535,In_624,In_374);
or U4536 (N_4536,In_15,In_1486);
and U4537 (N_4537,In_393,In_543);
or U4538 (N_4538,In_741,In_962);
nor U4539 (N_4539,In_419,In_696);
nand U4540 (N_4540,In_223,In_1021);
nor U4541 (N_4541,In_922,In_1386);
nor U4542 (N_4542,In_518,In_497);
nor U4543 (N_4543,In_839,In_1087);
nor U4544 (N_4544,In_511,In_1412);
nor U4545 (N_4545,In_898,In_694);
nor U4546 (N_4546,In_112,In_597);
nand U4547 (N_4547,In_157,In_771);
xnor U4548 (N_4548,In_371,In_54);
nand U4549 (N_4549,In_803,In_422);
nor U4550 (N_4550,In_61,In_275);
and U4551 (N_4551,In_1452,In_1494);
nand U4552 (N_4552,In_156,In_782);
nand U4553 (N_4553,In_1085,In_158);
or U4554 (N_4554,In_1310,In_329);
and U4555 (N_4555,In_253,In_1097);
nand U4556 (N_4556,In_332,In_434);
nor U4557 (N_4557,In_929,In_407);
nor U4558 (N_4558,In_607,In_1181);
xor U4559 (N_4559,In_553,In_1351);
or U4560 (N_4560,In_52,In_1094);
or U4561 (N_4561,In_8,In_1117);
and U4562 (N_4562,In_829,In_898);
nand U4563 (N_4563,In_723,In_1115);
or U4564 (N_4564,In_1274,In_662);
nand U4565 (N_4565,In_1051,In_774);
xor U4566 (N_4566,In_1232,In_215);
and U4567 (N_4567,In_699,In_665);
nand U4568 (N_4568,In_92,In_87);
or U4569 (N_4569,In_1135,In_1061);
xor U4570 (N_4570,In_93,In_287);
or U4571 (N_4571,In_226,In_1185);
or U4572 (N_4572,In_1142,In_410);
nor U4573 (N_4573,In_935,In_45);
nor U4574 (N_4574,In_1271,In_1026);
and U4575 (N_4575,In_643,In_594);
or U4576 (N_4576,In_791,In_1002);
xor U4577 (N_4577,In_920,In_291);
xor U4578 (N_4578,In_220,In_1361);
xnor U4579 (N_4579,In_1453,In_1231);
xnor U4580 (N_4580,In_392,In_1149);
and U4581 (N_4581,In_249,In_305);
xnor U4582 (N_4582,In_507,In_487);
nand U4583 (N_4583,In_942,In_653);
or U4584 (N_4584,In_408,In_960);
and U4585 (N_4585,In_77,In_833);
nand U4586 (N_4586,In_136,In_160);
nand U4587 (N_4587,In_718,In_861);
and U4588 (N_4588,In_1188,In_683);
and U4589 (N_4589,In_211,In_247);
nand U4590 (N_4590,In_53,In_879);
and U4591 (N_4591,In_128,In_365);
and U4592 (N_4592,In_28,In_485);
nor U4593 (N_4593,In_450,In_1073);
xor U4594 (N_4594,In_1021,In_1238);
nor U4595 (N_4595,In_751,In_1325);
or U4596 (N_4596,In_901,In_1061);
xnor U4597 (N_4597,In_407,In_1070);
nand U4598 (N_4598,In_938,In_611);
xor U4599 (N_4599,In_1355,In_1001);
nand U4600 (N_4600,In_279,In_788);
nor U4601 (N_4601,In_236,In_1433);
or U4602 (N_4602,In_317,In_798);
and U4603 (N_4603,In_1212,In_1256);
and U4604 (N_4604,In_694,In_339);
or U4605 (N_4605,In_1086,In_1457);
nand U4606 (N_4606,In_1166,In_920);
and U4607 (N_4607,In_881,In_1073);
nand U4608 (N_4608,In_1425,In_587);
xnor U4609 (N_4609,In_1209,In_168);
nand U4610 (N_4610,In_243,In_204);
xnor U4611 (N_4611,In_966,In_415);
nor U4612 (N_4612,In_686,In_511);
or U4613 (N_4613,In_889,In_803);
or U4614 (N_4614,In_224,In_236);
nand U4615 (N_4615,In_744,In_72);
xnor U4616 (N_4616,In_1052,In_1068);
or U4617 (N_4617,In_905,In_313);
xnor U4618 (N_4618,In_103,In_489);
xnor U4619 (N_4619,In_91,In_1189);
and U4620 (N_4620,In_1282,In_644);
nor U4621 (N_4621,In_619,In_1335);
nand U4622 (N_4622,In_1182,In_1377);
and U4623 (N_4623,In_1275,In_1353);
or U4624 (N_4624,In_249,In_268);
xor U4625 (N_4625,In_17,In_56);
or U4626 (N_4626,In_618,In_277);
or U4627 (N_4627,In_821,In_1170);
nor U4628 (N_4628,In_617,In_162);
nand U4629 (N_4629,In_14,In_265);
nor U4630 (N_4630,In_1297,In_59);
nand U4631 (N_4631,In_496,In_520);
and U4632 (N_4632,In_374,In_385);
xnor U4633 (N_4633,In_525,In_120);
nand U4634 (N_4634,In_1201,In_1013);
xnor U4635 (N_4635,In_740,In_772);
and U4636 (N_4636,In_1047,In_543);
nor U4637 (N_4637,In_255,In_900);
and U4638 (N_4638,In_1471,In_272);
nand U4639 (N_4639,In_1454,In_774);
or U4640 (N_4640,In_850,In_1353);
and U4641 (N_4641,In_402,In_286);
xor U4642 (N_4642,In_554,In_708);
nand U4643 (N_4643,In_989,In_451);
nand U4644 (N_4644,In_1266,In_354);
and U4645 (N_4645,In_565,In_1427);
nor U4646 (N_4646,In_922,In_986);
nor U4647 (N_4647,In_1379,In_1423);
and U4648 (N_4648,In_58,In_848);
and U4649 (N_4649,In_703,In_338);
and U4650 (N_4650,In_262,In_561);
nand U4651 (N_4651,In_996,In_791);
nand U4652 (N_4652,In_276,In_731);
and U4653 (N_4653,In_581,In_688);
nor U4654 (N_4654,In_883,In_698);
xor U4655 (N_4655,In_1202,In_984);
or U4656 (N_4656,In_314,In_1457);
and U4657 (N_4657,In_1144,In_1199);
nor U4658 (N_4658,In_281,In_467);
xor U4659 (N_4659,In_3,In_166);
xnor U4660 (N_4660,In_1404,In_589);
nand U4661 (N_4661,In_1320,In_1136);
and U4662 (N_4662,In_437,In_1214);
nor U4663 (N_4663,In_240,In_41);
xor U4664 (N_4664,In_1475,In_676);
or U4665 (N_4665,In_937,In_1024);
or U4666 (N_4666,In_1132,In_126);
nor U4667 (N_4667,In_647,In_1375);
or U4668 (N_4668,In_1070,In_458);
xnor U4669 (N_4669,In_378,In_1310);
and U4670 (N_4670,In_753,In_1367);
nor U4671 (N_4671,In_146,In_807);
and U4672 (N_4672,In_1115,In_1172);
xnor U4673 (N_4673,In_960,In_1385);
or U4674 (N_4674,In_615,In_161);
nor U4675 (N_4675,In_365,In_3);
nand U4676 (N_4676,In_786,In_58);
and U4677 (N_4677,In_1100,In_632);
and U4678 (N_4678,In_257,In_1320);
and U4679 (N_4679,In_1136,In_932);
nand U4680 (N_4680,In_1014,In_881);
xnor U4681 (N_4681,In_103,In_301);
nand U4682 (N_4682,In_6,In_729);
and U4683 (N_4683,In_1475,In_586);
or U4684 (N_4684,In_1359,In_244);
and U4685 (N_4685,In_531,In_208);
xnor U4686 (N_4686,In_434,In_1414);
and U4687 (N_4687,In_1374,In_694);
and U4688 (N_4688,In_24,In_1391);
and U4689 (N_4689,In_552,In_635);
nand U4690 (N_4690,In_1352,In_864);
nor U4691 (N_4691,In_560,In_1331);
xnor U4692 (N_4692,In_1049,In_1345);
xnor U4693 (N_4693,In_1096,In_563);
nor U4694 (N_4694,In_592,In_477);
or U4695 (N_4695,In_223,In_636);
or U4696 (N_4696,In_140,In_596);
or U4697 (N_4697,In_743,In_1295);
and U4698 (N_4698,In_138,In_161);
nand U4699 (N_4699,In_227,In_803);
xor U4700 (N_4700,In_555,In_900);
and U4701 (N_4701,In_362,In_1231);
xor U4702 (N_4702,In_150,In_1384);
nor U4703 (N_4703,In_668,In_755);
xor U4704 (N_4704,In_1098,In_582);
nor U4705 (N_4705,In_956,In_736);
nor U4706 (N_4706,In_326,In_857);
nand U4707 (N_4707,In_109,In_128);
nor U4708 (N_4708,In_572,In_385);
nand U4709 (N_4709,In_141,In_36);
nor U4710 (N_4710,In_642,In_1333);
nand U4711 (N_4711,In_86,In_487);
or U4712 (N_4712,In_1433,In_1462);
xor U4713 (N_4713,In_1281,In_1412);
xor U4714 (N_4714,In_557,In_356);
nor U4715 (N_4715,In_1281,In_266);
and U4716 (N_4716,In_877,In_483);
xnor U4717 (N_4717,In_202,In_379);
or U4718 (N_4718,In_1017,In_236);
or U4719 (N_4719,In_1076,In_1358);
xnor U4720 (N_4720,In_526,In_373);
xor U4721 (N_4721,In_1378,In_309);
and U4722 (N_4722,In_412,In_665);
nand U4723 (N_4723,In_693,In_967);
or U4724 (N_4724,In_1127,In_473);
or U4725 (N_4725,In_1373,In_253);
nor U4726 (N_4726,In_580,In_428);
or U4727 (N_4727,In_645,In_1449);
xnor U4728 (N_4728,In_447,In_123);
nor U4729 (N_4729,In_730,In_701);
or U4730 (N_4730,In_139,In_1310);
nand U4731 (N_4731,In_9,In_807);
nor U4732 (N_4732,In_308,In_323);
nand U4733 (N_4733,In_1360,In_552);
xor U4734 (N_4734,In_45,In_307);
nor U4735 (N_4735,In_377,In_1036);
nor U4736 (N_4736,In_252,In_107);
or U4737 (N_4737,In_1469,In_175);
xor U4738 (N_4738,In_693,In_828);
and U4739 (N_4739,In_1167,In_644);
and U4740 (N_4740,In_994,In_579);
xor U4741 (N_4741,In_1270,In_1065);
and U4742 (N_4742,In_554,In_813);
nor U4743 (N_4743,In_459,In_611);
nand U4744 (N_4744,In_1090,In_206);
nor U4745 (N_4745,In_1051,In_76);
xor U4746 (N_4746,In_709,In_644);
xnor U4747 (N_4747,In_621,In_855);
nor U4748 (N_4748,In_1275,In_382);
and U4749 (N_4749,In_1477,In_834);
nor U4750 (N_4750,In_367,In_517);
nand U4751 (N_4751,In_961,In_1132);
xnor U4752 (N_4752,In_367,In_1050);
and U4753 (N_4753,In_474,In_769);
xnor U4754 (N_4754,In_1395,In_813);
xor U4755 (N_4755,In_887,In_1053);
and U4756 (N_4756,In_726,In_553);
or U4757 (N_4757,In_1230,In_186);
nand U4758 (N_4758,In_1185,In_97);
nor U4759 (N_4759,In_569,In_1131);
xor U4760 (N_4760,In_725,In_689);
or U4761 (N_4761,In_1399,In_751);
or U4762 (N_4762,In_474,In_1000);
and U4763 (N_4763,In_899,In_1198);
xor U4764 (N_4764,In_1043,In_1052);
and U4765 (N_4765,In_1461,In_60);
and U4766 (N_4766,In_921,In_1195);
xnor U4767 (N_4767,In_766,In_574);
nor U4768 (N_4768,In_1386,In_588);
and U4769 (N_4769,In_112,In_557);
and U4770 (N_4770,In_3,In_902);
nor U4771 (N_4771,In_1073,In_235);
nand U4772 (N_4772,In_146,In_462);
nor U4773 (N_4773,In_659,In_195);
nand U4774 (N_4774,In_784,In_1000);
xor U4775 (N_4775,In_117,In_104);
and U4776 (N_4776,In_232,In_1136);
xnor U4777 (N_4777,In_468,In_1131);
or U4778 (N_4778,In_303,In_726);
nand U4779 (N_4779,In_1406,In_634);
or U4780 (N_4780,In_759,In_346);
xnor U4781 (N_4781,In_156,In_888);
xor U4782 (N_4782,In_975,In_1257);
or U4783 (N_4783,In_18,In_1401);
or U4784 (N_4784,In_1128,In_1122);
or U4785 (N_4785,In_924,In_971);
or U4786 (N_4786,In_56,In_1101);
or U4787 (N_4787,In_842,In_1312);
nor U4788 (N_4788,In_769,In_1103);
or U4789 (N_4789,In_945,In_1083);
xor U4790 (N_4790,In_1109,In_1396);
nor U4791 (N_4791,In_951,In_882);
nor U4792 (N_4792,In_1223,In_1477);
nor U4793 (N_4793,In_901,In_111);
and U4794 (N_4794,In_544,In_983);
and U4795 (N_4795,In_563,In_89);
or U4796 (N_4796,In_801,In_1381);
and U4797 (N_4797,In_1194,In_84);
nand U4798 (N_4798,In_1080,In_1356);
xnor U4799 (N_4799,In_437,In_1017);
nor U4800 (N_4800,In_1024,In_608);
nor U4801 (N_4801,In_1124,In_995);
and U4802 (N_4802,In_712,In_1008);
nand U4803 (N_4803,In_1012,In_1459);
xor U4804 (N_4804,In_333,In_780);
xor U4805 (N_4805,In_1245,In_168);
nand U4806 (N_4806,In_1066,In_987);
or U4807 (N_4807,In_1406,In_1366);
or U4808 (N_4808,In_787,In_148);
and U4809 (N_4809,In_1097,In_187);
nand U4810 (N_4810,In_1334,In_892);
and U4811 (N_4811,In_1408,In_14);
nand U4812 (N_4812,In_524,In_98);
and U4813 (N_4813,In_301,In_449);
nand U4814 (N_4814,In_605,In_1118);
xnor U4815 (N_4815,In_243,In_239);
or U4816 (N_4816,In_1491,In_216);
nand U4817 (N_4817,In_590,In_558);
xor U4818 (N_4818,In_389,In_331);
nor U4819 (N_4819,In_584,In_811);
nand U4820 (N_4820,In_1154,In_926);
xor U4821 (N_4821,In_391,In_512);
and U4822 (N_4822,In_491,In_432);
and U4823 (N_4823,In_1012,In_1337);
or U4824 (N_4824,In_37,In_1331);
nor U4825 (N_4825,In_868,In_776);
nor U4826 (N_4826,In_930,In_692);
and U4827 (N_4827,In_491,In_754);
nor U4828 (N_4828,In_1383,In_203);
or U4829 (N_4829,In_1210,In_1190);
or U4830 (N_4830,In_1396,In_1464);
nor U4831 (N_4831,In_9,In_221);
nand U4832 (N_4832,In_1014,In_1231);
nand U4833 (N_4833,In_487,In_1257);
xor U4834 (N_4834,In_315,In_487);
or U4835 (N_4835,In_1027,In_1370);
xnor U4836 (N_4836,In_246,In_560);
and U4837 (N_4837,In_1048,In_212);
xnor U4838 (N_4838,In_188,In_1458);
or U4839 (N_4839,In_865,In_17);
xnor U4840 (N_4840,In_142,In_875);
nor U4841 (N_4841,In_234,In_473);
and U4842 (N_4842,In_76,In_50);
nor U4843 (N_4843,In_319,In_61);
xnor U4844 (N_4844,In_673,In_46);
xnor U4845 (N_4845,In_649,In_1152);
or U4846 (N_4846,In_1222,In_1189);
nor U4847 (N_4847,In_641,In_712);
or U4848 (N_4848,In_709,In_977);
and U4849 (N_4849,In_749,In_229);
nand U4850 (N_4850,In_1083,In_568);
and U4851 (N_4851,In_914,In_1392);
and U4852 (N_4852,In_924,In_893);
or U4853 (N_4853,In_741,In_1234);
xnor U4854 (N_4854,In_980,In_505);
xor U4855 (N_4855,In_866,In_978);
xor U4856 (N_4856,In_650,In_285);
xor U4857 (N_4857,In_1259,In_1185);
xor U4858 (N_4858,In_153,In_766);
xor U4859 (N_4859,In_693,In_542);
and U4860 (N_4860,In_351,In_0);
nor U4861 (N_4861,In_39,In_442);
xnor U4862 (N_4862,In_1175,In_930);
or U4863 (N_4863,In_1082,In_1113);
nand U4864 (N_4864,In_339,In_1187);
nand U4865 (N_4865,In_394,In_845);
and U4866 (N_4866,In_830,In_1286);
or U4867 (N_4867,In_28,In_456);
or U4868 (N_4868,In_1209,In_907);
nor U4869 (N_4869,In_1463,In_875);
nand U4870 (N_4870,In_686,In_777);
xnor U4871 (N_4871,In_1417,In_266);
nor U4872 (N_4872,In_568,In_497);
xor U4873 (N_4873,In_859,In_420);
and U4874 (N_4874,In_844,In_475);
and U4875 (N_4875,In_1447,In_848);
nand U4876 (N_4876,In_546,In_1195);
xor U4877 (N_4877,In_917,In_1456);
or U4878 (N_4878,In_748,In_327);
or U4879 (N_4879,In_1142,In_323);
nor U4880 (N_4880,In_1353,In_1438);
and U4881 (N_4881,In_1471,In_5);
or U4882 (N_4882,In_1443,In_1123);
xnor U4883 (N_4883,In_1082,In_689);
nand U4884 (N_4884,In_1305,In_431);
nor U4885 (N_4885,In_1045,In_172);
or U4886 (N_4886,In_650,In_1450);
xor U4887 (N_4887,In_1034,In_1324);
nand U4888 (N_4888,In_77,In_880);
and U4889 (N_4889,In_1257,In_354);
nand U4890 (N_4890,In_801,In_972);
or U4891 (N_4891,In_1327,In_481);
nand U4892 (N_4892,In_1122,In_263);
and U4893 (N_4893,In_716,In_479);
nand U4894 (N_4894,In_618,In_1416);
or U4895 (N_4895,In_183,In_134);
nor U4896 (N_4896,In_22,In_1369);
or U4897 (N_4897,In_525,In_170);
nor U4898 (N_4898,In_1129,In_65);
nand U4899 (N_4899,In_891,In_1079);
xor U4900 (N_4900,In_1084,In_798);
nand U4901 (N_4901,In_268,In_895);
nand U4902 (N_4902,In_63,In_1439);
nand U4903 (N_4903,In_1269,In_1047);
nand U4904 (N_4904,In_399,In_592);
nand U4905 (N_4905,In_1163,In_488);
and U4906 (N_4906,In_1189,In_1228);
nor U4907 (N_4907,In_650,In_446);
nor U4908 (N_4908,In_1473,In_37);
xnor U4909 (N_4909,In_1189,In_765);
and U4910 (N_4910,In_1327,In_289);
xor U4911 (N_4911,In_894,In_132);
nor U4912 (N_4912,In_1020,In_412);
nand U4913 (N_4913,In_533,In_717);
nor U4914 (N_4914,In_124,In_1148);
xnor U4915 (N_4915,In_715,In_406);
or U4916 (N_4916,In_16,In_957);
nand U4917 (N_4917,In_577,In_730);
xor U4918 (N_4918,In_810,In_224);
nor U4919 (N_4919,In_265,In_700);
nor U4920 (N_4920,In_58,In_394);
or U4921 (N_4921,In_670,In_1093);
or U4922 (N_4922,In_863,In_1379);
or U4923 (N_4923,In_474,In_1124);
xnor U4924 (N_4924,In_493,In_12);
or U4925 (N_4925,In_1353,In_957);
nor U4926 (N_4926,In_50,In_470);
and U4927 (N_4927,In_1272,In_218);
nand U4928 (N_4928,In_464,In_214);
nand U4929 (N_4929,In_377,In_9);
and U4930 (N_4930,In_29,In_19);
and U4931 (N_4931,In_14,In_1415);
and U4932 (N_4932,In_1450,In_1140);
nor U4933 (N_4933,In_1368,In_579);
nor U4934 (N_4934,In_1366,In_726);
xnor U4935 (N_4935,In_412,In_1422);
nand U4936 (N_4936,In_686,In_1329);
and U4937 (N_4937,In_1269,In_462);
or U4938 (N_4938,In_505,In_934);
nand U4939 (N_4939,In_99,In_882);
xnor U4940 (N_4940,In_16,In_32);
or U4941 (N_4941,In_1082,In_37);
nand U4942 (N_4942,In_349,In_130);
and U4943 (N_4943,In_1149,In_1495);
or U4944 (N_4944,In_57,In_731);
nand U4945 (N_4945,In_190,In_1125);
or U4946 (N_4946,In_1044,In_258);
nor U4947 (N_4947,In_23,In_253);
or U4948 (N_4948,In_309,In_583);
and U4949 (N_4949,In_443,In_774);
and U4950 (N_4950,In_442,In_530);
nand U4951 (N_4951,In_354,In_130);
or U4952 (N_4952,In_721,In_1333);
nor U4953 (N_4953,In_1441,In_721);
and U4954 (N_4954,In_666,In_1276);
or U4955 (N_4955,In_287,In_1498);
and U4956 (N_4956,In_1363,In_105);
nor U4957 (N_4957,In_1310,In_771);
or U4958 (N_4958,In_1149,In_638);
nand U4959 (N_4959,In_1250,In_894);
xnor U4960 (N_4960,In_692,In_659);
nand U4961 (N_4961,In_1013,In_390);
nor U4962 (N_4962,In_231,In_1355);
nand U4963 (N_4963,In_932,In_1108);
nor U4964 (N_4964,In_1136,In_266);
nand U4965 (N_4965,In_351,In_1192);
xor U4966 (N_4966,In_522,In_1074);
nor U4967 (N_4967,In_333,In_705);
or U4968 (N_4968,In_1406,In_1156);
nor U4969 (N_4969,In_123,In_1289);
nand U4970 (N_4970,In_1416,In_1273);
or U4971 (N_4971,In_314,In_223);
and U4972 (N_4972,In_1343,In_38);
or U4973 (N_4973,In_581,In_821);
or U4974 (N_4974,In_1002,In_449);
nor U4975 (N_4975,In_738,In_155);
or U4976 (N_4976,In_872,In_257);
nand U4977 (N_4977,In_903,In_1203);
and U4978 (N_4978,In_1023,In_55);
xnor U4979 (N_4979,In_733,In_17);
nor U4980 (N_4980,In_499,In_55);
nand U4981 (N_4981,In_176,In_1134);
nand U4982 (N_4982,In_835,In_829);
and U4983 (N_4983,In_1238,In_927);
or U4984 (N_4984,In_472,In_1282);
and U4985 (N_4985,In_1365,In_239);
or U4986 (N_4986,In_907,In_184);
nand U4987 (N_4987,In_839,In_23);
and U4988 (N_4988,In_1458,In_816);
and U4989 (N_4989,In_975,In_1200);
nand U4990 (N_4990,In_275,In_1046);
nor U4991 (N_4991,In_407,In_639);
xnor U4992 (N_4992,In_1186,In_998);
and U4993 (N_4993,In_551,In_1127);
nor U4994 (N_4994,In_760,In_596);
or U4995 (N_4995,In_765,In_805);
xor U4996 (N_4996,In_457,In_553);
and U4997 (N_4997,In_527,In_566);
nor U4998 (N_4998,In_462,In_197);
nor U4999 (N_4999,In_9,In_1079);
and U5000 (N_5000,N_1598,N_494);
nand U5001 (N_5001,N_3512,N_375);
xnor U5002 (N_5002,N_1496,N_4904);
xor U5003 (N_5003,N_1851,N_1241);
xor U5004 (N_5004,N_1015,N_3539);
or U5005 (N_5005,N_43,N_3404);
and U5006 (N_5006,N_919,N_187);
nor U5007 (N_5007,N_735,N_965);
or U5008 (N_5008,N_1893,N_736);
xor U5009 (N_5009,N_3050,N_3556);
nand U5010 (N_5010,N_221,N_3949);
and U5011 (N_5011,N_1172,N_1468);
nor U5012 (N_5012,N_365,N_4873);
xor U5013 (N_5013,N_1880,N_2833);
xnor U5014 (N_5014,N_2382,N_3397);
nand U5015 (N_5015,N_1407,N_4265);
nand U5016 (N_5016,N_4200,N_2027);
nor U5017 (N_5017,N_9,N_742);
or U5018 (N_5018,N_3762,N_4411);
nor U5019 (N_5019,N_2050,N_2423);
xnor U5020 (N_5020,N_605,N_3578);
xnor U5021 (N_5021,N_4569,N_2767);
nand U5022 (N_5022,N_4857,N_4050);
xnor U5023 (N_5023,N_416,N_3016);
xnor U5024 (N_5024,N_1891,N_4881);
nor U5025 (N_5025,N_153,N_912);
nand U5026 (N_5026,N_4827,N_4193);
nand U5027 (N_5027,N_3612,N_578);
nor U5028 (N_5028,N_422,N_1109);
xor U5029 (N_5029,N_3433,N_2712);
xor U5030 (N_5030,N_1984,N_1961);
xor U5031 (N_5031,N_2340,N_2751);
nand U5032 (N_5032,N_4006,N_1579);
xnor U5033 (N_5033,N_2037,N_4263);
xor U5034 (N_5034,N_1458,N_3571);
nor U5035 (N_5035,N_4514,N_1261);
xnor U5036 (N_5036,N_2555,N_1383);
nor U5037 (N_5037,N_284,N_4964);
nand U5038 (N_5038,N_2719,N_32);
or U5039 (N_5039,N_2856,N_1113);
nor U5040 (N_5040,N_3113,N_2465);
nand U5041 (N_5041,N_3255,N_400);
and U5042 (N_5042,N_413,N_2764);
or U5043 (N_5043,N_606,N_800);
nor U5044 (N_5044,N_1382,N_3664);
and U5045 (N_5045,N_3020,N_3817);
or U5046 (N_5046,N_3650,N_4536);
nor U5047 (N_5047,N_1174,N_2273);
xnor U5048 (N_5048,N_1536,N_2511);
nand U5049 (N_5049,N_4093,N_4190);
and U5050 (N_5050,N_4042,N_3291);
and U5051 (N_5051,N_3683,N_3701);
nand U5052 (N_5052,N_4935,N_4224);
and U5053 (N_5053,N_2016,N_686);
nor U5054 (N_5054,N_3148,N_1732);
and U5055 (N_5055,N_500,N_3111);
nand U5056 (N_5056,N_841,N_1747);
nand U5057 (N_5057,N_3479,N_3848);
or U5058 (N_5058,N_2663,N_2035);
nor U5059 (N_5059,N_183,N_4153);
xnor U5060 (N_5060,N_1527,N_2725);
xnor U5061 (N_5061,N_3800,N_1127);
nand U5062 (N_5062,N_562,N_4926);
and U5063 (N_5063,N_4388,N_2627);
nor U5064 (N_5064,N_381,N_1288);
xnor U5065 (N_5065,N_53,N_1473);
xnor U5066 (N_5066,N_4324,N_2752);
xnor U5067 (N_5067,N_2458,N_2595);
nand U5068 (N_5068,N_456,N_3424);
and U5069 (N_5069,N_517,N_4933);
xor U5070 (N_5070,N_2641,N_780);
or U5071 (N_5071,N_2900,N_1665);
nor U5072 (N_5072,N_61,N_1583);
or U5073 (N_5073,N_4898,N_488);
and U5074 (N_5074,N_1006,N_3724);
xnor U5075 (N_5075,N_1378,N_4296);
xnor U5076 (N_5076,N_4977,N_2017);
xnor U5077 (N_5077,N_1460,N_3373);
and U5078 (N_5078,N_4094,N_3934);
nor U5079 (N_5079,N_3205,N_810);
nand U5080 (N_5080,N_4567,N_1103);
or U5081 (N_5081,N_1727,N_2957);
xor U5082 (N_5082,N_21,N_4192);
nand U5083 (N_5083,N_480,N_678);
nor U5084 (N_5084,N_4782,N_3064);
or U5085 (N_5085,N_175,N_4652);
nand U5086 (N_5086,N_672,N_1303);
and U5087 (N_5087,N_4290,N_4323);
and U5088 (N_5088,N_1795,N_1718);
or U5089 (N_5089,N_3428,N_425);
and U5090 (N_5090,N_1150,N_2443);
or U5091 (N_5091,N_4763,N_1039);
nand U5092 (N_5092,N_1020,N_4829);
and U5093 (N_5093,N_891,N_2987);
or U5094 (N_5094,N_1441,N_1203);
nand U5095 (N_5095,N_3352,N_3543);
nor U5096 (N_5096,N_4412,N_1495);
xnor U5097 (N_5097,N_110,N_1521);
nand U5098 (N_5098,N_3114,N_3210);
xor U5099 (N_5099,N_3450,N_1141);
xnor U5100 (N_5100,N_2055,N_1206);
nand U5101 (N_5101,N_3857,N_3915);
nand U5102 (N_5102,N_2177,N_1531);
xor U5103 (N_5103,N_99,N_3334);
nor U5104 (N_5104,N_4463,N_3906);
xnor U5105 (N_5105,N_254,N_2560);
nor U5106 (N_5106,N_201,N_4996);
and U5107 (N_5107,N_3407,N_493);
nor U5108 (N_5108,N_3832,N_3858);
and U5109 (N_5109,N_4951,N_979);
and U5110 (N_5110,N_1021,N_893);
nand U5111 (N_5111,N_3598,N_3788);
and U5112 (N_5112,N_2248,N_2876);
and U5113 (N_5113,N_3624,N_632);
nor U5114 (N_5114,N_184,N_726);
xor U5115 (N_5115,N_4397,N_1721);
xor U5116 (N_5116,N_2284,N_1632);
nor U5117 (N_5117,N_536,N_3487);
xnor U5118 (N_5118,N_2429,N_1777);
xnor U5119 (N_5119,N_2271,N_1275);
or U5120 (N_5120,N_333,N_4440);
or U5121 (N_5121,N_4171,N_3994);
and U5122 (N_5122,N_4267,N_4545);
xnor U5123 (N_5123,N_4141,N_4436);
and U5124 (N_5124,N_2233,N_4633);
nor U5125 (N_5125,N_1522,N_3620);
and U5126 (N_5126,N_3575,N_2899);
or U5127 (N_5127,N_4308,N_642);
and U5128 (N_5128,N_4096,N_302);
or U5129 (N_5129,N_395,N_424);
nor U5130 (N_5130,N_3583,N_2694);
nand U5131 (N_5131,N_854,N_3546);
and U5132 (N_5132,N_4066,N_2845);
nand U5133 (N_5133,N_4475,N_4466);
nand U5134 (N_5134,N_1101,N_4616);
nor U5135 (N_5135,N_4896,N_181);
nand U5136 (N_5136,N_3340,N_234);
and U5137 (N_5137,N_2625,N_3121);
or U5138 (N_5138,N_1041,N_3787);
or U5139 (N_5139,N_794,N_2777);
and U5140 (N_5140,N_1225,N_4973);
xor U5141 (N_5141,N_1847,N_4194);
nor U5142 (N_5142,N_2231,N_4457);
or U5143 (N_5143,N_2968,N_4826);
nor U5144 (N_5144,N_3072,N_3110);
or U5145 (N_5145,N_1106,N_1293);
and U5146 (N_5146,N_4086,N_3025);
and U5147 (N_5147,N_3715,N_2474);
and U5148 (N_5148,N_2519,N_1869);
nand U5149 (N_5149,N_1565,N_120);
or U5150 (N_5150,N_3029,N_2006);
nand U5151 (N_5151,N_1988,N_1262);
or U5152 (N_5152,N_348,N_1080);
and U5153 (N_5153,N_1230,N_1852);
and U5154 (N_5154,N_2144,N_3609);
xnor U5155 (N_5155,N_3347,N_2374);
nand U5156 (N_5156,N_4478,N_665);
nand U5157 (N_5157,N_4586,N_4554);
and U5158 (N_5158,N_906,N_762);
and U5159 (N_5159,N_4434,N_3507);
xnor U5160 (N_5160,N_1554,N_1641);
nor U5161 (N_5161,N_1363,N_3923);
and U5162 (N_5162,N_3948,N_2657);
nand U5163 (N_5163,N_2163,N_3458);
or U5164 (N_5164,N_740,N_1729);
nand U5165 (N_5165,N_689,N_4158);
or U5166 (N_5166,N_1821,N_3357);
nor U5167 (N_5167,N_2780,N_4980);
xnor U5168 (N_5168,N_265,N_4078);
and U5169 (N_5169,N_4049,N_2930);
or U5170 (N_5170,N_3386,N_3966);
nor U5171 (N_5171,N_353,N_2317);
nand U5172 (N_5172,N_2416,N_1047);
or U5173 (N_5173,N_2695,N_531);
and U5174 (N_5174,N_35,N_4753);
nand U5175 (N_5175,N_3851,N_1760);
and U5176 (N_5176,N_1018,N_802);
xnor U5177 (N_5177,N_3123,N_1836);
xor U5178 (N_5178,N_2138,N_2091);
or U5179 (N_5179,N_2524,N_4026);
nor U5180 (N_5180,N_2483,N_2387);
nor U5181 (N_5181,N_1714,N_4261);
nor U5182 (N_5182,N_3881,N_4936);
nor U5183 (N_5183,N_3807,N_1208);
xor U5184 (N_5184,N_2165,N_877);
or U5185 (N_5185,N_1350,N_2187);
and U5186 (N_5186,N_36,N_1387);
nor U5187 (N_5187,N_1181,N_4344);
xnor U5188 (N_5188,N_2424,N_3815);
nor U5189 (N_5189,N_237,N_3070);
or U5190 (N_5190,N_4143,N_1265);
xnor U5191 (N_5191,N_4556,N_297);
nand U5192 (N_5192,N_2958,N_2026);
and U5193 (N_5193,N_3738,N_2604);
or U5194 (N_5194,N_4840,N_481);
nor U5195 (N_5195,N_3155,N_2605);
xnor U5196 (N_5196,N_445,N_1909);
or U5197 (N_5197,N_871,N_2064);
nor U5198 (N_5198,N_1928,N_335);
and U5199 (N_5199,N_103,N_322);
nor U5200 (N_5200,N_1001,N_3495);
or U5201 (N_5201,N_1312,N_307);
nor U5202 (N_5202,N_573,N_4680);
nand U5203 (N_5203,N_4748,N_1576);
and U5204 (N_5204,N_2991,N_1846);
or U5205 (N_5205,N_2812,N_3860);
nand U5206 (N_5206,N_171,N_2012);
and U5207 (N_5207,N_1863,N_2320);
xnor U5208 (N_5208,N_2209,N_3791);
xor U5209 (N_5209,N_2115,N_3459);
and U5210 (N_5210,N_2992,N_783);
xor U5211 (N_5211,N_4963,N_2646);
xor U5212 (N_5212,N_3106,N_3721);
nand U5213 (N_5213,N_72,N_4882);
or U5214 (N_5214,N_2288,N_3378);
or U5215 (N_5215,N_4538,N_2307);
nor U5216 (N_5216,N_4288,N_4540);
or U5217 (N_5217,N_3117,N_805);
nand U5218 (N_5218,N_1032,N_4914);
xor U5219 (N_5219,N_1211,N_2183);
or U5220 (N_5220,N_4978,N_758);
nor U5221 (N_5221,N_1814,N_4467);
and U5222 (N_5222,N_4136,N_1072);
xor U5223 (N_5223,N_1175,N_435);
nor U5224 (N_5224,N_2167,N_1306);
or U5225 (N_5225,N_806,N_3538);
xnor U5226 (N_5226,N_4164,N_1200);
or U5227 (N_5227,N_3193,N_3919);
nand U5228 (N_5228,N_2190,N_1499);
or U5229 (N_5229,N_4894,N_3607);
or U5230 (N_5230,N_4019,N_3244);
and U5231 (N_5231,N_113,N_2832);
nor U5232 (N_5232,N_2457,N_1471);
xor U5233 (N_5233,N_403,N_2829);
nor U5234 (N_5234,N_308,N_3635);
nand U5235 (N_5235,N_420,N_186);
nor U5236 (N_5236,N_4565,N_2745);
or U5237 (N_5237,N_903,N_3831);
and U5238 (N_5238,N_639,N_6);
or U5239 (N_5239,N_693,N_4345);
or U5240 (N_5240,N_1298,N_4132);
xnor U5241 (N_5241,N_1385,N_1586);
nand U5242 (N_5242,N_660,N_895);
or U5243 (N_5243,N_1281,N_3931);
or U5244 (N_5244,N_3998,N_204);
xor U5245 (N_5245,N_1227,N_1853);
and U5246 (N_5246,N_3754,N_3035);
or U5247 (N_5247,N_303,N_4778);
xor U5248 (N_5248,N_467,N_2594);
and U5249 (N_5249,N_1201,N_4989);
nand U5250 (N_5250,N_916,N_3565);
xor U5251 (N_5251,N_2391,N_2974);
or U5252 (N_5252,N_3501,N_1987);
or U5253 (N_5253,N_1135,N_3587);
xor U5254 (N_5254,N_4295,N_1702);
nor U5255 (N_5255,N_939,N_4924);
nor U5256 (N_5256,N_1611,N_4728);
and U5257 (N_5257,N_4529,N_798);
and U5258 (N_5258,N_3989,N_4407);
nand U5259 (N_5259,N_2470,N_31);
or U5260 (N_5260,N_2372,N_3441);
and U5261 (N_5261,N_2994,N_2467);
and U5262 (N_5262,N_613,N_3585);
nor U5263 (N_5263,N_3263,N_2923);
nand U5264 (N_5264,N_1314,N_719);
or U5265 (N_5265,N_1654,N_957);
or U5266 (N_5266,N_3149,N_4819);
nor U5267 (N_5267,N_3038,N_1519);
nor U5268 (N_5268,N_464,N_2041);
nand U5269 (N_5269,N_4286,N_3276);
and U5270 (N_5270,N_4823,N_2668);
or U5271 (N_5271,N_2888,N_4161);
xor U5272 (N_5272,N_190,N_4689);
or U5273 (N_5273,N_3339,N_259);
or U5274 (N_5274,N_882,N_1011);
nor U5275 (N_5275,N_1986,N_4177);
or U5276 (N_5276,N_2619,N_2);
or U5277 (N_5277,N_1389,N_3653);
or U5278 (N_5278,N_3756,N_615);
nor U5279 (N_5279,N_4834,N_1341);
and U5280 (N_5280,N_2323,N_3734);
nor U5281 (N_5281,N_3658,N_1526);
xnor U5282 (N_5282,N_1927,N_4770);
nand U5283 (N_5283,N_1592,N_4719);
nor U5284 (N_5284,N_2475,N_534);
or U5285 (N_5285,N_3015,N_2097);
xor U5286 (N_5286,N_246,N_4932);
or U5287 (N_5287,N_1709,N_1449);
and U5288 (N_5288,N_2438,N_2312);
xor U5289 (N_5289,N_3160,N_700);
nand U5290 (N_5290,N_3173,N_3328);
nor U5291 (N_5291,N_71,N_4532);
and U5292 (N_5292,N_1299,N_875);
nor U5293 (N_5293,N_4034,N_385);
or U5294 (N_5294,N_857,N_1384);
nor U5295 (N_5295,N_202,N_1770);
nor U5296 (N_5296,N_4651,N_2535);
nor U5297 (N_5297,N_3592,N_2514);
nand U5298 (N_5298,N_272,N_631);
nand U5299 (N_5299,N_4509,N_4983);
nand U5300 (N_5300,N_3388,N_730);
nor U5301 (N_5301,N_1398,N_10);
or U5302 (N_5302,N_2543,N_3876);
nand U5303 (N_5303,N_2069,N_1983);
or U5304 (N_5304,N_2655,N_4931);
xnor U5305 (N_5305,N_1824,N_62);
nand U5306 (N_5306,N_4612,N_2647);
and U5307 (N_5307,N_3885,N_3518);
and U5308 (N_5308,N_4012,N_1036);
nor U5309 (N_5309,N_650,N_2274);
and U5310 (N_5310,N_1942,N_4106);
nor U5311 (N_5311,N_1994,N_3889);
xor U5312 (N_5312,N_2173,N_2858);
nand U5313 (N_5313,N_3890,N_807);
xor U5314 (N_5314,N_929,N_3985);
or U5315 (N_5315,N_941,N_2867);
nand U5316 (N_5316,N_4822,N_711);
nand U5317 (N_5317,N_2067,N_412);
or U5318 (N_5318,N_761,N_3238);
or U5319 (N_5319,N_2756,N_256);
nand U5320 (N_5320,N_3427,N_1662);
xnor U5321 (N_5321,N_3903,N_3248);
or U5322 (N_5322,N_1163,N_4154);
xor U5323 (N_5323,N_1152,N_940);
xnor U5324 (N_5324,N_1491,N_3437);
xor U5325 (N_5325,N_1883,N_3590);
or U5326 (N_5326,N_1012,N_2853);
nand U5327 (N_5327,N_2345,N_4000);
xnor U5328 (N_5328,N_4442,N_3709);
xor U5329 (N_5329,N_4886,N_2447);
and U5330 (N_5330,N_2418,N_3765);
nand U5331 (N_5331,N_824,N_155);
and U5332 (N_5332,N_2328,N_3820);
nand U5333 (N_5333,N_4516,N_4614);
nand U5334 (N_5334,N_831,N_4927);
or U5335 (N_5335,N_3484,N_718);
nor U5336 (N_5336,N_1631,N_737);
xnor U5337 (N_5337,N_775,N_2331);
xor U5338 (N_5338,N_123,N_1348);
or U5339 (N_5339,N_988,N_2341);
nor U5340 (N_5340,N_1764,N_1450);
and U5341 (N_5341,N_2815,N_3879);
nand U5342 (N_5342,N_1180,N_1255);
nand U5343 (N_5343,N_549,N_2473);
nand U5344 (N_5344,N_3203,N_4371);
nand U5345 (N_5345,N_2671,N_2682);
or U5346 (N_5346,N_1660,N_3391);
nor U5347 (N_5347,N_3936,N_2194);
nand U5348 (N_5348,N_4076,N_402);
nor U5349 (N_5349,N_4310,N_320);
nand U5350 (N_5350,N_253,N_1622);
or U5351 (N_5351,N_2077,N_70);
and U5352 (N_5352,N_4459,N_586);
and U5353 (N_5353,N_4937,N_2824);
nor U5354 (N_5354,N_3637,N_2933);
nor U5355 (N_5355,N_47,N_1695);
xnor U5356 (N_5356,N_3714,N_1750);
xnor U5357 (N_5357,N_599,N_2720);
nor U5358 (N_5358,N_812,N_2439);
xor U5359 (N_5359,N_670,N_4080);
nor U5360 (N_5360,N_3941,N_3237);
nor U5361 (N_5361,N_4287,N_3584);
and U5362 (N_5362,N_1748,N_2684);
nor U5363 (N_5363,N_2754,N_2609);
xnor U5364 (N_5364,N_3896,N_4868);
or U5365 (N_5365,N_2005,N_3892);
or U5366 (N_5366,N_1877,N_4798);
xor U5367 (N_5367,N_1758,N_1974);
nor U5368 (N_5368,N_250,N_679);
and U5369 (N_5369,N_1919,N_3104);
or U5370 (N_5370,N_2600,N_4752);
nand U5371 (N_5371,N_2488,N_1528);
nand U5372 (N_5372,N_1254,N_4421);
and U5373 (N_5373,N_727,N_1157);
nand U5374 (N_5374,N_4229,N_4302);
and U5375 (N_5375,N_1584,N_3644);
nor U5376 (N_5376,N_4750,N_4588);
nand U5377 (N_5377,N_4054,N_2112);
nand U5378 (N_5378,N_3400,N_2532);
or U5379 (N_5379,N_227,N_4941);
xnor U5380 (N_5380,N_4734,N_111);
and U5381 (N_5381,N_3116,N_1515);
and U5382 (N_5382,N_1644,N_2464);
nor U5383 (N_5383,N_1887,N_3991);
or U5384 (N_5384,N_1646,N_2141);
or U5385 (N_5385,N_3555,N_2364);
nand U5386 (N_5386,N_3986,N_1618);
and U5387 (N_5387,N_898,N_2776);
or U5388 (N_5388,N_3748,N_3535);
nand U5389 (N_5389,N_2969,N_682);
nand U5390 (N_5390,N_4995,N_1982);
or U5391 (N_5391,N_1464,N_3071);
or U5392 (N_5392,N_4115,N_3812);
xnor U5393 (N_5393,N_3201,N_4852);
and U5394 (N_5394,N_55,N_4965);
and U5395 (N_5395,N_3579,N_2260);
nor U5396 (N_5396,N_3321,N_2461);
or U5397 (N_5397,N_1235,N_1962);
xnor U5398 (N_5398,N_911,N_4550);
and U5399 (N_5399,N_4742,N_4640);
nor U5400 (N_5400,N_4490,N_1289);
or U5401 (N_5401,N_2807,N_2135);
and U5402 (N_5402,N_1486,N_1182);
and U5403 (N_5403,N_2285,N_1107);
nor U5404 (N_5404,N_4400,N_3976);
nor U5405 (N_5405,N_927,N_1674);
or U5406 (N_5406,N_3520,N_1892);
nor U5407 (N_5407,N_3599,N_236);
or U5408 (N_5408,N_3981,N_1765);
nor U5409 (N_5409,N_4124,N_1093);
xor U5410 (N_5410,N_1810,N_3646);
nand U5411 (N_5411,N_326,N_2820);
nand U5412 (N_5412,N_1420,N_661);
and U5413 (N_5413,N_3972,N_3383);
nand U5414 (N_5414,N_1297,N_4646);
nand U5415 (N_5415,N_458,N_2040);
nand U5416 (N_5416,N_2182,N_3181);
nor U5417 (N_5417,N_89,N_971);
or U5418 (N_5418,N_1691,N_721);
nor U5419 (N_5419,N_1086,N_3654);
xor U5420 (N_5420,N_1566,N_923);
nor U5421 (N_5421,N_4594,N_4038);
or U5422 (N_5422,N_1049,N_3527);
and U5423 (N_5423,N_2018,N_1381);
nor U5424 (N_5424,N_720,N_1530);
xor U5425 (N_5425,N_729,N_908);
and U5426 (N_5426,N_3220,N_4555);
nor U5427 (N_5427,N_2228,N_3743);
nand U5428 (N_5428,N_1899,N_79);
or U5429 (N_5429,N_2822,N_4417);
and U5430 (N_5430,N_3212,N_2197);
and U5431 (N_5431,N_3953,N_4568);
or U5432 (N_5432,N_949,N_3368);
nor U5433 (N_5433,N_2889,N_3872);
nand U5434 (N_5434,N_2536,N_2977);
and U5435 (N_5435,N_3303,N_2327);
nand U5436 (N_5436,N_3486,N_4386);
and U5437 (N_5437,N_4473,N_1040);
and U5438 (N_5438,N_3301,N_4211);
or U5439 (N_5439,N_280,N_2512);
and U5440 (N_5440,N_4667,N_3611);
and U5441 (N_5441,N_1075,N_4892);
nand U5442 (N_5442,N_4830,N_1508);
nor U5443 (N_5443,N_4291,N_4711);
or U5444 (N_5444,N_1483,N_1397);
or U5445 (N_5445,N_508,N_2564);
xor U5446 (N_5446,N_3156,N_3514);
nor U5447 (N_5447,N_4376,N_172);
nor U5448 (N_5448,N_3752,N_3408);
xnor U5449 (N_5449,N_4990,N_310);
and U5450 (N_5450,N_2166,N_1014);
or U5451 (N_5451,N_4333,N_1713);
nand U5452 (N_5452,N_3943,N_1689);
nand U5453 (N_5453,N_2490,N_3447);
nor U5454 (N_5454,N_3708,N_522);
or U5455 (N_5455,N_1309,N_3463);
nor U5456 (N_5456,N_1470,N_4183);
and U5457 (N_5457,N_2943,N_2466);
and U5458 (N_5458,N_2353,N_3137);
or U5459 (N_5459,N_3362,N_4727);
xor U5460 (N_5460,N_4890,N_4833);
and U5461 (N_5461,N_585,N_1775);
nor U5462 (N_5462,N_478,N_4530);
nor U5463 (N_5463,N_2015,N_471);
nor U5464 (N_5464,N_797,N_878);
nand U5465 (N_5465,N_3521,N_1875);
or U5466 (N_5466,N_2683,N_1533);
nor U5467 (N_5467,N_3629,N_3506);
or U5468 (N_5468,N_830,N_1831);
xnor U5469 (N_5469,N_3651,N_2747);
nand U5470 (N_5470,N_415,N_2314);
or U5471 (N_5471,N_4595,N_938);
and U5472 (N_5472,N_4648,N_2551);
nand U5473 (N_5473,N_1790,N_1068);
and U5474 (N_5474,N_1687,N_2582);
nand U5475 (N_5475,N_3060,N_2476);
nand U5476 (N_5476,N_2226,N_3382);
and U5477 (N_5477,N_610,N_2665);
nand U5478 (N_5478,N_4367,N_2243);
nand U5479 (N_5479,N_2351,N_1003);
nor U5480 (N_5480,N_4,N_3097);
and U5481 (N_5481,N_261,N_3547);
or U5482 (N_5482,N_2207,N_2222);
and U5483 (N_5483,N_2024,N_2614);
nor U5484 (N_5484,N_1567,N_3824);
and U5485 (N_5485,N_1484,N_2517);
and U5486 (N_5486,N_4972,N_3859);
and U5487 (N_5487,N_4653,N_2980);
xnor U5488 (N_5488,N_490,N_3026);
nand U5489 (N_5489,N_4630,N_1796);
nor U5490 (N_5490,N_1902,N_1881);
nor U5491 (N_5491,N_1791,N_3713);
nand U5492 (N_5492,N_767,N_2696);
nand U5493 (N_5493,N_2495,N_1812);
nor U5494 (N_5494,N_283,N_2905);
xnor U5495 (N_5495,N_1417,N_3829);
nand U5496 (N_5496,N_2076,N_2450);
xor U5497 (N_5497,N_3369,N_3451);
xnor U5498 (N_5498,N_2998,N_4395);
or U5499 (N_5499,N_185,N_3319);
or U5500 (N_5500,N_3318,N_867);
xor U5501 (N_5501,N_2471,N_2573);
nor U5502 (N_5502,N_2151,N_1870);
and U5503 (N_5503,N_315,N_2283);
nor U5504 (N_5504,N_3154,N_3268);
nand U5505 (N_5505,N_4844,N_4250);
and U5506 (N_5506,N_3870,N_431);
or U5507 (N_5507,N_3726,N_1835);
or U5508 (N_5508,N_2405,N_3842);
nor U5509 (N_5509,N_4611,N_2375);
nor U5510 (N_5510,N_260,N_2132);
xor U5511 (N_5511,N_816,N_1061);
nor U5512 (N_5512,N_4524,N_1188);
nor U5513 (N_5513,N_609,N_4351);
nand U5514 (N_5514,N_2926,N_2245);
xor U5515 (N_5515,N_4399,N_1453);
xor U5516 (N_5516,N_2852,N_378);
and U5517 (N_5517,N_548,N_4848);
nand U5518 (N_5518,N_1751,N_3917);
nor U5519 (N_5519,N_1443,N_746);
or U5520 (N_5520,N_788,N_793);
xor U5521 (N_5521,N_154,N_2057);
nand U5522 (N_5522,N_2419,N_3498);
or U5523 (N_5523,N_972,N_888);
or U5524 (N_5524,N_1154,N_2702);
or U5525 (N_5525,N_4498,N_352);
xnor U5526 (N_5526,N_4317,N_2116);
or U5527 (N_5527,N_3241,N_2721);
nand U5528 (N_5528,N_1668,N_1391);
nand U5529 (N_5529,N_1763,N_1210);
and U5530 (N_5530,N_441,N_3690);
and U5531 (N_5531,N_2541,N_1903);
nand U5532 (N_5532,N_2109,N_1252);
and U5533 (N_5533,N_2848,N_1324);
xor U5534 (N_5534,N_981,N_3452);
nand U5535 (N_5535,N_1755,N_3847);
or U5536 (N_5536,N_1167,N_4180);
or U5537 (N_5537,N_4637,N_228);
xor U5538 (N_5538,N_982,N_2603);
or U5539 (N_5539,N_4357,N_3908);
xor U5540 (N_5540,N_252,N_1954);
nor U5541 (N_5541,N_4878,N_1797);
or U5542 (N_5542,N_54,N_4913);
xor U5543 (N_5543,N_1432,N_4850);
nor U5544 (N_5544,N_3862,N_716);
xor U5545 (N_5545,N_2454,N_2139);
or U5546 (N_5546,N_3354,N_581);
or U5547 (N_5547,N_3226,N_712);
xnor U5548 (N_5548,N_1245,N_3942);
nand U5549 (N_5549,N_3780,N_4419);
or U5550 (N_5550,N_1487,N_2818);
nor U5551 (N_5551,N_3134,N_3613);
nor U5552 (N_5552,N_334,N_2389);
or U5553 (N_5553,N_2781,N_3775);
and U5554 (N_5554,N_3457,N_575);
nor U5555 (N_5555,N_1151,N_3833);
xnor U5556 (N_5556,N_1939,N_3040);
and U5557 (N_5557,N_3128,N_2066);
xnor U5558 (N_5558,N_3905,N_3115);
or U5559 (N_5559,N_4805,N_2347);
xnor U5560 (N_5560,N_864,N_2074);
nor U5561 (N_5561,N_2303,N_2584);
or U5562 (N_5562,N_274,N_282);
and U5563 (N_5563,N_4271,N_2585);
and U5564 (N_5564,N_3667,N_4361);
xnor U5565 (N_5565,N_779,N_3855);
nand U5566 (N_5566,N_1540,N_4974);
nor U5567 (N_5567,N_4025,N_2558);
nand U5568 (N_5568,N_2379,N_4451);
and U5569 (N_5569,N_950,N_733);
xnor U5570 (N_5570,N_1331,N_1590);
or U5571 (N_5571,N_1630,N_484);
nand U5572 (N_5572,N_4997,N_3865);
or U5573 (N_5573,N_1278,N_1216);
nor U5574 (N_5574,N_3993,N_4665);
nand U5575 (N_5575,N_4121,N_3251);
xnor U5576 (N_5576,N_3496,N_827);
and U5577 (N_5577,N_2596,N_2482);
nand U5578 (N_5578,N_4944,N_97);
nor U5579 (N_5579,N_2492,N_3099);
nor U5580 (N_5580,N_4401,N_3090);
and U5581 (N_5581,N_2048,N_2060);
and U5582 (N_5582,N_1502,N_4029);
nor U5583 (N_5583,N_2346,N_4606);
or U5584 (N_5584,N_29,N_2298);
nor U5585 (N_5585,N_3952,N_4301);
nand U5586 (N_5586,N_774,N_1307);
nand U5587 (N_5587,N_688,N_2268);
and U5588 (N_5588,N_1145,N_612);
or U5589 (N_5589,N_2153,N_1964);
nand U5590 (N_5590,N_1160,N_3494);
xnor U5591 (N_5591,N_2550,N_1558);
nand U5592 (N_5592,N_2644,N_389);
or U5593 (N_5593,N_676,N_3483);
xnor U5594 (N_5594,N_901,N_411);
nor U5595 (N_5595,N_1239,N_152);
and U5596 (N_5596,N_4358,N_3327);
or U5597 (N_5597,N_479,N_1007);
and U5598 (N_5598,N_3877,N_2962);
nor U5599 (N_5599,N_4175,N_1600);
xnor U5600 (N_5600,N_2131,N_3795);
or U5601 (N_5601,N_3302,N_1229);
nand U5602 (N_5602,N_541,N_502);
nor U5603 (N_5603,N_3967,N_4262);
and U5604 (N_5604,N_2927,N_473);
or U5605 (N_5605,N_3586,N_1130);
nand U5606 (N_5606,N_4618,N_2894);
nor U5607 (N_5607,N_1393,N_3228);
or U5608 (N_5608,N_23,N_2746);
nor U5609 (N_5609,N_3171,N_3662);
nand U5610 (N_5610,N_2875,N_2616);
nor U5611 (N_5611,N_4073,N_2844);
xnor U5612 (N_5612,N_4170,N_295);
and U5613 (N_5613,N_625,N_844);
nand U5614 (N_5614,N_2723,N_3088);
nand U5615 (N_5615,N_2469,N_2480);
or U5616 (N_5616,N_452,N_1058);
xor U5617 (N_5617,N_3356,N_2533);
xnor U5618 (N_5618,N_3074,N_1128);
xor U5619 (N_5619,N_2096,N_3010);
nor U5620 (N_5620,N_3315,N_4859);
or U5621 (N_5621,N_1941,N_3602);
or U5622 (N_5622,N_2506,N_4845);
or U5623 (N_5623,N_4704,N_2065);
nand U5624 (N_5624,N_3147,N_2310);
nand U5625 (N_5625,N_1728,N_423);
and U5626 (N_5626,N_1427,N_2983);
and U5627 (N_5627,N_3704,N_1682);
nand U5628 (N_5628,N_1051,N_2870);
nor U5629 (N_5629,N_4740,N_3329);
and U5630 (N_5630,N_3309,N_4129);
or U5631 (N_5631,N_3348,N_2749);
nand U5632 (N_5632,N_1168,N_2843);
nor U5633 (N_5633,N_4336,N_1901);
nor U5634 (N_5634,N_552,N_2762);
nand U5635 (N_5635,N_3898,N_2354);
and U5636 (N_5636,N_3262,N_2373);
nor U5637 (N_5637,N_2549,N_330);
and U5638 (N_5638,N_248,N_537);
nor U5639 (N_5639,N_3814,N_57);
nand U5640 (N_5640,N_822,N_311);
and U5641 (N_5641,N_4801,N_3840);
or U5642 (N_5642,N_2019,N_963);
and U5643 (N_5643,N_371,N_3677);
and U5644 (N_5644,N_4671,N_3359);
or U5645 (N_5645,N_557,N_3051);
and U5646 (N_5646,N_772,N_592);
and U5647 (N_5647,N_3465,N_4792);
and U5648 (N_5648,N_4240,N_3502);
and U5649 (N_5649,N_92,N_638);
nor U5650 (N_5650,N_19,N_4938);
nor U5651 (N_5651,N_2935,N_2638);
nor U5652 (N_5652,N_3034,N_2119);
nand U5653 (N_5653,N_367,N_4252);
xor U5654 (N_5654,N_414,N_4731);
xnor U5655 (N_5655,N_2145,N_3642);
and U5656 (N_5656,N_2785,N_1782);
xnor U5657 (N_5657,N_1349,N_3109);
nand U5658 (N_5658,N_630,N_139);
nand U5659 (N_5659,N_1480,N_3282);
and U5660 (N_5660,N_3711,N_108);
nor U5661 (N_5661,N_3413,N_951);
nand U5662 (N_5662,N_3723,N_2576);
nand U5663 (N_5663,N_2892,N_1937);
nand U5664 (N_5664,N_646,N_2256);
nor U5665 (N_5665,N_3673,N_4131);
and U5666 (N_5666,N_3381,N_2000);
or U5667 (N_5667,N_1056,N_2501);
or U5668 (N_5668,N_1082,N_754);
or U5669 (N_5669,N_1799,N_4761);
nand U5670 (N_5670,N_3092,N_2462);
and U5671 (N_5671,N_920,N_2437);
nand U5672 (N_5672,N_2122,N_4577);
nand U5673 (N_5673,N_396,N_2662);
xnor U5674 (N_5674,N_4910,N_2896);
and U5675 (N_5675,N_521,N_861);
xnor U5676 (N_5676,N_2787,N_225);
nand U5677 (N_5677,N_2525,N_1832);
and U5678 (N_5678,N_1411,N_4494);
xnor U5679 (N_5679,N_20,N_4404);
or U5680 (N_5680,N_4365,N_4694);
or U5681 (N_5681,N_278,N_1771);
and U5682 (N_5682,N_887,N_3473);
or U5683 (N_5683,N_741,N_1457);
nand U5684 (N_5684,N_3947,N_2493);
nor U5685 (N_5685,N_1308,N_4098);
nand U5686 (N_5686,N_2054,N_1435);
and U5687 (N_5687,N_1738,N_4605);
nand U5688 (N_5688,N_1136,N_1066);
and U5689 (N_5689,N_2681,N_1500);
nor U5690 (N_5690,N_2022,N_88);
nor U5691 (N_5691,N_2859,N_2409);
or U5692 (N_5692,N_4284,N_1222);
and U5693 (N_5693,N_2874,N_4418);
or U5694 (N_5694,N_1929,N_4318);
nor U5695 (N_5695,N_2956,N_316);
xor U5696 (N_5696,N_1089,N_760);
or U5697 (N_5697,N_2004,N_67);
nand U5698 (N_5698,N_1026,N_1376);
nand U5699 (N_5699,N_2453,N_1259);
nor U5700 (N_5700,N_4741,N_482);
and U5701 (N_5701,N_4236,N_4070);
nor U5702 (N_5702,N_3478,N_4448);
nand U5703 (N_5703,N_4055,N_2857);
and U5704 (N_5704,N_2629,N_3528);
or U5705 (N_5705,N_2615,N_865);
xnor U5706 (N_5706,N_2042,N_4380);
nand U5707 (N_5707,N_2846,N_4645);
xnor U5708 (N_5708,N_2691,N_34);
nand U5709 (N_5709,N_1640,N_3431);
xnor U5710 (N_5710,N_1429,N_3652);
nand U5711 (N_5711,N_1756,N_4837);
xnor U5712 (N_5712,N_4735,N_4866);
nor U5713 (N_5713,N_3188,N_2979);
nor U5714 (N_5714,N_4970,N_1400);
nand U5715 (N_5715,N_2329,N_3202);
xnor U5716 (N_5716,N_223,N_1827);
xor U5717 (N_5717,N_4638,N_4107);
or U5718 (N_5718,N_1196,N_4341);
and U5719 (N_5719,N_2940,N_2321);
and U5720 (N_5720,N_2513,N_980);
or U5721 (N_5721,N_1838,N_4888);
xnor U5722 (N_5722,N_4692,N_4708);
and U5723 (N_5723,N_328,N_2208);
and U5724 (N_5724,N_523,N_4533);
xor U5725 (N_5725,N_3779,N_127);
nand U5726 (N_5726,N_1615,N_3567);
nand U5727 (N_5727,N_1930,N_4945);
or U5728 (N_5728,N_1759,N_4396);
nand U5729 (N_5729,N_3838,N_4908);
nand U5730 (N_5730,N_1117,N_4228);
nor U5731 (N_5731,N_607,N_565);
or U5732 (N_5732,N_15,N_4634);
and U5733 (N_5733,N_1680,N_2124);
nand U5734 (N_5734,N_3474,N_4214);
or U5735 (N_5735,N_4522,N_3561);
nand U5736 (N_5736,N_818,N_4311);
nor U5737 (N_5737,N_2945,N_4063);
nand U5738 (N_5738,N_2736,N_1842);
xor U5739 (N_5739,N_2704,N_858);
nor U5740 (N_5740,N_388,N_3793);
nand U5741 (N_5741,N_3138,N_4369);
and U5742 (N_5742,N_1310,N_4201);
nor U5743 (N_5743,N_1138,N_3996);
xnor U5744 (N_5744,N_3298,N_2147);
and U5745 (N_5745,N_4930,N_3678);
xnor U5746 (N_5746,N_2922,N_3141);
and U5747 (N_5747,N_4013,N_1266);
nor U5748 (N_5748,N_4342,N_195);
nand U5749 (N_5749,N_3213,N_2701);
and U5750 (N_5750,N_76,N_3605);
xnor U5751 (N_5751,N_1701,N_782);
or U5752 (N_5752,N_1826,N_4221);
and U5753 (N_5753,N_2790,N_2880);
xnor U5754 (N_5754,N_1591,N_1588);
or U5755 (N_5755,N_1090,N_3267);
nand U5756 (N_5756,N_3977,N_2739);
nand U5757 (N_5757,N_3122,N_4383);
and U5758 (N_5758,N_466,N_4220);
or U5759 (N_5759,N_2143,N_1192);
nand U5760 (N_5760,N_1976,N_2380);
nand U5761 (N_5761,N_1535,N_2397);
nor U5762 (N_5762,N_2242,N_2158);
xnor U5763 (N_5763,N_983,N_2775);
or U5764 (N_5764,N_991,N_1616);
xnor U5765 (N_5765,N_4144,N_4870);
and U5766 (N_5766,N_4458,N_555);
nand U5767 (N_5767,N_1772,N_934);
and U5768 (N_5768,N_1274,N_2239);
nor U5769 (N_5769,N_3564,N_1744);
nand U5770 (N_5770,N_4590,N_5);
or U5771 (N_5771,N_3760,N_3254);
nor U5772 (N_5772,N_4804,N_1663);
or U5773 (N_5773,N_539,N_3508);
and U5774 (N_5774,N_4853,N_2254);
nand U5775 (N_5775,N_904,N_109);
nor U5776 (N_5776,N_2823,N_4915);
nand U5777 (N_5777,N_1031,N_475);
and U5778 (N_5778,N_1409,N_1573);
or U5779 (N_5779,N_2431,N_3694);
nor U5780 (N_5780,N_3211,N_4790);
nand U5781 (N_5781,N_777,N_1510);
nor U5782 (N_5782,N_4674,N_2199);
and U5783 (N_5783,N_684,N_314);
and U5784 (N_5784,N_2626,N_4531);
nor U5785 (N_5785,N_4068,N_3406);
and U5786 (N_5786,N_749,N_3194);
and U5787 (N_5787,N_3028,N_3265);
xor U5788 (N_5788,N_652,N_1076);
and U5789 (N_5789,N_3367,N_969);
xor U5790 (N_5790,N_1108,N_996);
or U5791 (N_5791,N_1712,N_738);
nand U5792 (N_5792,N_2496,N_2225);
nand U5793 (N_5793,N_886,N_3945);
and U5794 (N_5794,N_3819,N_2579);
nor U5795 (N_5795,N_2881,N_2967);
and U5796 (N_5796,N_4991,N_1898);
nand U5797 (N_5797,N_4897,N_1700);
or U5798 (N_5798,N_2631,N_224);
or U5799 (N_5799,N_1762,N_4736);
or U5800 (N_5800,N_1194,N_1577);
nand U5801 (N_5801,N_4373,N_3396);
nand U5802 (N_5802,N_1932,N_1465);
xnor U5803 (N_5803,N_2518,N_470);
xor U5804 (N_5804,N_2342,N_2673);
nor U5805 (N_5805,N_725,N_4867);
and U5806 (N_5806,N_3744,N_417);
nand U5807 (N_5807,N_300,N_4709);
xor U5808 (N_5808,N_3163,N_2649);
nor U5809 (N_5809,N_1178,N_817);
nand U5810 (N_5810,N_2965,N_3289);
nand U5811 (N_5811,N_4981,N_1494);
xnor U5812 (N_5812,N_2305,N_4402);
xor U5813 (N_5813,N_4135,N_116);
xnor U5814 (N_5814,N_4701,N_975);
or U5815 (N_5815,N_4552,N_931);
or U5816 (N_5816,N_469,N_1784);
and U5817 (N_5817,N_4542,N_465);
nor U5818 (N_5818,N_1318,N_2386);
and U5819 (N_5819,N_3180,N_1830);
nor U5820 (N_5820,N_2272,N_1008);
nor U5821 (N_5821,N_1872,N_3541);
and U5822 (N_5822,N_4209,N_2302);
xor U5823 (N_5823,N_3983,N_3971);
nand U5824 (N_5824,N_1708,N_4314);
or U5825 (N_5825,N_1095,N_2033);
and U5826 (N_5826,N_4040,N_4036);
nor U5827 (N_5827,N_3618,N_4700);
nor U5828 (N_5828,N_668,N_3951);
xnor U5829 (N_5829,N_1120,N_1704);
or U5830 (N_5830,N_2581,N_3270);
or U5831 (N_5831,N_203,N_3052);
or U5832 (N_5832,N_745,N_3706);
xor U5833 (N_5833,N_2110,N_3648);
nor U5834 (N_5834,N_2909,N_4703);
and U5835 (N_5835,N_2422,N_358);
xnor U5836 (N_5836,N_2087,N_87);
or U5837 (N_5837,N_3534,N_4007);
or U5838 (N_5838,N_2538,N_1099);
or U5839 (N_5839,N_359,N_3692);
xnor U5840 (N_5840,N_4716,N_305);
and U5841 (N_5841,N_4484,N_2258);
nand U5842 (N_5842,N_100,N_1340);
nand U5843 (N_5843,N_4001,N_2861);
nand U5844 (N_5844,N_2703,N_3119);
nand U5845 (N_5845,N_4686,N_3231);
or U5846 (N_5846,N_3191,N_3867);
nand U5847 (N_5847,N_472,N_4347);
or U5848 (N_5848,N_239,N_4503);
xor U5849 (N_5849,N_1647,N_1276);
and U5850 (N_5850,N_3974,N_4492);
nand U5851 (N_5851,N_164,N_1326);
xor U5852 (N_5852,N_4005,N_404);
and U5853 (N_5853,N_1419,N_25);
nand U5854 (N_5854,N_3661,N_1970);
nand U5855 (N_5855,N_4069,N_550);
nor U5856 (N_5856,N_2366,N_50);
nor U5857 (N_5857,N_1509,N_3434);
or U5858 (N_5858,N_2643,N_1544);
or U5859 (N_5859,N_2914,N_917);
or U5860 (N_5860,N_4572,N_2942);
nand U5861 (N_5861,N_1907,N_4075);
nand U5862 (N_5862,N_176,N_93);
nand U5863 (N_5863,N_4309,N_1905);
nor U5864 (N_5864,N_444,N_3403);
xor U5865 (N_5865,N_1067,N_528);
nand U5866 (N_5866,N_1710,N_1915);
xnor U5867 (N_5867,N_1859,N_582);
or U5868 (N_5868,N_3279,N_2319);
nor U5869 (N_5869,N_1884,N_4507);
or U5870 (N_5870,N_4045,N_4722);
nand U5871 (N_5871,N_48,N_3676);
xnor U5872 (N_5872,N_2651,N_4900);
or U5873 (N_5873,N_3655,N_4539);
or U5874 (N_5874,N_2877,N_497);
nor U5875 (N_5875,N_3086,N_3783);
xnor U5876 (N_5876,N_3513,N_998);
or U5877 (N_5877,N_4593,N_3557);
and U5878 (N_5878,N_2191,N_2677);
nand U5879 (N_5879,N_1060,N_3728);
xnor U5880 (N_5880,N_4172,N_1822);
nand U5881 (N_5881,N_436,N_900);
xor U5882 (N_5882,N_757,N_1676);
nor U5883 (N_5883,N_2851,N_4663);
or U5884 (N_5884,N_394,N_2697);
nor U5885 (N_5885,N_645,N_1319);
xnor U5886 (N_5886,N_4008,N_3718);
and U5887 (N_5887,N_3853,N_4168);
and U5888 (N_5888,N_961,N_3236);
xnor U5889 (N_5889,N_1639,N_3956);
nor U5890 (N_5890,N_2007,N_3595);
nor U5891 (N_5891,N_3275,N_1620);
and U5892 (N_5892,N_4403,N_2455);
nor U5893 (N_5893,N_4669,N_2193);
or U5894 (N_5894,N_2916,N_3846);
nor U5895 (N_5895,N_2137,N_2063);
nand U5896 (N_5896,N_2179,N_64);
nand U5897 (N_5897,N_3146,N_932);
nor U5898 (N_5898,N_850,N_2803);
nor U5899 (N_5899,N_658,N_1971);
and U5900 (N_5900,N_856,N_1645);
and U5901 (N_5901,N_242,N_1815);
or U5902 (N_5902,N_4176,N_2817);
and U5903 (N_5903,N_3370,N_407);
nand U5904 (N_5904,N_2174,N_1793);
or U5905 (N_5905,N_2919,N_1774);
and U5906 (N_5906,N_2280,N_3054);
nand U5907 (N_5907,N_3687,N_1652);
nor U5908 (N_5908,N_3959,N_1115);
or U5909 (N_5909,N_134,N_3940);
xnor U5910 (N_5910,N_3178,N_4389);
or U5911 (N_5911,N_1503,N_1693);
or U5912 (N_5912,N_1557,N_2508);
xnor U5913 (N_5913,N_4902,N_4518);
xor U5914 (N_5914,N_1968,N_4658);
nand U5915 (N_5915,N_2318,N_1034);
and U5916 (N_5916,N_4059,N_3429);
or U5917 (N_5917,N_1162,N_1943);
or U5918 (N_5918,N_3563,N_199);
nor U5919 (N_5919,N_4508,N_1856);
or U5920 (N_5920,N_1321,N_3505);
or U5921 (N_5921,N_3133,N_4133);
nand U5922 (N_5922,N_289,N_4786);
or U5923 (N_5923,N_2062,N_4282);
or U5924 (N_5924,N_2939,N_1742);
nand U5925 (N_5925,N_2505,N_1656);
nor U5926 (N_5926,N_2589,N_1949);
nor U5927 (N_5927,N_4023,N_1092);
or U5928 (N_5928,N_3699,N_3792);
nor U5929 (N_5929,N_674,N_4491);
xor U5930 (N_5930,N_1582,N_410);
nor U5931 (N_5931,N_2654,N_1896);
xor U5932 (N_5932,N_1910,N_1187);
xnor U5933 (N_5933,N_1786,N_331);
or U5934 (N_5934,N_39,N_4368);
nor U5935 (N_5935,N_106,N_4226);
nor U5936 (N_5936,N_4247,N_269);
or U5937 (N_5937,N_3189,N_2489);
or U5938 (N_5938,N_1604,N_4880);
or U5939 (N_5939,N_4039,N_2953);
and U5940 (N_5940,N_68,N_2808);
or U5941 (N_5941,N_1918,N_4928);
xnor U5942 (N_5942,N_4757,N_791);
or U5943 (N_5943,N_3307,N_2491);
xnor U5944 (N_5944,N_1542,N_3278);
and U5945 (N_5945,N_4181,N_4656);
and U5946 (N_5946,N_4292,N_814);
and U5947 (N_5947,N_2809,N_4120);
or U5948 (N_5948,N_2255,N_60);
xnor U5949 (N_5949,N_3910,N_1780);
nand U5950 (N_5950,N_2370,N_1659);
xnor U5951 (N_5951,N_1379,N_63);
xor U5952 (N_5952,N_45,N_1358);
xor U5953 (N_5953,N_1956,N_1282);
nand U5954 (N_5954,N_3544,N_3358);
nand U5955 (N_5955,N_1811,N_3384);
nor U5956 (N_5956,N_1218,N_4784);
and U5957 (N_5957,N_2842,N_232);
xnor U5958 (N_5958,N_3196,N_2836);
nand U5959 (N_5959,N_1841,N_3594);
xnor U5960 (N_5960,N_3125,N_1179);
nand U5961 (N_5961,N_212,N_477);
xnor U5962 (N_5962,N_11,N_4955);
nor U5963 (N_5963,N_2918,N_3509);
and U5964 (N_5964,N_3632,N_3438);
and U5965 (N_5965,N_2300,N_1532);
nand U5966 (N_5966,N_2290,N_3963);
and U5967 (N_5967,N_4195,N_4721);
nor U5968 (N_5968,N_1198,N_1238);
or U5969 (N_5969,N_2499,N_2178);
and U5970 (N_5970,N_1507,N_3094);
xor U5971 (N_5971,N_4796,N_244);
nand U5972 (N_5972,N_1785,N_18);
nor U5973 (N_5973,N_1757,N_498);
and U5974 (N_5974,N_1633,N_1922);
nor U5975 (N_5975,N_629,N_2414);
and U5976 (N_5976,N_869,N_2073);
xor U5977 (N_5977,N_3918,N_2211);
nand U5978 (N_5978,N_1323,N_4623);
or U5979 (N_5979,N_570,N_4780);
and U5980 (N_5980,N_3336,N_438);
nand U5981 (N_5981,N_1525,N_936);
xnor U5982 (N_5982,N_2442,N_3045);
nor U5983 (N_5983,N_255,N_1189);
nand U5984 (N_5984,N_41,N_126);
nand U5985 (N_5985,N_3707,N_2292);
or U5986 (N_5986,N_1963,N_2883);
or U5987 (N_5987,N_2399,N_715);
and U5988 (N_5988,N_4520,N_3753);
xnor U5989 (N_5989,N_3084,N_462);
and U5990 (N_5990,N_4788,N_3471);
and U5991 (N_5991,N_1129,N_3304);
xor U5992 (N_5992,N_2171,N_3553);
and U5993 (N_5993,N_3415,N_3574);
nand U5994 (N_5994,N_2989,N_451);
nor U5995 (N_5995,N_317,N_4387);
nand U5996 (N_5996,N_1125,N_2656);
nor U5997 (N_5997,N_4217,N_4815);
and U5998 (N_5998,N_4469,N_1873);
or U5999 (N_5999,N_1054,N_1079);
and U6000 (N_6000,N_2794,N_4566);
or U6001 (N_6001,N_2154,N_2755);
and U6002 (N_6002,N_1670,N_4052);
xor U6003 (N_6003,N_1935,N_3776);
nor U6004 (N_6004,N_114,N_3705);
or U6005 (N_6005,N_3355,N_2598);
xor U6006 (N_6006,N_3849,N_4994);
and U6007 (N_6007,N_182,N_2220);
nand U6008 (N_6008,N_1865,N_2456);
nand U6009 (N_6009,N_4398,N_4431);
or U6010 (N_6010,N_2825,N_4083);
and U6011 (N_6011,N_743,N_924);
nand U6012 (N_6012,N_1320,N_3572);
nand U6013 (N_6013,N_608,N_976);
and U6014 (N_6014,N_4751,N_701);
nand U6015 (N_6015,N_690,N_1408);
xnor U6016 (N_6016,N_2412,N_2344);
nand U6017 (N_6017,N_1071,N_2032);
and U6018 (N_6018,N_3409,N_2552);
nand U6019 (N_6019,N_634,N_3394);
nor U6020 (N_6020,N_2999,N_4832);
and U6021 (N_6021,N_3145,N_510);
and U6022 (N_6022,N_3670,N_853);
nor U6023 (N_6023,N_3011,N_4949);
and U6024 (N_6024,N_4084,N_4281);
nand U6025 (N_6025,N_4954,N_1171);
nand U6026 (N_6026,N_2827,N_1232);
xor U6027 (N_6027,N_3766,N_3797);
nor U6028 (N_6028,N_4125,N_249);
xor U6029 (N_6029,N_602,N_4670);
xor U6030 (N_6030,N_2334,N_928);
and U6031 (N_6031,N_2686,N_1908);
xor U6032 (N_6032,N_2103,N_2043);
xnor U6033 (N_6033,N_3198,N_1140);
xnor U6034 (N_6034,N_1388,N_2970);
and U6035 (N_6035,N_855,N_243);
or U6036 (N_6036,N_3308,N_4020);
or U6037 (N_6037,N_2500,N_579);
nand U6038 (N_6038,N_3988,N_1743);
or U6039 (N_6039,N_1916,N_2411);
or U6040 (N_6040,N_847,N_691);
and U6041 (N_6041,N_507,N_3617);
nand U6042 (N_6042,N_4015,N_3243);
xor U6043 (N_6043,N_1455,N_3679);
xor U6044 (N_6044,N_2238,N_2937);
nor U6045 (N_6045,N_1993,N_1005);
or U6046 (N_6046,N_2262,N_2140);
xor U6047 (N_6047,N_935,N_2792);
or U6048 (N_6048,N_17,N_2136);
or U6049 (N_6049,N_2013,N_1343);
and U6050 (N_6050,N_3854,N_3997);
or U6051 (N_6051,N_226,N_512);
nand U6052 (N_6052,N_2932,N_3630);
nor U6053 (N_6053,N_2912,N_3175);
and U6054 (N_6054,N_576,N_3069);
or U6055 (N_6055,N_1062,N_3897);
nand U6056 (N_6056,N_1116,N_808);
or U6057 (N_6057,N_1737,N_1110);
nor U6058 (N_6058,N_2218,N_4730);
xor U6059 (N_6059,N_454,N_3741);
nand U6060 (N_6060,N_1190,N_1);
nand U6061 (N_6061,N_4081,N_4666);
xor U6062 (N_6062,N_1834,N_4647);
nand U6063 (N_6063,N_1396,N_3187);
or U6064 (N_6064,N_457,N_2613);
nand U6065 (N_6065,N_4909,N_4327);
xor U6066 (N_6066,N_3423,N_2478);
nand U6067 (N_6067,N_4338,N_4116);
or U6068 (N_6068,N_4839,N_3317);
and U6069 (N_6069,N_3246,N_2544);
nand U6070 (N_6070,N_2797,N_1977);
and U6071 (N_6071,N_3803,N_4329);
nor U6072 (N_6072,N_3560,N_4602);
and U6073 (N_6073,N_3063,N_2960);
and U6074 (N_6074,N_876,N_4461);
nand U6075 (N_6075,N_2046,N_3295);
nor U6076 (N_6076,N_1860,N_463);
nand U6077 (N_6077,N_2769,N_1094);
or U6078 (N_6078,N_2650,N_1339);
nor U6079 (N_6079,N_2247,N_1037);
nand U6080 (N_6080,N_4472,N_1677);
and U6081 (N_6081,N_2250,N_3522);
nand U6082 (N_6082,N_3089,N_3827);
or U6083 (N_6083,N_2772,N_1596);
or U6084 (N_6084,N_621,N_1776);
xnor U6085 (N_6085,N_4726,N_4824);
nor U6086 (N_6086,N_3135,N_1541);
nor U6087 (N_6087,N_4806,N_657);
or U6088 (N_6088,N_4197,N_16);
nand U6089 (N_6089,N_1599,N_1642);
nand U6090 (N_6090,N_2494,N_483);
nor U6091 (N_6091,N_499,N_4356);
and U6092 (N_6092,N_4456,N_2884);
nor U6093 (N_6093,N_987,N_2531);
nor U6094 (N_6094,N_3042,N_1948);
and U6095 (N_6095,N_4627,N_2964);
and U6096 (N_6096,N_1267,N_1482);
or U6097 (N_6097,N_1176,N_4381);
or U6098 (N_6098,N_2460,N_4745);
nor U6099 (N_6099,N_2561,N_732);
xor U6100 (N_6100,N_3095,N_2948);
xor U6101 (N_6101,N_4838,N_4774);
or U6102 (N_6102,N_4321,N_2811);
or U6103 (N_6103,N_509,N_1933);
xnor U6104 (N_6104,N_2717,N_1371);
nand U6105 (N_6105,N_2692,N_1368);
and U6106 (N_6106,N_1953,N_3682);
nor U6107 (N_6107,N_2707,N_1059);
or U6108 (N_6108,N_4099,N_583);
or U6109 (N_6109,N_3374,N_1798);
nor U6110 (N_6110,N_1121,N_3468);
xor U6111 (N_6111,N_899,N_1224);
and U6112 (N_6112,N_3481,N_3895);
nor U6113 (N_6113,N_3271,N_2590);
xor U6114 (N_6114,N_301,N_3165);
xnor U6115 (N_6115,N_46,N_2913);
or U6116 (N_6116,N_1057,N_1147);
or U6117 (N_6117,N_1885,N_3816);
nor U6118 (N_6118,N_69,N_4439);
nor U6119 (N_6119,N_784,N_2034);
and U6120 (N_6120,N_2227,N_946);
and U6121 (N_6121,N_4769,N_3103);
nand U6122 (N_6122,N_2402,N_4043);
xor U6123 (N_6123,N_4122,N_355);
xnor U6124 (N_6124,N_3821,N_194);
xor U6125 (N_6125,N_2546,N_4505);
nor U6126 (N_6126,N_4650,N_2152);
or U6127 (N_6127,N_2996,N_1978);
xor U6128 (N_6128,N_3430,N_4348);
xor U6129 (N_6129,N_2118,N_1698);
nor U6130 (N_6130,N_1451,N_3965);
or U6131 (N_6131,N_1155,N_2734);
and U6132 (N_6132,N_401,N_3174);
and U6133 (N_6133,N_3640,N_910);
xor U6134 (N_6134,N_3868,N_3747);
and U6135 (N_6135,N_3684,N_4325);
or U6136 (N_6136,N_4179,N_4957);
xnor U6137 (N_6137,N_543,N_105);
nor U6138 (N_6138,N_4793,N_4416);
xor U6139 (N_6139,N_2316,N_755);
xor U6140 (N_6140,N_4062,N_3675);
nand U6141 (N_6141,N_4100,N_4268);
or U6142 (N_6142,N_3001,N_3195);
nand U6143 (N_6143,N_2330,N_3372);
and U6144 (N_6144,N_1874,N_4668);
nand U6145 (N_6145,N_2766,N_1818);
and U6146 (N_6146,N_4760,N_1706);
and U6147 (N_6147,N_3614,N_2868);
nand U6148 (N_6148,N_4596,N_4248);
nor U6149 (N_6149,N_2934,N_1084);
nand U6150 (N_6150,N_2301,N_3933);
nor U6151 (N_6151,N_984,N_3647);
xor U6152 (N_6152,N_2085,N_4581);
or U6153 (N_6153,N_1366,N_2133);
nor U6154 (N_6154,N_192,N_3671);
xor U6155 (N_6155,N_2872,N_3130);
xnor U6156 (N_6156,N_1637,N_4085);
or U6157 (N_6157,N_1185,N_4335);
nand U6158 (N_6158,N_1477,N_1735);
nand U6159 (N_6159,N_38,N_637);
nand U6160 (N_6160,N_1463,N_3825);
xnor U6161 (N_6161,N_357,N_2959);
nor U6162 (N_6162,N_1019,N_4953);
nand U6163 (N_6163,N_2885,N_4189);
nor U6164 (N_6164,N_4425,N_2636);
and U6165 (N_6165,N_1703,N_3786);
xnor U6166 (N_6166,N_1726,N_1719);
xnor U6167 (N_6167,N_1304,N_1864);
or U6168 (N_6168,N_2793,N_3108);
or U6169 (N_6169,N_4958,N_4010);
nand U6170 (N_6170,N_2408,N_3393);
and U6171 (N_6171,N_2477,N_580);
nand U6172 (N_6172,N_2587,N_4108);
nand U6173 (N_6173,N_836,N_2791);
and U6174 (N_6174,N_1925,N_617);
nor U6175 (N_6175,N_4187,N_2404);
or U6176 (N_6176,N_1214,N_4749);
xor U6177 (N_6177,N_1991,N_778);
or U6178 (N_6178,N_4800,N_1913);
or U6179 (N_6179,N_872,N_4114);
nand U6180 (N_6180,N_4863,N_1876);
or U6181 (N_6181,N_4130,N_2264);
nor U6182 (N_6182,N_4849,N_703);
and U6183 (N_6183,N_1819,N_918);
and U6184 (N_6184,N_4423,N_2403);
xnor U6185 (N_6185,N_1111,N_2622);
and U6186 (N_6186,N_1169,N_4808);
and U6187 (N_6187,N_1574,N_2393);
nand U6188 (N_6188,N_1805,N_3581);
nand U6189 (N_6189,N_3037,N_4041);
xor U6190 (N_6190,N_2056,N_1279);
or U6191 (N_6191,N_985,N_2947);
or U6192 (N_6192,N_426,N_1459);
and U6193 (N_6193,N_1534,N_3568);
nor U6194 (N_6194,N_4213,N_3511);
and U6195 (N_6195,N_4764,N_1390);
xnor U6196 (N_6196,N_2588,N_1917);
xor U6197 (N_6197,N_372,N_2572);
and U6198 (N_6198,N_1562,N_1270);
xnor U6199 (N_6199,N_4374,N_4767);
nor U6200 (N_6200,N_766,N_4551);
xnor U6201 (N_6201,N_1555,N_383);
nor U6202 (N_6202,N_4676,N_2805);
nor U6203 (N_6203,N_3100,N_1717);
or U6204 (N_6204,N_1286,N_773);
or U6205 (N_6205,N_1029,N_1362);
xor U6206 (N_6206,N_4390,N_2708);
xnor U6207 (N_6207,N_863,N_382);
nand U6208 (N_6208,N_4737,N_3475);
or U6209 (N_6209,N_2952,N_312);
nor U6210 (N_6210,N_4009,N_160);
and U6211 (N_6211,N_1434,N_4424);
or U6212 (N_6212,N_1931,N_3472);
nand U6213 (N_6213,N_1219,N_3176);
nor U6214 (N_6214,N_694,N_419);
xnor U6215 (N_6215,N_937,N_1447);
nor U6216 (N_6216,N_3245,N_1754);
and U6217 (N_6217,N_1437,N_1448);
xor U6218 (N_6218,N_1243,N_4723);
nand U6219 (N_6219,N_2061,N_838);
or U6220 (N_6220,N_1580,N_3491);
nor U6221 (N_6221,N_3297,N_374);
or U6222 (N_6222,N_157,N_4907);
nor U6223 (N_6223,N_3810,N_974);
nand U6224 (N_6224,N_3597,N_1624);
nor U6225 (N_6225,N_163,N_3420);
nor U6226 (N_6226,N_2902,N_3660);
xnor U6227 (N_6227,N_4090,N_4825);
or U6228 (N_6228,N_4821,N_3476);
nor U6229 (N_6229,N_4349,N_2426);
xor U6230 (N_6230,N_3041,N_3250);
nor U6231 (N_6231,N_3525,N_4275);
and U6232 (N_6232,N_3158,N_3672);
xor U6233 (N_6233,N_4048,N_2451);
nor U6234 (N_6234,N_2356,N_4264);
xor U6235 (N_6235,N_2107,N_968);
nand U6236 (N_6236,N_4985,N_2159);
nand U6237 (N_6237,N_4969,N_1529);
and U6238 (N_6238,N_4624,N_1990);
nor U6239 (N_6239,N_3342,N_4984);
xor U6240 (N_6240,N_4160,N_4919);
xor U6241 (N_6241,N_3120,N_4428);
nand U6242 (N_6242,N_1328,N_1431);
xor U6243 (N_6243,N_350,N_286);
nand U6244 (N_6244,N_3863,N_296);
or U6245 (N_6245,N_4243,N_1404);
xor U6246 (N_6246,N_3335,N_3260);
xnor U6247 (N_6247,N_4065,N_3938);
nor U6248 (N_6248,N_102,N_2634);
nor U6249 (N_6249,N_159,N_319);
nand U6250 (N_6250,N_257,N_3252);
or U6251 (N_6251,N_3177,N_4673);
nand U6252 (N_6252,N_3767,N_544);
nor U6253 (N_6253,N_4636,N_3536);
nand U6254 (N_6254,N_3621,N_4151);
and U6255 (N_6255,N_952,N_4662);
nor U6256 (N_6256,N_792,N_3999);
nor U6257 (N_6257,N_3221,N_514);
and U6258 (N_6258,N_3873,N_4759);
nor U6259 (N_6259,N_947,N_3542);
and U6260 (N_6260,N_1697,N_4580);
nor U6261 (N_6261,N_3014,N_1501);
xor U6262 (N_6262,N_1619,N_1370);
and U6263 (N_6263,N_129,N_448);
nor U6264 (N_6264,N_3049,N_4032);
nand U6265 (N_6265,N_4257,N_3880);
nand U6266 (N_6266,N_1209,N_4392);
or U6267 (N_6267,N_2398,N_3710);
or U6268 (N_6268,N_4225,N_4999);
and U6269 (N_6269,N_495,N_1801);
or U6270 (N_6270,N_3697,N_4699);
xnor U6271 (N_6271,N_4410,N_4372);
xor U6272 (N_6272,N_4305,N_3390);
and U6273 (N_6273,N_4432,N_1123);
and U6274 (N_6274,N_4346,N_2556);
and U6275 (N_6275,N_2148,N_98);
nor U6276 (N_6276,N_2931,N_84);
and U6277 (N_6277,N_1955,N_1924);
nand U6278 (N_6278,N_4468,N_2308);
nand U6279 (N_6279,N_433,N_1972);
nor U6280 (N_6280,N_2782,N_2425);
and U6281 (N_6281,N_287,N_4843);
nor U6282 (N_6282,N_4011,N_2309);
nor U6283 (N_6283,N_2821,N_3843);
and U6284 (N_6284,N_992,N_3470);
xor U6285 (N_6285,N_1412,N_4639);
xnor U6286 (N_6286,N_3957,N_4146);
nand U6287 (N_6287,N_3258,N_3046);
nor U6288 (N_6288,N_4102,N_1351);
xnor U6289 (N_6289,N_3338,N_180);
and U6290 (N_6290,N_4445,N_3492);
or U6291 (N_6291,N_1505,N_3217);
nor U6292 (N_6292,N_168,N_3206);
or U6293 (N_6293,N_166,N_763);
nand U6294 (N_6294,N_2601,N_1996);
nand U6295 (N_6295,N_4150,N_1257);
nand U6296 (N_6296,N_4858,N_4232);
and U6297 (N_6297,N_839,N_59);
xnor U6298 (N_6298,N_104,N_673);
or U6299 (N_6299,N_2679,N_1231);
xnor U6300 (N_6300,N_4810,N_2071);
xnor U6301 (N_6301,N_1356,N_406);
xor U6302 (N_6302,N_1564,N_1361);
nor U6303 (N_6303,N_1879,N_83);
or U6304 (N_6304,N_4198,N_3314);
nor U6305 (N_6305,N_1967,N_4865);
xor U6306 (N_6306,N_3875,N_3385);
or U6307 (N_6307,N_3425,N_4413);
xnor U6308 (N_6308,N_4147,N_4051);
nand U6309 (N_6309,N_3771,N_1078);
and U6310 (N_6310,N_4587,N_3091);
nor U6311 (N_6311,N_439,N_4776);
and U6312 (N_6312,N_3861,N_675);
nand U6313 (N_6313,N_3603,N_3401);
or U6314 (N_6314,N_4409,N_4797);
nand U6315 (N_6315,N_2800,N_2599);
nor U6316 (N_6316,N_4452,N_3076);
nand U6317 (N_6317,N_4664,N_1476);
and U6318 (N_6318,N_2891,N_3466);
nand U6319 (N_6319,N_78,N_4269);
xor U6320 (N_6320,N_4320,N_3524);
xnor U6321 (N_6321,N_3469,N_3969);
nand U6322 (N_6322,N_1516,N_3802);
nand U6323 (N_6323,N_1260,N_4112);
nor U6324 (N_6324,N_4097,N_4510);
and U6325 (N_6325,N_268,N_4259);
nor U6326 (N_6326,N_3341,N_1401);
nand U6327 (N_6327,N_3272,N_4298);
xor U6328 (N_6328,N_4574,N_4405);
and U6329 (N_6329,N_2897,N_3588);
or U6330 (N_6330,N_1207,N_4523);
nand U6331 (N_6331,N_4921,N_1575);
and U6332 (N_6332,N_3256,N_4330);
xnor U6333 (N_6333,N_2946,N_3975);
and U6334 (N_6334,N_4622,N_2565);
xor U6335 (N_6335,N_1716,N_3454);
and U6336 (N_6336,N_2732,N_3216);
nor U6337 (N_6337,N_2410,N_4477);
or U6338 (N_6338,N_2121,N_2864);
nor U6339 (N_6339,N_4313,N_4101);
and U6340 (N_6340,N_2289,N_3292);
and U6341 (N_6341,N_2214,N_7);
or U6342 (N_6342,N_2357,N_4621);
and U6343 (N_6343,N_4899,N_2716);
and U6344 (N_6344,N_594,N_4184);
nor U6345 (N_6345,N_4435,N_173);
nand U6346 (N_6346,N_590,N_1556);
nand U6347 (N_6347,N_3691,N_4174);
and U6348 (N_6348,N_518,N_2653);
nor U6349 (N_6349,N_1655,N_1895);
nand U6350 (N_6350,N_2548,N_1569);
nor U6351 (N_6351,N_4724,N_2571);
and U6352 (N_6352,N_391,N_4943);
xor U6353 (N_6353,N_567,N_3657);
nor U6354 (N_6354,N_1184,N_146);
nand U6355 (N_6355,N_277,N_4649);
nor U6356 (N_6356,N_66,N_130);
xnor U6357 (N_6357,N_450,N_14);
and U6358 (N_6358,N_4681,N_2763);
xnor U6359 (N_6359,N_4297,N_4560);
and U6360 (N_6360,N_3685,N_3774);
xnor U6361 (N_6361,N_4732,N_4573);
nor U6362 (N_6362,N_1514,N_4237);
xnor U6363 (N_6363,N_1675,N_826);
and U6364 (N_6364,N_3954,N_989);
nand U6365 (N_6365,N_2304,N_1973);
nand U6366 (N_6366,N_324,N_1634);
or U6367 (N_6367,N_525,N_4441);
xor U6368 (N_6368,N_1365,N_1440);
and U6369 (N_6369,N_3665,N_2295);
nor U6370 (N_6370,N_1921,N_2487);
nor U6371 (N_6371,N_4169,N_3519);
or U6372 (N_6372,N_2205,N_515);
xnor U6373 (N_6373,N_2637,N_3222);
nor U6374 (N_6374,N_294,N_3523);
and U6375 (N_6375,N_3737,N_2232);
nor U6376 (N_6376,N_4304,N_1837);
or U6377 (N_6377,N_2075,N_2430);
and U6378 (N_6378,N_2114,N_44);
xnor U6379 (N_6379,N_3839,N_141);
nand U6380 (N_6380,N_1570,N_4835);
and U6381 (N_6381,N_251,N_4642);
nor U6382 (N_6382,N_1246,N_3182);
xnor U6383 (N_6383,N_3078,N_1593);
xnor U6384 (N_6384,N_3127,N_3909);
nand U6385 (N_6385,N_2840,N_85);
xor U6386 (N_6386,N_1539,N_2224);
xnor U6387 (N_6387,N_647,N_3446);
or U6388 (N_6388,N_1118,N_1767);
or U6389 (N_6389,N_2961,N_803);
or U6390 (N_6390,N_3894,N_3240);
nor U6391 (N_6391,N_151,N_2528);
nand U6392 (N_6392,N_4057,N_340);
xnor U6393 (N_6393,N_1890,N_2984);
xnor U6394 (N_6394,N_2903,N_2415);
xor U6395 (N_6395,N_4105,N_795);
xor U6396 (N_6396,N_3891,N_211);
nor U6397 (N_6397,N_973,N_4218);
and U6398 (N_6398,N_4655,N_1733);
nor U6399 (N_6399,N_804,N_3018);
or U6400 (N_6400,N_2537,N_4856);
and U6401 (N_6401,N_1399,N_3500);
and U6402 (N_6402,N_3102,N_3549);
and U6403 (N_6403,N_2080,N_2507);
nand U6404 (N_6404,N_3636,N_4155);
and U6405 (N_6405,N_1191,N_3773);
and U6406 (N_6406,N_4256,N_809);
nor U6407 (N_6407,N_776,N_1287);
xnor U6408 (N_6408,N_1498,N_1344);
or U6409 (N_6409,N_74,N_649);
xor U6410 (N_6410,N_3921,N_2652);
xnor U6411 (N_6411,N_4860,N_73);
nor U6412 (N_6412,N_697,N_4702);
or U6413 (N_6413,N_959,N_4884);
nand U6414 (N_6414,N_2384,N_1673);
nor U6415 (N_6415,N_4163,N_4626);
nand U6416 (N_6416,N_1868,N_3551);
and U6417 (N_6417,N_2123,N_3312);
xor U6418 (N_6418,N_1817,N_3689);
or U6419 (N_6419,N_1653,N_3749);
nand U6420 (N_6420,N_3573,N_4239);
or U6421 (N_6421,N_709,N_3828);
or U6422 (N_6422,N_2203,N_285);
or U6423 (N_6423,N_2502,N_3361);
or U6424 (N_6424,N_4274,N_955);
xor U6425 (N_6425,N_220,N_4809);
nand U6426 (N_6426,N_4079,N_635);
nand U6427 (N_6427,N_4364,N_680);
or U6428 (N_6428,N_1923,N_2440);
and U6429 (N_6429,N_1602,N_2799);
and U6430 (N_6430,N_2126,N_1979);
or U6431 (N_6431,N_2484,N_2049);
and U6432 (N_6432,N_1134,N_535);
and U6433 (N_6433,N_1549,N_4481);
xor U6434 (N_6434,N_4535,N_1418);
nand U6435 (N_6435,N_3320,N_4947);
xnor U6436 (N_6436,N_588,N_3809);
and U6437 (N_6437,N_571,N_4903);
nor U6438 (N_6438,N_2783,N_4082);
nand U6439 (N_6439,N_1024,N_2893);
xor U6440 (N_6440,N_1046,N_2950);
and U6441 (N_6441,N_533,N_4988);
nor U6442 (N_6442,N_1256,N_273);
and U6443 (N_6443,N_4315,N_2090);
xnor U6444 (N_6444,N_1551,N_2395);
nand U6445 (N_6445,N_3242,N_2099);
or U6446 (N_6446,N_213,N_3784);
xor U6447 (N_6447,N_3866,N_2841);
or U6448 (N_6448,N_3266,N_834);
nor U6449 (N_6449,N_2929,N_3961);
nand U6450 (N_6450,N_2771,N_2774);
and U6451 (N_6451,N_3032,N_2570);
or U6452 (N_6452,N_309,N_2545);
nand U6453 (N_6453,N_2816,N_279);
nor U6454 (N_6454,N_4869,N_2216);
and U6455 (N_6455,N_1028,N_3461);
and U6456 (N_6456,N_1523,N_1952);
nor U6457 (N_6457,N_2523,N_2949);
or U6458 (N_6458,N_4450,N_1651);
nor U6459 (N_6459,N_1085,N_4064);
xor U6460 (N_6460,N_1550,N_329);
xnor U6461 (N_6461,N_3830,N_4799);
and U6462 (N_6462,N_921,N_978);
xnor U6463 (N_6463,N_325,N_1428);
nand U6464 (N_6464,N_4251,N_620);
or U6465 (N_6465,N_137,N_3591);
xor U6466 (N_6466,N_3224,N_4438);
xor U6467 (N_6467,N_3055,N_627);
and U6468 (N_6468,N_3631,N_345);
nand U6469 (N_6469,N_4739,N_3777);
and U6470 (N_6470,N_2819,N_3615);
nor U6471 (N_6471,N_1280,N_1284);
nand U6472 (N_6472,N_1561,N_4871);
or U6473 (N_6473,N_1985,N_3462);
and U6474 (N_6474,N_1669,N_1969);
nor U6475 (N_6475,N_2569,N_3725);
nand U6476 (N_6476,N_3331,N_3596);
and U6477 (N_6477,N_966,N_4382);
nand U6478 (N_6478,N_3980,N_4319);
nand U6479 (N_6479,N_393,N_2185);
or U6480 (N_6480,N_566,N_12);
and U6481 (N_6481,N_4643,N_3417);
nand U6482 (N_6482,N_344,N_506);
nand U6483 (N_6483,N_2169,N_4846);
nor U6484 (N_6484,N_2898,N_4887);
or U6485 (N_6485,N_90,N_4705);
or U6486 (N_6486,N_4030,N_1244);
and U6487 (N_6487,N_1273,N_2039);
or U6488 (N_6488,N_2072,N_2200);
nor U6489 (N_6489,N_4199,N_1684);
or U6490 (N_6490,N_1707,N_2724);
and U6491 (N_6491,N_2051,N_3343);
nand U6492 (N_6492,N_1300,N_3962);
and U6493 (N_6493,N_271,N_3722);
or U6494 (N_6494,N_3515,N_2911);
nand U6495 (N_6495,N_913,N_3727);
nand U6496 (N_6496,N_4447,N_3416);
xor U6497 (N_6497,N_2789,N_2212);
xnor U6498 (N_6498,N_4196,N_759);
xnor U6499 (N_6499,N_3142,N_292);
xor U6500 (N_6500,N_4166,N_2428);
nand U6501 (N_6501,N_1844,N_210);
nor U6502 (N_6502,N_3987,N_2401);
nand U6503 (N_6503,N_1294,N_2530);
xor U6504 (N_6504,N_2553,N_2854);
nor U6505 (N_6505,N_568,N_1325);
nand U6506 (N_6506,N_1626,N_2813);
nand U6507 (N_6507,N_748,N_3324);
nor U6508 (N_6508,N_3887,N_3310);
or U6509 (N_6509,N_2890,N_925);
and U6510 (N_6510,N_4003,N_2658);
xnor U6511 (N_6511,N_245,N_2838);
xor U6512 (N_6512,N_198,N_405);
xor U6513 (N_6513,N_3935,N_753);
nand U6514 (N_6514,N_2156,N_2002);
nor U6515 (N_6515,N_3696,N_669);
xnor U6516 (N_6516,N_2690,N_1936);
and U6517 (N_6517,N_1692,N_1614);
nor U6518 (N_6518,N_4644,N_1850);
or U6519 (N_6519,N_4738,N_486);
nor U6520 (N_6520,N_94,N_3085);
or U6521 (N_6521,N_4553,N_4127);
nor U6522 (N_6522,N_3330,N_3259);
nand U6523 (N_6523,N_1722,N_4293);
xnor U6524 (N_6524,N_4018,N_386);
and U6525 (N_6525,N_3499,N_2612);
nand U6526 (N_6526,N_3926,N_2693);
nand U6527 (N_6527,N_42,N_4775);
nand U6528 (N_6528,N_65,N_574);
nand U6529 (N_6529,N_2648,N_2761);
nand U6530 (N_6530,N_4743,N_3964);
or U6531 (N_6531,N_2795,N_3281);
xnor U6532 (N_6532,N_369,N_3674);
or U6533 (N_6533,N_2750,N_1966);
xnor U6534 (N_6534,N_698,N_4851);
xor U6535 (N_6535,N_4548,N_1594);
xnor U6536 (N_6536,N_2713,N_1367);
nor U6537 (N_6537,N_2279,N_304);
xor U6538 (N_6538,N_1685,N_2058);
xnor U6539 (N_6539,N_785,N_2406);
or U6540 (N_6540,N_1000,N_30);
nor U6541 (N_6541,N_598,N_2740);
nand U6542 (N_6542,N_4496,N_4526);
or U6543 (N_6543,N_4444,N_207);
and U6544 (N_6544,N_2672,N_1263);
and U6545 (N_6545,N_1960,N_1489);
and U6546 (N_6546,N_362,N_2070);
nor U6547 (N_6547,N_3731,N_4613);
nand U6548 (N_6548,N_2079,N_3274);
nor U6549 (N_6549,N_1959,N_1804);
xor U6550 (N_6550,N_1603,N_169);
nor U6551 (N_6551,N_2350,N_1165);
or U6552 (N_6552,N_4414,N_162);
nor U6553 (N_6553,N_1965,N_4210);
xor U6554 (N_6554,N_3763,N_82);
xnor U6555 (N_6555,N_3904,N_4185);
or U6556 (N_6556,N_135,N_692);
or U6557 (N_6557,N_4758,N_2990);
and U6558 (N_6558,N_739,N_4712);
nor U6559 (N_6559,N_4483,N_3845);
nand U6560 (N_6560,N_1889,N_558);
xor U6561 (N_6561,N_75,N_905);
nor U6562 (N_6562,N_1862,N_3172);
or U6563 (N_6563,N_4609,N_4047);
nand U6564 (N_6564,N_643,N_4306);
or U6565 (N_6565,N_3412,N_1568);
xor U6566 (N_6566,N_1237,N_2168);
and U6567 (N_6567,N_3770,N_1223);
nand U6568 (N_6568,N_2966,N_3190);
nand U6569 (N_6569,N_1334,N_3081);
and U6570 (N_6570,N_1359,N_3794);
nor U6571 (N_6571,N_1301,N_2362);
nand U6572 (N_6572,N_1589,N_3349);
nand U6573 (N_6573,N_3410,N_1809);
or U6574 (N_6574,N_2925,N_943);
nor U6575 (N_6575,N_3422,N_1621);
nand U6576 (N_6576,N_611,N_3759);
xor U6577 (N_6577,N_3157,N_3033);
xnor U6578 (N_6578,N_4230,N_2997);
nor U6579 (N_6579,N_165,N_4599);
or U6580 (N_6580,N_2325,N_2098);
xor U6581 (N_6581,N_3365,N_1436);
nor U6582 (N_6582,N_3185,N_349);
nand U6583 (N_6583,N_1228,N_2743);
nand U6584 (N_6584,N_4446,N_4922);
and U6585 (N_6585,N_200,N_4755);
nor U6586 (N_6586,N_2908,N_3209);
and U6587 (N_6587,N_618,N_1866);
nor U6588 (N_6588,N_2369,N_379);
xor U6589 (N_6589,N_2871,N_3214);
xor U6590 (N_6590,N_3083,N_1248);
xor U6591 (N_6591,N_3558,N_2368);
nand U6592 (N_6592,N_3517,N_1871);
and U6593 (N_6593,N_1013,N_217);
xor U6594 (N_6594,N_1517,N_663);
nor U6595 (N_6595,N_781,N_1920);
nand U6596 (N_6596,N_3253,N_119);
nand U6597 (N_6597,N_485,N_1083);
and U6598 (N_6598,N_3360,N_3455);
nor U6599 (N_6599,N_633,N_170);
xnor U6600 (N_6600,N_397,N_1945);
nor U6601 (N_6601,N_193,N_3280);
and U6602 (N_6602,N_829,N_1422);
or U6603 (N_6603,N_3623,N_4744);
or U6604 (N_6604,N_342,N_132);
xor U6605 (N_6605,N_1649,N_4889);
or U6606 (N_6606,N_1617,N_1010);
and U6607 (N_6607,N_2452,N_2420);
xor U6608 (N_6608,N_1158,N_1610);
and U6609 (N_6609,N_1212,N_124);
nand U6610 (N_6610,N_4628,N_4109);
or U6611 (N_6611,N_149,N_1524);
or U6612 (N_6612,N_2941,N_1048);
nand U6613 (N_6613,N_2479,N_3);
xor U6614 (N_6614,N_4891,N_2349);
and U6615 (N_6615,N_150,N_429);
and U6616 (N_6616,N_2886,N_1938);
or U6617 (N_6617,N_3978,N_3239);
and U6618 (N_6618,N_667,N_1285);
nor U6619 (N_6619,N_4549,N_4993);
and U6620 (N_6620,N_2125,N_2236);
xor U6621 (N_6621,N_1052,N_708);
xor U6622 (N_6622,N_4359,N_2093);
nand U6623 (N_6623,N_1546,N_1490);
and U6624 (N_6624,N_828,N_3277);
nand U6625 (N_6625,N_147,N_4534);
or U6626 (N_6626,N_2660,N_1042);
nor U6627 (N_6627,N_2102,N_3808);
nand U6628 (N_6628,N_156,N_449);
or U6629 (N_6629,N_4578,N_2278);
or U6630 (N_6630,N_3604,N_1088);
xor U6631 (N_6631,N_944,N_3232);
nand U6632 (N_6632,N_1734,N_2737);
and U6633 (N_6633,N_885,N_491);
or U6634 (N_6634,N_1803,N_2270);
and U6635 (N_6635,N_1355,N_2509);
and U6636 (N_6636,N_4355,N_2481);
or U6637 (N_6637,N_235,N_1808);
and U6638 (N_6638,N_3628,N_3712);
and U6639 (N_6639,N_2130,N_474);
xnor U6640 (N_6640,N_118,N_4816);
and U6641 (N_6641,N_948,N_3798);
and U6642 (N_6642,N_1126,N_3323);
and U6643 (N_6643,N_3769,N_3504);
and U6644 (N_6644,N_206,N_4204);
nor U6645 (N_6645,N_4714,N_880);
and U6646 (N_6646,N_3337,N_889);
nand U6647 (N_6647,N_2786,N_2181);
or U6648 (N_6648,N_4660,N_4033);
and U6649 (N_6649,N_1251,N_1202);
nor U6650 (N_6650,N_3057,N_3285);
nor U6651 (N_6651,N_4426,N_2162);
nor U6652 (N_6652,N_2045,N_4906);
xnor U6653 (N_6653,N_2241,N_293);
xnor U6654 (N_6654,N_1104,N_1139);
or U6655 (N_6655,N_4802,N_4497);
nand U6656 (N_6656,N_851,N_3118);
nor U6657 (N_6657,N_3973,N_4971);
nand U6658 (N_6658,N_1472,N_1694);
nor U6659 (N_6659,N_1258,N_3261);
nor U6660 (N_6660,N_1520,N_2869);
xor U6661 (N_6661,N_1357,N_3669);
nand U6662 (N_6662,N_1761,N_3166);
xnor U6663 (N_6663,N_655,N_3056);
nand U6664 (N_6664,N_178,N_197);
nand U6665 (N_6665,N_2828,N_361);
nor U6666 (N_6666,N_3790,N_4354);
nor U6667 (N_6667,N_1377,N_1030);
or U6668 (N_6668,N_2315,N_262);
xnor U6669 (N_6669,N_4110,N_695);
or U6670 (N_6670,N_3902,N_3152);
xor U6671 (N_6671,N_1346,N_722);
xnor U6672 (N_6672,N_3970,N_37);
or U6673 (N_6673,N_4583,N_4615);
xor U6674 (N_6674,N_101,N_4474);
nand U6675 (N_6675,N_3332,N_2297);
nand U6676 (N_6676,N_3757,N_4717);
xor U6677 (N_6677,N_299,N_3022);
nor U6678 (N_6678,N_4684,N_648);
and U6679 (N_6679,N_2082,N_1724);
or U6680 (N_6680,N_4519,N_2388);
nor U6681 (N_6681,N_527,N_3414);
or U6682 (N_6682,N_4162,N_1518);
nand U6683 (N_6683,N_1302,N_4234);
and U6684 (N_6684,N_1740,N_4579);
nor U6685 (N_6685,N_1369,N_770);
xnor U6686 (N_6686,N_3826,N_4562);
or U6687 (N_6687,N_4942,N_2294);
xnor U6688 (N_6688,N_1696,N_4682);
nor U6689 (N_6689,N_3432,N_3294);
or U6690 (N_6690,N_4619,N_2866);
xor U6691 (N_6691,N_2129,N_3659);
and U6692 (N_6692,N_3497,N_3688);
nor U6693 (N_6693,N_2001,N_3136);
or U6694 (N_6694,N_4547,N_1144);
xor U6695 (N_6695,N_1800,N_1461);
nand U6696 (N_6696,N_2664,N_258);
or U6697 (N_6697,N_1424,N_3772);
xor U6698 (N_6698,N_4462,N_4360);
or U6699 (N_6699,N_4148,N_2593);
nand U6700 (N_6700,N_1488,N_1242);
and U6701 (N_6701,N_2332,N_3363);
nand U6702 (N_6702,N_1283,N_4756);
nand U6703 (N_6703,N_3529,N_3306);
nand U6704 (N_6704,N_1806,N_2865);
nand U6705 (N_6705,N_1678,N_2029);
nor U6706 (N_6706,N_1688,N_3161);
and U6707 (N_6707,N_3371,N_4920);
nand U6708 (N_6708,N_922,N_3345);
nor U6709 (N_6709,N_3065,N_4558);
nor U6710 (N_6710,N_2675,N_399);
nand U6711 (N_6711,N_3299,N_4095);
xnor U6712 (N_6712,N_96,N_2435);
xnor U6713 (N_6713,N_4929,N_2286);
or U6714 (N_6714,N_641,N_214);
or U6715 (N_6715,N_1271,N_3925);
or U6716 (N_6716,N_4188,N_597);
or U6717 (N_6717,N_4182,N_1779);
xnor U6718 (N_6718,N_4137,N_4092);
nand U6719 (N_6719,N_3616,N_811);
xor U6720 (N_6720,N_2175,N_986);
nand U6721 (N_6721,N_4339,N_870);
and U6722 (N_6722,N_3225,N_744);
or U6723 (N_6723,N_614,N_1886);
nor U6724 (N_6724,N_1456,N_832);
nand U6725 (N_6725,N_4455,N_409);
nand U6726 (N_6726,N_4841,N_95);
xor U6727 (N_6727,N_121,N_1445);
or U6728 (N_6728,N_0,N_1975);
and U6729 (N_6729,N_3449,N_363);
nand U6730 (N_6730,N_56,N_1999);
and U6731 (N_6731,N_843,N_1720);
xnor U6732 (N_6732,N_3589,N_2921);
or U6733 (N_6733,N_3444,N_487);
nor U6734 (N_6734,N_2376,N_4454);
or U6735 (N_6735,N_492,N_820);
or U6736 (N_6736,N_860,N_890);
nand U6737 (N_6737,N_4449,N_2459);
nor U6738 (N_6738,N_4119,N_323);
or U6739 (N_6739,N_4014,N_1137);
nand U6740 (N_6740,N_4597,N_3227);
xnor U6741 (N_6741,N_1998,N_3900);
nor U6742 (N_6742,N_1940,N_2355);
nand U6743 (N_6743,N_2568,N_3663);
nand U6744 (N_6744,N_3007,N_2688);
xnor U6745 (N_6745,N_115,N_2192);
xor U6746 (N_6746,N_4517,N_3006);
or U6747 (N_6747,N_1572,N_1553);
nor U6748 (N_6748,N_4331,N_4546);
nor U6749 (N_6749,N_1547,N_2920);
nor U6750 (N_6750,N_28,N_3601);
and U6751 (N_6751,N_2539,N_2759);
and U6752 (N_6752,N_2306,N_769);
and U6753 (N_6753,N_1446,N_1296);
xor U6754 (N_6754,N_953,N_2611);
or U6755 (N_6755,N_327,N_4813);
nand U6756 (N_6756,N_3739,N_1829);
xnor U6757 (N_6757,N_80,N_977);
or U6758 (N_6758,N_752,N_3464);
xor U6759 (N_6759,N_1878,N_3958);
nand U6760 (N_6760,N_4208,N_3435);
or U6761 (N_6761,N_3344,N_2244);
nor U6762 (N_6762,N_907,N_4632);
nor U6763 (N_6763,N_4377,N_713);
xor U6764 (N_6764,N_3287,N_2715);
or U6765 (N_6765,N_604,N_4771);
or U6766 (N_6766,N_4216,N_4876);
or U6767 (N_6767,N_3167,N_3806);
nor U6768 (N_6768,N_2149,N_442);
nand U6769 (N_6769,N_1781,N_2337);
nand U6770 (N_6770,N_4877,N_545);
xnor U6771 (N_6771,N_3761,N_4883);
and U6772 (N_6772,N_1170,N_4544);
nand U6773 (N_6773,N_2753,N_3928);
and U6774 (N_6774,N_4429,N_3017);
or U6775 (N_6775,N_2230,N_4635);
or U6776 (N_6776,N_4152,N_3482);
and U6777 (N_6777,N_2044,N_4071);
nand U6778 (N_6778,N_653,N_3112);
nor U6779 (N_6779,N_3871,N_2150);
and U6780 (N_6780,N_3946,N_2383);
xor U6781 (N_6781,N_2540,N_4254);
nand U6782 (N_6782,N_540,N_993);
nor U6783 (N_6783,N_2659,N_3649);
and U6784 (N_6784,N_291,N_933);
and U6785 (N_6785,N_2714,N_1683);
and U6786 (N_6786,N_3477,N_91);
nand U6787 (N_6787,N_1332,N_3533);
xor U6788 (N_6788,N_4610,N_2527);
xor U6789 (N_6789,N_1739,N_3700);
or U6790 (N_6790,N_321,N_27);
nor U6791 (N_6791,N_2534,N_241);
or U6792 (N_6792,N_2639,N_849);
nand U6793 (N_6793,N_107,N_4576);
nor U6794 (N_6794,N_380,N_4303);
xnor U6795 (N_6795,N_569,N_3316);
nand U6796 (N_6796,N_2385,N_4046);
nor U6797 (N_6797,N_1405,N_526);
or U6798 (N_6798,N_1149,N_3645);
xnor U6799 (N_6799,N_4379,N_1064);
or U6800 (N_6800,N_13,N_3932);
nor U6801 (N_6801,N_1193,N_2266);
nor U6802 (N_6802,N_4912,N_819);
nand U6803 (N_6803,N_4718,N_677);
nor U6804 (N_6804,N_1627,N_2574);
xnor U6805 (N_6805,N_4901,N_2432);
nor U6806 (N_6806,N_556,N_4811);
or U6807 (N_6807,N_768,N_2669);
xor U6808 (N_6808,N_3698,N_2566);
and U6809 (N_6809,N_2882,N_368);
xnor U6810 (N_6810,N_2760,N_275);
or U6811 (N_6811,N_40,N_117);
xnor U6812 (N_6812,N_2973,N_2972);
nand U6813 (N_6813,N_1133,N_3013);
nand U6814 (N_6814,N_4279,N_4501);
or U6815 (N_6815,N_3290,N_4088);
xnor U6816 (N_6816,N_1394,N_1017);
xor U6817 (N_6817,N_4659,N_2448);
or U6818 (N_6818,N_3377,N_1912);
xor U6819 (N_6819,N_4253,N_2311);
xnor U6820 (N_6820,N_2434,N_58);
or U6821 (N_6821,N_2441,N_2976);
nand U6822 (N_6822,N_4482,N_1741);
nand U6823 (N_6823,N_1571,N_4480);
xnor U6824 (N_6824,N_1406,N_3082);
or U6825 (N_6825,N_81,N_4202);
or U6826 (N_6826,N_1854,N_3379);
or U6827 (N_6827,N_4720,N_3570);
and U6828 (N_6828,N_4294,N_1392);
xnor U6829 (N_6829,N_3531,N_2618);
xnor U6830 (N_6830,N_339,N_2400);
and U6831 (N_6831,N_4022,N_2709);
and U6832 (N_6832,N_2261,N_4787);
or U6833 (N_6833,N_4021,N_2726);
xnor U6834 (N_6834,N_584,N_3883);
nand U6835 (N_6835,N_2768,N_125);
xor U6836 (N_6836,N_1711,N_1438);
and U6837 (N_6837,N_2249,N_1690);
or U6838 (N_6838,N_2936,N_4433);
nor U6839 (N_6839,N_4683,N_3229);
nor U6840 (N_6840,N_4111,N_2757);
and U6841 (N_6841,N_2806,N_3510);
xnor U6842 (N_6842,N_4241,N_2860);
and U6843 (N_6843,N_1372,N_2365);
xnor U6844 (N_6844,N_1045,N_1658);
and U6845 (N_6845,N_656,N_1845);
xor U6846 (N_6846,N_430,N_3736);
or U6847 (N_6847,N_1607,N_4488);
and U6848 (N_6848,N_3566,N_2718);
nand U6849 (N_6849,N_2326,N_3695);
nor U6850 (N_6850,N_2951,N_1250);
nor U6851 (N_6851,N_3979,N_2014);
nor U6852 (N_6852,N_4363,N_1944);
xor U6853 (N_6853,N_2092,N_1402);
and U6854 (N_6854,N_2313,N_1423);
xor U6855 (N_6855,N_994,N_2678);
nor U6856 (N_6856,N_2100,N_4968);
and U6857 (N_6857,N_2904,N_2358);
xor U6858 (N_6858,N_1951,N_2269);
or U6859 (N_6859,N_813,N_4246);
xnor U6860 (N_6860,N_3799,N_3730);
and U6861 (N_6861,N_4027,N_476);
nand U6862 (N_6862,N_3593,N_3096);
xnor U6863 (N_6863,N_2765,N_1119);
or U6864 (N_6864,N_4479,N_427);
nor U6865 (N_6865,N_561,N_4471);
or U6866 (N_6866,N_4512,N_4842);
and U6867 (N_6867,N_1316,N_2221);
nor U6868 (N_6868,N_2336,N_3562);
xor U6869 (N_6869,N_3823,N_143);
and U6870 (N_6870,N_1087,N_1329);
nor U6871 (N_6871,N_3066,N_4543);
xor U6872 (N_6872,N_1234,N_3411);
xor U6873 (N_6873,N_4299,N_1858);
xnor U6874 (N_6874,N_4603,N_1403);
or U6875 (N_6875,N_902,N_554);
xnor U6876 (N_6876,N_4893,N_2666);
or U6877 (N_6877,N_999,N_3002);
and U6878 (N_6878,N_2486,N_2632);
nor U6879 (N_6879,N_4058,N_3019);
nor U6880 (N_6880,N_884,N_1897);
xnor U6881 (N_6881,N_4982,N_503);
nand U6882 (N_6882,N_1469,N_3008);
and U6883 (N_6883,N_2580,N_2578);
and U6884 (N_6884,N_3204,N_593);
nor U6885 (N_6885,N_4608,N_1268);
nand U6886 (N_6886,N_288,N_3493);
nor U6887 (N_6887,N_2554,N_1233);
nand U6888 (N_6888,N_4212,N_364);
nor U6889 (N_6889,N_3351,N_1511);
nand U6890 (N_6890,N_2277,N_2981);
nand U6891 (N_6891,N_247,N_3257);
or U6892 (N_6892,N_2711,N_2252);
or U6893 (N_6893,N_4521,N_3681);
nor U6894 (N_6894,N_4222,N_4513);
and U6895 (N_6895,N_4205,N_2602);
nand U6896 (N_6896,N_2597,N_2253);
nand U6897 (N_6897,N_3554,N_4582);
nand U6898 (N_6898,N_3835,N_4219);
or U6899 (N_6899,N_4885,N_4925);
nor U6900 (N_6900,N_2215,N_2003);
and U6901 (N_6901,N_1025,N_2106);
nand U6902 (N_6902,N_3080,N_1249);
nor U6903 (N_6903,N_2698,N_3249);
and U6904 (N_6904,N_3552,N_1648);
nor U6905 (N_6905,N_2985,N_3750);
nor U6906 (N_6906,N_2586,N_2485);
nor U6907 (N_6907,N_4249,N_2407);
or U6908 (N_6908,N_563,N_4916);
and U6909 (N_6909,N_4366,N_2030);
or U6910 (N_6910,N_1100,N_1813);
and U6911 (N_6911,N_3643,N_2710);
xor U6912 (N_6912,N_4698,N_4495);
xnor U6913 (N_6913,N_1752,N_460);
nor U6914 (N_6914,N_4004,N_3703);
nor U6915 (N_6915,N_2390,N_2468);
nor U6916 (N_6916,N_3418,N_3375);
and U6917 (N_6917,N_4312,N_1439);
nor U6918 (N_6918,N_2229,N_2522);
and U6919 (N_6919,N_2727,N_3311);
xor U6920 (N_6920,N_3680,N_2810);
or U6921 (N_6921,N_22,N_360);
nor U6922 (N_6922,N_2705,N_542);
and U6923 (N_6923,N_628,N_2104);
and U6924 (N_6924,N_1492,N_2463);
nand U6925 (N_6925,N_3882,N_4280);
nor U6926 (N_6926,N_366,N_3233);
nor U6927 (N_6927,N_3087,N_2575);
nand U6928 (N_6928,N_2562,N_1433);
or U6929 (N_6929,N_3850,N_3625);
nor U6930 (N_6930,N_1608,N_896);
and U6931 (N_6931,N_3764,N_2020);
nor U6932 (N_6932,N_1004,N_1264);
nor U6933 (N_6933,N_2608,N_747);
nor U6934 (N_6934,N_3192,N_267);
or U6935 (N_6935,N_418,N_4729);
xnor U6936 (N_6936,N_4803,N_705);
nand U6937 (N_6937,N_1002,N_1197);
and U6938 (N_6938,N_2503,N_596);
xnor U6939 (N_6939,N_790,N_3439);
nand U6940 (N_6940,N_443,N_2516);
nand U6941 (N_6941,N_3907,N_4629);
or U6942 (N_6942,N_4895,N_2955);
and U6943 (N_6943,N_4443,N_1290);
nand U6944 (N_6944,N_2010,N_343);
nor U6945 (N_6945,N_3716,N_1327);
nand U6946 (N_6946,N_1681,N_3929);
and U6947 (N_6947,N_3639,N_3399);
or U6948 (N_6948,N_3313,N_1543);
or U6949 (N_6949,N_3577,N_1221);
and U6950 (N_6950,N_731,N_1360);
nor U6951 (N_6951,N_4657,N_3419);
xor U6952 (N_6952,N_1217,N_1671);
or U6953 (N_6953,N_2689,N_2394);
or U6954 (N_6954,N_351,N_1091);
nand U6955 (N_6955,N_4362,N_408);
nor U6956 (N_6956,N_338,N_3627);
xor U6957 (N_6957,N_2617,N_848);
and U6958 (N_6958,N_868,N_3200);
nor U6959 (N_6959,N_4939,N_3456);
or U6960 (N_6960,N_3608,N_4173);
xor U6961 (N_6961,N_4795,N_4515);
xnor U6962 (N_6962,N_3924,N_4353);
and U6963 (N_6963,N_4631,N_4601);
nor U6964 (N_6964,N_3150,N_3207);
or U6965 (N_6965,N_1112,N_564);
nor U6966 (N_6966,N_2101,N_591);
and U6967 (N_6967,N_1475,N_144);
nand U6968 (N_6968,N_894,N_799);
nor U6969 (N_6969,N_2633,N_3380);
nor U6970 (N_6970,N_840,N_4044);
nand U6971 (N_6971,N_835,N_997);
xor U6972 (N_6972,N_683,N_2281);
nor U6973 (N_6973,N_1723,N_2729);
or U6974 (N_6974,N_2188,N_3269);
and U6975 (N_6975,N_4104,N_3686);
and U6976 (N_6976,N_133,N_233);
and U6977 (N_6977,N_3044,N_336);
nand U6978 (N_6978,N_1199,N_3169);
nor U6979 (N_6979,N_685,N_724);
xor U6980 (N_6980,N_3392,N_2201);
xnor U6981 (N_6981,N_3124,N_2161);
xnor U6982 (N_6982,N_3922,N_4233);
nor U6983 (N_6983,N_3068,N_2521);
xor U6984 (N_6984,N_2542,N_4511);
nor U6985 (N_6985,N_1513,N_687);
or U6986 (N_6986,N_1506,N_626);
nand U6987 (N_6987,N_4685,N_833);
nor U6988 (N_6988,N_3914,N_1166);
or U6989 (N_6989,N_4976,N_623);
nand U6990 (N_6990,N_2180,N_332);
xnor U6991 (N_6991,N_390,N_1462);
nor U6992 (N_6992,N_3075,N_2873);
nor U6993 (N_6993,N_3350,N_4589);
or U6994 (N_6994,N_2741,N_3162);
xor U6995 (N_6995,N_4861,N_1650);
nand U6996 (N_6996,N_266,N_706);
xor U6997 (N_6997,N_2265,N_2804);
xor U6998 (N_6998,N_3488,N_4818);
nand U6999 (N_6999,N_263,N_4998);
xor U7000 (N_7000,N_765,N_2023);
nor U7001 (N_7001,N_142,N_4028);
and U7002 (N_7002,N_4675,N_1055);
nor U7003 (N_7003,N_3537,N_2172);
and U7004 (N_7004,N_1415,N_4289);
xor U7005 (N_7005,N_4814,N_4872);
nor U7006 (N_7006,N_2237,N_3151);
nor U7007 (N_7007,N_1291,N_3886);
or U7008 (N_7008,N_3920,N_4328);
and U7009 (N_7009,N_2083,N_3024);
and U7010 (N_7010,N_2381,N_496);
and U7011 (N_7011,N_2674,N_1313);
nor U7012 (N_7012,N_4270,N_3834);
xor U7013 (N_7013,N_2796,N_216);
and U7014 (N_7014,N_2621,N_4923);
or U7015 (N_7015,N_1783,N_3789);
or U7016 (N_7016,N_1773,N_4747);
and U7017 (N_7017,N_3027,N_883);
or U7018 (N_7018,N_3569,N_2421);
or U7019 (N_7019,N_1177,N_2667);
and U7020 (N_7020,N_4772,N_2915);
and U7021 (N_7021,N_4500,N_1322);
and U7022 (N_7022,N_3582,N_2472);
nand U7023 (N_7023,N_2773,N_3950);
nor U7024 (N_7024,N_167,N_3186);
nand U7025 (N_7025,N_2176,N_4060);
nand U7026 (N_7026,N_2642,N_398);
nor U7027 (N_7027,N_2246,N_3530);
and U7028 (N_7028,N_3283,N_1807);
nand U7029 (N_7029,N_2047,N_2623);
or U7030 (N_7030,N_3526,N_3939);
nor U7031 (N_7031,N_2449,N_4427);
and U7032 (N_7032,N_4273,N_1900);
or U7033 (N_7033,N_1904,N_3405);
nor U7034 (N_7034,N_3366,N_4661);
xor U7035 (N_7035,N_771,N_2577);
xor U7036 (N_7036,N_3009,N_945);
and U7037 (N_7037,N_3467,N_4178);
and U7038 (N_7038,N_1105,N_4591);
or U7039 (N_7039,N_1253,N_3742);
and U7040 (N_7040,N_2839,N_2028);
nor U7041 (N_7041,N_4620,N_2078);
nor U7042 (N_7042,N_2863,N_3778);
nor U7043 (N_7043,N_1374,N_4203);
and U7044 (N_7044,N_2607,N_4053);
and U7045 (N_7045,N_1820,N_4165);
nor U7046 (N_7046,N_4975,N_4244);
and U7047 (N_7047,N_1787,N_1077);
nor U7048 (N_7048,N_3053,N_2184);
nand U7049 (N_7049,N_3023,N_624);
or U7050 (N_7050,N_122,N_174);
and U7051 (N_7051,N_4035,N_2210);
and U7052 (N_7052,N_572,N_4126);
and U7053 (N_7053,N_1778,N_1065);
or U7054 (N_7054,N_3325,N_2170);
nand U7055 (N_7055,N_4453,N_930);
nor U7056 (N_7056,N_24,N_520);
nor U7057 (N_7057,N_2117,N_2591);
and U7058 (N_7058,N_3048,N_4332);
nor U7059 (N_7059,N_710,N_222);
and U7060 (N_7060,N_1474,N_2134);
and U7061 (N_7061,N_1478,N_4992);
or U7062 (N_7062,N_3606,N_926);
or U7063 (N_7063,N_4504,N_3445);
and U7064 (N_7064,N_699,N_4186);
nand U7065 (N_7065,N_1430,N_3841);
nor U7066 (N_7066,N_995,N_3140);
xor U7067 (N_7067,N_1183,N_440);
nand U7068 (N_7068,N_1142,N_2676);
nand U7069 (N_7069,N_4918,N_3864);
and U7070 (N_7070,N_2887,N_2640);
or U7071 (N_7071,N_954,N_3702);
nand U7072 (N_7072,N_4502,N_651);
and U7073 (N_7073,N_1493,N_821);
nand U7074 (N_7074,N_538,N_2722);
nand U7075 (N_7075,N_128,N_3485);
and U7076 (N_7076,N_1195,N_2735);
xor U7077 (N_7077,N_4285,N_1679);
nor U7078 (N_7078,N_2975,N_4959);
nand U7079 (N_7079,N_3333,N_1612);
nor U7080 (N_7080,N_501,N_1364);
nand U7081 (N_7081,N_3982,N_4828);
and U7082 (N_7082,N_3235,N_2113);
nand U7083 (N_7083,N_2901,N_589);
xor U7084 (N_7084,N_2202,N_2730);
and U7085 (N_7085,N_1421,N_1906);
and U7086 (N_7086,N_3532,N_2089);
xnor U7087 (N_7087,N_4420,N_4149);
or U7088 (N_7088,N_370,N_4283);
or U7089 (N_7089,N_595,N_1035);
and U7090 (N_7090,N_145,N_3031);
xor U7091 (N_7091,N_1597,N_33);
nor U7092 (N_7092,N_4206,N_3580);
and U7093 (N_7093,N_4952,N_4557);
xnor U7094 (N_7094,N_4074,N_489);
or U7095 (N_7095,N_1629,N_2798);
nand U7096 (N_7096,N_3916,N_4258);
or U7097 (N_7097,N_600,N_1073);
and U7098 (N_7098,N_2504,N_640);
nand U7099 (N_7099,N_3836,N_4617);
and U7100 (N_7100,N_51,N_3720);
nor U7101 (N_7101,N_3326,N_3719);
and U7102 (N_7102,N_3101,N_4499);
or U7103 (N_7103,N_2744,N_2847);
nand U7104 (N_7104,N_387,N_2563);
and U7105 (N_7105,N_1497,N_1947);
and U7106 (N_7106,N_2223,N_796);
and U7107 (N_7107,N_873,N_4966);
and U7108 (N_7108,N_547,N_4960);
xor U7109 (N_7109,N_77,N_4862);
nor U7110 (N_7110,N_4598,N_3818);
or U7111 (N_7111,N_1613,N_4123);
and U7112 (N_7112,N_2779,N_4561);
nor U7113 (N_7113,N_1788,N_879);
and U7114 (N_7114,N_4167,N_4570);
or U7115 (N_7115,N_3804,N_3610);
nand U7116 (N_7116,N_1911,N_1636);
xor U7117 (N_7117,N_4307,N_1153);
xor U7118 (N_7118,N_2343,N_3199);
xnor U7119 (N_7119,N_4278,N_3927);
or U7120 (N_7120,N_4875,N_1186);
xor U7121 (N_7121,N_1292,N_2758);
or U7122 (N_7122,N_1643,N_881);
or U7123 (N_7123,N_3768,N_846);
or U7124 (N_7124,N_2567,N_3215);
nand U7125 (N_7125,N_4695,N_2392);
xnor U7126 (N_7126,N_1548,N_3844);
nor U7127 (N_7127,N_4156,N_2954);
or U7128 (N_7128,N_516,N_4794);
or U7129 (N_7129,N_1426,N_2360);
and U7130 (N_7130,N_4067,N_1467);
or U7131 (N_7131,N_1981,N_3098);
or U7132 (N_7132,N_4391,N_4017);
nor U7133 (N_7133,N_2333,N_4950);
xnor U7134 (N_7134,N_1601,N_1849);
nor U7135 (N_7135,N_616,N_702);
and U7136 (N_7136,N_4159,N_1625);
and U7137 (N_7137,N_337,N_3300);
and U7138 (N_7138,N_2928,N_1414);
nor U7139 (N_7139,N_4528,N_4592);
xnor U7140 (N_7140,N_2128,N_1305);
or U7141 (N_7141,N_2728,N_461);
nand U7142 (N_7142,N_3234,N_4697);
nor U7143 (N_7143,N_4563,N_3751);
or U7144 (N_7144,N_1454,N_960);
nand U7145 (N_7145,N_4791,N_3395);
nor U7146 (N_7146,N_4559,N_577);
or U7147 (N_7147,N_4688,N_892);
xnor U7148 (N_7148,N_1159,N_4393);
or U7149 (N_7149,N_4537,N_161);
and U7150 (N_7150,N_1699,N_4693);
nor U7151 (N_7151,N_1769,N_3012);
or U7152 (N_7152,N_1749,N_874);
xor U7153 (N_7153,N_4422,N_4002);
and U7154 (N_7154,N_696,N_2835);
nor U7155 (N_7155,N_2529,N_764);
nand U7156 (N_7156,N_3995,N_1672);
or U7157 (N_7157,N_1124,N_1894);
and U7158 (N_7158,N_354,N_4031);
nand U7159 (N_7159,N_2826,N_4128);
and U7160 (N_7160,N_4207,N_1538);
and U7161 (N_7161,N_1009,N_3218);
and U7162 (N_7162,N_4715,N_3874);
nor U7163 (N_7163,N_3426,N_815);
nor U7164 (N_7164,N_4489,N_3480);
xnor U7165 (N_7165,N_4987,N_2251);
nor U7166 (N_7166,N_4255,N_3634);
nand U7167 (N_7167,N_3930,N_2971);
xnor U7168 (N_7168,N_4113,N_205);
and U7169 (N_7169,N_4527,N_2322);
nor U7170 (N_7170,N_4238,N_3168);
nor U7171 (N_7171,N_3745,N_3619);
nor U7172 (N_7172,N_2988,N_3656);
nor U7173 (N_7173,N_1934,N_1843);
nor U7174 (N_7174,N_1016,N_644);
and U7175 (N_7175,N_845,N_4272);
or U7176 (N_7176,N_3740,N_1413);
nor U7177 (N_7177,N_4157,N_3805);
nand U7178 (N_7178,N_3073,N_2038);
nand U7179 (N_7179,N_751,N_270);
or U7180 (N_7180,N_3735,N_4746);
nor U7181 (N_7181,N_4117,N_3296);
nor U7182 (N_7182,N_4911,N_3811);
or U7183 (N_7183,N_4487,N_671);
nand U7184 (N_7184,N_4820,N_2731);
and U7185 (N_7185,N_8,N_2127);
nor U7186 (N_7186,N_3059,N_897);
xor U7187 (N_7187,N_4600,N_1070);
xnor U7188 (N_7188,N_2661,N_2738);
nor U7189 (N_7189,N_3668,N_1857);
nand U7190 (N_7190,N_347,N_3548);
or U7191 (N_7191,N_4460,N_4812);
nand U7192 (N_7192,N_2510,N_2195);
nand U7193 (N_7193,N_1802,N_1958);
xnor U7194 (N_7194,N_1333,N_3641);
nand U7195 (N_7195,N_622,N_2198);
and U7196 (N_7196,N_2498,N_2788);
or U7197 (N_7197,N_2120,N_4072);
nand U7198 (N_7198,N_1317,N_4242);
xor U7199 (N_7199,N_2189,N_189);
nor U7200 (N_7200,N_2862,N_2906);
nor U7201 (N_7201,N_3139,N_2282);
nor U7202 (N_7202,N_3955,N_1926);
and U7203 (N_7203,N_188,N_3884);
or U7204 (N_7204,N_1205,N_3490);
or U7205 (N_7205,N_4485,N_2396);
nand U7206 (N_7206,N_1989,N_4962);
or U7207 (N_7207,N_4370,N_3129);
nor U7208 (N_7208,N_3442,N_1882);
and U7209 (N_7209,N_86,N_3460);
xor U7210 (N_7210,N_2628,N_3288);
and U7211 (N_7211,N_2635,N_2801);
nand U7212 (N_7212,N_2978,N_2291);
or U7213 (N_7213,N_140,N_3837);
xnor U7214 (N_7214,N_1277,N_4486);
nand U7215 (N_7215,N_191,N_1053);
and U7216 (N_7216,N_1664,N_2878);
or U7217 (N_7217,N_468,N_4754);
and U7218 (N_7218,N_4394,N_958);
and U7219 (N_7219,N_4375,N_3453);
nor U7220 (N_7220,N_915,N_546);
nand U7221 (N_7221,N_2259,N_3869);
or U7222 (N_7222,N_1132,N_447);
and U7223 (N_7223,N_3755,N_4235);
and U7224 (N_7224,N_4118,N_209);
and U7225 (N_7225,N_1995,N_2583);
xnor U7226 (N_7226,N_1731,N_4986);
nand U7227 (N_7227,N_504,N_3443);
xnor U7228 (N_7228,N_3638,N_4785);
nand U7229 (N_7229,N_1746,N_2059);
and U7230 (N_7230,N_4089,N_3402);
or U7231 (N_7231,N_519,N_4138);
xnor U7232 (N_7232,N_131,N_4476);
nor U7233 (N_7233,N_662,N_4506);
xor U7234 (N_7234,N_341,N_2830);
or U7235 (N_7235,N_3184,N_2146);
xor U7236 (N_7236,N_2371,N_4227);
and U7237 (N_7237,N_1950,N_1220);
xnor U7238 (N_7238,N_1833,N_2547);
nor U7239 (N_7239,N_559,N_1730);
nand U7240 (N_7240,N_2624,N_2700);
or U7241 (N_7241,N_2217,N_513);
xor U7242 (N_7242,N_2084,N_158);
or U7243 (N_7243,N_215,N_231);
and U7244 (N_7244,N_2748,N_1311);
and U7245 (N_7245,N_4687,N_3284);
nor U7246 (N_7246,N_2433,N_3448);
nor U7247 (N_7247,N_4934,N_392);
nand U7248 (N_7248,N_3305,N_218);
xnor U7249 (N_7249,N_4077,N_4276);
nand U7250 (N_7250,N_1143,N_3911);
nor U7251 (N_7251,N_3733,N_4352);
or U7252 (N_7252,N_3852,N_2592);
xnor U7253 (N_7253,N_2982,N_3944);
xor U7254 (N_7254,N_2895,N_3516);
or U7255 (N_7255,N_4300,N_2993);
and U7256 (N_7256,N_1096,N_3813);
nor U7257 (N_7257,N_3912,N_437);
nand U7258 (N_7258,N_4940,N_2094);
xor U7259 (N_7259,N_4337,N_2497);
and U7260 (N_7260,N_1715,N_2742);
nor U7261 (N_7261,N_524,N_1353);
or U7262 (N_7262,N_3183,N_1609);
and U7263 (N_7263,N_3899,N_3179);
nand U7264 (N_7264,N_1380,N_2963);
nor U7265 (N_7265,N_1395,N_4493);
or U7266 (N_7266,N_2068,N_4917);
and U7267 (N_7267,N_4134,N_4140);
nor U7268 (N_7268,N_1148,N_377);
or U7269 (N_7269,N_4575,N_3878);
or U7270 (N_7270,N_1164,N_4807);
and U7271 (N_7271,N_1354,N_2234);
nor U7272 (N_7272,N_2359,N_3322);
nand U7273 (N_7273,N_2557,N_942);
and U7274 (N_7274,N_1466,N_654);
or U7275 (N_7275,N_4215,N_4672);
nand U7276 (N_7276,N_3197,N_4465);
xnor U7277 (N_7277,N_723,N_3247);
or U7278 (N_7278,N_4905,N_2520);
and U7279 (N_7279,N_346,N_4385);
xnor U7280 (N_7280,N_553,N_1023);
or U7281 (N_7281,N_3550,N_4564);
or U7282 (N_7282,N_3984,N_4725);
nor U7283 (N_7283,N_2338,N_428);
nor U7284 (N_7284,N_2837,N_3717);
or U7285 (N_7285,N_619,N_4525);
or U7286 (N_7286,N_2263,N_2879);
and U7287 (N_7287,N_659,N_1479);
xnor U7288 (N_7288,N_1022,N_1537);
nor U7289 (N_7289,N_4946,N_1560);
nor U7290 (N_7290,N_2850,N_859);
and U7291 (N_7291,N_3219,N_3782);
nor U7292 (N_7292,N_2111,N_1452);
nor U7293 (N_7293,N_2088,N_909);
nor U7294 (N_7294,N_1667,N_1657);
nand U7295 (N_7295,N_825,N_3421);
and U7296 (N_7296,N_1768,N_3062);
or U7297 (N_7297,N_3264,N_2413);
or U7298 (N_7298,N_3079,N_1825);
and U7299 (N_7299,N_750,N_1097);
xnor U7300 (N_7300,N_956,N_3153);
nor U7301 (N_7301,N_4847,N_1442);
or U7302 (N_7302,N_636,N_1336);
nand U7303 (N_7303,N_4874,N_3067);
nor U7304 (N_7304,N_4340,N_4678);
or U7305 (N_7305,N_666,N_3208);
and U7306 (N_7306,N_2276,N_4679);
or U7307 (N_7307,N_4016,N_3781);
xor U7308 (N_7308,N_4690,N_1605);
and U7309 (N_7309,N_2206,N_2526);
xor U7310 (N_7310,N_1587,N_1033);
and U7311 (N_7311,N_1840,N_4266);
nand U7312 (N_7312,N_384,N_704);
xnor U7313 (N_7313,N_1766,N_2687);
or U7314 (N_7314,N_1027,N_4231);
and U7315 (N_7315,N_3093,N_2053);
and U7316 (N_7316,N_1623,N_1410);
and U7317 (N_7317,N_1861,N_2834);
nand U7318 (N_7318,N_2784,N_2378);
or U7319 (N_7319,N_4779,N_3732);
or U7320 (N_7320,N_3159,N_3376);
nor U7321 (N_7321,N_2699,N_264);
xnor U7322 (N_7322,N_4765,N_3968);
or U7323 (N_7323,N_2938,N_4350);
nand U7324 (N_7324,N_1050,N_4691);
xnor U7325 (N_7325,N_4408,N_4773);
nor U7326 (N_7326,N_3901,N_3043);
and U7327 (N_7327,N_1375,N_356);
xnor U7328 (N_7328,N_1946,N_2296);
xor U7329 (N_7329,N_3387,N_1444);
nand U7330 (N_7330,N_3440,N_4091);
xnor U7331 (N_7331,N_2436,N_4604);
or U7332 (N_7332,N_4677,N_3131);
xnor U7333 (N_7333,N_3105,N_1745);
and U7334 (N_7334,N_801,N_1753);
xnor U7335 (N_7335,N_4139,N_2361);
nand U7336 (N_7336,N_148,N_3039);
or U7337 (N_7337,N_1794,N_138);
nor U7338 (N_7338,N_4854,N_2257);
nand U7339 (N_7339,N_786,N_2352);
or U7340 (N_7340,N_3293,N_3992);
nor U7341 (N_7341,N_1236,N_4056);
nor U7342 (N_7342,N_4142,N_52);
nand U7343 (N_7343,N_2339,N_1816);
or U7344 (N_7344,N_1295,N_3785);
or U7345 (N_7345,N_4415,N_1789);
nor U7346 (N_7346,N_529,N_4707);
nand U7347 (N_7347,N_3126,N_1074);
or U7348 (N_7348,N_511,N_1563);
and U7349 (N_7349,N_4766,N_177);
and U7350 (N_7350,N_1792,N_4277);
nor U7351 (N_7351,N_4607,N_3540);
nand U7352 (N_7352,N_1686,N_4625);
nor U7353 (N_7353,N_1512,N_1855);
or U7354 (N_7354,N_3559,N_4733);
and U7355 (N_7355,N_2052,N_1736);
xor U7356 (N_7356,N_1131,N_3888);
nand U7357 (N_7357,N_230,N_2995);
xnor U7358 (N_7358,N_4384,N_4781);
xor U7359 (N_7359,N_4768,N_4145);
and U7360 (N_7360,N_1069,N_4191);
nor U7361 (N_7361,N_2417,N_3273);
xor U7362 (N_7362,N_714,N_2009);
xor U7363 (N_7363,N_1504,N_2986);
nand U7364 (N_7364,N_3223,N_1545);
nand U7365 (N_7365,N_3693,N_962);
or U7366 (N_7366,N_2917,N_3576);
xor U7367 (N_7367,N_2036,N_1595);
xnor U7368 (N_7368,N_4322,N_728);
nor U7369 (N_7369,N_1272,N_3913);
nand U7370 (N_7370,N_3364,N_2770);
xor U7371 (N_7371,N_4103,N_3047);
nor U7372 (N_7372,N_3960,N_1425);
nor U7373 (N_7373,N_1226,N_2924);
nand U7374 (N_7374,N_1578,N_3077);
nand U7375 (N_7375,N_2515,N_837);
and U7376 (N_7376,N_4789,N_717);
nand U7377 (N_7377,N_432,N_238);
nand U7378 (N_7378,N_2275,N_2025);
xor U7379 (N_7379,N_1828,N_4855);
nor U7380 (N_7380,N_2855,N_4260);
or U7381 (N_7381,N_2219,N_3058);
nor U7382 (N_7382,N_4541,N_4706);
nand U7383 (N_7383,N_2108,N_1997);
or U7384 (N_7384,N_459,N_421);
nand U7385 (N_7385,N_664,N_4762);
xor U7386 (N_7386,N_560,N_2680);
and U7387 (N_7387,N_2907,N_505);
and U7388 (N_7388,N_4696,N_4967);
or U7389 (N_7389,N_1173,N_1481);
or U7390 (N_7390,N_2287,N_4979);
nor U7391 (N_7391,N_1204,N_3822);
nor U7392 (N_7392,N_376,N_26);
and U7393 (N_7393,N_2155,N_1114);
and U7394 (N_7394,N_2008,N_2021);
xor U7395 (N_7395,N_3353,N_3005);
or U7396 (N_7396,N_4836,N_2645);
and U7397 (N_7397,N_4831,N_4783);
xnor U7398 (N_7398,N_1098,N_373);
or U7399 (N_7399,N_313,N_3230);
nand U7400 (N_7400,N_3000,N_2240);
nor U7401 (N_7401,N_842,N_2802);
and U7402 (N_7402,N_3801,N_967);
nor U7403 (N_7403,N_3170,N_2031);
nor U7404 (N_7404,N_990,N_1914);
nor U7405 (N_7405,N_1240,N_2160);
or U7406 (N_7406,N_2142,N_2559);
or U7407 (N_7407,N_970,N_823);
nor U7408 (N_7408,N_3937,N_3489);
or U7409 (N_7409,N_1606,N_112);
xnor U7410 (N_7410,N_2630,N_2367);
nand U7411 (N_7411,N_306,N_3622);
or U7412 (N_7412,N_2444,N_281);
or U7413 (N_7413,N_3796,N_3746);
or U7414 (N_7414,N_1102,N_4879);
nand U7415 (N_7415,N_2204,N_1957);
or U7416 (N_7416,N_2081,N_2335);
xor U7417 (N_7417,N_3107,N_4378);
or U7418 (N_7418,N_2086,N_3666);
xor U7419 (N_7419,N_4470,N_3545);
or U7420 (N_7420,N_3758,N_1063);
xnor U7421 (N_7421,N_2944,N_2620);
nor U7422 (N_7422,N_681,N_1342);
nand U7423 (N_7423,N_2348,N_3143);
or U7424 (N_7424,N_707,N_4464);
xor U7425 (N_7425,N_2196,N_587);
xor U7426 (N_7426,N_4571,N_3856);
nor U7427 (N_7427,N_3503,N_4245);
and U7428 (N_7428,N_1585,N_229);
nand U7429 (N_7429,N_4654,N_787);
xor U7430 (N_7430,N_4777,N_756);
and U7431 (N_7431,N_208,N_4334);
or U7432 (N_7432,N_1666,N_551);
nand U7433 (N_7433,N_4584,N_3633);
xor U7434 (N_7434,N_219,N_2849);
xor U7435 (N_7435,N_3398,N_3626);
nor U7436 (N_7436,N_2157,N_2706);
or U7437 (N_7437,N_290,N_3132);
xnor U7438 (N_7438,N_603,N_1661);
and U7439 (N_7439,N_4864,N_1215);
and U7440 (N_7440,N_1485,N_4948);
nor U7441 (N_7441,N_2778,N_1839);
nand U7442 (N_7442,N_862,N_4024);
nor U7443 (N_7443,N_1247,N_1416);
xnor U7444 (N_7444,N_852,N_3436);
and U7445 (N_7445,N_4316,N_1352);
nand U7446 (N_7446,N_530,N_446);
or U7447 (N_7447,N_1725,N_1635);
nand U7448 (N_7448,N_4641,N_2299);
and U7449 (N_7449,N_4087,N_4710);
nand U7450 (N_7450,N_1386,N_2814);
nand U7451 (N_7451,N_2445,N_1043);
nand U7452 (N_7452,N_2011,N_2670);
nor U7453 (N_7453,N_2606,N_1581);
nand U7454 (N_7454,N_1330,N_4817);
xnor U7455 (N_7455,N_789,N_1269);
xor U7456 (N_7456,N_1638,N_2831);
xnor U7457 (N_7457,N_3144,N_2164);
nand U7458 (N_7458,N_2186,N_298);
nand U7459 (N_7459,N_3893,N_49);
xor U7460 (N_7460,N_3021,N_196);
nand U7461 (N_7461,N_3003,N_2733);
nor U7462 (N_7462,N_3346,N_240);
nor U7463 (N_7463,N_4061,N_1628);
xor U7464 (N_7464,N_2267,N_4585);
nor U7465 (N_7465,N_2324,N_2610);
nor U7466 (N_7466,N_2293,N_4437);
and U7467 (N_7467,N_4223,N_2685);
nor U7468 (N_7468,N_1347,N_136);
or U7469 (N_7469,N_4343,N_1992);
or U7470 (N_7470,N_4406,N_3004);
nor U7471 (N_7471,N_3164,N_1552);
xor U7472 (N_7472,N_3061,N_4326);
nand U7473 (N_7473,N_1161,N_4713);
or U7474 (N_7474,N_3990,N_3030);
or U7475 (N_7475,N_318,N_1122);
xor U7476 (N_7476,N_3729,N_3389);
or U7477 (N_7477,N_1867,N_2105);
or U7478 (N_7478,N_1705,N_4037);
nor U7479 (N_7479,N_1315,N_1373);
nand U7480 (N_7480,N_1038,N_2377);
or U7481 (N_7481,N_866,N_734);
nand U7482 (N_7482,N_2363,N_1044);
or U7483 (N_7483,N_1980,N_453);
and U7484 (N_7484,N_1337,N_1338);
or U7485 (N_7485,N_434,N_1888);
nor U7486 (N_7486,N_276,N_601);
nor U7487 (N_7487,N_1848,N_3036);
nor U7488 (N_7488,N_1146,N_2213);
nor U7489 (N_7489,N_3600,N_2095);
xnor U7490 (N_7490,N_532,N_1823);
nand U7491 (N_7491,N_2446,N_4430);
or U7492 (N_7492,N_179,N_964);
and U7493 (N_7493,N_3286,N_4956);
and U7494 (N_7494,N_1559,N_2235);
nand U7495 (N_7495,N_1335,N_1081);
nand U7496 (N_7496,N_1213,N_455);
xor U7497 (N_7497,N_2910,N_1156);
or U7498 (N_7498,N_1345,N_2427);
and U7499 (N_7499,N_4961,N_914);
nor U7500 (N_7500,N_1174,N_3719);
and U7501 (N_7501,N_3624,N_622);
nor U7502 (N_7502,N_4703,N_1282);
nand U7503 (N_7503,N_2791,N_2313);
and U7504 (N_7504,N_863,N_1747);
xor U7505 (N_7505,N_3978,N_4788);
or U7506 (N_7506,N_939,N_1324);
nand U7507 (N_7507,N_2826,N_4195);
or U7508 (N_7508,N_567,N_2770);
or U7509 (N_7509,N_203,N_3896);
or U7510 (N_7510,N_3125,N_3292);
and U7511 (N_7511,N_319,N_3588);
nor U7512 (N_7512,N_126,N_64);
xor U7513 (N_7513,N_123,N_256);
nor U7514 (N_7514,N_4380,N_2782);
and U7515 (N_7515,N_581,N_2921);
nand U7516 (N_7516,N_839,N_3125);
nand U7517 (N_7517,N_2913,N_1199);
and U7518 (N_7518,N_886,N_4061);
nand U7519 (N_7519,N_366,N_2822);
nand U7520 (N_7520,N_2394,N_4618);
and U7521 (N_7521,N_2627,N_646);
xor U7522 (N_7522,N_871,N_1930);
nor U7523 (N_7523,N_2937,N_3353);
nand U7524 (N_7524,N_2943,N_2687);
xnor U7525 (N_7525,N_1560,N_3218);
or U7526 (N_7526,N_102,N_1811);
nand U7527 (N_7527,N_3397,N_430);
or U7528 (N_7528,N_3306,N_144);
and U7529 (N_7529,N_1135,N_1810);
nand U7530 (N_7530,N_894,N_3953);
and U7531 (N_7531,N_4553,N_4191);
xor U7532 (N_7532,N_3824,N_4886);
or U7533 (N_7533,N_4545,N_1272);
or U7534 (N_7534,N_3303,N_4144);
and U7535 (N_7535,N_464,N_4078);
xnor U7536 (N_7536,N_4748,N_1462);
nor U7537 (N_7537,N_1704,N_139);
nor U7538 (N_7538,N_4065,N_2455);
or U7539 (N_7539,N_2865,N_2270);
nor U7540 (N_7540,N_3437,N_3015);
nand U7541 (N_7541,N_762,N_581);
nor U7542 (N_7542,N_4648,N_2646);
nor U7543 (N_7543,N_1320,N_759);
or U7544 (N_7544,N_2460,N_1247);
and U7545 (N_7545,N_4852,N_2548);
or U7546 (N_7546,N_2896,N_3525);
nor U7547 (N_7547,N_462,N_3810);
nand U7548 (N_7548,N_3205,N_2324);
or U7549 (N_7549,N_3298,N_163);
nand U7550 (N_7550,N_1454,N_3162);
or U7551 (N_7551,N_108,N_11);
and U7552 (N_7552,N_915,N_2354);
xor U7553 (N_7553,N_2951,N_693);
nor U7554 (N_7554,N_3429,N_4213);
xnor U7555 (N_7555,N_346,N_3939);
nor U7556 (N_7556,N_2006,N_1977);
xnor U7557 (N_7557,N_4120,N_1944);
nand U7558 (N_7558,N_277,N_4149);
and U7559 (N_7559,N_3006,N_2183);
nand U7560 (N_7560,N_1524,N_340);
nor U7561 (N_7561,N_4353,N_3929);
and U7562 (N_7562,N_1275,N_4049);
and U7563 (N_7563,N_1124,N_4649);
and U7564 (N_7564,N_2791,N_919);
nand U7565 (N_7565,N_3577,N_1495);
xnor U7566 (N_7566,N_4645,N_2285);
or U7567 (N_7567,N_2146,N_42);
or U7568 (N_7568,N_4448,N_1859);
nand U7569 (N_7569,N_1648,N_3768);
or U7570 (N_7570,N_3892,N_3076);
xor U7571 (N_7571,N_1858,N_2331);
and U7572 (N_7572,N_2235,N_3552);
nor U7573 (N_7573,N_730,N_2613);
or U7574 (N_7574,N_2956,N_3804);
or U7575 (N_7575,N_349,N_30);
and U7576 (N_7576,N_1817,N_1158);
nor U7577 (N_7577,N_175,N_2576);
or U7578 (N_7578,N_2337,N_4519);
xnor U7579 (N_7579,N_4938,N_948);
nor U7580 (N_7580,N_973,N_4151);
nor U7581 (N_7581,N_1423,N_2520);
and U7582 (N_7582,N_1219,N_4817);
and U7583 (N_7583,N_4687,N_694);
or U7584 (N_7584,N_996,N_1248);
nand U7585 (N_7585,N_3483,N_2519);
or U7586 (N_7586,N_2221,N_4841);
nor U7587 (N_7587,N_3326,N_2831);
and U7588 (N_7588,N_2689,N_793);
or U7589 (N_7589,N_3064,N_2938);
and U7590 (N_7590,N_4983,N_3701);
or U7591 (N_7591,N_1199,N_719);
or U7592 (N_7592,N_4229,N_4504);
nor U7593 (N_7593,N_2809,N_1725);
nor U7594 (N_7594,N_4280,N_1217);
or U7595 (N_7595,N_1375,N_2698);
and U7596 (N_7596,N_1991,N_937);
and U7597 (N_7597,N_4198,N_1787);
nand U7598 (N_7598,N_4896,N_4883);
and U7599 (N_7599,N_1906,N_295);
nor U7600 (N_7600,N_3188,N_4414);
or U7601 (N_7601,N_3021,N_2655);
and U7602 (N_7602,N_4194,N_1537);
nor U7603 (N_7603,N_4900,N_31);
xnor U7604 (N_7604,N_3292,N_2627);
xnor U7605 (N_7605,N_3401,N_1242);
and U7606 (N_7606,N_2776,N_566);
nand U7607 (N_7607,N_4887,N_2359);
and U7608 (N_7608,N_3668,N_556);
and U7609 (N_7609,N_408,N_42);
nand U7610 (N_7610,N_73,N_4893);
nor U7611 (N_7611,N_3506,N_3598);
nand U7612 (N_7612,N_4593,N_4187);
nand U7613 (N_7613,N_4122,N_654);
or U7614 (N_7614,N_2530,N_2448);
or U7615 (N_7615,N_4974,N_861);
or U7616 (N_7616,N_1034,N_4588);
or U7617 (N_7617,N_2653,N_1041);
nor U7618 (N_7618,N_1566,N_2683);
nor U7619 (N_7619,N_444,N_1931);
and U7620 (N_7620,N_4099,N_391);
xnor U7621 (N_7621,N_591,N_1612);
and U7622 (N_7622,N_1497,N_1160);
or U7623 (N_7623,N_2682,N_706);
nor U7624 (N_7624,N_434,N_3230);
or U7625 (N_7625,N_2562,N_1929);
and U7626 (N_7626,N_4810,N_544);
xor U7627 (N_7627,N_3955,N_1128);
xnor U7628 (N_7628,N_1038,N_4628);
xnor U7629 (N_7629,N_59,N_606);
nand U7630 (N_7630,N_771,N_1596);
or U7631 (N_7631,N_4880,N_4511);
xor U7632 (N_7632,N_3590,N_2317);
nand U7633 (N_7633,N_2258,N_2947);
xor U7634 (N_7634,N_3645,N_3853);
nand U7635 (N_7635,N_4546,N_1066);
nor U7636 (N_7636,N_233,N_3216);
and U7637 (N_7637,N_4819,N_250);
nand U7638 (N_7638,N_2232,N_1922);
or U7639 (N_7639,N_2477,N_765);
nand U7640 (N_7640,N_347,N_1454);
nor U7641 (N_7641,N_4952,N_984);
xnor U7642 (N_7642,N_4817,N_2970);
and U7643 (N_7643,N_1907,N_1454);
xnor U7644 (N_7644,N_4111,N_2054);
and U7645 (N_7645,N_3699,N_3711);
nor U7646 (N_7646,N_1535,N_1793);
and U7647 (N_7647,N_2345,N_1920);
xnor U7648 (N_7648,N_628,N_1559);
nor U7649 (N_7649,N_1800,N_3673);
and U7650 (N_7650,N_2746,N_2409);
or U7651 (N_7651,N_390,N_2169);
and U7652 (N_7652,N_1551,N_2895);
nor U7653 (N_7653,N_2177,N_1561);
or U7654 (N_7654,N_1346,N_3926);
and U7655 (N_7655,N_1911,N_3992);
xor U7656 (N_7656,N_2683,N_817);
nor U7657 (N_7657,N_61,N_1090);
xnor U7658 (N_7658,N_3849,N_3689);
or U7659 (N_7659,N_3824,N_201);
nand U7660 (N_7660,N_1316,N_3628);
xor U7661 (N_7661,N_3773,N_567);
nor U7662 (N_7662,N_1140,N_3900);
and U7663 (N_7663,N_4639,N_1762);
xor U7664 (N_7664,N_2718,N_4237);
or U7665 (N_7665,N_2102,N_2851);
xor U7666 (N_7666,N_2150,N_3859);
nor U7667 (N_7667,N_1869,N_4701);
and U7668 (N_7668,N_2606,N_4913);
nand U7669 (N_7669,N_2816,N_882);
xor U7670 (N_7670,N_3286,N_3884);
or U7671 (N_7671,N_1549,N_1066);
xor U7672 (N_7672,N_3906,N_215);
or U7673 (N_7673,N_3119,N_2981);
and U7674 (N_7674,N_3598,N_2622);
or U7675 (N_7675,N_3840,N_2961);
nor U7676 (N_7676,N_3869,N_4881);
xor U7677 (N_7677,N_4374,N_639);
xor U7678 (N_7678,N_2896,N_921);
or U7679 (N_7679,N_802,N_2428);
and U7680 (N_7680,N_851,N_4498);
and U7681 (N_7681,N_2472,N_2359);
nand U7682 (N_7682,N_1950,N_3807);
nand U7683 (N_7683,N_2488,N_966);
nor U7684 (N_7684,N_1098,N_650);
nor U7685 (N_7685,N_2384,N_1914);
nand U7686 (N_7686,N_1428,N_2685);
nand U7687 (N_7687,N_2063,N_824);
nor U7688 (N_7688,N_2592,N_1750);
xnor U7689 (N_7689,N_156,N_1127);
nand U7690 (N_7690,N_36,N_297);
and U7691 (N_7691,N_1685,N_2017);
or U7692 (N_7692,N_2218,N_4546);
xnor U7693 (N_7693,N_4998,N_2866);
or U7694 (N_7694,N_2889,N_512);
nor U7695 (N_7695,N_1158,N_1840);
or U7696 (N_7696,N_217,N_3654);
and U7697 (N_7697,N_3879,N_2101);
and U7698 (N_7698,N_3522,N_4926);
xnor U7699 (N_7699,N_2721,N_1714);
or U7700 (N_7700,N_4678,N_1093);
xnor U7701 (N_7701,N_1410,N_4211);
and U7702 (N_7702,N_4091,N_2927);
nor U7703 (N_7703,N_2432,N_888);
or U7704 (N_7704,N_3775,N_2749);
or U7705 (N_7705,N_22,N_24);
nor U7706 (N_7706,N_3986,N_1231);
or U7707 (N_7707,N_4481,N_298);
or U7708 (N_7708,N_1501,N_2643);
and U7709 (N_7709,N_3764,N_4951);
nand U7710 (N_7710,N_3640,N_256);
or U7711 (N_7711,N_2472,N_4303);
and U7712 (N_7712,N_1219,N_2811);
nor U7713 (N_7713,N_3497,N_3761);
xnor U7714 (N_7714,N_4249,N_4184);
nor U7715 (N_7715,N_4802,N_3624);
xor U7716 (N_7716,N_4428,N_2023);
nor U7717 (N_7717,N_1370,N_2757);
or U7718 (N_7718,N_3758,N_3233);
xnor U7719 (N_7719,N_4686,N_1838);
nor U7720 (N_7720,N_3534,N_2624);
or U7721 (N_7721,N_4355,N_545);
nand U7722 (N_7722,N_376,N_2838);
nor U7723 (N_7723,N_603,N_2772);
nor U7724 (N_7724,N_1965,N_62);
nor U7725 (N_7725,N_3477,N_3544);
nand U7726 (N_7726,N_3432,N_2270);
or U7727 (N_7727,N_2242,N_2021);
nor U7728 (N_7728,N_2320,N_795);
xor U7729 (N_7729,N_3082,N_3627);
xnor U7730 (N_7730,N_3597,N_2697);
nor U7731 (N_7731,N_3484,N_4982);
nor U7732 (N_7732,N_4961,N_3290);
nand U7733 (N_7733,N_1104,N_1033);
xor U7734 (N_7734,N_4975,N_1007);
nor U7735 (N_7735,N_3379,N_4860);
xor U7736 (N_7736,N_1309,N_4914);
and U7737 (N_7737,N_39,N_3271);
nor U7738 (N_7738,N_3252,N_1298);
or U7739 (N_7739,N_1448,N_1632);
or U7740 (N_7740,N_2487,N_4145);
xor U7741 (N_7741,N_301,N_3305);
nor U7742 (N_7742,N_1131,N_2486);
nor U7743 (N_7743,N_3089,N_1881);
nand U7744 (N_7744,N_2088,N_1905);
and U7745 (N_7745,N_3149,N_1472);
nor U7746 (N_7746,N_1071,N_2610);
nor U7747 (N_7747,N_94,N_3677);
nand U7748 (N_7748,N_2581,N_1221);
nor U7749 (N_7749,N_1703,N_1674);
nand U7750 (N_7750,N_1704,N_727);
xor U7751 (N_7751,N_1592,N_4493);
xor U7752 (N_7752,N_3395,N_3661);
or U7753 (N_7753,N_4286,N_4211);
and U7754 (N_7754,N_3769,N_664);
nor U7755 (N_7755,N_3194,N_1707);
and U7756 (N_7756,N_2986,N_525);
nand U7757 (N_7757,N_1103,N_4591);
or U7758 (N_7758,N_1508,N_1899);
or U7759 (N_7759,N_238,N_1852);
nand U7760 (N_7760,N_848,N_2095);
nor U7761 (N_7761,N_3940,N_3572);
and U7762 (N_7762,N_1166,N_4921);
and U7763 (N_7763,N_3212,N_111);
xnor U7764 (N_7764,N_4104,N_2164);
xor U7765 (N_7765,N_1326,N_4147);
nand U7766 (N_7766,N_848,N_3104);
nand U7767 (N_7767,N_258,N_1543);
or U7768 (N_7768,N_2027,N_3428);
nand U7769 (N_7769,N_1515,N_3346);
nor U7770 (N_7770,N_2611,N_2399);
nand U7771 (N_7771,N_4767,N_1267);
or U7772 (N_7772,N_2460,N_3097);
and U7773 (N_7773,N_1782,N_3656);
nor U7774 (N_7774,N_907,N_4528);
xnor U7775 (N_7775,N_1747,N_1622);
or U7776 (N_7776,N_3618,N_4196);
and U7777 (N_7777,N_2663,N_281);
and U7778 (N_7778,N_1067,N_2314);
or U7779 (N_7779,N_4766,N_4491);
xnor U7780 (N_7780,N_1758,N_1629);
or U7781 (N_7781,N_2048,N_3228);
or U7782 (N_7782,N_1541,N_207);
xnor U7783 (N_7783,N_4399,N_3261);
nand U7784 (N_7784,N_1412,N_4861);
nor U7785 (N_7785,N_3818,N_1691);
nor U7786 (N_7786,N_422,N_679);
nand U7787 (N_7787,N_115,N_1836);
and U7788 (N_7788,N_3329,N_2074);
nand U7789 (N_7789,N_3021,N_2484);
nor U7790 (N_7790,N_257,N_3125);
nor U7791 (N_7791,N_4975,N_2829);
and U7792 (N_7792,N_3540,N_4829);
nor U7793 (N_7793,N_637,N_3765);
and U7794 (N_7794,N_2490,N_2318);
and U7795 (N_7795,N_1442,N_4230);
or U7796 (N_7796,N_2120,N_4323);
nor U7797 (N_7797,N_643,N_288);
nor U7798 (N_7798,N_4326,N_3577);
and U7799 (N_7799,N_1964,N_4544);
xor U7800 (N_7800,N_466,N_4769);
nand U7801 (N_7801,N_221,N_1199);
xor U7802 (N_7802,N_1274,N_1296);
nand U7803 (N_7803,N_1708,N_1208);
and U7804 (N_7804,N_2473,N_4266);
nor U7805 (N_7805,N_3579,N_2900);
nand U7806 (N_7806,N_316,N_2060);
nor U7807 (N_7807,N_3502,N_1128);
nand U7808 (N_7808,N_3162,N_2042);
and U7809 (N_7809,N_1000,N_4081);
nand U7810 (N_7810,N_3986,N_2458);
and U7811 (N_7811,N_3267,N_4296);
or U7812 (N_7812,N_2006,N_2707);
xnor U7813 (N_7813,N_3894,N_4455);
or U7814 (N_7814,N_526,N_2072);
nand U7815 (N_7815,N_3418,N_936);
nor U7816 (N_7816,N_4309,N_4527);
and U7817 (N_7817,N_4927,N_3296);
nor U7818 (N_7818,N_731,N_2571);
and U7819 (N_7819,N_3705,N_2440);
and U7820 (N_7820,N_4541,N_3333);
nand U7821 (N_7821,N_4521,N_1709);
xnor U7822 (N_7822,N_3709,N_1035);
nor U7823 (N_7823,N_1769,N_2395);
and U7824 (N_7824,N_1741,N_4529);
nand U7825 (N_7825,N_4903,N_4851);
nor U7826 (N_7826,N_1493,N_4683);
nand U7827 (N_7827,N_1381,N_4630);
nor U7828 (N_7828,N_3361,N_3087);
or U7829 (N_7829,N_2648,N_1835);
or U7830 (N_7830,N_217,N_270);
and U7831 (N_7831,N_3799,N_2133);
or U7832 (N_7832,N_1696,N_1752);
xor U7833 (N_7833,N_3543,N_2806);
or U7834 (N_7834,N_967,N_2182);
or U7835 (N_7835,N_3444,N_3496);
or U7836 (N_7836,N_2708,N_4055);
and U7837 (N_7837,N_3338,N_3807);
nand U7838 (N_7838,N_1570,N_3498);
or U7839 (N_7839,N_82,N_4530);
xnor U7840 (N_7840,N_847,N_2418);
or U7841 (N_7841,N_256,N_389);
nand U7842 (N_7842,N_2170,N_3166);
nand U7843 (N_7843,N_2425,N_4825);
and U7844 (N_7844,N_4515,N_2298);
and U7845 (N_7845,N_2913,N_2034);
or U7846 (N_7846,N_1579,N_2479);
nor U7847 (N_7847,N_4072,N_4442);
or U7848 (N_7848,N_4961,N_1910);
nand U7849 (N_7849,N_3651,N_1976);
nand U7850 (N_7850,N_3001,N_2103);
nand U7851 (N_7851,N_2084,N_179);
nand U7852 (N_7852,N_750,N_478);
and U7853 (N_7853,N_2921,N_3497);
and U7854 (N_7854,N_1158,N_1889);
xnor U7855 (N_7855,N_4109,N_3555);
and U7856 (N_7856,N_410,N_129);
or U7857 (N_7857,N_3888,N_3444);
nor U7858 (N_7858,N_3746,N_2341);
xor U7859 (N_7859,N_4583,N_4015);
or U7860 (N_7860,N_2041,N_2939);
or U7861 (N_7861,N_1535,N_1324);
or U7862 (N_7862,N_807,N_3037);
nand U7863 (N_7863,N_4651,N_3042);
xor U7864 (N_7864,N_830,N_4852);
and U7865 (N_7865,N_3714,N_2752);
or U7866 (N_7866,N_4724,N_1990);
nor U7867 (N_7867,N_1438,N_3575);
nor U7868 (N_7868,N_925,N_4244);
nor U7869 (N_7869,N_4699,N_134);
and U7870 (N_7870,N_4920,N_3736);
xor U7871 (N_7871,N_1398,N_940);
xor U7872 (N_7872,N_556,N_3087);
or U7873 (N_7873,N_2465,N_1129);
or U7874 (N_7874,N_1769,N_2422);
nor U7875 (N_7875,N_3804,N_3820);
nand U7876 (N_7876,N_4094,N_3528);
nand U7877 (N_7877,N_4090,N_1214);
nor U7878 (N_7878,N_4558,N_4663);
and U7879 (N_7879,N_975,N_1433);
or U7880 (N_7880,N_3691,N_3102);
or U7881 (N_7881,N_3670,N_145);
nand U7882 (N_7882,N_298,N_2694);
nand U7883 (N_7883,N_3846,N_4199);
nor U7884 (N_7884,N_59,N_2253);
and U7885 (N_7885,N_2342,N_4853);
nor U7886 (N_7886,N_3425,N_4218);
nor U7887 (N_7887,N_2050,N_4676);
or U7888 (N_7888,N_725,N_462);
and U7889 (N_7889,N_2816,N_69);
xnor U7890 (N_7890,N_4909,N_1399);
nand U7891 (N_7891,N_924,N_3499);
and U7892 (N_7892,N_3623,N_2644);
nor U7893 (N_7893,N_4731,N_3240);
xnor U7894 (N_7894,N_3446,N_3911);
nor U7895 (N_7895,N_1864,N_1279);
nand U7896 (N_7896,N_2720,N_3679);
and U7897 (N_7897,N_581,N_408);
nor U7898 (N_7898,N_3205,N_731);
and U7899 (N_7899,N_4658,N_1998);
or U7900 (N_7900,N_2491,N_85);
nor U7901 (N_7901,N_2117,N_1860);
and U7902 (N_7902,N_837,N_4190);
nor U7903 (N_7903,N_2058,N_1714);
and U7904 (N_7904,N_782,N_19);
and U7905 (N_7905,N_2281,N_4267);
xnor U7906 (N_7906,N_461,N_964);
or U7907 (N_7907,N_2848,N_908);
xnor U7908 (N_7908,N_863,N_3796);
and U7909 (N_7909,N_1808,N_2139);
and U7910 (N_7910,N_719,N_1249);
nor U7911 (N_7911,N_3687,N_2952);
nor U7912 (N_7912,N_4097,N_1285);
xor U7913 (N_7913,N_4645,N_1095);
nand U7914 (N_7914,N_3756,N_3037);
or U7915 (N_7915,N_3347,N_1957);
nor U7916 (N_7916,N_2385,N_4637);
nand U7917 (N_7917,N_2793,N_3199);
and U7918 (N_7918,N_2753,N_2609);
nand U7919 (N_7919,N_4792,N_4160);
xnor U7920 (N_7920,N_3121,N_837);
and U7921 (N_7921,N_4110,N_490);
xnor U7922 (N_7922,N_3921,N_312);
and U7923 (N_7923,N_2890,N_2928);
or U7924 (N_7924,N_365,N_2049);
xor U7925 (N_7925,N_2686,N_1534);
nor U7926 (N_7926,N_2997,N_4725);
nand U7927 (N_7927,N_4852,N_1702);
nor U7928 (N_7928,N_1665,N_1836);
nor U7929 (N_7929,N_3606,N_1879);
nor U7930 (N_7930,N_1771,N_670);
nor U7931 (N_7931,N_4190,N_2811);
nand U7932 (N_7932,N_3176,N_3518);
nand U7933 (N_7933,N_3693,N_820);
and U7934 (N_7934,N_2486,N_1967);
or U7935 (N_7935,N_2882,N_4419);
xor U7936 (N_7936,N_2972,N_4817);
xor U7937 (N_7937,N_2072,N_2917);
nand U7938 (N_7938,N_2691,N_4162);
or U7939 (N_7939,N_557,N_3066);
xor U7940 (N_7940,N_1333,N_4837);
nand U7941 (N_7941,N_3200,N_2531);
or U7942 (N_7942,N_381,N_1832);
and U7943 (N_7943,N_2621,N_509);
nor U7944 (N_7944,N_2958,N_2122);
nand U7945 (N_7945,N_3068,N_989);
nor U7946 (N_7946,N_461,N_2077);
xnor U7947 (N_7947,N_1090,N_4606);
or U7948 (N_7948,N_3699,N_602);
xnor U7949 (N_7949,N_612,N_18);
or U7950 (N_7950,N_1040,N_868);
nand U7951 (N_7951,N_1713,N_167);
or U7952 (N_7952,N_2386,N_4451);
xnor U7953 (N_7953,N_1892,N_4901);
nor U7954 (N_7954,N_4310,N_2662);
nor U7955 (N_7955,N_1226,N_357);
nand U7956 (N_7956,N_4029,N_1958);
nand U7957 (N_7957,N_1830,N_4503);
nor U7958 (N_7958,N_4370,N_1956);
or U7959 (N_7959,N_471,N_2683);
nand U7960 (N_7960,N_4186,N_4940);
nand U7961 (N_7961,N_1793,N_2747);
or U7962 (N_7962,N_4054,N_2050);
and U7963 (N_7963,N_1779,N_4509);
nand U7964 (N_7964,N_1629,N_3306);
xnor U7965 (N_7965,N_4731,N_1807);
nand U7966 (N_7966,N_800,N_3094);
xor U7967 (N_7967,N_166,N_2897);
xnor U7968 (N_7968,N_3435,N_19);
or U7969 (N_7969,N_237,N_1066);
nand U7970 (N_7970,N_3015,N_3003);
or U7971 (N_7971,N_599,N_2305);
xnor U7972 (N_7972,N_860,N_4893);
and U7973 (N_7973,N_1368,N_1899);
xnor U7974 (N_7974,N_97,N_248);
nand U7975 (N_7975,N_792,N_4303);
nor U7976 (N_7976,N_4140,N_3166);
xor U7977 (N_7977,N_4236,N_1015);
xor U7978 (N_7978,N_1835,N_2662);
or U7979 (N_7979,N_967,N_964);
nand U7980 (N_7980,N_2594,N_2858);
and U7981 (N_7981,N_464,N_2024);
nand U7982 (N_7982,N_4876,N_1502);
and U7983 (N_7983,N_529,N_569);
and U7984 (N_7984,N_372,N_1080);
or U7985 (N_7985,N_4787,N_1303);
or U7986 (N_7986,N_4771,N_4682);
xor U7987 (N_7987,N_4452,N_3201);
nand U7988 (N_7988,N_2677,N_3627);
nand U7989 (N_7989,N_2791,N_943);
and U7990 (N_7990,N_1538,N_1262);
and U7991 (N_7991,N_3014,N_3631);
or U7992 (N_7992,N_4235,N_806);
xor U7993 (N_7993,N_1488,N_3202);
or U7994 (N_7994,N_4276,N_265);
and U7995 (N_7995,N_1927,N_4867);
nor U7996 (N_7996,N_1495,N_4102);
nor U7997 (N_7997,N_2727,N_86);
or U7998 (N_7998,N_3632,N_2359);
xor U7999 (N_7999,N_4784,N_3305);
and U8000 (N_8000,N_1574,N_1682);
or U8001 (N_8001,N_3748,N_2494);
nand U8002 (N_8002,N_1973,N_4969);
and U8003 (N_8003,N_3462,N_1551);
nand U8004 (N_8004,N_4808,N_1223);
or U8005 (N_8005,N_247,N_971);
or U8006 (N_8006,N_4165,N_4707);
nor U8007 (N_8007,N_689,N_4840);
nand U8008 (N_8008,N_2128,N_3962);
nor U8009 (N_8009,N_1052,N_2042);
nand U8010 (N_8010,N_4926,N_1514);
nor U8011 (N_8011,N_2677,N_1810);
xor U8012 (N_8012,N_3894,N_205);
and U8013 (N_8013,N_2457,N_2845);
nand U8014 (N_8014,N_622,N_2339);
xor U8015 (N_8015,N_2391,N_4208);
and U8016 (N_8016,N_3930,N_2277);
and U8017 (N_8017,N_65,N_3975);
and U8018 (N_8018,N_2140,N_3845);
nand U8019 (N_8019,N_301,N_756);
or U8020 (N_8020,N_3758,N_2053);
xor U8021 (N_8021,N_3183,N_463);
or U8022 (N_8022,N_1035,N_2845);
or U8023 (N_8023,N_1333,N_4923);
xnor U8024 (N_8024,N_3671,N_1379);
xnor U8025 (N_8025,N_3833,N_1853);
or U8026 (N_8026,N_4415,N_254);
nand U8027 (N_8027,N_2899,N_1043);
or U8028 (N_8028,N_2789,N_4728);
and U8029 (N_8029,N_2209,N_4251);
or U8030 (N_8030,N_756,N_1529);
nand U8031 (N_8031,N_3721,N_365);
xor U8032 (N_8032,N_1309,N_2631);
or U8033 (N_8033,N_504,N_3609);
or U8034 (N_8034,N_252,N_825);
or U8035 (N_8035,N_1071,N_4033);
xnor U8036 (N_8036,N_861,N_835);
or U8037 (N_8037,N_3770,N_2277);
and U8038 (N_8038,N_3049,N_464);
nor U8039 (N_8039,N_420,N_1193);
nor U8040 (N_8040,N_3719,N_3151);
nand U8041 (N_8041,N_4697,N_3252);
nand U8042 (N_8042,N_1018,N_240);
nor U8043 (N_8043,N_2622,N_2316);
and U8044 (N_8044,N_2964,N_535);
nor U8045 (N_8045,N_838,N_2245);
nor U8046 (N_8046,N_3900,N_2044);
xnor U8047 (N_8047,N_4756,N_2069);
nor U8048 (N_8048,N_4792,N_1170);
xor U8049 (N_8049,N_101,N_3572);
or U8050 (N_8050,N_1212,N_2593);
or U8051 (N_8051,N_2561,N_3883);
nor U8052 (N_8052,N_1425,N_3821);
xor U8053 (N_8053,N_959,N_3807);
nor U8054 (N_8054,N_3367,N_3639);
xor U8055 (N_8055,N_4561,N_264);
or U8056 (N_8056,N_549,N_2610);
xnor U8057 (N_8057,N_3867,N_967);
xor U8058 (N_8058,N_3281,N_1801);
and U8059 (N_8059,N_2292,N_71);
or U8060 (N_8060,N_1617,N_3203);
xor U8061 (N_8061,N_2057,N_4517);
xor U8062 (N_8062,N_4516,N_1644);
xnor U8063 (N_8063,N_2437,N_4430);
nand U8064 (N_8064,N_2139,N_228);
and U8065 (N_8065,N_243,N_2863);
or U8066 (N_8066,N_814,N_1051);
nand U8067 (N_8067,N_3605,N_3271);
xor U8068 (N_8068,N_1201,N_2620);
and U8069 (N_8069,N_3146,N_4620);
xnor U8070 (N_8070,N_4453,N_991);
and U8071 (N_8071,N_803,N_3397);
and U8072 (N_8072,N_752,N_2374);
xnor U8073 (N_8073,N_4744,N_1842);
or U8074 (N_8074,N_1524,N_4735);
xor U8075 (N_8075,N_251,N_369);
and U8076 (N_8076,N_3008,N_2741);
and U8077 (N_8077,N_721,N_3960);
nor U8078 (N_8078,N_2506,N_1790);
or U8079 (N_8079,N_3170,N_30);
and U8080 (N_8080,N_2011,N_2424);
and U8081 (N_8081,N_7,N_474);
nand U8082 (N_8082,N_1016,N_3705);
xor U8083 (N_8083,N_2559,N_1209);
and U8084 (N_8084,N_1815,N_1921);
and U8085 (N_8085,N_1068,N_4382);
nor U8086 (N_8086,N_4325,N_417);
or U8087 (N_8087,N_3634,N_4986);
xor U8088 (N_8088,N_3899,N_1255);
nor U8089 (N_8089,N_2568,N_3218);
and U8090 (N_8090,N_2424,N_3455);
and U8091 (N_8091,N_3224,N_2217);
nand U8092 (N_8092,N_994,N_208);
nor U8093 (N_8093,N_2070,N_4840);
nor U8094 (N_8094,N_1383,N_3647);
and U8095 (N_8095,N_889,N_759);
and U8096 (N_8096,N_2074,N_4638);
and U8097 (N_8097,N_2755,N_4326);
or U8098 (N_8098,N_4834,N_4579);
and U8099 (N_8099,N_3886,N_2425);
nor U8100 (N_8100,N_821,N_887);
nand U8101 (N_8101,N_2304,N_3452);
nor U8102 (N_8102,N_4977,N_1423);
or U8103 (N_8103,N_4189,N_1171);
nand U8104 (N_8104,N_2432,N_1972);
xor U8105 (N_8105,N_3169,N_4671);
or U8106 (N_8106,N_2393,N_4855);
xor U8107 (N_8107,N_4354,N_3551);
nand U8108 (N_8108,N_1069,N_3524);
or U8109 (N_8109,N_4754,N_2476);
nand U8110 (N_8110,N_1014,N_759);
or U8111 (N_8111,N_2459,N_1577);
nand U8112 (N_8112,N_602,N_2759);
and U8113 (N_8113,N_1751,N_3624);
or U8114 (N_8114,N_1011,N_1322);
nand U8115 (N_8115,N_2988,N_2243);
or U8116 (N_8116,N_1571,N_4163);
or U8117 (N_8117,N_606,N_498);
nand U8118 (N_8118,N_4238,N_1302);
nand U8119 (N_8119,N_1621,N_2659);
xnor U8120 (N_8120,N_3554,N_419);
or U8121 (N_8121,N_1870,N_1688);
nand U8122 (N_8122,N_4995,N_3846);
xnor U8123 (N_8123,N_4490,N_2323);
nor U8124 (N_8124,N_1245,N_2547);
nor U8125 (N_8125,N_4857,N_4230);
nand U8126 (N_8126,N_3065,N_1584);
and U8127 (N_8127,N_4466,N_2702);
and U8128 (N_8128,N_3034,N_2076);
or U8129 (N_8129,N_1122,N_460);
xor U8130 (N_8130,N_3251,N_2392);
xor U8131 (N_8131,N_437,N_472);
nand U8132 (N_8132,N_1150,N_223);
or U8133 (N_8133,N_1748,N_2878);
xnor U8134 (N_8134,N_449,N_541);
and U8135 (N_8135,N_4019,N_1505);
nor U8136 (N_8136,N_2709,N_780);
xnor U8137 (N_8137,N_4101,N_3297);
or U8138 (N_8138,N_2173,N_3014);
nor U8139 (N_8139,N_3838,N_2269);
nor U8140 (N_8140,N_4323,N_4830);
nor U8141 (N_8141,N_2002,N_4375);
or U8142 (N_8142,N_2846,N_200);
or U8143 (N_8143,N_1352,N_4905);
and U8144 (N_8144,N_921,N_2913);
or U8145 (N_8145,N_3588,N_986);
or U8146 (N_8146,N_3744,N_1489);
nand U8147 (N_8147,N_2410,N_335);
and U8148 (N_8148,N_276,N_3022);
and U8149 (N_8149,N_388,N_2964);
nor U8150 (N_8150,N_1320,N_301);
or U8151 (N_8151,N_709,N_962);
nor U8152 (N_8152,N_2666,N_494);
or U8153 (N_8153,N_1513,N_3642);
or U8154 (N_8154,N_4269,N_571);
xnor U8155 (N_8155,N_843,N_4288);
nor U8156 (N_8156,N_445,N_2029);
nor U8157 (N_8157,N_4963,N_2040);
nor U8158 (N_8158,N_817,N_137);
nor U8159 (N_8159,N_1385,N_37);
and U8160 (N_8160,N_4766,N_4176);
and U8161 (N_8161,N_1411,N_1384);
nor U8162 (N_8162,N_912,N_1634);
nand U8163 (N_8163,N_1375,N_4394);
or U8164 (N_8164,N_1212,N_3779);
and U8165 (N_8165,N_3178,N_1761);
nor U8166 (N_8166,N_2343,N_2851);
nand U8167 (N_8167,N_1404,N_3760);
xor U8168 (N_8168,N_793,N_4283);
nand U8169 (N_8169,N_3904,N_1670);
xor U8170 (N_8170,N_1226,N_1007);
and U8171 (N_8171,N_2061,N_325);
xnor U8172 (N_8172,N_2165,N_1591);
nand U8173 (N_8173,N_2024,N_2707);
nand U8174 (N_8174,N_4550,N_680);
and U8175 (N_8175,N_4617,N_1188);
and U8176 (N_8176,N_4809,N_1041);
nor U8177 (N_8177,N_1703,N_1590);
nor U8178 (N_8178,N_4529,N_2534);
nor U8179 (N_8179,N_4269,N_2130);
or U8180 (N_8180,N_688,N_2608);
and U8181 (N_8181,N_4352,N_4975);
nand U8182 (N_8182,N_699,N_4890);
nor U8183 (N_8183,N_4612,N_3686);
or U8184 (N_8184,N_2346,N_2961);
nand U8185 (N_8185,N_2850,N_2573);
nor U8186 (N_8186,N_4608,N_4638);
xor U8187 (N_8187,N_1729,N_2652);
nor U8188 (N_8188,N_2733,N_38);
nand U8189 (N_8189,N_402,N_3885);
xor U8190 (N_8190,N_1993,N_4223);
and U8191 (N_8191,N_2058,N_3545);
xor U8192 (N_8192,N_1053,N_357);
xnor U8193 (N_8193,N_2533,N_2727);
xnor U8194 (N_8194,N_2087,N_1532);
and U8195 (N_8195,N_3630,N_639);
and U8196 (N_8196,N_2043,N_517);
or U8197 (N_8197,N_3116,N_516);
nand U8198 (N_8198,N_4834,N_3493);
or U8199 (N_8199,N_1649,N_2491);
xnor U8200 (N_8200,N_2945,N_3489);
or U8201 (N_8201,N_193,N_3936);
and U8202 (N_8202,N_4051,N_2025);
xor U8203 (N_8203,N_4513,N_543);
or U8204 (N_8204,N_2841,N_2714);
nor U8205 (N_8205,N_2165,N_3716);
or U8206 (N_8206,N_3495,N_4653);
or U8207 (N_8207,N_1403,N_3895);
or U8208 (N_8208,N_4034,N_2363);
nor U8209 (N_8209,N_1271,N_988);
xor U8210 (N_8210,N_4915,N_1885);
nor U8211 (N_8211,N_4323,N_4683);
xor U8212 (N_8212,N_1360,N_1475);
nor U8213 (N_8213,N_4115,N_3249);
xor U8214 (N_8214,N_978,N_3111);
or U8215 (N_8215,N_4542,N_2885);
or U8216 (N_8216,N_2042,N_4817);
xnor U8217 (N_8217,N_2369,N_232);
and U8218 (N_8218,N_1729,N_2811);
nor U8219 (N_8219,N_4369,N_3407);
nand U8220 (N_8220,N_4228,N_3522);
xnor U8221 (N_8221,N_1062,N_4112);
or U8222 (N_8222,N_4620,N_707);
nor U8223 (N_8223,N_3657,N_290);
nor U8224 (N_8224,N_4817,N_650);
and U8225 (N_8225,N_4198,N_2152);
nor U8226 (N_8226,N_3779,N_3891);
or U8227 (N_8227,N_4482,N_3548);
and U8228 (N_8228,N_755,N_3173);
or U8229 (N_8229,N_832,N_1078);
or U8230 (N_8230,N_1962,N_4182);
or U8231 (N_8231,N_4779,N_790);
nand U8232 (N_8232,N_1831,N_686);
nand U8233 (N_8233,N_1455,N_3650);
xnor U8234 (N_8234,N_4986,N_587);
or U8235 (N_8235,N_3522,N_763);
and U8236 (N_8236,N_4444,N_2221);
or U8237 (N_8237,N_358,N_3759);
or U8238 (N_8238,N_166,N_2443);
and U8239 (N_8239,N_4979,N_2854);
and U8240 (N_8240,N_4651,N_2576);
or U8241 (N_8241,N_2375,N_1879);
nand U8242 (N_8242,N_3445,N_2394);
xor U8243 (N_8243,N_4503,N_128);
nand U8244 (N_8244,N_1844,N_3057);
nand U8245 (N_8245,N_1820,N_3326);
nor U8246 (N_8246,N_954,N_1307);
or U8247 (N_8247,N_2724,N_3071);
xnor U8248 (N_8248,N_3653,N_1507);
xnor U8249 (N_8249,N_669,N_3196);
nor U8250 (N_8250,N_3585,N_1376);
xnor U8251 (N_8251,N_2307,N_4021);
or U8252 (N_8252,N_3341,N_3551);
nand U8253 (N_8253,N_1723,N_2090);
or U8254 (N_8254,N_4534,N_3137);
nand U8255 (N_8255,N_2263,N_1034);
nand U8256 (N_8256,N_307,N_1011);
and U8257 (N_8257,N_3157,N_4276);
or U8258 (N_8258,N_3585,N_1968);
xor U8259 (N_8259,N_4488,N_268);
xnor U8260 (N_8260,N_3381,N_4571);
xnor U8261 (N_8261,N_2491,N_3225);
nor U8262 (N_8262,N_4152,N_687);
xor U8263 (N_8263,N_2369,N_4861);
xor U8264 (N_8264,N_4921,N_3947);
nand U8265 (N_8265,N_2255,N_4733);
nand U8266 (N_8266,N_322,N_2460);
or U8267 (N_8267,N_392,N_4768);
xnor U8268 (N_8268,N_2275,N_2483);
xnor U8269 (N_8269,N_1441,N_1693);
xor U8270 (N_8270,N_828,N_3696);
or U8271 (N_8271,N_4327,N_2273);
nand U8272 (N_8272,N_3497,N_4818);
and U8273 (N_8273,N_1929,N_1338);
nor U8274 (N_8274,N_1320,N_2528);
xnor U8275 (N_8275,N_1073,N_2302);
xor U8276 (N_8276,N_390,N_2469);
or U8277 (N_8277,N_4667,N_1193);
and U8278 (N_8278,N_3673,N_4780);
and U8279 (N_8279,N_1381,N_3724);
or U8280 (N_8280,N_1919,N_3659);
and U8281 (N_8281,N_2744,N_1237);
xor U8282 (N_8282,N_2662,N_389);
nand U8283 (N_8283,N_2294,N_2174);
nor U8284 (N_8284,N_4213,N_1435);
or U8285 (N_8285,N_191,N_396);
nor U8286 (N_8286,N_4920,N_4704);
nor U8287 (N_8287,N_2586,N_1686);
nand U8288 (N_8288,N_4449,N_3616);
nand U8289 (N_8289,N_1327,N_3282);
and U8290 (N_8290,N_3041,N_2955);
nor U8291 (N_8291,N_650,N_3782);
xor U8292 (N_8292,N_2053,N_4815);
or U8293 (N_8293,N_2526,N_2416);
nor U8294 (N_8294,N_2221,N_2418);
xor U8295 (N_8295,N_505,N_2442);
and U8296 (N_8296,N_2019,N_442);
and U8297 (N_8297,N_743,N_296);
and U8298 (N_8298,N_3517,N_1316);
or U8299 (N_8299,N_2272,N_644);
nor U8300 (N_8300,N_4978,N_1118);
xor U8301 (N_8301,N_4638,N_902);
or U8302 (N_8302,N_4297,N_2986);
nand U8303 (N_8303,N_11,N_2536);
nor U8304 (N_8304,N_4752,N_30);
and U8305 (N_8305,N_3381,N_1470);
xnor U8306 (N_8306,N_3969,N_1990);
nor U8307 (N_8307,N_900,N_2541);
or U8308 (N_8308,N_454,N_3625);
or U8309 (N_8309,N_1662,N_442);
and U8310 (N_8310,N_770,N_798);
xor U8311 (N_8311,N_3623,N_1122);
nor U8312 (N_8312,N_647,N_3061);
nand U8313 (N_8313,N_1732,N_1561);
and U8314 (N_8314,N_216,N_3208);
xor U8315 (N_8315,N_264,N_4513);
or U8316 (N_8316,N_4928,N_3862);
nand U8317 (N_8317,N_3596,N_127);
or U8318 (N_8318,N_3266,N_677);
nor U8319 (N_8319,N_4447,N_2680);
or U8320 (N_8320,N_147,N_1025);
nor U8321 (N_8321,N_15,N_501);
or U8322 (N_8322,N_995,N_1647);
or U8323 (N_8323,N_3470,N_348);
nor U8324 (N_8324,N_3397,N_2003);
xor U8325 (N_8325,N_3978,N_502);
and U8326 (N_8326,N_1438,N_4116);
or U8327 (N_8327,N_3831,N_786);
and U8328 (N_8328,N_3719,N_1749);
nand U8329 (N_8329,N_3637,N_1545);
nand U8330 (N_8330,N_633,N_3840);
nor U8331 (N_8331,N_2730,N_691);
or U8332 (N_8332,N_4119,N_3969);
nor U8333 (N_8333,N_4364,N_1473);
nor U8334 (N_8334,N_2648,N_848);
and U8335 (N_8335,N_774,N_176);
nor U8336 (N_8336,N_2656,N_3759);
nor U8337 (N_8337,N_1197,N_2958);
or U8338 (N_8338,N_207,N_1192);
xor U8339 (N_8339,N_2666,N_2946);
nor U8340 (N_8340,N_3241,N_1263);
nand U8341 (N_8341,N_1777,N_1096);
and U8342 (N_8342,N_1797,N_1608);
xnor U8343 (N_8343,N_3488,N_1406);
nand U8344 (N_8344,N_1897,N_1109);
and U8345 (N_8345,N_1952,N_43);
or U8346 (N_8346,N_3333,N_2139);
nand U8347 (N_8347,N_4523,N_3780);
xnor U8348 (N_8348,N_1971,N_1935);
nand U8349 (N_8349,N_3569,N_2718);
and U8350 (N_8350,N_3683,N_2666);
nand U8351 (N_8351,N_1239,N_982);
xnor U8352 (N_8352,N_1826,N_1860);
nor U8353 (N_8353,N_2380,N_764);
or U8354 (N_8354,N_2402,N_2298);
or U8355 (N_8355,N_2115,N_4359);
xnor U8356 (N_8356,N_1820,N_2207);
nor U8357 (N_8357,N_181,N_3807);
or U8358 (N_8358,N_1292,N_4531);
nand U8359 (N_8359,N_490,N_2589);
nand U8360 (N_8360,N_4027,N_4352);
or U8361 (N_8361,N_2082,N_1582);
nand U8362 (N_8362,N_3182,N_4505);
nor U8363 (N_8363,N_1274,N_3263);
xor U8364 (N_8364,N_378,N_99);
nand U8365 (N_8365,N_4260,N_506);
nand U8366 (N_8366,N_2891,N_4789);
or U8367 (N_8367,N_1630,N_2934);
or U8368 (N_8368,N_4362,N_4850);
and U8369 (N_8369,N_790,N_35);
nand U8370 (N_8370,N_4591,N_301);
nor U8371 (N_8371,N_3402,N_4876);
xnor U8372 (N_8372,N_689,N_4623);
nand U8373 (N_8373,N_4317,N_2022);
xor U8374 (N_8374,N_9,N_836);
xor U8375 (N_8375,N_4245,N_3632);
nor U8376 (N_8376,N_342,N_4931);
xor U8377 (N_8377,N_3129,N_4503);
nor U8378 (N_8378,N_2471,N_2307);
nand U8379 (N_8379,N_4950,N_3629);
nand U8380 (N_8380,N_3966,N_2190);
and U8381 (N_8381,N_2275,N_2716);
or U8382 (N_8382,N_3133,N_2952);
and U8383 (N_8383,N_69,N_1382);
nand U8384 (N_8384,N_4139,N_4009);
or U8385 (N_8385,N_710,N_4589);
nor U8386 (N_8386,N_3979,N_4938);
nor U8387 (N_8387,N_3101,N_4116);
nand U8388 (N_8388,N_738,N_4504);
and U8389 (N_8389,N_456,N_1602);
and U8390 (N_8390,N_338,N_689);
xor U8391 (N_8391,N_4310,N_1177);
nor U8392 (N_8392,N_1094,N_2483);
or U8393 (N_8393,N_1878,N_1982);
nand U8394 (N_8394,N_773,N_1231);
nand U8395 (N_8395,N_505,N_861);
or U8396 (N_8396,N_4238,N_2170);
nor U8397 (N_8397,N_3556,N_4461);
and U8398 (N_8398,N_3762,N_993);
and U8399 (N_8399,N_2068,N_4084);
nand U8400 (N_8400,N_4760,N_294);
xnor U8401 (N_8401,N_1869,N_1162);
and U8402 (N_8402,N_132,N_989);
and U8403 (N_8403,N_1181,N_4651);
nand U8404 (N_8404,N_2658,N_1289);
nor U8405 (N_8405,N_33,N_125);
or U8406 (N_8406,N_329,N_2840);
or U8407 (N_8407,N_2678,N_4653);
or U8408 (N_8408,N_1949,N_2856);
and U8409 (N_8409,N_2402,N_1744);
nor U8410 (N_8410,N_3035,N_4769);
nand U8411 (N_8411,N_4067,N_936);
xor U8412 (N_8412,N_2165,N_4702);
xnor U8413 (N_8413,N_852,N_480);
or U8414 (N_8414,N_1517,N_4780);
nand U8415 (N_8415,N_4173,N_2770);
and U8416 (N_8416,N_662,N_400);
xor U8417 (N_8417,N_3448,N_3496);
or U8418 (N_8418,N_3525,N_1741);
or U8419 (N_8419,N_715,N_1640);
or U8420 (N_8420,N_2501,N_1325);
and U8421 (N_8421,N_2585,N_2798);
nor U8422 (N_8422,N_2300,N_4140);
and U8423 (N_8423,N_4242,N_3488);
and U8424 (N_8424,N_1966,N_4843);
nor U8425 (N_8425,N_3171,N_1647);
nand U8426 (N_8426,N_1953,N_2353);
or U8427 (N_8427,N_1032,N_4753);
nor U8428 (N_8428,N_2131,N_3945);
xor U8429 (N_8429,N_2828,N_4645);
and U8430 (N_8430,N_3505,N_18);
nor U8431 (N_8431,N_2983,N_4068);
and U8432 (N_8432,N_1505,N_927);
and U8433 (N_8433,N_1732,N_1554);
nand U8434 (N_8434,N_1457,N_264);
and U8435 (N_8435,N_1444,N_4579);
or U8436 (N_8436,N_414,N_3592);
nor U8437 (N_8437,N_4495,N_3056);
xor U8438 (N_8438,N_1271,N_2922);
or U8439 (N_8439,N_2957,N_4996);
nand U8440 (N_8440,N_4103,N_1991);
and U8441 (N_8441,N_1674,N_4503);
or U8442 (N_8442,N_4258,N_1994);
nor U8443 (N_8443,N_2988,N_474);
and U8444 (N_8444,N_2913,N_4069);
or U8445 (N_8445,N_396,N_4546);
and U8446 (N_8446,N_933,N_5);
nand U8447 (N_8447,N_4523,N_1721);
and U8448 (N_8448,N_2014,N_2611);
or U8449 (N_8449,N_3421,N_1734);
and U8450 (N_8450,N_2705,N_1669);
or U8451 (N_8451,N_76,N_1110);
nand U8452 (N_8452,N_2539,N_1043);
nand U8453 (N_8453,N_3957,N_2292);
nor U8454 (N_8454,N_1285,N_2161);
or U8455 (N_8455,N_1648,N_4545);
nor U8456 (N_8456,N_557,N_3759);
or U8457 (N_8457,N_3904,N_3992);
nand U8458 (N_8458,N_1970,N_4461);
nor U8459 (N_8459,N_1935,N_351);
nor U8460 (N_8460,N_4104,N_2253);
or U8461 (N_8461,N_1410,N_3450);
xor U8462 (N_8462,N_3980,N_150);
nor U8463 (N_8463,N_1665,N_1006);
xnor U8464 (N_8464,N_321,N_2758);
or U8465 (N_8465,N_2018,N_4550);
nor U8466 (N_8466,N_4363,N_839);
and U8467 (N_8467,N_2949,N_3738);
nand U8468 (N_8468,N_3492,N_3532);
xor U8469 (N_8469,N_3616,N_2164);
nor U8470 (N_8470,N_4382,N_4438);
xnor U8471 (N_8471,N_1774,N_4469);
xnor U8472 (N_8472,N_215,N_4895);
or U8473 (N_8473,N_3296,N_3165);
or U8474 (N_8474,N_587,N_633);
nor U8475 (N_8475,N_2458,N_22);
nand U8476 (N_8476,N_25,N_3566);
nor U8477 (N_8477,N_4171,N_1294);
and U8478 (N_8478,N_2420,N_3599);
or U8479 (N_8479,N_1102,N_4358);
and U8480 (N_8480,N_976,N_2946);
or U8481 (N_8481,N_1932,N_1701);
nand U8482 (N_8482,N_3098,N_77);
or U8483 (N_8483,N_609,N_498);
or U8484 (N_8484,N_4400,N_4965);
nor U8485 (N_8485,N_2533,N_4099);
nand U8486 (N_8486,N_2833,N_2066);
nand U8487 (N_8487,N_3411,N_2198);
nor U8488 (N_8488,N_872,N_1283);
and U8489 (N_8489,N_2087,N_2328);
nor U8490 (N_8490,N_2615,N_3160);
nand U8491 (N_8491,N_1670,N_368);
xor U8492 (N_8492,N_3867,N_4522);
nor U8493 (N_8493,N_3823,N_2104);
and U8494 (N_8494,N_2909,N_4377);
nor U8495 (N_8495,N_3677,N_3158);
nand U8496 (N_8496,N_3196,N_39);
nand U8497 (N_8497,N_3569,N_464);
xor U8498 (N_8498,N_374,N_1119);
nand U8499 (N_8499,N_1433,N_2810);
xor U8500 (N_8500,N_2815,N_2157);
xnor U8501 (N_8501,N_708,N_4434);
nor U8502 (N_8502,N_888,N_537);
nor U8503 (N_8503,N_4795,N_2179);
nor U8504 (N_8504,N_655,N_1400);
or U8505 (N_8505,N_1840,N_2487);
or U8506 (N_8506,N_606,N_4006);
nor U8507 (N_8507,N_4522,N_1757);
nand U8508 (N_8508,N_2732,N_2727);
or U8509 (N_8509,N_3304,N_1520);
nor U8510 (N_8510,N_2971,N_3349);
nor U8511 (N_8511,N_1143,N_3361);
xnor U8512 (N_8512,N_465,N_3723);
or U8513 (N_8513,N_3106,N_729);
nand U8514 (N_8514,N_4636,N_1455);
or U8515 (N_8515,N_4179,N_3319);
nor U8516 (N_8516,N_733,N_3072);
xnor U8517 (N_8517,N_1629,N_2349);
nand U8518 (N_8518,N_879,N_1836);
nand U8519 (N_8519,N_2499,N_2978);
nand U8520 (N_8520,N_3883,N_2570);
or U8521 (N_8521,N_2810,N_1075);
or U8522 (N_8522,N_2901,N_4903);
or U8523 (N_8523,N_2802,N_1472);
nor U8524 (N_8524,N_4096,N_1880);
nor U8525 (N_8525,N_4306,N_627);
nand U8526 (N_8526,N_1095,N_2471);
and U8527 (N_8527,N_1151,N_286);
xor U8528 (N_8528,N_3570,N_3671);
or U8529 (N_8529,N_3252,N_696);
or U8530 (N_8530,N_3366,N_100);
or U8531 (N_8531,N_3487,N_4550);
and U8532 (N_8532,N_3548,N_3905);
and U8533 (N_8533,N_3518,N_1412);
or U8534 (N_8534,N_721,N_1945);
and U8535 (N_8535,N_1535,N_3534);
or U8536 (N_8536,N_365,N_970);
and U8537 (N_8537,N_2684,N_3868);
nand U8538 (N_8538,N_2941,N_2807);
nor U8539 (N_8539,N_3697,N_115);
nand U8540 (N_8540,N_1705,N_3442);
nand U8541 (N_8541,N_3582,N_865);
nand U8542 (N_8542,N_854,N_3049);
nand U8543 (N_8543,N_3640,N_2333);
or U8544 (N_8544,N_4035,N_1484);
nand U8545 (N_8545,N_4217,N_1952);
nor U8546 (N_8546,N_3755,N_3224);
or U8547 (N_8547,N_855,N_3604);
xnor U8548 (N_8548,N_1489,N_3279);
nor U8549 (N_8549,N_3552,N_3443);
or U8550 (N_8550,N_3123,N_779);
or U8551 (N_8551,N_3619,N_1137);
xor U8552 (N_8552,N_2072,N_3276);
or U8553 (N_8553,N_2982,N_4262);
nand U8554 (N_8554,N_518,N_575);
nand U8555 (N_8555,N_2894,N_4171);
or U8556 (N_8556,N_1143,N_4605);
nor U8557 (N_8557,N_4820,N_1514);
xnor U8558 (N_8558,N_2899,N_2665);
nor U8559 (N_8559,N_3074,N_4);
nor U8560 (N_8560,N_1961,N_71);
and U8561 (N_8561,N_2566,N_771);
xor U8562 (N_8562,N_1959,N_2839);
or U8563 (N_8563,N_2147,N_1552);
and U8564 (N_8564,N_147,N_2996);
or U8565 (N_8565,N_4861,N_4541);
nor U8566 (N_8566,N_1698,N_1708);
nand U8567 (N_8567,N_701,N_1288);
or U8568 (N_8568,N_1425,N_1840);
and U8569 (N_8569,N_1278,N_3710);
xor U8570 (N_8570,N_4469,N_465);
nand U8571 (N_8571,N_4491,N_52);
xor U8572 (N_8572,N_240,N_4742);
nand U8573 (N_8573,N_684,N_2987);
or U8574 (N_8574,N_684,N_4685);
nor U8575 (N_8575,N_1519,N_1697);
nor U8576 (N_8576,N_3606,N_1172);
xor U8577 (N_8577,N_3699,N_4868);
or U8578 (N_8578,N_4388,N_1679);
and U8579 (N_8579,N_1115,N_2668);
xor U8580 (N_8580,N_707,N_317);
and U8581 (N_8581,N_4071,N_1504);
xnor U8582 (N_8582,N_4473,N_515);
nor U8583 (N_8583,N_664,N_3500);
xnor U8584 (N_8584,N_2258,N_808);
or U8585 (N_8585,N_3820,N_634);
nand U8586 (N_8586,N_3335,N_4754);
xnor U8587 (N_8587,N_4441,N_1016);
and U8588 (N_8588,N_275,N_790);
xnor U8589 (N_8589,N_3275,N_114);
and U8590 (N_8590,N_614,N_3918);
xnor U8591 (N_8591,N_1391,N_4549);
nand U8592 (N_8592,N_4744,N_977);
nor U8593 (N_8593,N_2999,N_615);
and U8594 (N_8594,N_1620,N_2940);
nor U8595 (N_8595,N_80,N_2831);
xnor U8596 (N_8596,N_4907,N_3726);
xor U8597 (N_8597,N_3631,N_3203);
or U8598 (N_8598,N_778,N_3360);
nand U8599 (N_8599,N_4424,N_2746);
and U8600 (N_8600,N_4107,N_2215);
nand U8601 (N_8601,N_3259,N_1620);
or U8602 (N_8602,N_3983,N_4702);
nor U8603 (N_8603,N_771,N_4810);
and U8604 (N_8604,N_4316,N_2492);
xnor U8605 (N_8605,N_544,N_138);
nand U8606 (N_8606,N_3709,N_4972);
or U8607 (N_8607,N_3576,N_2243);
nand U8608 (N_8608,N_749,N_2002);
and U8609 (N_8609,N_2916,N_1522);
xnor U8610 (N_8610,N_420,N_2163);
nand U8611 (N_8611,N_198,N_796);
nor U8612 (N_8612,N_3624,N_2372);
nor U8613 (N_8613,N_880,N_1005);
nor U8614 (N_8614,N_1387,N_337);
nand U8615 (N_8615,N_1799,N_1198);
nor U8616 (N_8616,N_4350,N_2604);
nor U8617 (N_8617,N_4089,N_976);
nor U8618 (N_8618,N_1635,N_829);
and U8619 (N_8619,N_4879,N_2861);
nor U8620 (N_8620,N_712,N_3009);
xor U8621 (N_8621,N_200,N_2474);
or U8622 (N_8622,N_689,N_1325);
xor U8623 (N_8623,N_4984,N_749);
xor U8624 (N_8624,N_429,N_188);
xnor U8625 (N_8625,N_1446,N_2223);
nand U8626 (N_8626,N_4453,N_1838);
nand U8627 (N_8627,N_2148,N_90);
and U8628 (N_8628,N_2264,N_386);
nor U8629 (N_8629,N_1136,N_3691);
nand U8630 (N_8630,N_3652,N_4772);
nor U8631 (N_8631,N_3054,N_2330);
and U8632 (N_8632,N_3563,N_63);
xor U8633 (N_8633,N_4644,N_8);
xnor U8634 (N_8634,N_2168,N_2367);
and U8635 (N_8635,N_295,N_100);
or U8636 (N_8636,N_4109,N_359);
and U8637 (N_8637,N_2831,N_1556);
xor U8638 (N_8638,N_3121,N_1199);
nand U8639 (N_8639,N_1317,N_1523);
nor U8640 (N_8640,N_2957,N_4517);
nor U8641 (N_8641,N_4435,N_1684);
nor U8642 (N_8642,N_2967,N_2002);
xnor U8643 (N_8643,N_2020,N_1222);
or U8644 (N_8644,N_4057,N_1708);
or U8645 (N_8645,N_4810,N_3546);
nor U8646 (N_8646,N_2769,N_1532);
or U8647 (N_8647,N_1889,N_2942);
xor U8648 (N_8648,N_826,N_2797);
xor U8649 (N_8649,N_3766,N_2938);
xor U8650 (N_8650,N_3308,N_3430);
and U8651 (N_8651,N_263,N_3718);
and U8652 (N_8652,N_21,N_1459);
and U8653 (N_8653,N_4330,N_184);
and U8654 (N_8654,N_4014,N_2921);
nand U8655 (N_8655,N_4053,N_4309);
nor U8656 (N_8656,N_2357,N_3567);
xor U8657 (N_8657,N_993,N_583);
nand U8658 (N_8658,N_4510,N_1840);
xnor U8659 (N_8659,N_2177,N_1194);
nor U8660 (N_8660,N_3885,N_4304);
nor U8661 (N_8661,N_2301,N_1231);
and U8662 (N_8662,N_3007,N_3304);
nor U8663 (N_8663,N_1968,N_1359);
and U8664 (N_8664,N_2687,N_3284);
or U8665 (N_8665,N_3546,N_3008);
and U8666 (N_8666,N_3021,N_2414);
nor U8667 (N_8667,N_2410,N_3204);
nand U8668 (N_8668,N_4021,N_4688);
nand U8669 (N_8669,N_4368,N_2420);
xnor U8670 (N_8670,N_4490,N_2188);
nor U8671 (N_8671,N_3231,N_3009);
and U8672 (N_8672,N_4372,N_4244);
nor U8673 (N_8673,N_3196,N_2592);
nor U8674 (N_8674,N_4701,N_4017);
xor U8675 (N_8675,N_2316,N_100);
and U8676 (N_8676,N_3492,N_3486);
or U8677 (N_8677,N_4857,N_1756);
or U8678 (N_8678,N_2873,N_646);
xnor U8679 (N_8679,N_2727,N_266);
xnor U8680 (N_8680,N_2794,N_3296);
nand U8681 (N_8681,N_806,N_1642);
or U8682 (N_8682,N_3625,N_3260);
and U8683 (N_8683,N_345,N_599);
xor U8684 (N_8684,N_96,N_2333);
xnor U8685 (N_8685,N_1750,N_501);
nor U8686 (N_8686,N_1652,N_24);
and U8687 (N_8687,N_1598,N_139);
xnor U8688 (N_8688,N_379,N_851);
or U8689 (N_8689,N_161,N_1033);
xor U8690 (N_8690,N_979,N_4874);
nand U8691 (N_8691,N_1292,N_4536);
nor U8692 (N_8692,N_4613,N_261);
xnor U8693 (N_8693,N_3171,N_2431);
nor U8694 (N_8694,N_2110,N_21);
and U8695 (N_8695,N_4091,N_4481);
or U8696 (N_8696,N_3418,N_3512);
xor U8697 (N_8697,N_759,N_3007);
nor U8698 (N_8698,N_2814,N_3020);
or U8699 (N_8699,N_1721,N_3002);
xnor U8700 (N_8700,N_4716,N_1582);
and U8701 (N_8701,N_2336,N_2212);
or U8702 (N_8702,N_2643,N_358);
or U8703 (N_8703,N_1914,N_1357);
xor U8704 (N_8704,N_4244,N_4633);
or U8705 (N_8705,N_4452,N_1679);
nand U8706 (N_8706,N_3000,N_2197);
xor U8707 (N_8707,N_1985,N_3590);
nor U8708 (N_8708,N_4745,N_1310);
nand U8709 (N_8709,N_1358,N_1228);
and U8710 (N_8710,N_2644,N_480);
and U8711 (N_8711,N_902,N_1685);
nand U8712 (N_8712,N_155,N_4622);
nor U8713 (N_8713,N_3601,N_1767);
nand U8714 (N_8714,N_191,N_1820);
nand U8715 (N_8715,N_4090,N_3752);
or U8716 (N_8716,N_3460,N_2243);
and U8717 (N_8717,N_2154,N_2930);
nor U8718 (N_8718,N_4427,N_1490);
xor U8719 (N_8719,N_4388,N_3964);
and U8720 (N_8720,N_3826,N_89);
nand U8721 (N_8721,N_4178,N_117);
xor U8722 (N_8722,N_70,N_4120);
and U8723 (N_8723,N_2072,N_3003);
xor U8724 (N_8724,N_3407,N_3740);
and U8725 (N_8725,N_2700,N_3965);
or U8726 (N_8726,N_4814,N_2849);
or U8727 (N_8727,N_93,N_1994);
or U8728 (N_8728,N_2015,N_293);
and U8729 (N_8729,N_1095,N_3102);
and U8730 (N_8730,N_4363,N_2323);
nand U8731 (N_8731,N_2554,N_2234);
or U8732 (N_8732,N_2839,N_2467);
and U8733 (N_8733,N_2183,N_3159);
or U8734 (N_8734,N_447,N_2716);
nor U8735 (N_8735,N_3261,N_1718);
xor U8736 (N_8736,N_3782,N_817);
and U8737 (N_8737,N_572,N_3612);
xor U8738 (N_8738,N_1217,N_436);
nand U8739 (N_8739,N_4216,N_1676);
xor U8740 (N_8740,N_4004,N_3981);
nor U8741 (N_8741,N_4651,N_1449);
nand U8742 (N_8742,N_864,N_3269);
nor U8743 (N_8743,N_4253,N_1449);
nor U8744 (N_8744,N_3774,N_3418);
and U8745 (N_8745,N_1480,N_2520);
and U8746 (N_8746,N_2445,N_4486);
or U8747 (N_8747,N_4464,N_925);
nor U8748 (N_8748,N_1450,N_4979);
or U8749 (N_8749,N_1190,N_95);
nand U8750 (N_8750,N_285,N_2752);
nand U8751 (N_8751,N_3602,N_2237);
xor U8752 (N_8752,N_3162,N_632);
or U8753 (N_8753,N_3649,N_2042);
nand U8754 (N_8754,N_817,N_1353);
nor U8755 (N_8755,N_654,N_2804);
xnor U8756 (N_8756,N_1897,N_1753);
nor U8757 (N_8757,N_2191,N_1534);
nor U8758 (N_8758,N_43,N_4963);
and U8759 (N_8759,N_4032,N_3891);
nand U8760 (N_8760,N_1912,N_4538);
nor U8761 (N_8761,N_1252,N_3128);
xnor U8762 (N_8762,N_4237,N_3333);
or U8763 (N_8763,N_1769,N_1762);
nor U8764 (N_8764,N_1292,N_366);
and U8765 (N_8765,N_1291,N_1474);
nor U8766 (N_8766,N_564,N_2079);
xnor U8767 (N_8767,N_3009,N_3767);
or U8768 (N_8768,N_2807,N_3487);
nand U8769 (N_8769,N_4161,N_204);
nand U8770 (N_8770,N_644,N_1326);
and U8771 (N_8771,N_4929,N_1312);
or U8772 (N_8772,N_2981,N_2569);
xor U8773 (N_8773,N_4015,N_3177);
and U8774 (N_8774,N_2393,N_346);
and U8775 (N_8775,N_4803,N_2467);
or U8776 (N_8776,N_2858,N_3745);
nand U8777 (N_8777,N_1077,N_3990);
and U8778 (N_8778,N_95,N_2330);
nand U8779 (N_8779,N_2854,N_670);
nor U8780 (N_8780,N_736,N_2461);
nor U8781 (N_8781,N_2154,N_1377);
xor U8782 (N_8782,N_4654,N_1654);
or U8783 (N_8783,N_2731,N_4116);
nor U8784 (N_8784,N_949,N_3310);
nor U8785 (N_8785,N_262,N_1270);
nor U8786 (N_8786,N_3775,N_3969);
and U8787 (N_8787,N_2208,N_338);
or U8788 (N_8788,N_3074,N_3844);
xor U8789 (N_8789,N_4891,N_3402);
xor U8790 (N_8790,N_4415,N_1579);
and U8791 (N_8791,N_2334,N_4196);
and U8792 (N_8792,N_3298,N_4954);
nand U8793 (N_8793,N_1254,N_174);
nand U8794 (N_8794,N_3934,N_946);
nand U8795 (N_8795,N_3432,N_4040);
or U8796 (N_8796,N_1635,N_1034);
and U8797 (N_8797,N_4315,N_4119);
or U8798 (N_8798,N_3104,N_2752);
nor U8799 (N_8799,N_3587,N_1812);
and U8800 (N_8800,N_3614,N_3882);
or U8801 (N_8801,N_998,N_2895);
and U8802 (N_8802,N_745,N_4307);
or U8803 (N_8803,N_769,N_3109);
and U8804 (N_8804,N_3492,N_1375);
and U8805 (N_8805,N_3416,N_2864);
nor U8806 (N_8806,N_3444,N_4520);
nor U8807 (N_8807,N_3028,N_690);
xnor U8808 (N_8808,N_2753,N_1214);
xnor U8809 (N_8809,N_2409,N_913);
nand U8810 (N_8810,N_323,N_2500);
xnor U8811 (N_8811,N_2681,N_2549);
and U8812 (N_8812,N_1065,N_1463);
and U8813 (N_8813,N_3578,N_4298);
nor U8814 (N_8814,N_2602,N_2960);
xnor U8815 (N_8815,N_3735,N_3912);
xor U8816 (N_8816,N_789,N_4364);
or U8817 (N_8817,N_3543,N_4790);
or U8818 (N_8818,N_4058,N_2143);
nor U8819 (N_8819,N_4682,N_3110);
and U8820 (N_8820,N_3228,N_2018);
nor U8821 (N_8821,N_513,N_2198);
or U8822 (N_8822,N_1262,N_4129);
or U8823 (N_8823,N_1690,N_3929);
or U8824 (N_8824,N_942,N_2709);
nor U8825 (N_8825,N_686,N_2820);
and U8826 (N_8826,N_3614,N_3056);
xor U8827 (N_8827,N_1925,N_3886);
or U8828 (N_8828,N_4264,N_3269);
xnor U8829 (N_8829,N_2760,N_4961);
xor U8830 (N_8830,N_775,N_1343);
xor U8831 (N_8831,N_1887,N_1483);
nand U8832 (N_8832,N_4384,N_3779);
or U8833 (N_8833,N_3452,N_720);
or U8834 (N_8834,N_715,N_1975);
and U8835 (N_8835,N_3164,N_4796);
nor U8836 (N_8836,N_3230,N_2832);
and U8837 (N_8837,N_327,N_2956);
nand U8838 (N_8838,N_4806,N_344);
xnor U8839 (N_8839,N_3596,N_3734);
nand U8840 (N_8840,N_2589,N_2839);
nand U8841 (N_8841,N_2694,N_1728);
and U8842 (N_8842,N_3319,N_4609);
or U8843 (N_8843,N_2545,N_4517);
nor U8844 (N_8844,N_2274,N_715);
nand U8845 (N_8845,N_1272,N_4990);
xor U8846 (N_8846,N_1527,N_3143);
or U8847 (N_8847,N_2547,N_625);
or U8848 (N_8848,N_3500,N_3057);
nor U8849 (N_8849,N_158,N_3971);
and U8850 (N_8850,N_3755,N_2056);
nand U8851 (N_8851,N_3870,N_507);
nand U8852 (N_8852,N_816,N_1516);
or U8853 (N_8853,N_3836,N_1410);
and U8854 (N_8854,N_2689,N_3821);
xnor U8855 (N_8855,N_4201,N_4657);
or U8856 (N_8856,N_4182,N_2071);
and U8857 (N_8857,N_2941,N_2637);
xnor U8858 (N_8858,N_4376,N_769);
and U8859 (N_8859,N_4849,N_3508);
or U8860 (N_8860,N_2256,N_4490);
nand U8861 (N_8861,N_2096,N_2434);
and U8862 (N_8862,N_3782,N_1046);
and U8863 (N_8863,N_4559,N_4588);
xnor U8864 (N_8864,N_2868,N_425);
nand U8865 (N_8865,N_3673,N_1641);
and U8866 (N_8866,N_1879,N_272);
nor U8867 (N_8867,N_69,N_1022);
or U8868 (N_8868,N_3870,N_4251);
and U8869 (N_8869,N_1885,N_3617);
nand U8870 (N_8870,N_2801,N_891);
nand U8871 (N_8871,N_1034,N_3063);
and U8872 (N_8872,N_4356,N_1938);
and U8873 (N_8873,N_3902,N_2441);
xnor U8874 (N_8874,N_1039,N_4110);
nor U8875 (N_8875,N_3851,N_529);
and U8876 (N_8876,N_3921,N_2488);
and U8877 (N_8877,N_4982,N_3365);
nand U8878 (N_8878,N_1882,N_246);
and U8879 (N_8879,N_3176,N_4532);
nand U8880 (N_8880,N_4102,N_473);
or U8881 (N_8881,N_4465,N_2835);
or U8882 (N_8882,N_567,N_1748);
nor U8883 (N_8883,N_4916,N_136);
nor U8884 (N_8884,N_1849,N_4765);
or U8885 (N_8885,N_2286,N_2);
or U8886 (N_8886,N_1592,N_1011);
and U8887 (N_8887,N_2450,N_4927);
or U8888 (N_8888,N_888,N_2821);
xnor U8889 (N_8889,N_3471,N_2186);
and U8890 (N_8890,N_2315,N_23);
xnor U8891 (N_8891,N_4981,N_4368);
and U8892 (N_8892,N_3338,N_4434);
and U8893 (N_8893,N_2949,N_2314);
xor U8894 (N_8894,N_191,N_4230);
nand U8895 (N_8895,N_3042,N_4431);
nand U8896 (N_8896,N_2961,N_698);
xnor U8897 (N_8897,N_808,N_2546);
and U8898 (N_8898,N_4283,N_3719);
or U8899 (N_8899,N_2408,N_256);
nand U8900 (N_8900,N_3341,N_774);
or U8901 (N_8901,N_1521,N_3805);
or U8902 (N_8902,N_4523,N_592);
and U8903 (N_8903,N_1051,N_3567);
nand U8904 (N_8904,N_3126,N_504);
nand U8905 (N_8905,N_1666,N_2381);
or U8906 (N_8906,N_2231,N_4236);
nand U8907 (N_8907,N_3546,N_2364);
and U8908 (N_8908,N_0,N_2309);
xnor U8909 (N_8909,N_1245,N_1428);
or U8910 (N_8910,N_1415,N_31);
or U8911 (N_8911,N_3240,N_3919);
nand U8912 (N_8912,N_503,N_4627);
or U8913 (N_8913,N_2822,N_779);
xnor U8914 (N_8914,N_1548,N_221);
nand U8915 (N_8915,N_4348,N_4223);
nand U8916 (N_8916,N_4815,N_304);
nand U8917 (N_8917,N_1668,N_699);
and U8918 (N_8918,N_4874,N_3987);
nor U8919 (N_8919,N_1573,N_674);
and U8920 (N_8920,N_3438,N_3306);
xnor U8921 (N_8921,N_3163,N_2292);
xnor U8922 (N_8922,N_4029,N_4429);
or U8923 (N_8923,N_2871,N_4139);
nand U8924 (N_8924,N_2475,N_766);
or U8925 (N_8925,N_4730,N_3676);
or U8926 (N_8926,N_3797,N_4120);
nor U8927 (N_8927,N_4239,N_107);
and U8928 (N_8928,N_2852,N_1645);
nand U8929 (N_8929,N_872,N_4012);
or U8930 (N_8930,N_4494,N_4483);
or U8931 (N_8931,N_4050,N_1836);
nand U8932 (N_8932,N_904,N_746);
and U8933 (N_8933,N_1023,N_4590);
nand U8934 (N_8934,N_2532,N_2823);
or U8935 (N_8935,N_2711,N_211);
nor U8936 (N_8936,N_4568,N_2055);
nor U8937 (N_8937,N_4334,N_4688);
nor U8938 (N_8938,N_2820,N_3839);
and U8939 (N_8939,N_4328,N_4571);
and U8940 (N_8940,N_4820,N_4606);
or U8941 (N_8941,N_827,N_3384);
and U8942 (N_8942,N_4203,N_1485);
nand U8943 (N_8943,N_3671,N_1308);
and U8944 (N_8944,N_3631,N_301);
nand U8945 (N_8945,N_2440,N_3267);
nor U8946 (N_8946,N_3648,N_4370);
nor U8947 (N_8947,N_2133,N_3142);
nor U8948 (N_8948,N_1382,N_440);
or U8949 (N_8949,N_4310,N_2813);
xnor U8950 (N_8950,N_1049,N_2441);
or U8951 (N_8951,N_2259,N_3414);
nand U8952 (N_8952,N_3770,N_2942);
nand U8953 (N_8953,N_4805,N_4581);
or U8954 (N_8954,N_267,N_1851);
nor U8955 (N_8955,N_1127,N_3280);
nor U8956 (N_8956,N_1890,N_3562);
nor U8957 (N_8957,N_4309,N_67);
and U8958 (N_8958,N_4273,N_1838);
or U8959 (N_8959,N_3614,N_898);
nor U8960 (N_8960,N_2497,N_3823);
nand U8961 (N_8961,N_4237,N_2123);
and U8962 (N_8962,N_807,N_2541);
and U8963 (N_8963,N_756,N_2854);
and U8964 (N_8964,N_2705,N_1222);
and U8965 (N_8965,N_1864,N_20);
and U8966 (N_8966,N_4137,N_2128);
nor U8967 (N_8967,N_915,N_1254);
and U8968 (N_8968,N_523,N_1235);
nor U8969 (N_8969,N_3850,N_343);
nor U8970 (N_8970,N_64,N_4841);
xnor U8971 (N_8971,N_2016,N_2777);
xor U8972 (N_8972,N_3858,N_3132);
xor U8973 (N_8973,N_1693,N_3595);
and U8974 (N_8974,N_116,N_188);
and U8975 (N_8975,N_1666,N_3599);
xnor U8976 (N_8976,N_952,N_824);
nand U8977 (N_8977,N_4767,N_1016);
or U8978 (N_8978,N_3694,N_1785);
or U8979 (N_8979,N_818,N_4292);
nand U8980 (N_8980,N_2912,N_415);
xor U8981 (N_8981,N_3440,N_3065);
xnor U8982 (N_8982,N_3443,N_3275);
nor U8983 (N_8983,N_2954,N_1654);
and U8984 (N_8984,N_1208,N_3629);
nand U8985 (N_8985,N_3661,N_3034);
or U8986 (N_8986,N_2527,N_4396);
nor U8987 (N_8987,N_3829,N_4716);
or U8988 (N_8988,N_4222,N_85);
nand U8989 (N_8989,N_42,N_3039);
nor U8990 (N_8990,N_4635,N_730);
nand U8991 (N_8991,N_2550,N_1110);
nor U8992 (N_8992,N_4479,N_4843);
and U8993 (N_8993,N_4181,N_3239);
or U8994 (N_8994,N_4757,N_1057);
nor U8995 (N_8995,N_2101,N_3258);
nand U8996 (N_8996,N_4234,N_1515);
and U8997 (N_8997,N_1378,N_1346);
nand U8998 (N_8998,N_4054,N_926);
or U8999 (N_8999,N_1257,N_1624);
or U9000 (N_9000,N_1444,N_4347);
xnor U9001 (N_9001,N_1852,N_3205);
nor U9002 (N_9002,N_984,N_4154);
xnor U9003 (N_9003,N_3214,N_1495);
nand U9004 (N_9004,N_3272,N_3411);
and U9005 (N_9005,N_4281,N_3705);
or U9006 (N_9006,N_73,N_2866);
nor U9007 (N_9007,N_650,N_3474);
xor U9008 (N_9008,N_1121,N_1844);
or U9009 (N_9009,N_2403,N_1602);
or U9010 (N_9010,N_1813,N_269);
nand U9011 (N_9011,N_2975,N_4269);
or U9012 (N_9012,N_3414,N_678);
nand U9013 (N_9013,N_435,N_2830);
nor U9014 (N_9014,N_57,N_3448);
nand U9015 (N_9015,N_2543,N_2028);
nor U9016 (N_9016,N_3679,N_1704);
nand U9017 (N_9017,N_440,N_3453);
nor U9018 (N_9018,N_4900,N_4019);
and U9019 (N_9019,N_3324,N_1629);
xor U9020 (N_9020,N_2474,N_4313);
and U9021 (N_9021,N_913,N_1809);
xor U9022 (N_9022,N_3654,N_3172);
nand U9023 (N_9023,N_1322,N_3875);
nor U9024 (N_9024,N_3035,N_1281);
or U9025 (N_9025,N_1294,N_1228);
nand U9026 (N_9026,N_4133,N_430);
xor U9027 (N_9027,N_1805,N_2597);
or U9028 (N_9028,N_4573,N_4112);
xnor U9029 (N_9029,N_1628,N_3599);
nor U9030 (N_9030,N_3486,N_1824);
or U9031 (N_9031,N_2430,N_4942);
nand U9032 (N_9032,N_4046,N_4835);
or U9033 (N_9033,N_4672,N_132);
or U9034 (N_9034,N_1366,N_3887);
and U9035 (N_9035,N_2197,N_4335);
nor U9036 (N_9036,N_4365,N_620);
or U9037 (N_9037,N_1591,N_1545);
and U9038 (N_9038,N_385,N_574);
nor U9039 (N_9039,N_1300,N_905);
xor U9040 (N_9040,N_2826,N_3215);
and U9041 (N_9041,N_1139,N_2328);
and U9042 (N_9042,N_3127,N_1937);
xnor U9043 (N_9043,N_2902,N_4939);
xor U9044 (N_9044,N_4271,N_679);
nor U9045 (N_9045,N_3915,N_996);
nor U9046 (N_9046,N_4215,N_4818);
xor U9047 (N_9047,N_4307,N_2156);
nor U9048 (N_9048,N_3745,N_4427);
or U9049 (N_9049,N_3033,N_1232);
and U9050 (N_9050,N_1963,N_2400);
nor U9051 (N_9051,N_3492,N_3227);
or U9052 (N_9052,N_606,N_1497);
xor U9053 (N_9053,N_3740,N_2115);
xnor U9054 (N_9054,N_2868,N_2606);
nor U9055 (N_9055,N_3863,N_4069);
nor U9056 (N_9056,N_4868,N_1621);
nand U9057 (N_9057,N_3474,N_1194);
or U9058 (N_9058,N_1525,N_4);
and U9059 (N_9059,N_4035,N_3128);
and U9060 (N_9060,N_4153,N_188);
xnor U9061 (N_9061,N_1774,N_3986);
or U9062 (N_9062,N_4305,N_1559);
and U9063 (N_9063,N_4064,N_3787);
or U9064 (N_9064,N_4898,N_1832);
xnor U9065 (N_9065,N_672,N_590);
or U9066 (N_9066,N_3586,N_1014);
nand U9067 (N_9067,N_3303,N_3064);
xnor U9068 (N_9068,N_1883,N_4151);
xnor U9069 (N_9069,N_4779,N_4066);
nor U9070 (N_9070,N_1000,N_3575);
or U9071 (N_9071,N_3018,N_4657);
or U9072 (N_9072,N_4679,N_4035);
or U9073 (N_9073,N_3900,N_729);
nand U9074 (N_9074,N_4181,N_3579);
and U9075 (N_9075,N_4182,N_2654);
and U9076 (N_9076,N_341,N_486);
and U9077 (N_9077,N_1175,N_1726);
xor U9078 (N_9078,N_4605,N_1358);
nand U9079 (N_9079,N_3610,N_138);
nand U9080 (N_9080,N_2119,N_2251);
nand U9081 (N_9081,N_4028,N_2634);
or U9082 (N_9082,N_652,N_4467);
or U9083 (N_9083,N_2615,N_284);
or U9084 (N_9084,N_3124,N_4212);
nand U9085 (N_9085,N_634,N_4859);
nand U9086 (N_9086,N_1321,N_3476);
and U9087 (N_9087,N_3773,N_4621);
or U9088 (N_9088,N_1188,N_607);
and U9089 (N_9089,N_3683,N_1877);
nor U9090 (N_9090,N_134,N_3980);
nor U9091 (N_9091,N_2759,N_967);
or U9092 (N_9092,N_3674,N_157);
and U9093 (N_9093,N_2216,N_2440);
or U9094 (N_9094,N_819,N_1149);
nand U9095 (N_9095,N_1735,N_1710);
and U9096 (N_9096,N_3710,N_3274);
xnor U9097 (N_9097,N_2323,N_267);
or U9098 (N_9098,N_3208,N_77);
and U9099 (N_9099,N_1067,N_73);
nor U9100 (N_9100,N_4699,N_2450);
xor U9101 (N_9101,N_638,N_722);
xor U9102 (N_9102,N_1868,N_324);
nand U9103 (N_9103,N_4561,N_414);
or U9104 (N_9104,N_1826,N_1641);
nor U9105 (N_9105,N_1387,N_3117);
and U9106 (N_9106,N_4876,N_1668);
xor U9107 (N_9107,N_3660,N_2978);
or U9108 (N_9108,N_4806,N_1769);
and U9109 (N_9109,N_3336,N_3061);
nor U9110 (N_9110,N_2194,N_54);
and U9111 (N_9111,N_1504,N_2413);
or U9112 (N_9112,N_298,N_3236);
xor U9113 (N_9113,N_3742,N_2094);
and U9114 (N_9114,N_258,N_2277);
xor U9115 (N_9115,N_1901,N_1487);
and U9116 (N_9116,N_2453,N_4106);
or U9117 (N_9117,N_150,N_2339);
nor U9118 (N_9118,N_2811,N_1699);
or U9119 (N_9119,N_4329,N_4294);
and U9120 (N_9120,N_2548,N_4021);
nand U9121 (N_9121,N_3301,N_407);
or U9122 (N_9122,N_464,N_2842);
or U9123 (N_9123,N_667,N_2095);
or U9124 (N_9124,N_336,N_3793);
xor U9125 (N_9125,N_303,N_1437);
nor U9126 (N_9126,N_2975,N_2556);
nand U9127 (N_9127,N_2692,N_3275);
or U9128 (N_9128,N_2205,N_3380);
nand U9129 (N_9129,N_1568,N_4931);
xnor U9130 (N_9130,N_2105,N_4762);
nor U9131 (N_9131,N_2029,N_1766);
nor U9132 (N_9132,N_3193,N_1623);
xnor U9133 (N_9133,N_4085,N_2740);
and U9134 (N_9134,N_2285,N_4909);
or U9135 (N_9135,N_4790,N_3113);
nand U9136 (N_9136,N_15,N_1832);
nand U9137 (N_9137,N_1973,N_2149);
and U9138 (N_9138,N_3771,N_448);
nor U9139 (N_9139,N_3480,N_775);
or U9140 (N_9140,N_4023,N_1269);
xor U9141 (N_9141,N_2821,N_1016);
nor U9142 (N_9142,N_1515,N_327);
nand U9143 (N_9143,N_463,N_2771);
nand U9144 (N_9144,N_2163,N_3667);
nand U9145 (N_9145,N_704,N_2226);
and U9146 (N_9146,N_455,N_3343);
nor U9147 (N_9147,N_2653,N_541);
nand U9148 (N_9148,N_4003,N_896);
nor U9149 (N_9149,N_2145,N_90);
nand U9150 (N_9150,N_4928,N_102);
and U9151 (N_9151,N_4142,N_3950);
xor U9152 (N_9152,N_1811,N_2901);
nor U9153 (N_9153,N_4637,N_4859);
nand U9154 (N_9154,N_4504,N_1883);
or U9155 (N_9155,N_417,N_2202);
and U9156 (N_9156,N_3227,N_2893);
nand U9157 (N_9157,N_3467,N_2942);
xor U9158 (N_9158,N_1847,N_4134);
or U9159 (N_9159,N_3793,N_2077);
nor U9160 (N_9160,N_2836,N_451);
nand U9161 (N_9161,N_1424,N_1947);
nand U9162 (N_9162,N_3851,N_1411);
nand U9163 (N_9163,N_1114,N_1937);
or U9164 (N_9164,N_2664,N_4277);
or U9165 (N_9165,N_993,N_222);
xnor U9166 (N_9166,N_74,N_2223);
or U9167 (N_9167,N_4016,N_2870);
xor U9168 (N_9168,N_1957,N_870);
nor U9169 (N_9169,N_397,N_2970);
or U9170 (N_9170,N_4033,N_94);
nand U9171 (N_9171,N_2684,N_2068);
nand U9172 (N_9172,N_3984,N_2551);
and U9173 (N_9173,N_4252,N_4439);
or U9174 (N_9174,N_3336,N_552);
nand U9175 (N_9175,N_4277,N_56);
and U9176 (N_9176,N_810,N_4318);
nand U9177 (N_9177,N_1435,N_4625);
or U9178 (N_9178,N_4630,N_3811);
nand U9179 (N_9179,N_4571,N_2298);
or U9180 (N_9180,N_2338,N_1818);
or U9181 (N_9181,N_3336,N_550);
and U9182 (N_9182,N_4702,N_4135);
and U9183 (N_9183,N_2655,N_894);
xnor U9184 (N_9184,N_4692,N_4254);
and U9185 (N_9185,N_4607,N_1310);
or U9186 (N_9186,N_830,N_2037);
xnor U9187 (N_9187,N_1240,N_1809);
nor U9188 (N_9188,N_3529,N_3866);
nand U9189 (N_9189,N_520,N_383);
or U9190 (N_9190,N_920,N_3837);
or U9191 (N_9191,N_2229,N_2594);
and U9192 (N_9192,N_3429,N_3073);
and U9193 (N_9193,N_3323,N_2912);
or U9194 (N_9194,N_3424,N_1410);
xnor U9195 (N_9195,N_1444,N_2525);
nor U9196 (N_9196,N_3782,N_1640);
nand U9197 (N_9197,N_3879,N_3085);
nor U9198 (N_9198,N_4635,N_1784);
nand U9199 (N_9199,N_2476,N_3129);
nor U9200 (N_9200,N_1163,N_4298);
xor U9201 (N_9201,N_269,N_1039);
xor U9202 (N_9202,N_2416,N_857);
and U9203 (N_9203,N_560,N_948);
or U9204 (N_9204,N_3470,N_2589);
and U9205 (N_9205,N_33,N_666);
xor U9206 (N_9206,N_211,N_3534);
and U9207 (N_9207,N_161,N_1902);
xnor U9208 (N_9208,N_2279,N_2876);
nand U9209 (N_9209,N_188,N_2890);
or U9210 (N_9210,N_2599,N_4150);
and U9211 (N_9211,N_2543,N_3431);
or U9212 (N_9212,N_2241,N_2015);
nor U9213 (N_9213,N_1931,N_2667);
nor U9214 (N_9214,N_2114,N_302);
or U9215 (N_9215,N_3991,N_4755);
nand U9216 (N_9216,N_3862,N_4501);
or U9217 (N_9217,N_3189,N_146);
and U9218 (N_9218,N_2049,N_338);
nand U9219 (N_9219,N_4286,N_3697);
xor U9220 (N_9220,N_1511,N_1623);
or U9221 (N_9221,N_1972,N_1283);
and U9222 (N_9222,N_2338,N_2079);
or U9223 (N_9223,N_1805,N_1469);
nor U9224 (N_9224,N_2511,N_3310);
nand U9225 (N_9225,N_897,N_2899);
xor U9226 (N_9226,N_2487,N_2222);
nand U9227 (N_9227,N_2307,N_1911);
nand U9228 (N_9228,N_1137,N_1797);
and U9229 (N_9229,N_3530,N_1975);
xor U9230 (N_9230,N_2891,N_3806);
nor U9231 (N_9231,N_4551,N_4624);
nand U9232 (N_9232,N_488,N_457);
nand U9233 (N_9233,N_4321,N_4615);
nor U9234 (N_9234,N_83,N_2936);
and U9235 (N_9235,N_169,N_3552);
and U9236 (N_9236,N_271,N_2587);
nand U9237 (N_9237,N_3324,N_3086);
nor U9238 (N_9238,N_4772,N_615);
nor U9239 (N_9239,N_4434,N_1495);
nor U9240 (N_9240,N_118,N_3379);
nor U9241 (N_9241,N_2951,N_1789);
nor U9242 (N_9242,N_1916,N_2057);
nand U9243 (N_9243,N_1514,N_4257);
xor U9244 (N_9244,N_1091,N_1044);
nand U9245 (N_9245,N_4706,N_1711);
xnor U9246 (N_9246,N_2912,N_2830);
nand U9247 (N_9247,N_4708,N_2240);
and U9248 (N_9248,N_309,N_4896);
xor U9249 (N_9249,N_831,N_3189);
xnor U9250 (N_9250,N_3570,N_4146);
xor U9251 (N_9251,N_4224,N_4577);
or U9252 (N_9252,N_3338,N_4761);
and U9253 (N_9253,N_4535,N_421);
nand U9254 (N_9254,N_4979,N_2949);
nor U9255 (N_9255,N_1837,N_2640);
xnor U9256 (N_9256,N_408,N_1936);
nor U9257 (N_9257,N_4365,N_2089);
nor U9258 (N_9258,N_234,N_2582);
or U9259 (N_9259,N_4472,N_2517);
xnor U9260 (N_9260,N_4083,N_860);
xor U9261 (N_9261,N_4313,N_2710);
xnor U9262 (N_9262,N_4896,N_3204);
and U9263 (N_9263,N_2776,N_832);
xor U9264 (N_9264,N_2443,N_1602);
xnor U9265 (N_9265,N_3169,N_3554);
nor U9266 (N_9266,N_3258,N_1311);
or U9267 (N_9267,N_3682,N_826);
nor U9268 (N_9268,N_4166,N_3554);
and U9269 (N_9269,N_3694,N_4981);
nor U9270 (N_9270,N_4155,N_2749);
xor U9271 (N_9271,N_4779,N_4028);
and U9272 (N_9272,N_1253,N_3573);
nand U9273 (N_9273,N_3364,N_3407);
nor U9274 (N_9274,N_3217,N_704);
nor U9275 (N_9275,N_2887,N_3500);
or U9276 (N_9276,N_2815,N_3647);
nand U9277 (N_9277,N_2165,N_2764);
nor U9278 (N_9278,N_1898,N_2873);
xnor U9279 (N_9279,N_3570,N_2723);
and U9280 (N_9280,N_1446,N_1930);
xnor U9281 (N_9281,N_1460,N_3200);
nor U9282 (N_9282,N_3813,N_4156);
nand U9283 (N_9283,N_2428,N_2281);
nor U9284 (N_9284,N_785,N_3894);
xnor U9285 (N_9285,N_2234,N_4918);
and U9286 (N_9286,N_563,N_3789);
and U9287 (N_9287,N_4406,N_584);
and U9288 (N_9288,N_4220,N_1706);
nand U9289 (N_9289,N_4442,N_1839);
nand U9290 (N_9290,N_1725,N_1066);
or U9291 (N_9291,N_4904,N_1502);
and U9292 (N_9292,N_4809,N_425);
xnor U9293 (N_9293,N_4399,N_1779);
and U9294 (N_9294,N_3326,N_1500);
or U9295 (N_9295,N_1199,N_301);
nand U9296 (N_9296,N_232,N_1885);
nand U9297 (N_9297,N_2968,N_546);
nor U9298 (N_9298,N_3978,N_1393);
or U9299 (N_9299,N_1641,N_646);
and U9300 (N_9300,N_392,N_2538);
nand U9301 (N_9301,N_1977,N_937);
and U9302 (N_9302,N_1410,N_3961);
nand U9303 (N_9303,N_2606,N_839);
xnor U9304 (N_9304,N_4994,N_1542);
and U9305 (N_9305,N_2542,N_4253);
nor U9306 (N_9306,N_3713,N_846);
and U9307 (N_9307,N_2362,N_4148);
and U9308 (N_9308,N_2288,N_3894);
xor U9309 (N_9309,N_1474,N_202);
and U9310 (N_9310,N_2018,N_530);
or U9311 (N_9311,N_2928,N_4170);
or U9312 (N_9312,N_1055,N_91);
or U9313 (N_9313,N_4313,N_4229);
xnor U9314 (N_9314,N_3528,N_329);
or U9315 (N_9315,N_821,N_551);
nor U9316 (N_9316,N_1254,N_428);
and U9317 (N_9317,N_4382,N_4672);
and U9318 (N_9318,N_3270,N_1799);
xor U9319 (N_9319,N_513,N_3243);
and U9320 (N_9320,N_720,N_2888);
and U9321 (N_9321,N_2825,N_1233);
xnor U9322 (N_9322,N_3084,N_664);
nor U9323 (N_9323,N_430,N_253);
nand U9324 (N_9324,N_2390,N_1612);
and U9325 (N_9325,N_3507,N_3350);
or U9326 (N_9326,N_353,N_2687);
xor U9327 (N_9327,N_925,N_3333);
nor U9328 (N_9328,N_1640,N_686);
or U9329 (N_9329,N_2913,N_2566);
nand U9330 (N_9330,N_1373,N_1511);
and U9331 (N_9331,N_80,N_2507);
xor U9332 (N_9332,N_3313,N_1435);
nand U9333 (N_9333,N_812,N_199);
and U9334 (N_9334,N_3713,N_576);
xor U9335 (N_9335,N_4670,N_299);
nand U9336 (N_9336,N_4400,N_2071);
xnor U9337 (N_9337,N_2255,N_899);
nor U9338 (N_9338,N_1128,N_3228);
xor U9339 (N_9339,N_2451,N_1425);
and U9340 (N_9340,N_1518,N_105);
or U9341 (N_9341,N_1089,N_2437);
xor U9342 (N_9342,N_208,N_655);
nand U9343 (N_9343,N_3057,N_472);
xnor U9344 (N_9344,N_3410,N_2389);
and U9345 (N_9345,N_2444,N_4331);
and U9346 (N_9346,N_226,N_1911);
and U9347 (N_9347,N_3605,N_4023);
nor U9348 (N_9348,N_3468,N_1765);
or U9349 (N_9349,N_607,N_775);
and U9350 (N_9350,N_4745,N_2576);
or U9351 (N_9351,N_1961,N_1376);
or U9352 (N_9352,N_3163,N_1460);
xor U9353 (N_9353,N_3264,N_4773);
nand U9354 (N_9354,N_3518,N_1635);
nand U9355 (N_9355,N_3894,N_2306);
xor U9356 (N_9356,N_111,N_3020);
and U9357 (N_9357,N_348,N_4720);
and U9358 (N_9358,N_4282,N_2597);
or U9359 (N_9359,N_3035,N_4465);
and U9360 (N_9360,N_641,N_3905);
nand U9361 (N_9361,N_3951,N_3616);
nor U9362 (N_9362,N_1039,N_2946);
nand U9363 (N_9363,N_2461,N_2054);
nor U9364 (N_9364,N_4313,N_3120);
and U9365 (N_9365,N_4467,N_3799);
nand U9366 (N_9366,N_684,N_2138);
or U9367 (N_9367,N_4740,N_1441);
nand U9368 (N_9368,N_3585,N_2763);
nand U9369 (N_9369,N_2908,N_27);
or U9370 (N_9370,N_4279,N_4189);
and U9371 (N_9371,N_897,N_1972);
xnor U9372 (N_9372,N_1517,N_1701);
or U9373 (N_9373,N_2612,N_2590);
or U9374 (N_9374,N_1288,N_3124);
nor U9375 (N_9375,N_4159,N_1986);
nor U9376 (N_9376,N_2056,N_1606);
nor U9377 (N_9377,N_942,N_733);
xor U9378 (N_9378,N_298,N_2972);
nor U9379 (N_9379,N_3866,N_4308);
xnor U9380 (N_9380,N_759,N_487);
or U9381 (N_9381,N_1486,N_849);
or U9382 (N_9382,N_4865,N_800);
nand U9383 (N_9383,N_4636,N_3645);
nand U9384 (N_9384,N_4336,N_748);
xor U9385 (N_9385,N_761,N_2285);
xnor U9386 (N_9386,N_1389,N_4844);
nand U9387 (N_9387,N_330,N_556);
or U9388 (N_9388,N_3781,N_765);
xnor U9389 (N_9389,N_3491,N_3432);
or U9390 (N_9390,N_593,N_1517);
nor U9391 (N_9391,N_3665,N_4221);
xor U9392 (N_9392,N_960,N_1327);
nor U9393 (N_9393,N_1944,N_2870);
nor U9394 (N_9394,N_974,N_963);
nand U9395 (N_9395,N_4487,N_2649);
xor U9396 (N_9396,N_3414,N_3293);
nor U9397 (N_9397,N_4837,N_3319);
and U9398 (N_9398,N_3079,N_1733);
and U9399 (N_9399,N_198,N_692);
xnor U9400 (N_9400,N_2937,N_2121);
nor U9401 (N_9401,N_553,N_1291);
nand U9402 (N_9402,N_3863,N_1959);
nand U9403 (N_9403,N_3726,N_3094);
xnor U9404 (N_9404,N_3909,N_2989);
xor U9405 (N_9405,N_1434,N_4164);
nand U9406 (N_9406,N_2841,N_2649);
nand U9407 (N_9407,N_4986,N_2425);
nor U9408 (N_9408,N_1228,N_3802);
nor U9409 (N_9409,N_4986,N_2145);
or U9410 (N_9410,N_1493,N_1173);
or U9411 (N_9411,N_582,N_2092);
and U9412 (N_9412,N_1793,N_3914);
nand U9413 (N_9413,N_252,N_2373);
nor U9414 (N_9414,N_3296,N_1725);
nand U9415 (N_9415,N_1791,N_783);
or U9416 (N_9416,N_3692,N_3141);
nand U9417 (N_9417,N_3363,N_4223);
xor U9418 (N_9418,N_2927,N_1778);
or U9419 (N_9419,N_3985,N_3581);
and U9420 (N_9420,N_2791,N_2824);
and U9421 (N_9421,N_948,N_4527);
and U9422 (N_9422,N_695,N_3543);
and U9423 (N_9423,N_2846,N_925);
and U9424 (N_9424,N_3436,N_1753);
xor U9425 (N_9425,N_4920,N_2010);
or U9426 (N_9426,N_4389,N_1034);
and U9427 (N_9427,N_4156,N_2633);
nor U9428 (N_9428,N_1826,N_161);
xor U9429 (N_9429,N_3109,N_1089);
nor U9430 (N_9430,N_622,N_816);
nor U9431 (N_9431,N_1633,N_3900);
nor U9432 (N_9432,N_2325,N_3794);
xor U9433 (N_9433,N_1243,N_281);
or U9434 (N_9434,N_487,N_2442);
and U9435 (N_9435,N_2689,N_4754);
nor U9436 (N_9436,N_4995,N_692);
and U9437 (N_9437,N_3683,N_4125);
or U9438 (N_9438,N_1878,N_4976);
nand U9439 (N_9439,N_3122,N_2229);
nand U9440 (N_9440,N_3319,N_3207);
nand U9441 (N_9441,N_3058,N_997);
nand U9442 (N_9442,N_3561,N_2206);
nor U9443 (N_9443,N_14,N_1253);
and U9444 (N_9444,N_3636,N_2059);
xnor U9445 (N_9445,N_2525,N_1070);
nand U9446 (N_9446,N_4552,N_1201);
nor U9447 (N_9447,N_2854,N_1356);
nand U9448 (N_9448,N_3017,N_1469);
xnor U9449 (N_9449,N_646,N_2462);
nand U9450 (N_9450,N_3521,N_987);
nor U9451 (N_9451,N_439,N_52);
and U9452 (N_9452,N_2804,N_4528);
or U9453 (N_9453,N_4964,N_2094);
xor U9454 (N_9454,N_2985,N_170);
xor U9455 (N_9455,N_3951,N_2370);
xor U9456 (N_9456,N_2057,N_3361);
nor U9457 (N_9457,N_3,N_1739);
nand U9458 (N_9458,N_2330,N_11);
and U9459 (N_9459,N_4123,N_3734);
xnor U9460 (N_9460,N_3795,N_1424);
nor U9461 (N_9461,N_2711,N_2575);
or U9462 (N_9462,N_1972,N_4001);
nand U9463 (N_9463,N_3604,N_2875);
nor U9464 (N_9464,N_1931,N_1783);
xor U9465 (N_9465,N_4560,N_4562);
or U9466 (N_9466,N_3152,N_1846);
and U9467 (N_9467,N_3222,N_2240);
xor U9468 (N_9468,N_3856,N_4411);
nor U9469 (N_9469,N_2478,N_1738);
nor U9470 (N_9470,N_709,N_4055);
nand U9471 (N_9471,N_498,N_3499);
nand U9472 (N_9472,N_1374,N_2577);
xor U9473 (N_9473,N_1019,N_4686);
xor U9474 (N_9474,N_2559,N_4883);
nand U9475 (N_9475,N_1188,N_4696);
nand U9476 (N_9476,N_4856,N_853);
nor U9477 (N_9477,N_1740,N_2558);
nand U9478 (N_9478,N_585,N_3059);
nand U9479 (N_9479,N_95,N_1208);
or U9480 (N_9480,N_603,N_4675);
or U9481 (N_9481,N_2400,N_3891);
and U9482 (N_9482,N_1150,N_2125);
nand U9483 (N_9483,N_4411,N_787);
nor U9484 (N_9484,N_3046,N_400);
xor U9485 (N_9485,N_2208,N_4529);
nand U9486 (N_9486,N_3650,N_2012);
and U9487 (N_9487,N_3544,N_3213);
nor U9488 (N_9488,N_846,N_1844);
nor U9489 (N_9489,N_2530,N_4087);
nor U9490 (N_9490,N_3860,N_2695);
nand U9491 (N_9491,N_3092,N_2668);
xor U9492 (N_9492,N_961,N_1045);
xnor U9493 (N_9493,N_263,N_4105);
nand U9494 (N_9494,N_3518,N_3351);
nor U9495 (N_9495,N_2805,N_984);
nor U9496 (N_9496,N_4958,N_3925);
nand U9497 (N_9497,N_1141,N_2820);
or U9498 (N_9498,N_1234,N_2803);
xor U9499 (N_9499,N_2082,N_3938);
nor U9500 (N_9500,N_4649,N_3479);
and U9501 (N_9501,N_2633,N_2877);
xnor U9502 (N_9502,N_3392,N_793);
or U9503 (N_9503,N_1455,N_4570);
or U9504 (N_9504,N_981,N_1352);
or U9505 (N_9505,N_497,N_4368);
or U9506 (N_9506,N_1248,N_641);
xnor U9507 (N_9507,N_1922,N_954);
nor U9508 (N_9508,N_1809,N_1301);
nor U9509 (N_9509,N_4011,N_4388);
nor U9510 (N_9510,N_2321,N_1259);
nor U9511 (N_9511,N_2117,N_592);
xnor U9512 (N_9512,N_110,N_4685);
nand U9513 (N_9513,N_401,N_2218);
and U9514 (N_9514,N_4363,N_2743);
and U9515 (N_9515,N_2458,N_1466);
nor U9516 (N_9516,N_4854,N_3206);
and U9517 (N_9517,N_3380,N_4260);
and U9518 (N_9518,N_1890,N_3699);
xor U9519 (N_9519,N_2057,N_2047);
nand U9520 (N_9520,N_895,N_4345);
nand U9521 (N_9521,N_2949,N_1822);
and U9522 (N_9522,N_4679,N_2046);
nand U9523 (N_9523,N_4422,N_923);
nor U9524 (N_9524,N_3690,N_2348);
nand U9525 (N_9525,N_4233,N_1896);
or U9526 (N_9526,N_1342,N_4427);
nor U9527 (N_9527,N_2714,N_3743);
or U9528 (N_9528,N_392,N_358);
and U9529 (N_9529,N_4512,N_4044);
nor U9530 (N_9530,N_562,N_1385);
and U9531 (N_9531,N_3002,N_3208);
or U9532 (N_9532,N_668,N_4621);
or U9533 (N_9533,N_3082,N_4592);
and U9534 (N_9534,N_4337,N_3455);
nor U9535 (N_9535,N_3320,N_2679);
or U9536 (N_9536,N_4052,N_2379);
and U9537 (N_9537,N_1204,N_4791);
or U9538 (N_9538,N_35,N_942);
and U9539 (N_9539,N_125,N_2005);
or U9540 (N_9540,N_1238,N_301);
or U9541 (N_9541,N_4509,N_4221);
and U9542 (N_9542,N_3517,N_4765);
and U9543 (N_9543,N_4135,N_4364);
nand U9544 (N_9544,N_1245,N_4392);
nand U9545 (N_9545,N_3414,N_2278);
nand U9546 (N_9546,N_999,N_4373);
or U9547 (N_9547,N_2132,N_2310);
and U9548 (N_9548,N_3593,N_2969);
and U9549 (N_9549,N_1525,N_681);
xor U9550 (N_9550,N_760,N_4363);
and U9551 (N_9551,N_2558,N_1642);
and U9552 (N_9552,N_4305,N_4447);
nor U9553 (N_9553,N_4030,N_984);
xnor U9554 (N_9554,N_1501,N_2022);
nor U9555 (N_9555,N_3941,N_3732);
and U9556 (N_9556,N_1232,N_4073);
or U9557 (N_9557,N_1941,N_1662);
or U9558 (N_9558,N_2062,N_57);
nor U9559 (N_9559,N_4638,N_115);
xor U9560 (N_9560,N_3460,N_966);
or U9561 (N_9561,N_2692,N_3063);
or U9562 (N_9562,N_373,N_4481);
or U9563 (N_9563,N_1034,N_3328);
xor U9564 (N_9564,N_3891,N_3325);
nor U9565 (N_9565,N_2245,N_2737);
nand U9566 (N_9566,N_1251,N_886);
nor U9567 (N_9567,N_4284,N_2350);
nor U9568 (N_9568,N_3275,N_3440);
nand U9569 (N_9569,N_3812,N_3560);
xnor U9570 (N_9570,N_2435,N_810);
nor U9571 (N_9571,N_3616,N_2511);
xor U9572 (N_9572,N_3526,N_2318);
nand U9573 (N_9573,N_3570,N_2144);
nand U9574 (N_9574,N_1427,N_2474);
xor U9575 (N_9575,N_3764,N_1031);
or U9576 (N_9576,N_4,N_1645);
nand U9577 (N_9577,N_4197,N_3146);
nor U9578 (N_9578,N_1560,N_4605);
xnor U9579 (N_9579,N_3182,N_1132);
nor U9580 (N_9580,N_6,N_3549);
or U9581 (N_9581,N_309,N_584);
or U9582 (N_9582,N_770,N_1572);
xor U9583 (N_9583,N_4753,N_4314);
or U9584 (N_9584,N_4247,N_2078);
xnor U9585 (N_9585,N_1259,N_1452);
nand U9586 (N_9586,N_2910,N_194);
xnor U9587 (N_9587,N_1391,N_3827);
nand U9588 (N_9588,N_2266,N_4644);
xnor U9589 (N_9589,N_3594,N_2913);
or U9590 (N_9590,N_1985,N_4806);
nand U9591 (N_9591,N_1360,N_265);
or U9592 (N_9592,N_2787,N_4930);
xnor U9593 (N_9593,N_3051,N_4689);
xor U9594 (N_9594,N_4302,N_616);
nor U9595 (N_9595,N_2422,N_4836);
nor U9596 (N_9596,N_1232,N_614);
nor U9597 (N_9597,N_264,N_1833);
nand U9598 (N_9598,N_4176,N_3967);
nor U9599 (N_9599,N_359,N_1378);
and U9600 (N_9600,N_39,N_538);
or U9601 (N_9601,N_2767,N_420);
and U9602 (N_9602,N_1435,N_1228);
or U9603 (N_9603,N_895,N_2739);
nor U9604 (N_9604,N_450,N_330);
and U9605 (N_9605,N_4401,N_4061);
xnor U9606 (N_9606,N_4022,N_1088);
and U9607 (N_9607,N_2633,N_332);
or U9608 (N_9608,N_4961,N_4846);
and U9609 (N_9609,N_3518,N_3482);
xnor U9610 (N_9610,N_2198,N_2115);
and U9611 (N_9611,N_1890,N_229);
or U9612 (N_9612,N_4243,N_3168);
or U9613 (N_9613,N_3781,N_3680);
nor U9614 (N_9614,N_4632,N_1694);
nand U9615 (N_9615,N_1951,N_2114);
xnor U9616 (N_9616,N_4167,N_3350);
or U9617 (N_9617,N_176,N_1935);
nand U9618 (N_9618,N_3338,N_3861);
or U9619 (N_9619,N_1106,N_2045);
nor U9620 (N_9620,N_4721,N_1047);
xnor U9621 (N_9621,N_2825,N_4874);
or U9622 (N_9622,N_3,N_2079);
nand U9623 (N_9623,N_2594,N_1507);
nand U9624 (N_9624,N_1751,N_3382);
and U9625 (N_9625,N_68,N_3394);
nor U9626 (N_9626,N_2020,N_1611);
xnor U9627 (N_9627,N_1538,N_370);
nand U9628 (N_9628,N_3440,N_1048);
xor U9629 (N_9629,N_1783,N_856);
and U9630 (N_9630,N_1850,N_1309);
nand U9631 (N_9631,N_3147,N_4616);
nor U9632 (N_9632,N_2696,N_4167);
xnor U9633 (N_9633,N_86,N_1493);
nand U9634 (N_9634,N_4024,N_1580);
nand U9635 (N_9635,N_3888,N_1494);
and U9636 (N_9636,N_2233,N_605);
and U9637 (N_9637,N_2689,N_1083);
nand U9638 (N_9638,N_4881,N_1);
nand U9639 (N_9639,N_3942,N_4307);
nor U9640 (N_9640,N_1032,N_4975);
and U9641 (N_9641,N_407,N_763);
nand U9642 (N_9642,N_556,N_1389);
and U9643 (N_9643,N_2059,N_2930);
and U9644 (N_9644,N_4040,N_3778);
and U9645 (N_9645,N_4642,N_1931);
and U9646 (N_9646,N_4913,N_1435);
nand U9647 (N_9647,N_2626,N_264);
or U9648 (N_9648,N_2257,N_4027);
nor U9649 (N_9649,N_1424,N_2256);
or U9650 (N_9650,N_3062,N_250);
nor U9651 (N_9651,N_1145,N_2273);
and U9652 (N_9652,N_1153,N_4809);
or U9653 (N_9653,N_4531,N_2646);
or U9654 (N_9654,N_4145,N_3691);
nor U9655 (N_9655,N_2769,N_26);
nor U9656 (N_9656,N_3066,N_3438);
and U9657 (N_9657,N_3009,N_3083);
nand U9658 (N_9658,N_3111,N_2328);
or U9659 (N_9659,N_3210,N_2821);
nand U9660 (N_9660,N_2196,N_3617);
xor U9661 (N_9661,N_402,N_2775);
nor U9662 (N_9662,N_4160,N_3834);
xor U9663 (N_9663,N_4529,N_593);
or U9664 (N_9664,N_2258,N_2541);
nor U9665 (N_9665,N_2024,N_4030);
xnor U9666 (N_9666,N_4250,N_4941);
nand U9667 (N_9667,N_38,N_2150);
nor U9668 (N_9668,N_4958,N_3499);
and U9669 (N_9669,N_4408,N_3125);
or U9670 (N_9670,N_806,N_4068);
nand U9671 (N_9671,N_3072,N_4918);
and U9672 (N_9672,N_2779,N_3726);
or U9673 (N_9673,N_4373,N_181);
and U9674 (N_9674,N_4799,N_573);
nor U9675 (N_9675,N_3435,N_2983);
nand U9676 (N_9676,N_3621,N_4320);
and U9677 (N_9677,N_852,N_4365);
or U9678 (N_9678,N_2300,N_1852);
nor U9679 (N_9679,N_2904,N_3765);
and U9680 (N_9680,N_3358,N_3049);
xnor U9681 (N_9681,N_3021,N_1659);
or U9682 (N_9682,N_2750,N_2072);
xnor U9683 (N_9683,N_4205,N_4677);
nor U9684 (N_9684,N_478,N_1886);
xnor U9685 (N_9685,N_3619,N_3770);
or U9686 (N_9686,N_3342,N_4369);
or U9687 (N_9687,N_3578,N_4435);
xor U9688 (N_9688,N_130,N_529);
xnor U9689 (N_9689,N_3992,N_1578);
xnor U9690 (N_9690,N_1977,N_4050);
xor U9691 (N_9691,N_104,N_3250);
xor U9692 (N_9692,N_3229,N_3398);
or U9693 (N_9693,N_3569,N_1945);
nand U9694 (N_9694,N_2826,N_1898);
or U9695 (N_9695,N_4020,N_46);
or U9696 (N_9696,N_2563,N_504);
nor U9697 (N_9697,N_2768,N_3222);
nand U9698 (N_9698,N_4110,N_2048);
nor U9699 (N_9699,N_2980,N_2856);
and U9700 (N_9700,N_4246,N_4184);
nand U9701 (N_9701,N_356,N_1827);
xor U9702 (N_9702,N_3182,N_4652);
nand U9703 (N_9703,N_2418,N_3219);
or U9704 (N_9704,N_3709,N_697);
nand U9705 (N_9705,N_4375,N_1783);
nand U9706 (N_9706,N_1920,N_2645);
and U9707 (N_9707,N_2447,N_4756);
and U9708 (N_9708,N_1816,N_73);
or U9709 (N_9709,N_3539,N_3458);
nor U9710 (N_9710,N_2975,N_1090);
or U9711 (N_9711,N_1783,N_2693);
nor U9712 (N_9712,N_347,N_3105);
nand U9713 (N_9713,N_786,N_4322);
nor U9714 (N_9714,N_3492,N_1605);
and U9715 (N_9715,N_4766,N_2384);
nand U9716 (N_9716,N_4074,N_4199);
or U9717 (N_9717,N_4901,N_3106);
or U9718 (N_9718,N_2191,N_4792);
and U9719 (N_9719,N_1407,N_4966);
xor U9720 (N_9720,N_3263,N_127);
nor U9721 (N_9721,N_4760,N_4572);
and U9722 (N_9722,N_3174,N_1301);
and U9723 (N_9723,N_1461,N_3334);
or U9724 (N_9724,N_1851,N_4842);
and U9725 (N_9725,N_3796,N_3434);
nand U9726 (N_9726,N_593,N_1532);
and U9727 (N_9727,N_425,N_2626);
xor U9728 (N_9728,N_1168,N_2993);
nor U9729 (N_9729,N_3193,N_2677);
nor U9730 (N_9730,N_3468,N_186);
nand U9731 (N_9731,N_3326,N_4307);
or U9732 (N_9732,N_661,N_4582);
or U9733 (N_9733,N_3703,N_839);
xnor U9734 (N_9734,N_1735,N_3209);
xnor U9735 (N_9735,N_1535,N_2527);
nand U9736 (N_9736,N_1284,N_2857);
or U9737 (N_9737,N_2555,N_4020);
nand U9738 (N_9738,N_3580,N_3695);
and U9739 (N_9739,N_237,N_4219);
nor U9740 (N_9740,N_3793,N_2948);
xnor U9741 (N_9741,N_105,N_117);
or U9742 (N_9742,N_3999,N_83);
or U9743 (N_9743,N_1692,N_3421);
nor U9744 (N_9744,N_1702,N_2885);
xnor U9745 (N_9745,N_3481,N_4644);
nor U9746 (N_9746,N_3633,N_4919);
and U9747 (N_9747,N_2427,N_1759);
nor U9748 (N_9748,N_476,N_575);
or U9749 (N_9749,N_1048,N_327);
xnor U9750 (N_9750,N_651,N_4734);
xor U9751 (N_9751,N_2118,N_3843);
nor U9752 (N_9752,N_3418,N_3974);
nor U9753 (N_9753,N_947,N_4989);
and U9754 (N_9754,N_1081,N_4430);
nor U9755 (N_9755,N_3787,N_1951);
xnor U9756 (N_9756,N_3317,N_3075);
nand U9757 (N_9757,N_3261,N_1189);
or U9758 (N_9758,N_3154,N_2037);
and U9759 (N_9759,N_1260,N_2249);
and U9760 (N_9760,N_467,N_1041);
and U9761 (N_9761,N_2429,N_459);
nand U9762 (N_9762,N_2819,N_3446);
and U9763 (N_9763,N_2332,N_3001);
xnor U9764 (N_9764,N_3109,N_1374);
nand U9765 (N_9765,N_2316,N_2079);
nand U9766 (N_9766,N_2334,N_2659);
nand U9767 (N_9767,N_1864,N_2610);
nand U9768 (N_9768,N_252,N_72);
nor U9769 (N_9769,N_2736,N_3148);
xnor U9770 (N_9770,N_4700,N_3981);
xor U9771 (N_9771,N_4172,N_3401);
nor U9772 (N_9772,N_3498,N_519);
nand U9773 (N_9773,N_3397,N_4625);
xor U9774 (N_9774,N_4276,N_1242);
nor U9775 (N_9775,N_172,N_1260);
or U9776 (N_9776,N_1063,N_3001);
xor U9777 (N_9777,N_3011,N_2731);
or U9778 (N_9778,N_4965,N_4799);
xnor U9779 (N_9779,N_1089,N_593);
or U9780 (N_9780,N_1466,N_650);
or U9781 (N_9781,N_2535,N_1802);
nor U9782 (N_9782,N_2291,N_3593);
xnor U9783 (N_9783,N_3857,N_1034);
xor U9784 (N_9784,N_1909,N_2148);
nor U9785 (N_9785,N_4257,N_1607);
or U9786 (N_9786,N_1146,N_2789);
nor U9787 (N_9787,N_318,N_3124);
xnor U9788 (N_9788,N_4810,N_3527);
nand U9789 (N_9789,N_1124,N_4287);
xnor U9790 (N_9790,N_2423,N_872);
nand U9791 (N_9791,N_2609,N_3082);
nor U9792 (N_9792,N_2841,N_4764);
nand U9793 (N_9793,N_2224,N_4548);
and U9794 (N_9794,N_773,N_2255);
and U9795 (N_9795,N_4921,N_4361);
xor U9796 (N_9796,N_2494,N_1839);
or U9797 (N_9797,N_773,N_4297);
nand U9798 (N_9798,N_2303,N_4841);
xor U9799 (N_9799,N_1163,N_2868);
nor U9800 (N_9800,N_657,N_2110);
and U9801 (N_9801,N_591,N_3930);
nor U9802 (N_9802,N_3017,N_698);
nor U9803 (N_9803,N_389,N_2242);
and U9804 (N_9804,N_2104,N_4069);
or U9805 (N_9805,N_2539,N_1342);
and U9806 (N_9806,N_199,N_1276);
nand U9807 (N_9807,N_3862,N_2208);
xor U9808 (N_9808,N_1209,N_1950);
nor U9809 (N_9809,N_4287,N_3222);
or U9810 (N_9810,N_2337,N_913);
or U9811 (N_9811,N_2303,N_4499);
nor U9812 (N_9812,N_3271,N_3760);
or U9813 (N_9813,N_4426,N_4412);
or U9814 (N_9814,N_3907,N_836);
nand U9815 (N_9815,N_2211,N_3673);
nor U9816 (N_9816,N_386,N_1572);
and U9817 (N_9817,N_4358,N_3356);
nor U9818 (N_9818,N_4122,N_557);
xnor U9819 (N_9819,N_1171,N_4772);
nor U9820 (N_9820,N_1828,N_178);
or U9821 (N_9821,N_2848,N_4829);
nor U9822 (N_9822,N_609,N_3496);
or U9823 (N_9823,N_1311,N_4657);
and U9824 (N_9824,N_4488,N_793);
nand U9825 (N_9825,N_4228,N_2837);
and U9826 (N_9826,N_3322,N_4067);
or U9827 (N_9827,N_4783,N_4656);
nor U9828 (N_9828,N_2290,N_3493);
or U9829 (N_9829,N_1247,N_1936);
and U9830 (N_9830,N_2655,N_3917);
xor U9831 (N_9831,N_475,N_2416);
or U9832 (N_9832,N_3466,N_303);
or U9833 (N_9833,N_1368,N_3087);
nor U9834 (N_9834,N_668,N_2881);
nor U9835 (N_9835,N_1011,N_837);
and U9836 (N_9836,N_596,N_3784);
or U9837 (N_9837,N_4394,N_3177);
xor U9838 (N_9838,N_2165,N_4076);
nor U9839 (N_9839,N_4031,N_2688);
xor U9840 (N_9840,N_3481,N_712);
xor U9841 (N_9841,N_4370,N_61);
or U9842 (N_9842,N_4107,N_4595);
nor U9843 (N_9843,N_4803,N_4981);
and U9844 (N_9844,N_1764,N_1717);
and U9845 (N_9845,N_3511,N_4158);
nor U9846 (N_9846,N_791,N_1207);
and U9847 (N_9847,N_3053,N_3526);
and U9848 (N_9848,N_384,N_2794);
or U9849 (N_9849,N_3874,N_2248);
nor U9850 (N_9850,N_176,N_4024);
or U9851 (N_9851,N_2887,N_4646);
nor U9852 (N_9852,N_297,N_2302);
nor U9853 (N_9853,N_4558,N_4865);
xnor U9854 (N_9854,N_2302,N_2913);
xnor U9855 (N_9855,N_2880,N_64);
or U9856 (N_9856,N_1729,N_188);
nand U9857 (N_9857,N_686,N_1524);
and U9858 (N_9858,N_1021,N_217);
or U9859 (N_9859,N_1887,N_2583);
xor U9860 (N_9860,N_1487,N_3015);
xnor U9861 (N_9861,N_2222,N_4483);
xnor U9862 (N_9862,N_1562,N_3460);
nor U9863 (N_9863,N_4657,N_613);
and U9864 (N_9864,N_3064,N_4792);
or U9865 (N_9865,N_4213,N_3723);
and U9866 (N_9866,N_815,N_691);
nor U9867 (N_9867,N_116,N_4659);
and U9868 (N_9868,N_3642,N_2125);
or U9869 (N_9869,N_2336,N_2878);
nor U9870 (N_9870,N_4220,N_2895);
xnor U9871 (N_9871,N_515,N_4978);
or U9872 (N_9872,N_1886,N_907);
xnor U9873 (N_9873,N_4897,N_4690);
nor U9874 (N_9874,N_24,N_826);
or U9875 (N_9875,N_2998,N_2592);
nor U9876 (N_9876,N_4053,N_2907);
xor U9877 (N_9877,N_2294,N_2188);
and U9878 (N_9878,N_4215,N_930);
or U9879 (N_9879,N_2828,N_372);
nand U9880 (N_9880,N_3225,N_4697);
nor U9881 (N_9881,N_4685,N_934);
nor U9882 (N_9882,N_15,N_145);
nand U9883 (N_9883,N_923,N_4056);
or U9884 (N_9884,N_3881,N_4543);
and U9885 (N_9885,N_3760,N_3362);
nand U9886 (N_9886,N_3321,N_1489);
xnor U9887 (N_9887,N_1426,N_2187);
nor U9888 (N_9888,N_4964,N_516);
or U9889 (N_9889,N_256,N_4550);
and U9890 (N_9890,N_483,N_77);
nand U9891 (N_9891,N_2690,N_2886);
and U9892 (N_9892,N_1253,N_495);
and U9893 (N_9893,N_4203,N_3395);
and U9894 (N_9894,N_1067,N_3984);
xor U9895 (N_9895,N_1858,N_4536);
and U9896 (N_9896,N_3894,N_4135);
or U9897 (N_9897,N_3461,N_1783);
and U9898 (N_9898,N_166,N_3841);
nand U9899 (N_9899,N_2501,N_4469);
nor U9900 (N_9900,N_4944,N_2252);
nand U9901 (N_9901,N_263,N_1928);
nor U9902 (N_9902,N_3768,N_2818);
or U9903 (N_9903,N_4150,N_3475);
xor U9904 (N_9904,N_4279,N_2642);
and U9905 (N_9905,N_1395,N_4456);
and U9906 (N_9906,N_996,N_4066);
nor U9907 (N_9907,N_1550,N_2430);
and U9908 (N_9908,N_636,N_3004);
or U9909 (N_9909,N_2194,N_1247);
nor U9910 (N_9910,N_3697,N_2041);
nor U9911 (N_9911,N_2732,N_391);
or U9912 (N_9912,N_374,N_1533);
and U9913 (N_9913,N_2632,N_914);
and U9914 (N_9914,N_2409,N_2415);
nand U9915 (N_9915,N_580,N_2167);
or U9916 (N_9916,N_237,N_3651);
or U9917 (N_9917,N_3146,N_1000);
and U9918 (N_9918,N_4916,N_2261);
nor U9919 (N_9919,N_274,N_4117);
nand U9920 (N_9920,N_2215,N_4053);
xnor U9921 (N_9921,N_1741,N_511);
or U9922 (N_9922,N_2069,N_1672);
nor U9923 (N_9923,N_1882,N_3605);
xnor U9924 (N_9924,N_3900,N_4272);
nand U9925 (N_9925,N_577,N_3539);
or U9926 (N_9926,N_3558,N_3197);
nand U9927 (N_9927,N_3108,N_3454);
or U9928 (N_9928,N_3716,N_1026);
or U9929 (N_9929,N_1436,N_414);
nand U9930 (N_9930,N_1284,N_3424);
nor U9931 (N_9931,N_4061,N_4045);
xnor U9932 (N_9932,N_1137,N_1431);
and U9933 (N_9933,N_4695,N_4704);
or U9934 (N_9934,N_673,N_3862);
xnor U9935 (N_9935,N_3887,N_2086);
nor U9936 (N_9936,N_4842,N_1471);
nor U9937 (N_9937,N_2405,N_1306);
or U9938 (N_9938,N_2265,N_3007);
nand U9939 (N_9939,N_125,N_2582);
xnor U9940 (N_9940,N_2730,N_2886);
xnor U9941 (N_9941,N_3963,N_538);
nand U9942 (N_9942,N_2420,N_4147);
xnor U9943 (N_9943,N_3232,N_3444);
and U9944 (N_9944,N_3460,N_1386);
xnor U9945 (N_9945,N_1772,N_615);
nand U9946 (N_9946,N_770,N_3096);
or U9947 (N_9947,N_1459,N_1635);
nor U9948 (N_9948,N_1407,N_3816);
or U9949 (N_9949,N_57,N_987);
nand U9950 (N_9950,N_2276,N_1165);
xnor U9951 (N_9951,N_3881,N_3780);
or U9952 (N_9952,N_1508,N_3660);
and U9953 (N_9953,N_4008,N_3452);
nand U9954 (N_9954,N_2587,N_2052);
nand U9955 (N_9955,N_1476,N_4262);
or U9956 (N_9956,N_2199,N_2172);
or U9957 (N_9957,N_2431,N_643);
or U9958 (N_9958,N_3348,N_3363);
nor U9959 (N_9959,N_2953,N_1079);
nand U9960 (N_9960,N_1253,N_677);
and U9961 (N_9961,N_3917,N_673);
xor U9962 (N_9962,N_4414,N_2359);
nor U9963 (N_9963,N_1540,N_4104);
and U9964 (N_9964,N_3794,N_3334);
xor U9965 (N_9965,N_4644,N_4378);
and U9966 (N_9966,N_4058,N_2165);
nand U9967 (N_9967,N_592,N_575);
nor U9968 (N_9968,N_2168,N_4884);
nand U9969 (N_9969,N_2251,N_1032);
nor U9970 (N_9970,N_1808,N_1625);
and U9971 (N_9971,N_1283,N_955);
and U9972 (N_9972,N_4078,N_720);
or U9973 (N_9973,N_20,N_1431);
nand U9974 (N_9974,N_2107,N_3604);
nor U9975 (N_9975,N_4340,N_1731);
or U9976 (N_9976,N_2800,N_1841);
or U9977 (N_9977,N_1083,N_1775);
nor U9978 (N_9978,N_33,N_2921);
or U9979 (N_9979,N_3248,N_1202);
and U9980 (N_9980,N_594,N_2537);
xnor U9981 (N_9981,N_1736,N_3787);
and U9982 (N_9982,N_991,N_3625);
nand U9983 (N_9983,N_3362,N_4173);
and U9984 (N_9984,N_1622,N_1873);
xnor U9985 (N_9985,N_2607,N_3100);
nor U9986 (N_9986,N_708,N_4196);
xnor U9987 (N_9987,N_3459,N_888);
nand U9988 (N_9988,N_2569,N_1217);
nor U9989 (N_9989,N_4553,N_3059);
nor U9990 (N_9990,N_3296,N_2378);
nor U9991 (N_9991,N_4236,N_1069);
xnor U9992 (N_9992,N_1966,N_3131);
nor U9993 (N_9993,N_857,N_447);
nor U9994 (N_9994,N_249,N_1884);
and U9995 (N_9995,N_3348,N_2679);
xor U9996 (N_9996,N_2038,N_2583);
xnor U9997 (N_9997,N_3000,N_3917);
and U9998 (N_9998,N_4663,N_72);
nand U9999 (N_9999,N_1525,N_4682);
and U10000 (N_10000,N_6203,N_8126);
nor U10001 (N_10001,N_6248,N_7561);
nor U10002 (N_10002,N_8202,N_8464);
nor U10003 (N_10003,N_8333,N_6014);
or U10004 (N_10004,N_6618,N_6988);
nand U10005 (N_10005,N_9260,N_6461);
xor U10006 (N_10006,N_5698,N_8011);
xor U10007 (N_10007,N_9710,N_9863);
nor U10008 (N_10008,N_8406,N_6929);
and U10009 (N_10009,N_7746,N_7801);
and U10010 (N_10010,N_5787,N_6730);
or U10011 (N_10011,N_5649,N_7444);
nor U10012 (N_10012,N_8878,N_9517);
nor U10013 (N_10013,N_5814,N_8695);
xor U10014 (N_10014,N_5143,N_9798);
and U10015 (N_10015,N_9227,N_8924);
nand U10016 (N_10016,N_7026,N_7550);
or U10017 (N_10017,N_6228,N_5511);
nor U10018 (N_10018,N_8873,N_6869);
nand U10019 (N_10019,N_5539,N_9459);
or U10020 (N_10020,N_8999,N_5528);
xnor U10021 (N_10021,N_7449,N_9480);
or U10022 (N_10022,N_6895,N_5777);
nor U10023 (N_10023,N_9874,N_5112);
nand U10024 (N_10024,N_6654,N_6061);
or U10025 (N_10025,N_5911,N_7773);
xnor U10026 (N_10026,N_9036,N_5750);
and U10027 (N_10027,N_8137,N_5653);
nor U10028 (N_10028,N_8714,N_6965);
nor U10029 (N_10029,N_7052,N_8972);
nand U10030 (N_10030,N_9443,N_7359);
or U10031 (N_10031,N_8483,N_9623);
xnor U10032 (N_10032,N_9085,N_9274);
or U10033 (N_10033,N_9921,N_5681);
nand U10034 (N_10034,N_8017,N_8396);
xor U10035 (N_10035,N_9140,N_9853);
nand U10036 (N_10036,N_6298,N_7689);
or U10037 (N_10037,N_5248,N_6712);
nor U10038 (N_10038,N_9157,N_5437);
nand U10039 (N_10039,N_8160,N_7518);
nand U10040 (N_10040,N_6714,N_8640);
xnor U10041 (N_10041,N_8095,N_7984);
or U10042 (N_10042,N_5860,N_8948);
nand U10043 (N_10043,N_9252,N_6900);
xnor U10044 (N_10044,N_9807,N_6257);
nor U10045 (N_10045,N_9888,N_6270);
or U10046 (N_10046,N_5493,N_7881);
nor U10047 (N_10047,N_8851,N_8470);
nand U10048 (N_10048,N_5565,N_9263);
nand U10049 (N_10049,N_9707,N_9027);
and U10050 (N_10050,N_7694,N_8225);
or U10051 (N_10051,N_9880,N_8284);
xnor U10052 (N_10052,N_7736,N_9005);
nor U10053 (N_10053,N_5224,N_6287);
and U10054 (N_10054,N_6790,N_9918);
nor U10055 (N_10055,N_8757,N_8957);
or U10056 (N_10056,N_7897,N_6375);
and U10057 (N_10057,N_8743,N_6097);
nor U10058 (N_10058,N_6514,N_5356);
nand U10059 (N_10059,N_9533,N_6453);
nand U10060 (N_10060,N_7265,N_9792);
xnor U10061 (N_10061,N_6944,N_9995);
nand U10062 (N_10062,N_5989,N_7584);
xor U10063 (N_10063,N_7218,N_6420);
and U10064 (N_10064,N_6671,N_8331);
nor U10065 (N_10065,N_6455,N_7139);
or U10066 (N_10066,N_7315,N_7662);
and U10067 (N_10067,N_6512,N_6362);
nand U10068 (N_10068,N_8986,N_7802);
nor U10069 (N_10069,N_6973,N_6488);
nor U10070 (N_10070,N_9300,N_7529);
nor U10071 (N_10071,N_8554,N_5587);
and U10072 (N_10072,N_9047,N_6577);
and U10073 (N_10073,N_8159,N_6625);
or U10074 (N_10074,N_6334,N_5991);
nor U10075 (N_10075,N_6767,N_7892);
nor U10076 (N_10076,N_7851,N_6725);
xnor U10077 (N_10077,N_9940,N_6414);
or U10078 (N_10078,N_8961,N_9887);
and U10079 (N_10079,N_9749,N_7551);
and U10080 (N_10080,N_5434,N_8089);
nand U10081 (N_10081,N_9708,N_9396);
xnor U10082 (N_10082,N_7304,N_9331);
nand U10083 (N_10083,N_6795,N_5669);
and U10084 (N_10084,N_5510,N_9923);
nand U10085 (N_10085,N_9595,N_8979);
nor U10086 (N_10086,N_8509,N_7752);
nand U10087 (N_10087,N_6152,N_9837);
or U10088 (N_10088,N_5870,N_6523);
xor U10089 (N_10089,N_8759,N_8492);
xnor U10090 (N_10090,N_6890,N_5223);
or U10091 (N_10091,N_5946,N_6893);
nand U10092 (N_10092,N_6506,N_8098);
or U10093 (N_10093,N_8270,N_9860);
nand U10094 (N_10094,N_5906,N_8609);
xnor U10095 (N_10095,N_8808,N_7691);
or U10096 (N_10096,N_9893,N_6398);
nand U10097 (N_10097,N_8591,N_6755);
or U10098 (N_10098,N_8477,N_6460);
or U10099 (N_10099,N_8033,N_9372);
and U10100 (N_10100,N_9366,N_8821);
and U10101 (N_10101,N_5430,N_7905);
nor U10102 (N_10102,N_7708,N_7739);
nand U10103 (N_10103,N_9123,N_8614);
nor U10104 (N_10104,N_7778,N_8970);
xnor U10105 (N_10105,N_7619,N_5772);
nor U10106 (N_10106,N_8361,N_5054);
nand U10107 (N_10107,N_8227,N_5426);
nand U10108 (N_10108,N_8858,N_6915);
nand U10109 (N_10109,N_6952,N_9230);
and U10110 (N_10110,N_8708,N_9993);
and U10111 (N_10111,N_7507,N_8579);
nor U10112 (N_10112,N_5109,N_9661);
xor U10113 (N_10113,N_8795,N_9314);
xor U10114 (N_10114,N_9079,N_9981);
and U10115 (N_10115,N_5723,N_5811);
or U10116 (N_10116,N_6439,N_9075);
or U10117 (N_10117,N_5280,N_6233);
or U10118 (N_10118,N_7781,N_6073);
xnor U10119 (N_10119,N_7384,N_7065);
and U10120 (N_10120,N_7213,N_5402);
xnor U10121 (N_10121,N_9838,N_9616);
nand U10122 (N_10122,N_7209,N_6210);
and U10123 (N_10123,N_8679,N_9135);
xnor U10124 (N_10124,N_7314,N_5775);
xor U10125 (N_10125,N_5214,N_7246);
and U10126 (N_10126,N_8032,N_8587);
nor U10127 (N_10127,N_8271,N_7625);
or U10128 (N_10128,N_8908,N_6080);
and U10129 (N_10129,N_8261,N_6614);
nand U10130 (N_10130,N_9392,N_7512);
and U10131 (N_10131,N_7942,N_5263);
or U10132 (N_10132,N_9345,N_8917);
xnor U10133 (N_10133,N_5862,N_5451);
and U10134 (N_10134,N_8001,N_9925);
or U10135 (N_10135,N_6074,N_8811);
nor U10136 (N_10136,N_9333,N_7981);
nand U10137 (N_10137,N_9769,N_5399);
nor U10138 (N_10138,N_6076,N_6591);
nand U10139 (N_10139,N_9060,N_6743);
or U10140 (N_10140,N_9698,N_5004);
nand U10141 (N_10141,N_6206,N_8845);
xor U10142 (N_10142,N_9412,N_5879);
nand U10143 (N_10143,N_6817,N_9729);
nand U10144 (N_10144,N_5216,N_6843);
xnor U10145 (N_10145,N_9719,N_9676);
or U10146 (N_10146,N_6813,N_9907);
xor U10147 (N_10147,N_7122,N_9960);
nor U10148 (N_10148,N_6505,N_6892);
or U10149 (N_10149,N_9321,N_8774);
xor U10150 (N_10150,N_6429,N_6150);
nor U10151 (N_10151,N_9267,N_5081);
nor U10152 (N_10152,N_6557,N_7903);
xor U10153 (N_10153,N_8481,N_6914);
xor U10154 (N_10154,N_6969,N_6905);
xnor U10155 (N_10155,N_9950,N_6217);
and U10156 (N_10156,N_7682,N_8253);
or U10157 (N_10157,N_5047,N_7254);
and U10158 (N_10158,N_7661,N_5377);
xnor U10159 (N_10159,N_7239,N_8930);
nor U10160 (N_10160,N_5741,N_5804);
nand U10161 (N_10161,N_6999,N_8398);
and U10162 (N_10162,N_7834,N_8728);
and U10163 (N_10163,N_5285,N_5984);
or U10164 (N_10164,N_8904,N_8628);
or U10165 (N_10165,N_7933,N_9695);
or U10166 (N_10166,N_6789,N_8560);
or U10167 (N_10167,N_7492,N_8316);
and U10168 (N_10168,N_9247,N_9696);
nor U10169 (N_10169,N_9814,N_5923);
xnor U10170 (N_10170,N_6432,N_5136);
xnor U10171 (N_10171,N_7135,N_9186);
and U10172 (N_10172,N_9813,N_6934);
and U10173 (N_10173,N_9091,N_5350);
nor U10174 (N_10174,N_9858,N_5190);
nand U10175 (N_10175,N_6943,N_8934);
and U10176 (N_10176,N_5931,N_8898);
or U10177 (N_10177,N_6612,N_5854);
nand U10178 (N_10178,N_9675,N_8019);
nor U10179 (N_10179,N_8935,N_6516);
nor U10180 (N_10180,N_6918,N_6205);
or U10181 (N_10181,N_8395,N_9919);
nand U10182 (N_10182,N_9354,N_6476);
nor U10183 (N_10183,N_8713,N_7402);
nor U10184 (N_10184,N_6631,N_7809);
nand U10185 (N_10185,N_8175,N_9532);
xnor U10186 (N_10186,N_7876,N_9519);
or U10187 (N_10187,N_5564,N_7210);
or U10188 (N_10188,N_9238,N_6531);
or U10189 (N_10189,N_7856,N_6345);
or U10190 (N_10190,N_6159,N_6397);
xnor U10191 (N_10191,N_5327,N_9967);
nand U10192 (N_10192,N_6665,N_5383);
xnor U10193 (N_10193,N_6288,N_7080);
or U10194 (N_10194,N_6953,N_5545);
and U10195 (N_10195,N_8684,N_8677);
nand U10196 (N_10196,N_9779,N_5781);
or U10197 (N_10197,N_9360,N_6197);
and U10198 (N_10198,N_6276,N_5494);
xor U10199 (N_10199,N_7282,N_6576);
nand U10200 (N_10200,N_6582,N_7362);
nor U10201 (N_10201,N_7760,N_8312);
or U10202 (N_10202,N_5160,N_6050);
xor U10203 (N_10203,N_8437,N_7249);
xnor U10204 (N_10204,N_9470,N_6481);
and U10205 (N_10205,N_8035,N_6387);
and U10206 (N_10206,N_5193,N_9545);
nand U10207 (N_10207,N_5287,N_9946);
and U10208 (N_10208,N_6682,N_6782);
or U10209 (N_10209,N_9100,N_6503);
xnor U10210 (N_10210,N_5941,N_7858);
nand U10211 (N_10211,N_9795,N_5101);
xor U10212 (N_10212,N_7496,N_7543);
nand U10213 (N_10213,N_9910,N_6381);
and U10214 (N_10214,N_5724,N_7458);
nand U10215 (N_10215,N_7462,N_6694);
nor U10216 (N_10216,N_7792,N_6449);
nand U10217 (N_10217,N_6143,N_5268);
and U10218 (N_10218,N_8540,N_8959);
nor U10219 (N_10219,N_9142,N_6799);
or U10220 (N_10220,N_9884,N_5291);
xor U10221 (N_10221,N_7953,N_9453);
xor U10222 (N_10222,N_6367,N_5255);
nor U10223 (N_10223,N_7436,N_8149);
and U10224 (N_10224,N_5466,N_9776);
nor U10225 (N_10225,N_5739,N_5914);
and U10226 (N_10226,N_9611,N_9662);
nor U10227 (N_10227,N_8615,N_6090);
and U10228 (N_10228,N_7889,N_7390);
nand U10229 (N_10229,N_9567,N_5512);
or U10230 (N_10230,N_8295,N_5122);
or U10231 (N_10231,N_8402,N_7419);
xor U10232 (N_10232,N_7959,N_5140);
nand U10233 (N_10233,N_7546,N_7335);
and U10234 (N_10234,N_9964,N_8324);
xnor U10235 (N_10235,N_6008,N_6685);
nor U10236 (N_10236,N_7750,N_8818);
or U10237 (N_10237,N_8231,N_8599);
nor U10238 (N_10238,N_6761,N_9515);
nand U10239 (N_10239,N_9777,N_8413);
nor U10240 (N_10240,N_6422,N_9020);
nand U10241 (N_10241,N_7958,N_9931);
and U10242 (N_10242,N_6489,N_8949);
and U10243 (N_10243,N_7755,N_6036);
nand U10244 (N_10244,N_7181,N_7464);
and U10245 (N_10245,N_7127,N_9098);
xor U10246 (N_10246,N_6332,N_5352);
nor U10247 (N_10247,N_5177,N_6348);
or U10248 (N_10248,N_6803,N_5533);
or U10249 (N_10249,N_6471,N_9117);
nand U10250 (N_10250,N_7114,N_6272);
and U10251 (N_10251,N_9229,N_5035);
and U10252 (N_10252,N_6964,N_5945);
nor U10253 (N_10253,N_9934,N_7311);
xor U10254 (N_10254,N_8860,N_8990);
nor U10255 (N_10255,N_6444,N_9574);
nor U10256 (N_10256,N_8163,N_7678);
and U10257 (N_10257,N_9589,N_8596);
nor U10258 (N_10258,N_5542,N_9996);
and U10259 (N_10259,N_7641,N_5876);
nand U10260 (N_10260,N_6095,N_8800);
xor U10261 (N_10261,N_5491,N_5992);
or U10262 (N_10262,N_7463,N_7993);
nor U10263 (N_10263,N_7544,N_5640);
nor U10264 (N_10264,N_7681,N_7130);
or U10265 (N_10265,N_6054,N_9320);
or U10266 (N_10266,N_9678,N_7124);
nor U10267 (N_10267,N_6148,N_5960);
or U10268 (N_10268,N_7805,N_9518);
and U10269 (N_10269,N_8381,N_6668);
nor U10270 (N_10270,N_5927,N_5784);
nor U10271 (N_10271,N_6509,N_6423);
xor U10272 (N_10272,N_5376,N_7638);
xor U10273 (N_10273,N_9865,N_5305);
nand U10274 (N_10274,N_9387,N_5389);
nand U10275 (N_10275,N_5387,N_7675);
or U10276 (N_10276,N_5676,N_8044);
nor U10277 (N_10277,N_5391,N_5487);
xnor U10278 (N_10278,N_9144,N_5056);
nand U10279 (N_10279,N_6294,N_7860);
nor U10280 (N_10280,N_9601,N_8134);
nand U10281 (N_10281,N_6924,N_6160);
nor U10282 (N_10282,N_5566,N_7669);
xor U10283 (N_10283,N_5887,N_6794);
or U10284 (N_10284,N_9531,N_5692);
and U10285 (N_10285,N_7298,N_9659);
or U10286 (N_10286,N_6747,N_5372);
and U10287 (N_10287,N_7278,N_8520);
and U10288 (N_10288,N_8584,N_6066);
nand U10289 (N_10289,N_9181,N_8450);
nand U10290 (N_10290,N_8940,N_7145);
or U10291 (N_10291,N_7407,N_5002);
and U10292 (N_10292,N_6847,N_6802);
or U10293 (N_10293,N_8519,N_9579);
xor U10294 (N_10294,N_5489,N_7457);
xnor U10295 (N_10295,N_8191,N_8275);
nor U10296 (N_10296,N_9861,N_6030);
nand U10297 (N_10297,N_9419,N_9906);
nand U10298 (N_10298,N_6570,N_7997);
or U10299 (N_10299,N_6251,N_5701);
or U10300 (N_10300,N_9492,N_9829);
xor U10301 (N_10301,N_9199,N_6109);
xor U10302 (N_10302,N_5294,N_6963);
or U10303 (N_10303,N_7872,N_9451);
nand U10304 (N_10304,N_7286,N_6114);
nor U10305 (N_10305,N_8418,N_6753);
xnor U10306 (N_10306,N_7144,N_9882);
nand U10307 (N_10307,N_7626,N_5668);
nand U10308 (N_10308,N_5475,N_9620);
xnor U10309 (N_10309,N_9179,N_7133);
xnor U10310 (N_10310,N_7799,N_5303);
xnor U10311 (N_10311,N_8844,N_9365);
xor U10312 (N_10312,N_5105,N_7992);
nor U10313 (N_10313,N_6209,N_9322);
and U10314 (N_10314,N_9872,N_6660);
nand U10315 (N_10315,N_7225,N_9954);
nor U10316 (N_10316,N_7814,N_5585);
nor U10317 (N_10317,N_8391,N_7508);
or U10318 (N_10318,N_6947,N_9415);
nor U10319 (N_10319,N_5218,N_6504);
nor U10320 (N_10320,N_8721,N_8829);
nor U10321 (N_10321,N_9767,N_9556);
or U10322 (N_10322,N_6039,N_6457);
nor U10323 (N_10323,N_8740,N_9414);
or U10324 (N_10324,N_9735,N_7058);
or U10325 (N_10325,N_6921,N_7164);
and U10326 (N_10326,N_5735,N_6325);
nand U10327 (N_10327,N_9163,N_6775);
or U10328 (N_10328,N_5357,N_6513);
nand U10329 (N_10329,N_8547,N_6472);
nor U10330 (N_10330,N_7329,N_9766);
and U10331 (N_10331,N_5265,N_5928);
xnor U10332 (N_10332,N_6780,N_7207);
nor U10333 (N_10333,N_7380,N_8238);
nor U10334 (N_10334,N_9422,N_9957);
nand U10335 (N_10335,N_5233,N_9189);
nor U10336 (N_10336,N_9525,N_6344);
and U10337 (N_10337,N_9466,N_6316);
nand U10338 (N_10338,N_5447,N_5791);
nand U10339 (N_10339,N_9430,N_9765);
nor U10340 (N_10340,N_9541,N_8248);
nand U10341 (N_10341,N_9210,N_7285);
xor U10342 (N_10342,N_5505,N_5410);
xnor U10343 (N_10343,N_6437,N_7924);
nor U10344 (N_10344,N_6385,N_5902);
nand U10345 (N_10345,N_7523,N_7715);
or U10346 (N_10346,N_6038,N_5824);
nor U10347 (N_10347,N_7623,N_7084);
xor U10348 (N_10348,N_9243,N_6163);
xnor U10349 (N_10349,N_8545,N_9512);
nand U10350 (N_10350,N_9702,N_9764);
nand U10351 (N_10351,N_9236,N_9001);
xor U10352 (N_10352,N_6335,N_6252);
nor U10353 (N_10353,N_6708,N_5604);
or U10354 (N_10354,N_6102,N_5881);
nand U10355 (N_10355,N_5625,N_6260);
and U10356 (N_10356,N_8621,N_8651);
xnor U10357 (N_10357,N_8265,N_8273);
nor U10358 (N_10358,N_6913,N_9019);
nor U10359 (N_10359,N_7979,N_7810);
nor U10360 (N_10360,N_5110,N_7969);
xnor U10361 (N_10361,N_6840,N_8296);
nor U10362 (N_10362,N_8931,N_8247);
or U10363 (N_10363,N_7852,N_8962);
or U10364 (N_10364,N_5253,N_6566);
or U10365 (N_10365,N_7838,N_8243);
or U10366 (N_10366,N_8896,N_7494);
or U10367 (N_10367,N_6604,N_8573);
or U10368 (N_10368,N_6555,N_9246);
nor U10369 (N_10369,N_6681,N_6589);
and U10370 (N_10370,N_8010,N_9832);
xor U10371 (N_10371,N_6907,N_5710);
and U10372 (N_10372,N_7790,N_9239);
xnor U10373 (N_10373,N_8868,N_7002);
and U10374 (N_10374,N_5012,N_7895);
nand U10375 (N_10375,N_6574,N_6154);
or U10376 (N_10376,N_6037,N_8981);
nor U10377 (N_10377,N_6010,N_7352);
or U10378 (N_10378,N_7046,N_7132);
xnor U10379 (N_10379,N_7393,N_7827);
or U10380 (N_10380,N_9277,N_7577);
nand U10381 (N_10381,N_6713,N_8392);
nand U10382 (N_10382,N_7977,N_9012);
xnor U10383 (N_10383,N_7811,N_6842);
xnor U10384 (N_10384,N_7261,N_7107);
and U10385 (N_10385,N_7535,N_9324);
or U10386 (N_10386,N_7610,N_7168);
or U10387 (N_10387,N_8143,N_6638);
or U10388 (N_10388,N_6527,N_7306);
or U10389 (N_10389,N_9706,N_5774);
nor U10390 (N_10390,N_5563,N_9418);
or U10391 (N_10391,N_7737,N_8498);
nor U10392 (N_10392,N_7845,N_8119);
nand U10393 (N_10393,N_6986,N_6897);
or U10394 (N_10394,N_8076,N_9894);
nor U10395 (N_10395,N_6408,N_9066);
or U10396 (N_10396,N_9619,N_8315);
or U10397 (N_10397,N_6331,N_6355);
nor U10398 (N_10398,N_8091,N_8796);
xnor U10399 (N_10399,N_8776,N_7121);
nor U10400 (N_10400,N_5022,N_6026);
nor U10401 (N_10401,N_5951,N_8195);
nand U10402 (N_10402,N_6166,N_6979);
or U10403 (N_10403,N_6369,N_7212);
nor U10404 (N_10404,N_5175,N_6278);
nor U10405 (N_10405,N_9849,N_7158);
and U10406 (N_10406,N_6827,N_6751);
nor U10407 (N_10407,N_9442,N_8720);
nor U10408 (N_10408,N_9737,N_8952);
nor U10409 (N_10409,N_6613,N_5599);
nor U10410 (N_10410,N_5773,N_8289);
nand U10411 (N_10411,N_5948,N_7795);
and U10412 (N_10412,N_7321,N_5152);
nor U10413 (N_10413,N_8342,N_6374);
and U10414 (N_10414,N_6139,N_7466);
nor U10415 (N_10415,N_5380,N_6891);
or U10416 (N_10416,N_8928,N_6884);
nand U10417 (N_10417,N_8699,N_9114);
and U10418 (N_10418,N_5544,N_9969);
or U10419 (N_10419,N_5456,N_7024);
and U10420 (N_10420,N_7461,N_8528);
nand U10421 (N_10421,N_8592,N_7732);
xnor U10422 (N_10422,N_6958,N_6939);
nor U10423 (N_10423,N_9353,N_7617);
or U10424 (N_10424,N_6974,N_8151);
or U10425 (N_10425,N_5379,N_9250);
nor U10426 (N_10426,N_6264,N_7653);
xnor U10427 (N_10427,N_7722,N_6018);
or U10428 (N_10428,N_9498,N_5815);
or U10429 (N_10429,N_7375,N_8964);
nor U10430 (N_10430,N_8777,N_5172);
nand U10431 (N_10431,N_9059,N_6350);
nand U10432 (N_10432,N_8881,N_8054);
and U10433 (N_10433,N_7235,N_7302);
or U10434 (N_10434,N_9602,N_7118);
xnor U10435 (N_10435,N_9680,N_8021);
and U10436 (N_10436,N_6399,N_9026);
nor U10437 (N_10437,N_9555,N_6838);
and U10438 (N_10438,N_7686,N_7408);
nand U10439 (N_10439,N_9118,N_9650);
or U10440 (N_10440,N_9069,N_7309);
and U10441 (N_10441,N_8337,N_5969);
and U10442 (N_10442,N_8320,N_8194);
xor U10443 (N_10443,N_7729,N_5219);
and U10444 (N_10444,N_5798,N_5188);
nor U10445 (N_10445,N_9063,N_5745);
or U10446 (N_10446,N_6550,N_8240);
or U10447 (N_10447,N_8394,N_7073);
and U10448 (N_10448,N_6722,N_9275);
or U10449 (N_10449,N_8114,N_7221);
or U10450 (N_10450,N_5716,N_5632);
or U10451 (N_10451,N_7774,N_5146);
nand U10452 (N_10452,N_6075,N_7763);
xnor U10453 (N_10453,N_9053,N_9130);
xnor U10454 (N_10454,N_6501,N_5994);
nand U10455 (N_10455,N_8988,N_8963);
xor U10456 (N_10456,N_9817,N_7287);
xor U10457 (N_10457,N_6729,N_6436);
and U10458 (N_10458,N_9024,N_9389);
nor U10459 (N_10459,N_8219,N_5976);
or U10460 (N_10460,N_7711,N_9987);
or U10461 (N_10461,N_9472,N_6519);
or U10462 (N_10462,N_7150,N_7602);
nor U10463 (N_10463,N_8830,N_6136);
nand U10464 (N_10464,N_8213,N_6749);
or U10465 (N_10465,N_5609,N_9639);
xnor U10466 (N_10466,N_6823,N_9337);
and U10467 (N_10467,N_7303,N_6330);
nand U10468 (N_10468,N_9298,N_9564);
and U10469 (N_10469,N_5405,N_6342);
xor U10470 (N_10470,N_8619,N_8132);
or U10471 (N_10471,N_6495,N_6368);
nand U10472 (N_10472,N_8729,N_7850);
xor U10473 (N_10473,N_7930,N_6889);
or U10474 (N_10474,N_8662,N_9883);
or U10475 (N_10475,N_6544,N_9788);
and U10476 (N_10476,N_9989,N_8526);
xnor U10477 (N_10477,N_5636,N_9093);
and U10478 (N_10478,N_9870,N_7070);
xor U10479 (N_10479,N_9568,N_8150);
nand U10480 (N_10480,N_6820,N_7477);
xnor U10481 (N_10481,N_5361,N_9688);
nor U10482 (N_10482,N_7651,N_5553);
or U10483 (N_10483,N_7358,N_7102);
nand U10484 (N_10484,N_9223,N_7049);
and U10485 (N_10485,N_5628,N_6565);
xnor U10486 (N_10486,N_6845,N_7497);
xnor U10487 (N_10487,N_5819,N_9618);
or U10488 (N_10488,N_8186,N_5334);
nor U10489 (N_10489,N_6882,N_7172);
xnor U10490 (N_10490,N_8086,N_5141);
and U10491 (N_10491,N_7009,N_7256);
nor U10492 (N_10492,N_9553,N_5232);
nand U10493 (N_10493,N_9222,N_8709);
nand U10494 (N_10494,N_8472,N_5316);
nor U10495 (N_10495,N_8521,N_8856);
or U10496 (N_10496,N_7332,N_6663);
or U10497 (N_10497,N_8926,N_6704);
and U10498 (N_10498,N_8070,N_7388);
or U10499 (N_10499,N_7775,N_8706);
xnor U10500 (N_10500,N_9203,N_5169);
and U10501 (N_10501,N_9625,N_9966);
or U10502 (N_10502,N_8081,N_7806);
nor U10503 (N_10503,N_5930,N_9850);
xnor U10504 (N_10504,N_5052,N_6189);
and U10505 (N_10505,N_7912,N_9032);
nor U10506 (N_10506,N_6617,N_9326);
nor U10507 (N_10507,N_6615,N_6868);
or U10508 (N_10508,N_9649,N_9171);
or U10509 (N_10509,N_5181,N_8358);
nor U10510 (N_10510,N_5418,N_9468);
nor U10511 (N_10511,N_6211,N_5973);
xnor U10512 (N_10512,N_9843,N_5850);
and U10513 (N_10513,N_5952,N_5807);
xnor U10514 (N_10514,N_8696,N_9065);
or U10515 (N_10515,N_8298,N_6942);
or U10516 (N_10516,N_7060,N_7989);
xnor U10517 (N_10517,N_6672,N_6475);
nand U10518 (N_10518,N_5166,N_6190);
xor U10519 (N_10519,N_6177,N_6563);
or U10520 (N_10520,N_5382,N_8008);
nor U10521 (N_10521,N_6232,N_9129);
xnor U10522 (N_10522,N_8744,N_7050);
nand U10523 (N_10523,N_8542,N_8200);
and U10524 (N_10524,N_8344,N_8003);
nand U10525 (N_10525,N_8672,N_8286);
and U10526 (N_10526,N_8326,N_9081);
nor U10527 (N_10527,N_7027,N_7945);
or U10528 (N_10528,N_9483,N_8386);
nor U10529 (N_10529,N_9428,N_8073);
or U10530 (N_10530,N_5220,N_7010);
xnor U10531 (N_10531,N_9319,N_5252);
nand U10532 (N_10532,N_9455,N_6901);
or U10533 (N_10533,N_6562,N_8837);
nand U10534 (N_10534,N_7898,N_7970);
or U10535 (N_10535,N_6490,N_6425);
xnor U10536 (N_10536,N_8383,N_5097);
nor U10537 (N_10537,N_7220,N_5856);
or U10538 (N_10538,N_8781,N_8550);
and U10539 (N_10539,N_6926,N_8690);
nor U10540 (N_10540,N_9244,N_9983);
nor U10541 (N_10541,N_5882,N_8890);
or U10542 (N_10542,N_6551,N_8182);
and U10543 (N_10543,N_5737,N_6434);
and U10544 (N_10544,N_9534,N_5579);
xor U10545 (N_10545,N_9701,N_8929);
and U10546 (N_10546,N_7326,N_6229);
nand U10547 (N_10547,N_7759,N_6534);
xor U10548 (N_10548,N_8042,N_5720);
nor U10549 (N_10549,N_6837,N_7170);
or U10550 (N_10550,N_6314,N_8434);
nor U10551 (N_10551,N_6226,N_5749);
xnor U10552 (N_10552,N_9693,N_8162);
nand U10553 (N_10553,N_7189,N_8511);
nor U10554 (N_10554,N_8185,N_5349);
and U10555 (N_10555,N_9824,N_9867);
nand U10556 (N_10556,N_8506,N_7267);
nor U10557 (N_10557,N_7453,N_8539);
xor U10558 (N_10558,N_7879,N_5568);
nand U10559 (N_10559,N_8115,N_8487);
nor U10560 (N_10560,N_9159,N_6435);
and U10561 (N_10561,N_6635,N_5032);
or U10562 (N_10562,N_8268,N_9770);
xnor U10563 (N_10563,N_7700,N_5453);
or U10564 (N_10564,N_8078,N_5445);
nor U10565 (N_10565,N_6029,N_5312);
xnor U10566 (N_10566,N_7500,N_5107);
nand U10567 (N_10567,N_7514,N_5179);
nor U10568 (N_10568,N_7893,N_6130);
nor U10569 (N_10569,N_8080,N_8495);
nor U10570 (N_10570,N_6880,N_5414);
nand U10571 (N_10571,N_7635,N_5757);
or U10572 (N_10572,N_9436,N_5550);
nor U10573 (N_10573,N_9092,N_8336);
nor U10574 (N_10574,N_5290,N_7428);
nor U10575 (N_10575,N_8339,N_5961);
xnor U10576 (N_10576,N_9138,N_9658);
xnor U10577 (N_10577,N_8120,N_7377);
or U10578 (N_10578,N_7126,N_8906);
and U10579 (N_10579,N_8180,N_9510);
or U10580 (N_10580,N_9963,N_9576);
nor U10581 (N_10581,N_8303,N_5726);
nand U10582 (N_10582,N_6923,N_9152);
and U10583 (N_10583,N_7202,N_8130);
and U10584 (N_10584,N_7016,N_9160);
nor U10585 (N_10585,N_7902,N_8401);
nor U10586 (N_10586,N_6839,N_7129);
and U10587 (N_10587,N_5892,N_9645);
xnor U10588 (N_10588,N_9635,N_5849);
and U10589 (N_10589,N_6581,N_6554);
nor U10590 (N_10590,N_7618,N_8892);
or U10591 (N_10591,N_5062,N_5159);
nor U10592 (N_10592,N_8864,N_8622);
xor U10593 (N_10593,N_5718,N_8364);
nor U10594 (N_10594,N_5988,N_6469);
nor U10595 (N_10595,N_5439,N_9221);
xnor U10596 (N_10596,N_8485,N_9057);
xnor U10597 (N_10597,N_6007,N_7075);
xnor U10598 (N_10598,N_7939,N_9477);
and U10599 (N_10599,N_9316,N_9232);
and U10600 (N_10600,N_6781,N_6225);
and U10601 (N_10601,N_9196,N_5603);
and U10602 (N_10602,N_7001,N_9871);
nor U10603 (N_10603,N_5957,N_5621);
nand U10604 (N_10604,N_9938,N_9476);
nand U10605 (N_10605,N_9040,N_9105);
xnor U10606 (N_10606,N_9962,N_5877);
xor U10607 (N_10607,N_6972,N_6904);
nor U10608 (N_10608,N_8482,N_8715);
xnor U10609 (N_10609,N_7644,N_6752);
nand U10610 (N_10610,N_6310,N_6874);
nand U10611 (N_10611,N_7859,N_8764);
or U10612 (N_10612,N_8531,N_6590);
and U10613 (N_10613,N_7855,N_8665);
nor U10614 (N_10614,N_9191,N_5693);
xnor U10615 (N_10615,N_8976,N_7908);
and U10616 (N_10616,N_8223,N_5407);
or U10617 (N_10617,N_5810,N_8474);
xnor U10618 (N_10618,N_8946,N_7968);
nand U10619 (N_10619,N_6289,N_9099);
or U10620 (N_10620,N_6140,N_8165);
xor U10621 (N_10621,N_7337,N_9329);
or U10622 (N_10622,N_8104,N_8356);
or U10623 (N_10623,N_7079,N_9381);
or U10624 (N_10624,N_5714,N_6001);
xor U10625 (N_10625,N_9304,N_8857);
nor U10626 (N_10626,N_9634,N_5435);
nor U10627 (N_10627,N_5488,N_8473);
nor U10628 (N_10628,N_8580,N_7068);
xnor U10629 (N_10629,N_8558,N_7655);
nor U10630 (N_10630,N_9150,N_8480);
or U10631 (N_10631,N_9254,N_6315);
nand U10632 (N_10632,N_7274,N_6311);
or U10633 (N_10633,N_8441,N_8711);
xor U10634 (N_10634,N_7308,N_7141);
or U10635 (N_10635,N_8431,N_9013);
and U10636 (N_10636,N_6156,N_5256);
or U10637 (N_10637,N_5011,N_7511);
xnor U10638 (N_10638,N_8887,N_7527);
and U10639 (N_10639,N_5027,N_5240);
and U10640 (N_10640,N_7777,N_5966);
and U10641 (N_10641,N_9755,N_5717);
xor U10642 (N_10642,N_7649,N_7100);
nor U10643 (N_10643,N_5178,N_5885);
nand U10644 (N_10644,N_5955,N_6022);
or U10645 (N_10645,N_6865,N_7331);
and U10646 (N_10646,N_8783,N_5345);
xor U10647 (N_10647,N_5574,N_6451);
xnor U10648 (N_10648,N_8772,N_9241);
xnor U10649 (N_10649,N_6982,N_7054);
xnor U10650 (N_10650,N_9043,N_9561);
nand U10651 (N_10651,N_7579,N_8748);
nor U10652 (N_10652,N_5129,N_5898);
nand U10653 (N_10653,N_9259,N_6520);
xor U10654 (N_10654,N_5520,N_6127);
and U10655 (N_10655,N_6473,N_5050);
or U10656 (N_10656,N_6376,N_8260);
and U10657 (N_10657,N_8282,N_5409);
nor U10658 (N_10658,N_6219,N_6677);
nand U10659 (N_10659,N_5838,N_9166);
nand U10660 (N_10660,N_8117,N_7825);
nand U10661 (N_10661,N_8912,N_9169);
xnor U10662 (N_10662,N_8751,N_9109);
and U10663 (N_10663,N_7648,N_9796);
or U10664 (N_10664,N_7340,N_6064);
or U10665 (N_10665,N_5215,N_6003);
nand U10666 (N_10666,N_7949,N_9432);
nor U10667 (N_10667,N_9313,N_8328);
xor U10668 (N_10668,N_8382,N_7187);
nand U10669 (N_10669,N_8886,N_6128);
and U10670 (N_10670,N_7350,N_5778);
or U10671 (N_10671,N_8832,N_5249);
and U10672 (N_10672,N_7467,N_7142);
xnor U10673 (N_10673,N_8734,N_6903);
nand U10674 (N_10674,N_7251,N_6100);
xor U10675 (N_10675,N_9575,N_9806);
nand U10676 (N_10676,N_9226,N_6249);
or U10677 (N_10677,N_7615,N_8467);
nor U10678 (N_10678,N_9056,N_9347);
nand U10679 (N_10679,N_6404,N_9738);
nand U10680 (N_10680,N_7117,N_7757);
xnor U10681 (N_10681,N_9790,N_7807);
nand U10682 (N_10682,N_8647,N_9640);
and U10683 (N_10683,N_7242,N_6881);
or U10684 (N_10684,N_9992,N_9523);
nor U10685 (N_10685,N_8214,N_9580);
nand U10686 (N_10686,N_7573,N_5163);
or U10687 (N_10687,N_8387,N_6807);
nor U10688 (N_10688,N_7833,N_5353);
or U10689 (N_10689,N_5483,N_5229);
nor U10690 (N_10690,N_7808,N_5119);
xor U10691 (N_10691,N_7784,N_8034);
nor U10692 (N_10692,N_5206,N_8861);
xor U10693 (N_10693,N_5589,N_7726);
xnor U10694 (N_10694,N_6906,N_7656);
nand U10695 (N_10695,N_7772,N_8673);
xor U10696 (N_10696,N_9070,N_9201);
nor U10697 (N_10697,N_9198,N_9953);
or U10698 (N_10698,N_5910,N_6624);
nor U10699 (N_10699,N_8155,N_8533);
or U10700 (N_10700,N_6588,N_5597);
and U10701 (N_10701,N_7112,N_5863);
xnor U10702 (N_10702,N_6950,N_6797);
nand U10703 (N_10703,N_7671,N_9615);
xnor U10704 (N_10704,N_9692,N_5051);
nor U10705 (N_10705,N_5534,N_8608);
xnor U10706 (N_10706,N_7751,N_9317);
or U10707 (N_10707,N_5421,N_8779);
nor U10708 (N_10708,N_9890,N_7109);
or U10709 (N_10709,N_5884,N_5748);
or U10710 (N_10710,N_9539,N_7575);
xor U10711 (N_10711,N_9335,N_6960);
or U10712 (N_10712,N_6370,N_6482);
nand U10713 (N_10713,N_7247,N_9375);
xnor U10714 (N_10714,N_6357,N_6405);
or U10715 (N_10715,N_7951,N_6186);
or U10716 (N_10716,N_9131,N_6221);
and U10717 (N_10717,N_7421,N_9301);
or U10718 (N_10718,N_6057,N_9978);
nand U10719 (N_10719,N_5087,N_8502);
nand U10720 (N_10720,N_5161,N_7175);
or U10721 (N_10721,N_6517,N_5010);
and U10722 (N_10722,N_7698,N_7670);
and U10723 (N_10723,N_7647,N_9281);
nand U10724 (N_10724,N_8043,N_9679);
xor U10725 (N_10725,N_5629,N_5576);
and U10726 (N_10726,N_7947,N_8604);
nand U10727 (N_10727,N_6785,N_6502);
xor U10728 (N_10728,N_5595,N_8183);
nor U10729 (N_10729,N_5654,N_5046);
nor U10730 (N_10730,N_7157,N_6157);
and U10731 (N_10731,N_7280,N_5733);
xor U10732 (N_10732,N_5438,N_7515);
or U10733 (N_10733,N_8201,N_8718);
nand U10734 (N_10734,N_9721,N_6059);
nand U10735 (N_10735,N_7622,N_7025);
and U10736 (N_10736,N_6546,N_9791);
and U10737 (N_10737,N_5156,N_6745);
nand U10738 (N_10738,N_7316,N_8913);
nand U10739 (N_10739,N_6430,N_7899);
nand U10740 (N_10740,N_7474,N_9450);
nor U10741 (N_10741,N_9905,N_8343);
xor U10742 (N_10742,N_8835,N_8793);
or U10743 (N_10743,N_7580,N_8206);
and U10744 (N_10744,N_8843,N_7232);
and U10745 (N_10745,N_8379,N_8925);
nor U10746 (N_10746,N_5947,N_5874);
nor U10747 (N_10747,N_9760,N_7273);
nand U10748 (N_10748,N_7151,N_5921);
and U10749 (N_10749,N_8146,N_7849);
xor U10750 (N_10750,N_7988,N_8824);
xnor U10751 (N_10751,N_9374,N_8637);
or U10752 (N_10752,N_8293,N_7926);
or U10753 (N_10753,N_7679,N_6170);
nor U10754 (N_10754,N_6935,N_5731);
or U10755 (N_10755,N_7843,N_5425);
nand U10756 (N_10756,N_5446,N_9599);
nor U10757 (N_10757,N_7472,N_8172);
and U10758 (N_10758,N_6698,N_8079);
or U10759 (N_10759,N_6680,N_6549);
or U10760 (N_10760,N_8576,N_5970);
xor U10761 (N_10761,N_5066,N_6858);
and U10762 (N_10762,N_7702,N_8850);
or U10763 (N_10763,N_8735,N_6237);
nand U10764 (N_10764,N_7103,N_6771);
nor U10765 (N_10765,N_7931,N_6770);
and U10766 (N_10766,N_6991,N_7513);
nor U10767 (N_10767,N_5531,N_5663);
nor U10768 (N_10768,N_9642,N_5170);
nand U10769 (N_10769,N_8582,N_8249);
or U10770 (N_10770,N_9452,N_5744);
nor U10771 (N_10771,N_6231,N_8258);
nor U10772 (N_10772,N_8517,N_6125);
xnor U10773 (N_10773,N_7768,N_7720);
xnor U10774 (N_10774,N_7620,N_5131);
or U10775 (N_10775,N_8006,N_9786);
or U10776 (N_10776,N_6002,N_6732);
nand U10777 (N_10777,N_5825,N_8313);
nor U10778 (N_10778,N_5106,N_7263);
and U10779 (N_10779,N_7687,N_7299);
and U10780 (N_10780,N_8152,N_8691);
xor U10781 (N_10781,N_9089,N_6220);
nor U10782 (N_10782,N_8507,N_7608);
nor U10783 (N_10783,N_7536,N_7520);
nand U10784 (N_10784,N_5326,N_5673);
nor U10785 (N_10785,N_6149,N_7487);
nor U10786 (N_10786,N_6898,N_9929);
nand U10787 (N_10787,N_7987,N_7290);
or U10788 (N_10788,N_7381,N_9608);
or U10789 (N_10789,N_5571,N_7704);
or U10790 (N_10790,N_8967,N_9280);
or U10791 (N_10791,N_5315,N_9578);
xnor U10792 (N_10792,N_9393,N_9127);
xnor U10793 (N_10793,N_9286,N_9988);
nand U10794 (N_10794,N_6746,N_8330);
xnor U10795 (N_10795,N_8047,N_8977);
or U10796 (N_10796,N_8118,N_7222);
or U10797 (N_10797,N_7666,N_5462);
xor U10798 (N_10798,N_5789,N_6360);
or U10799 (N_10799,N_5959,N_7611);
and U10800 (N_10800,N_6641,N_9058);
nor U10801 (N_10801,N_7006,N_7171);
and U10802 (N_10802,N_8508,N_6639);
or U10803 (N_10803,N_5443,N_9783);
and U10804 (N_10804,N_9610,N_7946);
xor U10805 (N_10805,N_5920,N_8681);
nand U10806 (N_10806,N_8668,N_6980);
or U10807 (N_10807,N_6303,N_9581);
or U10808 (N_10808,N_5795,N_5697);
nand U10809 (N_10809,N_9341,N_9664);
and U10810 (N_10810,N_5580,N_7727);
and U10811 (N_10811,N_8422,N_8697);
xor U10812 (N_10812,N_6968,N_7560);
xor U10813 (N_10813,N_5638,N_9268);
nor U10814 (N_10814,N_5554,N_7983);
nor U10815 (N_10815,N_8648,N_7243);
and U10816 (N_10816,N_7627,N_9306);
nand U10817 (N_10817,N_7660,N_5937);
nand U10818 (N_10818,N_9543,N_6793);
nand U10819 (N_10819,N_5467,N_5711);
and U10820 (N_10820,N_7643,N_9147);
nor U10821 (N_10821,N_9302,N_7713);
nor U10822 (N_10822,N_7252,N_6967);
or U10823 (N_10823,N_7250,N_6951);
nand U10824 (N_10824,N_8397,N_6162);
and U10825 (N_10825,N_5238,N_8670);
nor U10826 (N_10826,N_7753,N_6676);
or U10827 (N_10827,N_6280,N_9303);
nand U10828 (N_10828,N_6961,N_7771);
or U10829 (N_10829,N_8574,N_7307);
or U10830 (N_10830,N_9376,N_8083);
nor U10831 (N_10831,N_8525,N_5005);
nand U10832 (N_10832,N_5076,N_6811);
and U10833 (N_10833,N_8785,N_6135);
xnor U10834 (N_10834,N_9318,N_8128);
and U10835 (N_10835,N_7780,N_7980);
and U10836 (N_10836,N_9828,N_7389);
nand U10837 (N_10837,N_7676,N_8625);
and U10838 (N_10838,N_5828,N_7005);
xor U10839 (N_10839,N_6928,N_5208);
xnor U10840 (N_10840,N_6017,N_5540);
or U10841 (N_10841,N_8833,N_8605);
xor U10842 (N_10842,N_7837,N_9809);
nand U10843 (N_10843,N_8354,N_5647);
nand U10844 (N_10844,N_7839,N_9577);
and U10845 (N_10845,N_5644,N_8476);
nand U10846 (N_10846,N_8319,N_8203);
or U10847 (N_10847,N_6199,N_8263);
and U10848 (N_10848,N_8488,N_6180);
xnor U10849 (N_10849,N_8762,N_6620);
nor U10850 (N_10850,N_7224,N_6327);
nand U10851 (N_10851,N_5611,N_5982);
nor U10852 (N_10852,N_8110,N_6552);
xnor U10853 (N_10853,N_7938,N_7099);
or U10854 (N_10854,N_9473,N_9522);
and U10855 (N_10855,N_5818,N_7556);
and U10856 (N_10856,N_7257,N_5461);
xnor U10857 (N_10857,N_7416,N_6716);
and U10858 (N_10858,N_8329,N_7909);
and U10859 (N_10859,N_5396,N_5029);
nand U10860 (N_10860,N_6726,N_7363);
and U10861 (N_10861,N_5369,N_9039);
xnor U10862 (N_10862,N_9563,N_5788);
xnor U10863 (N_10863,N_9656,N_6670);
nand U10864 (N_10864,N_9461,N_5917);
and U10865 (N_10865,N_6353,N_8932);
and U10866 (N_10866,N_8029,N_7258);
nor U10867 (N_10867,N_8633,N_6372);
or U10868 (N_10868,N_8301,N_8875);
and U10869 (N_10869,N_9416,N_7517);
nor U10870 (N_10870,N_6389,N_8566);
nor U10871 (N_10871,N_8568,N_6695);
or U10872 (N_10872,N_6748,N_5643);
nor U10873 (N_10873,N_5670,N_8433);
nand U10874 (N_10874,N_9370,N_7818);
xor U10875 (N_10875,N_7519,N_8973);
xnor U10876 (N_10876,N_8366,N_5168);
nand U10877 (N_10877,N_6684,N_5513);
nand U10878 (N_10878,N_5230,N_6533);
or U10879 (N_10879,N_6479,N_8951);
or U10880 (N_10880,N_6312,N_7160);
nand U10881 (N_10881,N_6706,N_6564);
xnor U10882 (N_10882,N_7495,N_7219);
xnor U10883 (N_10883,N_9740,N_6886);
xor U10884 (N_10884,N_9622,N_9185);
and U10885 (N_10885,N_9819,N_5038);
xnor U10886 (N_10886,N_5978,N_5707);
nand U10887 (N_10887,N_7932,N_8048);
nor U10888 (N_10888,N_6224,N_8230);
nor U10889 (N_10889,N_7343,N_7628);
nand U10890 (N_10890,N_5064,N_9355);
xor U10891 (N_10891,N_9050,N_8613);
and U10892 (N_10892,N_8514,N_9090);
nor U10893 (N_10893,N_7654,N_9956);
nand U10894 (N_10894,N_5138,N_6025);
nor U10895 (N_10895,N_5043,N_7712);
nor U10896 (N_10896,N_8516,N_6833);
nor U10897 (N_10897,N_7297,N_5061);
or U10898 (N_10898,N_5135,N_5806);
nor U10899 (N_10899,N_6738,N_9899);
xnor U10900 (N_10900,N_5217,N_5460);
and U10901 (N_10901,N_6402,N_5840);
nand U10902 (N_10902,N_8463,N_8572);
nand U10903 (N_10903,N_9052,N_9279);
or U10904 (N_10904,N_7521,N_6593);
nor U10905 (N_10905,N_5333,N_7510);
or U10906 (N_10906,N_5114,N_8819);
nor U10907 (N_10907,N_6521,N_8466);
xor U10908 (N_10908,N_9346,N_8885);
xor U10909 (N_10909,N_6134,N_7430);
or U10910 (N_10910,N_5600,N_6822);
nor U10911 (N_10911,N_5411,N_7501);
xnor U10912 (N_10912,N_6111,N_7357);
xnor U10913 (N_10913,N_9624,N_8812);
xor U10914 (N_10914,N_7873,N_7169);
and U10915 (N_10915,N_8166,N_7403);
or U10916 (N_10916,N_5419,N_9889);
and U10917 (N_10917,N_6318,N_7067);
and U10918 (N_10918,N_6441,N_8874);
nor U10919 (N_10919,N_7057,N_7074);
and U10920 (N_10920,N_7910,N_8384);
nor U10921 (N_10921,N_7714,N_7578);
or U10922 (N_10922,N_6734,N_5269);
and U10923 (N_10923,N_7347,N_5696);
and U10924 (N_10924,N_5412,N_9216);
nand U10925 (N_10925,N_5675,N_5167);
or U10926 (N_10926,N_8232,N_9061);
nor U10927 (N_10927,N_8399,N_9514);
nor U10928 (N_10928,N_9031,N_6529);
nor U10929 (N_10929,N_7361,N_9491);
nor U10930 (N_10930,N_9739,N_6486);
nand U10931 (N_10931,N_6082,N_9405);
nand U10932 (N_10932,N_5627,N_5365);
and U10933 (N_10933,N_6333,N_7078);
nor U10934 (N_10934,N_7667,N_9666);
or U10935 (N_10935,N_9305,N_7204);
or U10936 (N_10936,N_5059,N_7441);
and U10937 (N_10937,N_5180,N_5492);
xnor U10938 (N_10938,N_9744,N_7123);
and U10939 (N_10939,N_5134,N_6540);
nand U10940 (N_10940,N_7206,N_5995);
nor U10941 (N_10941,N_9951,N_6167);
nor U10942 (N_10942,N_9276,N_8915);
nand U10943 (N_10943,N_9465,N_9038);
nand U10944 (N_10944,N_8869,N_6300);
nand U10945 (N_10945,N_9003,N_6442);
and U10946 (N_10946,N_5057,N_6971);
and U10947 (N_10947,N_5536,N_9248);
or U10948 (N_10948,N_5331,N_7966);
xor U10949 (N_10949,N_7935,N_8283);
nor U10950 (N_10950,N_6710,N_9175);
and U10951 (N_10951,N_8737,N_7925);
and U10952 (N_10952,N_8920,N_9023);
and U10953 (N_10953,N_8277,N_9891);
and U10954 (N_10954,N_9839,N_8512);
nand U10955 (N_10955,N_9509,N_5987);
nand U10956 (N_10956,N_9486,N_7216);
nor U10957 (N_10957,N_7592,N_5348);
xor U10958 (N_10958,N_9629,N_8601);
or U10959 (N_10959,N_5040,N_5276);
nor U10960 (N_10960,N_8046,N_7423);
and U10961 (N_10961,N_7526,N_9445);
nor U10962 (N_10962,N_6027,N_7554);
or U10963 (N_10963,N_9399,N_7813);
xnor U10964 (N_10964,N_5635,N_5783);
nor U10965 (N_10965,N_7226,N_6996);
nand U10966 (N_10966,N_8357,N_5104);
nand U10967 (N_10967,N_9357,N_7391);
or U10968 (N_10968,N_5477,N_8955);
xor U10969 (N_10969,N_8109,N_9261);
xnor U10970 (N_10970,N_9562,N_8061);
and U10971 (N_10971,N_8365,N_9048);
xnor U10972 (N_10972,N_7417,N_9854);
nor U10973 (N_10973,N_6678,N_6171);
and U10974 (N_10974,N_7197,N_6826);
and U10975 (N_10975,N_8376,N_7740);
nor U10976 (N_10976,N_9750,N_9985);
nand U10977 (N_10977,N_6878,N_6737);
and U10978 (N_10978,N_8769,N_5728);
nand U10979 (N_10979,N_6772,N_5709);
nor U10980 (N_10980,N_9524,N_8352);
xor U10981 (N_10981,N_6261,N_9778);
nor U10982 (N_10982,N_5763,N_8636);
nor U10983 (N_10983,N_8421,N_7438);
xnor U10984 (N_10984,N_6699,N_9590);
nor U10985 (N_10985,N_8650,N_6305);
nand U10986 (N_10986,N_6867,N_9536);
or U10987 (N_10987,N_9251,N_5154);
nor U10988 (N_10988,N_8009,N_9294);
xnor U10989 (N_10989,N_8902,N_8411);
nor U10990 (N_10990,N_9605,N_9000);
or U10991 (N_10991,N_8116,N_6198);
xor U10992 (N_10992,N_7087,N_9288);
nor U10993 (N_10993,N_5820,N_8020);
or U10994 (N_10994,N_9896,N_8716);
nor U10995 (N_10995,N_5626,N_7113);
and U10996 (N_10996,N_8363,N_7048);
and U10997 (N_10997,N_8755,N_7334);
or U10998 (N_10998,N_8235,N_7410);
nand U10999 (N_10999,N_7435,N_8405);
or U11000 (N_11000,N_9165,N_8106);
nor U11001 (N_11001,N_7880,N_9295);
nand U11002 (N_11002,N_8746,N_7767);
xor U11003 (N_11003,N_7665,N_7883);
or U11004 (N_11004,N_5853,N_7528);
nand U11005 (N_11005,N_7155,N_7323);
xnor U11006 (N_11006,N_5834,N_7125);
xnor U11007 (N_11007,N_5337,N_8028);
nor U11008 (N_11008,N_9511,N_5126);
nor U11009 (N_11009,N_6126,N_7223);
xnor U11010 (N_11010,N_8251,N_6493);
nand U11011 (N_11011,N_5441,N_9460);
or U11012 (N_11012,N_7844,N_7104);
nor U11013 (N_11013,N_7033,N_5659);
xor U11014 (N_11014,N_7835,N_7066);
xnor U11015 (N_11015,N_5296,N_6689);
or U11016 (N_11016,N_9644,N_9868);
xor U11017 (N_11017,N_5705,N_8088);
and U11018 (N_11018,N_6883,N_6196);
nand U11019 (N_11019,N_9566,N_7812);
xnor U11020 (N_11020,N_5759,N_9034);
and U11021 (N_11021,N_8719,N_8978);
and U11022 (N_11022,N_6524,N_8188);
or U11023 (N_11023,N_7245,N_6596);
nand U11024 (N_11024,N_5678,N_5164);
nand U11025 (N_11025,N_5373,N_9187);
xor U11026 (N_11026,N_8209,N_7919);
xor U11027 (N_11027,N_6659,N_6424);
nor U11028 (N_11028,N_9002,N_7995);
or U11029 (N_11029,N_7820,N_9213);
and U11030 (N_11030,N_6783,N_7174);
or U11031 (N_11031,N_8618,N_9731);
or U11032 (N_11032,N_5527,N_5416);
nand U11033 (N_11033,N_8798,N_5351);
nand U11034 (N_11034,N_9781,N_7096);
and U11035 (N_11035,N_9875,N_8589);
and U11036 (N_11036,N_7652,N_9774);
nand U11037 (N_11037,N_6652,N_7884);
or U11038 (N_11038,N_9759,N_5529);
xnor U11039 (N_11039,N_9836,N_7601);
nor U11040 (N_11040,N_9475,N_9864);
or U11041 (N_11041,N_7769,N_6019);
or U11042 (N_11042,N_9339,N_9811);
and U11043 (N_11043,N_8646,N_9386);
nor U11044 (N_11044,N_8055,N_5762);
xnor U11045 (N_11045,N_9840,N_6144);
xnor U11046 (N_11046,N_5321,N_8026);
or U11047 (N_11047,N_9030,N_7131);
nor U11048 (N_11048,N_9433,N_8415);
xor U11049 (N_11049,N_5650,N_8606);
nor U11050 (N_11050,N_5656,N_5346);
xnor U11051 (N_11051,N_7531,N_9217);
or U11052 (N_11052,N_6995,N_8077);
nand U11053 (N_11053,N_7558,N_6306);
nand U11054 (N_11054,N_9398,N_9018);
nor U11055 (N_11055,N_8168,N_9377);
or U11056 (N_11056,N_9587,N_8069);
xnor U11057 (N_11057,N_6079,N_5080);
and U11058 (N_11058,N_9877,N_8578);
and U11059 (N_11059,N_9984,N_7392);
xor U11060 (N_11060,N_8094,N_6788);
or U11061 (N_11061,N_9920,N_9560);
xor U11062 (N_11062,N_5524,N_7178);
nand U11063 (N_11063,N_8002,N_7193);
xor U11064 (N_11064,N_8880,N_8290);
nor U11065 (N_11065,N_5023,N_9273);
nor U11066 (N_11066,N_9192,N_8585);
xnor U11067 (N_11067,N_9421,N_8780);
or U11068 (N_11068,N_5821,N_6151);
and U11069 (N_11069,N_5974,N_7976);
and U11070 (N_11070,N_8448,N_9308);
nor U11071 (N_11071,N_5187,N_9818);
nor U11072 (N_11072,N_9609,N_7485);
and U11073 (N_11073,N_6428,N_7624);
or U11074 (N_11074,N_7059,N_8947);
nand U11075 (N_11075,N_8666,N_9961);
and U11076 (N_11076,N_5281,N_6941);
nand U11077 (N_11077,N_5896,N_9037);
nor U11078 (N_11078,N_8139,N_8870);
xor U11079 (N_11079,N_6110,N_9833);
xor U11080 (N_11080,N_7688,N_8423);
or U11081 (N_11081,N_5257,N_6661);
xnor U11082 (N_11082,N_9080,N_9686);
or U11083 (N_11083,N_8562,N_6443);
nand U11084 (N_11084,N_9797,N_5144);
or U11085 (N_11085,N_6587,N_5044);
and U11086 (N_11086,N_8649,N_9200);
and U11087 (N_11087,N_6688,N_7030);
and U11088 (N_11088,N_8754,N_6966);
nor U11089 (N_11089,N_6319,N_5127);
nand U11090 (N_11090,N_5413,N_6409);
nor U11091 (N_11091,N_8192,N_7022);
nor U11092 (N_11092,N_8752,N_9126);
xor U11093 (N_11093,N_7015,N_9369);
xnor U11094 (N_11094,N_6121,N_5588);
xor U11095 (N_11095,N_8439,N_6108);
and U11096 (N_11096,N_6778,N_6766);
nor U11097 (N_11097,N_9336,N_6719);
nor U11098 (N_11098,N_5171,N_5145);
or U11099 (N_11099,N_7043,N_6997);
nor U11100 (N_11100,N_6742,N_9952);
xor U11101 (N_11101,N_7596,N_5324);
or U11102 (N_11102,N_7208,N_7998);
nand U11103 (N_11103,N_8359,N_8565);
or U11104 (N_11104,N_9694,N_6352);
or U11105 (N_11105,N_8982,N_9846);
nand U11106 (N_11106,N_5388,N_9170);
and U11107 (N_11107,N_7031,N_9042);
or U11108 (N_11108,N_6086,N_6118);
xnor U11109 (N_11109,N_6138,N_8635);
nand U11110 (N_11110,N_7229,N_6798);
nor U11111 (N_11111,N_6132,N_5746);
nand U11112 (N_11112,N_5031,N_8465);
or U11113 (N_11113,N_9311,N_7532);
xor U11114 (N_11114,N_7488,N_7398);
xor U11115 (N_11115,N_7327,N_6055);
nand U11116 (N_11116,N_9782,N_6718);
and U11117 (N_11117,N_6356,N_6829);
nor U11118 (N_11118,N_8414,N_9497);
or U11119 (N_11119,N_5001,N_8127);
and U11120 (N_11120,N_7971,N_6020);
nor U11121 (N_11121,N_8987,N_6285);
nand U11122 (N_11122,N_9011,N_8491);
or U11123 (N_11123,N_8943,N_9773);
xnor U11124 (N_11124,N_9939,N_9916);
xor U11125 (N_11125,N_8831,N_7716);
nand U11126 (N_11126,N_6917,N_5436);
or U11127 (N_11127,N_5194,N_5120);
and U11128 (N_11128,N_8288,N_8058);
nor U11129 (N_11129,N_7957,N_6247);
xor U11130 (N_11130,N_8332,N_7183);
nor U11131 (N_11131,N_8996,N_5715);
nor U11132 (N_11132,N_7236,N_7539);
or U11133 (N_11133,N_6611,N_8872);
or U11134 (N_11134,N_6392,N_8794);
or U11135 (N_11135,N_7480,N_7325);
nor U11136 (N_11136,N_5295,N_8778);
nor U11137 (N_11137,N_7963,N_8905);
or U11138 (N_11138,N_8440,N_5342);
nor U11139 (N_11139,N_5090,N_5964);
or U11140 (N_11140,N_5859,N_8760);
xnor U11141 (N_11141,N_6948,N_6637);
and U11142 (N_11142,N_6200,N_7629);
nor U11143 (N_11143,N_5393,N_7961);
and U11144 (N_11144,N_7349,N_8535);
xnor U11145 (N_11145,N_9293,N_5189);
nand U11146 (N_11146,N_5234,N_7277);
nor U11147 (N_11147,N_9559,N_6131);
xor U11148 (N_11148,N_7344,N_8541);
and U11149 (N_11149,N_7724,N_6366);
nor U11150 (N_11150,N_9033,N_9633);
or U11151 (N_11151,N_8135,N_6263);
or U11152 (N_11152,N_7846,N_6015);
and U11153 (N_11153,N_6223,N_6879);
xor U11154 (N_11154,N_9958,N_5476);
and U11155 (N_11155,N_6407,N_5808);
nor U11156 (N_11156,N_5463,N_5197);
xor U11157 (N_11157,N_7305,N_5086);
nand U11158 (N_11158,N_5761,N_9586);
nand U11159 (N_11159,N_5118,N_7581);
nand U11160 (N_11160,N_6619,N_8167);
and U11161 (N_11161,N_6908,N_8210);
xor U11162 (N_11162,N_9426,N_5612);
or U11163 (N_11163,N_8971,N_5366);
nor U11164 (N_11164,N_6078,N_7706);
nand U11165 (N_11165,N_6494,N_6478);
nand U11166 (N_11166,N_9852,N_8660);
and U11167 (N_11167,N_5325,N_6246);
or U11168 (N_11168,N_7685,N_6433);
and U11169 (N_11169,N_6235,N_5271);
nand U11170 (N_11170,N_8763,N_6459);
nand U11171 (N_11171,N_7861,N_8189);
and U11172 (N_11172,N_7659,N_8322);
or U11173 (N_11173,N_9804,N_5738);
nor U11174 (N_11174,N_5690,N_8598);
or U11175 (N_11175,N_9438,N_7385);
and U11176 (N_11176,N_6341,N_6584);
nor U11177 (N_11177,N_5962,N_8307);
xnor U11178 (N_11178,N_9115,N_8369);
or U11179 (N_11179,N_8204,N_6595);
xor U11180 (N_11180,N_6431,N_8703);
or U11181 (N_11181,N_9862,N_6470);
nor U11182 (N_11182,N_6774,N_6243);
nand U11183 (N_11183,N_5958,N_8656);
nor U11184 (N_11184,N_5151,N_6860);
xnor U11185 (N_11185,N_8170,N_9121);
nor U11186 (N_11186,N_6575,N_5586);
and U11187 (N_11187,N_5481,N_9062);
and U11188 (N_11188,N_8643,N_5355);
and U11189 (N_11189,N_9110,N_5306);
nand U11190 (N_11190,N_8499,N_7616);
nand U11191 (N_11191,N_5578,N_9869);
nand U11192 (N_11192,N_9700,N_6141);
nand U11193 (N_11193,N_9082,N_5805);
and U11194 (N_11194,N_9641,N_9591);
and U11195 (N_11195,N_7683,N_6621);
nor U11196 (N_11196,N_8389,N_9373);
xor U11197 (N_11197,N_6916,N_5075);
or U11198 (N_11198,N_5686,N_9990);
nand U11199 (N_11199,N_5796,N_7275);
and U11200 (N_11200,N_8994,N_7077);
xor U11201 (N_11201,N_8122,N_9394);
and U11202 (N_11202,N_8177,N_5699);
nor U11203 (N_11203,N_5142,N_5639);
nand U11204 (N_11204,N_5800,N_7489);
nor U11205 (N_11205,N_9125,N_9648);
or U11206 (N_11206,N_6870,N_7941);
nand U11207 (N_11207,N_9292,N_5330);
xor U11208 (N_11208,N_6768,N_8921);
and U11209 (N_11209,N_8408,N_5176);
xnor U11210 (N_11210,N_9550,N_9651);
or U11211 (N_11211,N_9859,N_5065);
or U11212 (N_11212,N_5688,N_7188);
nor U11213 (N_11213,N_8974,N_8022);
xnor U11214 (N_11214,N_5085,N_5631);
nand U11215 (N_11215,N_7614,N_5015);
and U11216 (N_11216,N_8680,N_8317);
or U11217 (N_11217,N_7955,N_7636);
nor U11218 (N_11218,N_9718,N_7719);
xnor U11219 (N_11219,N_8171,N_9933);
and U11220 (N_11220,N_9262,N_8616);
and U11221 (N_11221,N_8676,N_6202);
nand U11222 (N_11222,N_8918,N_5518);
nor U11223 (N_11223,N_7165,N_6846);
nand U11224 (N_11224,N_5648,N_5843);
and U11225 (N_11225,N_7429,N_6792);
nand U11226 (N_11226,N_6291,N_7748);
or U11227 (N_11227,N_8153,N_5128);
or U11228 (N_11228,N_8775,N_6023);
and U11229 (N_11229,N_8594,N_6047);
or U11230 (N_11230,N_6072,N_5685);
nand U11231 (N_11231,N_8049,N_8883);
and U11232 (N_11232,N_9500,N_5014);
or U11233 (N_11233,N_5297,N_5719);
nor U11234 (N_11234,N_6643,N_7668);
xnor U11235 (N_11235,N_8348,N_8157);
or U11236 (N_11236,N_5662,N_7268);
xor U11237 (N_11237,N_7338,N_6009);
or U11238 (N_11238,N_7166,N_6183);
nor U11239 (N_11239,N_9535,N_9554);
nor U11240 (N_11240,N_8820,N_6667);
xor U11241 (N_11241,N_8877,N_6279);
nor U11242 (N_11242,N_7823,N_9206);
xor U11243 (N_11243,N_8855,N_8642);
or U11244 (N_11244,N_6586,N_6244);
nor U11245 (N_11245,N_8810,N_5890);
and U11246 (N_11246,N_8173,N_8553);
nor U11247 (N_11247,N_9878,N_6744);
or U11248 (N_11248,N_8484,N_8953);
nand U11249 (N_11249,N_5384,N_6222);
nand U11250 (N_11250,N_6717,N_8138);
or U11251 (N_11251,N_6885,N_9340);
nand U11252 (N_11252,N_7690,N_5894);
nor U11253 (N_11253,N_7721,N_7916);
and U11254 (N_11254,N_8367,N_6804);
xor U11255 (N_11255,N_9133,N_6569);
and U11256 (N_11256,N_9290,N_9655);
nor U11257 (N_11257,N_9297,N_5712);
and U11258 (N_11258,N_6087,N_6810);
nand U11259 (N_11259,N_7555,N_5204);
and U11260 (N_11260,N_5830,N_5736);
and U11261 (N_11261,N_8847,N_7468);
or U11262 (N_11262,N_6692,N_9712);
and U11263 (N_11263,N_7071,N_5555);
nand U11264 (N_11264,N_8093,N_5394);
xnor U11265 (N_11265,N_9271,N_5484);
xor U11266 (N_11266,N_5655,N_6707);
or U11267 (N_11267,N_6363,N_8698);
and U11268 (N_11268,N_6962,N_8455);
and U11269 (N_11269,N_8145,N_6894);
nor U11270 (N_11270,N_7865,N_5459);
nor U11271 (N_11271,N_9021,N_6011);
nand U11272 (N_11272,N_6088,N_8792);
and U11273 (N_11273,N_9385,N_7482);
xnor U11274 (N_11274,N_8350,N_9822);
nor U11275 (N_11275,N_8933,N_8309);
or U11276 (N_11276,N_9022,N_6255);
xor U11277 (N_11277,N_6594,N_8771);
nand U11278 (N_11278,N_8839,N_9367);
and U11279 (N_11279,N_6993,N_8228);
and U11280 (N_11280,N_7756,N_7680);
or U11281 (N_11281,N_9162,N_6507);
or U11282 (N_11282,N_8620,N_6089);
nor U11283 (N_11283,N_6750,N_8663);
nor U11284 (N_11284,N_8014,N_7821);
nor U11285 (N_11285,N_5695,N_5743);
or U11286 (N_11286,N_7779,N_6808);
xnor U11287 (N_11287,N_9391,N_7744);
or U11288 (N_11288,N_8279,N_6194);
nor U11289 (N_11289,N_5878,N_6779);
nor U11290 (N_11290,N_7826,N_7233);
and U11291 (N_11291,N_7875,N_6954);
nand U11292 (N_11292,N_8425,N_7056);
nor U11293 (N_11293,N_9488,N_6760);
nor U11294 (N_11294,N_8278,N_8853);
or U11295 (N_11295,N_9307,N_6218);
nand U11296 (N_11296,N_9106,N_9176);
xnor U11297 (N_11297,N_9427,N_8567);
nor U11298 (N_11298,N_7138,N_7097);
xnor U11299 (N_11299,N_5953,N_8828);
nand U11300 (N_11300,N_5851,N_5756);
nor U11301 (N_11301,N_5458,N_6975);
nor U11302 (N_11302,N_5981,N_9732);
nand U11303 (N_11303,N_9761,N_9727);
nand U11304 (N_11304,N_8969,N_8427);
xor U11305 (N_11305,N_5672,N_8954);
or U11306 (N_11306,N_8246,N_7140);
and U11307 (N_11307,N_5683,N_7791);
nor U11308 (N_11308,N_7264,N_7986);
nand U11309 (N_11309,N_7738,N_6656);
nor U11310 (N_11310,N_5034,N_5025);
or U11311 (N_11311,N_6024,N_6579);
and U11312 (N_11312,N_9726,N_8600);
xor U11313 (N_11313,N_8942,N_9237);
or U11314 (N_11314,N_6664,N_6395);
xor U11315 (N_11315,N_9359,N_9668);
xnor U11316 (N_11316,N_8355,N_9119);
xnor U11317 (N_11317,N_8712,N_7272);
xor U11318 (N_11318,N_6535,N_5833);
xor U11319 (N_11319,N_7538,N_5742);
xnor U11320 (N_11320,N_6877,N_8629);
nor U11321 (N_11321,N_8221,N_7585);
nor U11322 (N_11322,N_6990,N_6474);
and U11323 (N_11323,N_6391,N_5495);
xnor U11324 (N_11324,N_5336,N_5371);
nand U11325 (N_11325,N_7396,N_8393);
or U11326 (N_11326,N_5583,N_7952);
xor U11327 (N_11327,N_7345,N_8527);
and U11328 (N_11328,N_9717,N_6987);
nor U11329 (N_11329,N_8624,N_9168);
nand U11330 (N_11330,N_5702,N_5417);
nand U11331 (N_11331,N_7541,N_6184);
xnor U11332 (N_11332,N_9607,N_5270);
nor U11333 (N_11333,N_8164,N_5274);
nor U11334 (N_11334,N_6016,N_7650);
nand U11335 (N_11335,N_9816,N_9746);
xor U11336 (N_11336,N_9291,N_5517);
nand U11337 (N_11337,N_8907,N_9636);
nand U11338 (N_11338,N_9456,N_5048);
xnor U11339 (N_11339,N_5284,N_9084);
nand U11340 (N_11340,N_5003,N_9937);
or U11341 (N_11341,N_6989,N_8659);
and U11342 (N_11342,N_7887,N_5904);
or U11343 (N_11343,N_7735,N_8460);
xnor U11344 (N_11344,N_8004,N_5019);
and U11345 (N_11345,N_5226,N_8638);
xnor U11346 (N_11346,N_7564,N_5872);
and U11347 (N_11347,N_6871,N_7589);
nor U11348 (N_11348,N_8471,N_6844);
or U11349 (N_11349,N_8726,N_6697);
nor U11350 (N_11350,N_9603,N_7562);
xnor U11351 (N_11351,N_7481,N_5532);
nor U11352 (N_11352,N_7973,N_9914);
nor U11353 (N_11353,N_8603,N_9627);
nand U11354 (N_11354,N_9088,N_8859);
and U11355 (N_11355,N_5320,N_5868);
xnor U11356 (N_11356,N_7776,N_5464);
xnor U11357 (N_11357,N_7593,N_8803);
nand U11358 (N_11358,N_8148,N_7371);
nor U11359 (N_11359,N_7372,N_9979);
nand U11360 (N_11360,N_9404,N_5869);
nor U11361 (N_11361,N_6032,N_7534);
and U11362 (N_11362,N_8370,N_7470);
and U11363 (N_11363,N_6084,N_5258);
xnor U11364 (N_11364,N_6394,N_9264);
xnor U11365 (N_11365,N_5839,N_6830);
and U11366 (N_11366,N_9898,N_9826);
xnor U11367 (N_11367,N_6343,N_7864);
nand U11368 (N_11368,N_9879,N_6608);
xor U11369 (N_11369,N_5374,N_8815);
nor U11370 (N_11370,N_8866,N_7364);
nor U11371 (N_11371,N_7936,N_6123);
nand U11372 (N_11372,N_9287,N_6675);
and U11373 (N_11373,N_6462,N_9315);
nand U11374 (N_11374,N_7637,N_8469);
nand U11375 (N_11375,N_8939,N_7742);
and U11376 (N_11376,N_7259,N_8129);
nor U11377 (N_11377,N_9479,N_9516);
or U11378 (N_11378,N_8958,N_6258);
nor U11379 (N_11379,N_9148,N_5867);
or U11380 (N_11380,N_6004,N_7605);
nor U11381 (N_11381,N_8063,N_9108);
xor U11382 (N_11382,N_5752,N_6463);
nand U11383 (N_11383,N_9713,N_8442);
nor U11384 (N_11384,N_7831,N_9128);
or U11385 (N_11385,N_7498,N_6165);
nor U11386 (N_11386,N_8984,N_9046);
nor U11387 (N_11387,N_9598,N_7414);
xor U11388 (N_11388,N_7836,N_6012);
nor U11389 (N_11389,N_9420,N_5030);
or U11390 (N_11390,N_5278,N_5237);
or U11391 (N_11391,N_7874,N_7153);
nor U11392 (N_11392,N_7348,N_9076);
or U11393 (N_11393,N_5432,N_8380);
nor U11394 (N_11394,N_8552,N_5261);
nand U11395 (N_11395,N_8092,N_5809);
and U11396 (N_11396,N_6598,N_5516);
or U11397 (N_11397,N_7956,N_6242);
xor U11398 (N_11398,N_8016,N_9413);
nor U11399 (N_11399,N_5103,N_9256);
and U11400 (N_11400,N_6866,N_5347);
nand U11401 (N_11401,N_6585,N_9999);
xor U11402 (N_11402,N_6164,N_7530);
or U11403 (N_11403,N_6426,N_6477);
xnor U11404 (N_11404,N_9218,N_6105);
or U11405 (N_11405,N_6763,N_7913);
or U11406 (N_11406,N_5323,N_9667);
nand U11407 (N_11407,N_8723,N_8451);
and U11408 (N_11408,N_8285,N_7053);
and U11409 (N_11409,N_7915,N_5060);
or U11410 (N_11410,N_5691,N_9527);
or U11411 (N_11411,N_7828,N_8105);
nor U11412 (N_11412,N_5123,N_8992);
nor U11413 (N_11413,N_6537,N_7041);
nand U11414 (N_11414,N_5942,N_9733);
and U11415 (N_11415,N_9328,N_8453);
and U11416 (N_11416,N_7012,N_7699);
nor U11417 (N_11417,N_9449,N_7244);
nand U11418 (N_11418,N_8588,N_5950);
nor U11419 (N_11419,N_7974,N_9006);
nand U11420 (N_11420,N_5956,N_5766);
and U11421 (N_11421,N_5273,N_5497);
nor U11422 (N_11422,N_5133,N_5262);
xor U11423 (N_11423,N_6347,N_6539);
nor U11424 (N_11424,N_6116,N_5332);
or U11425 (N_11425,N_6045,N_6227);
or U11426 (N_11426,N_8158,N_8879);
or U11427 (N_11427,N_6307,N_9643);
xnor U11428 (N_11428,N_8687,N_8664);
nand U11429 (N_11429,N_8797,N_5033);
nand U11430 (N_11430,N_8702,N_5130);
and U11431 (N_11431,N_5861,N_7177);
nor U11432 (N_11432,N_9289,N_9356);
xnor U11433 (N_11433,N_5264,N_5200);
xor U11434 (N_11434,N_6956,N_8788);
or U11435 (N_11435,N_8532,N_8310);
nor U11436 (N_11436,N_8586,N_7954);
nor U11437 (N_11437,N_5725,N_5689);
nand U11438 (N_11438,N_5486,N_5173);
and U11439 (N_11439,N_5328,N_5801);
nor U11440 (N_11440,N_5272,N_8784);
nor U11441 (N_11441,N_8314,N_8995);
or U11442 (N_11442,N_5832,N_9378);
nand U11443 (N_11443,N_8555,N_7566);
and U11444 (N_11444,N_5185,N_8292);
xor U11445 (N_11445,N_8215,N_6735);
nor U11446 (N_11446,N_6985,N_9406);
and U11447 (N_11447,N_5786,N_8424);
nor U11448 (N_11448,N_5408,N_5390);
nand U11449 (N_11449,N_9754,N_9073);
nor U11450 (N_11450,N_5139,N_7609);
or U11451 (N_11451,N_9606,N_8123);
nand U11452 (N_11452,N_7545,N_6609);
and U11453 (N_11453,N_9401,N_9448);
xnor U11454 (N_11454,N_5979,N_6927);
and U11455 (N_11455,N_6468,N_6518);
or U11456 (N_11456,N_8187,N_7136);
xor U11457 (N_11457,N_8667,N_9924);
nor U11458 (N_11458,N_6526,N_7707);
or U11459 (N_11459,N_8701,N_8341);
nand U11460 (N_11460,N_9209,N_5472);
nor U11461 (N_11461,N_7848,N_7505);
nor U11462 (N_11462,N_7386,N_9017);
nor U11463 (N_11463,N_5581,N_5855);
nor U11464 (N_11464,N_9435,N_5474);
and U11465 (N_11465,N_9010,N_5301);
xor U11466 (N_11466,N_5888,N_8050);
xnor U11467 (N_11467,N_5277,N_9464);
or U11468 (N_11468,N_5573,N_9631);
xnor U11469 (N_11469,N_7948,N_6051);
nor U11470 (N_11470,N_7657,N_6304);
nor U11471 (N_11471,N_9380,N_6955);
nor U11472 (N_11472,N_8813,N_9723);
or U11473 (N_11473,N_9799,N_8051);
and U11474 (N_11474,N_5817,N_5213);
nand U11475 (N_11475,N_7524,N_8693);
or U11476 (N_11476,N_6919,N_5242);
and U11477 (N_11477,N_7296,N_7841);
xnor U11478 (N_11478,N_7176,N_6666);
nand U11479 (N_11479,N_8447,N_8854);
xnor U11480 (N_11480,N_8304,N_9193);
nand U11481 (N_11481,N_9312,N_5844);
nor U11482 (N_11482,N_6787,N_8903);
and U11483 (N_11483,N_9269,N_8297);
or U11484 (N_11484,N_8549,N_6275);
or U11485 (N_11485,N_8400,N_8863);
nand U11486 (N_11486,N_9425,N_5907);
nand U11487 (N_11487,N_8805,N_5899);
xor U11488 (N_11488,N_8753,N_6633);
or U11489 (N_11489,N_6484,N_8113);
nor U11490 (N_11490,N_9876,N_8220);
and U11491 (N_11491,N_8287,N_9211);
nand U11492 (N_11492,N_7425,N_6861);
nor U11493 (N_11493,N_5452,N_7901);
and U11494 (N_11494,N_6825,N_8281);
or U11495 (N_11495,N_9663,N_7289);
nand U11496 (N_11496,N_7162,N_9334);
or U11497 (N_11497,N_8443,N_5794);
xor U11498 (N_11498,N_6147,N_8321);
xor U11499 (N_11499,N_7597,N_8791);
or U11500 (N_11500,N_9188,N_8272);
and U11501 (N_11501,N_5864,N_5149);
nor U11502 (N_11502,N_9035,N_7922);
or U11503 (N_11503,N_5582,N_8252);
nand U11504 (N_11504,N_7537,N_6687);
and U11505 (N_11505,N_9278,N_7634);
or U11506 (N_11506,N_8725,N_6545);
nor U11507 (N_11507,N_6497,N_8688);
nand U11508 (N_11508,N_8561,N_6764);
xnor U11509 (N_11509,N_9139,N_8241);
nor U11510 (N_11510,N_6815,N_6896);
nor U11511 (N_11511,N_6378,N_8786);
nand U11512 (N_11512,N_7469,N_5674);
or U11513 (N_11513,N_6727,N_5111);
xnor U11514 (N_11514,N_9959,N_7120);
and U11515 (N_11515,N_7284,N_7190);
or U11516 (N_11516,N_6721,N_6268);
or U11517 (N_11517,N_8941,N_8597);
nand U11518 (N_11518,N_9671,N_5429);
and U11519 (N_11519,N_8950,N_7346);
and U11520 (N_11520,N_6580,N_7411);
nor U11521 (N_11521,N_9691,N_5522);
and U11522 (N_11522,N_9604,N_7281);
xor U11523 (N_11523,N_9283,N_8612);
or U11524 (N_11524,N_8264,N_5753);
nand U11525 (N_11525,N_8216,N_7928);
and U11526 (N_11526,N_6021,N_8475);
or U11527 (N_11527,N_6777,N_8244);
and U11528 (N_11528,N_9630,N_9546);
nor U11529 (N_11529,N_9660,N_9382);
and U11530 (N_11530,N_6290,N_8233);
nor U11531 (N_11531,N_9948,N_8694);
xnor U11532 (N_11532,N_9856,N_8224);
nor U11533 (N_11533,N_9368,N_5771);
and U11534 (N_11534,N_7062,N_5020);
nand U11535 (N_11535,N_9998,N_7789);
nand U11536 (N_11536,N_9520,N_8731);
and U11537 (N_11537,N_8968,N_9390);
nor U11538 (N_11538,N_5021,N_6806);
nand U11539 (N_11539,N_8888,N_5601);
and U11540 (N_11540,N_5400,N_5431);
nand U11541 (N_11541,N_6146,N_6172);
nor U11542 (N_11542,N_6857,N_8570);
or U11543 (N_11543,N_7035,N_5893);
nor U11544 (N_11544,N_9670,N_5972);
nor U11545 (N_11545,N_6686,N_5018);
nand U11546 (N_11546,N_6213,N_8335);
xor U11547 (N_11547,N_5490,N_8564);
nand U11548 (N_11548,N_8602,N_5468);
nor U11549 (N_11549,N_9549,N_8062);
nand U11550 (N_11550,N_8108,N_8617);
and U11551 (N_11551,N_9097,N_5370);
nand U11552 (N_11552,N_9265,N_5000);
nor U11553 (N_11553,N_8848,N_6850);
xnor U11554 (N_11554,N_9909,N_8438);
or U11555 (N_11555,N_8385,N_6709);
or U11556 (N_11556,N_8041,N_5496);
and U11557 (N_11557,N_6515,N_5993);
nand U11558 (N_11558,N_6864,N_7440);
and U11559 (N_11559,N_6083,N_9847);
nand U11560 (N_11560,N_7929,N_8468);
nor U11561 (N_11561,N_8515,N_8510);
nor U11562 (N_11562,N_6642,N_9758);
or U11563 (N_11563,N_6373,N_5153);
xor U11564 (N_11564,N_5916,N_5977);
xnor U11565 (N_11565,N_7758,N_9903);
nand U11566 (N_11566,N_6323,N_7559);
nand U11567 (N_11567,N_9682,N_5222);
nand U11568 (N_11568,N_8136,N_9507);
and U11569 (N_11569,N_8799,N_7318);
xor U11570 (N_11570,N_5116,N_8059);
xor U11571 (N_11571,N_5755,N_6340);
and U11572 (N_11572,N_9379,N_6875);
nand U11573 (N_11573,N_6724,N_8522);
or U11574 (N_11574,N_5471,N_7044);
nor U11575 (N_11575,N_9552,N_8478);
xnor U11576 (N_11576,N_7004,N_7567);
nor U11577 (N_11577,N_8403,N_8318);
or U11578 (N_11578,N_5998,N_7446);
nand U11579 (N_11579,N_6679,N_6571);
or U11580 (N_11580,N_8910,N_6556);
nand U11581 (N_11581,N_9310,N_8193);
xnor U11582 (N_11582,N_6636,N_7796);
xnor U11583 (N_11583,N_9495,N_6693);
or U11584 (N_11584,N_7854,N_5658);
nor U11585 (N_11585,N_5765,N_7406);
nor U11586 (N_11586,N_6651,N_6216);
nand U11587 (N_11587,N_5633,N_5228);
xnor U11588 (N_11588,N_5509,N_5192);
xnor U11589 (N_11589,N_6809,N_6762);
or U11590 (N_11590,N_7741,N_5058);
xnor U11591 (N_11591,N_8919,N_7310);
nand U11592 (N_11592,N_5102,N_8234);
and U11593 (N_11593,N_6630,N_5616);
or U11594 (N_11594,N_6271,N_7445);
nand U11595 (N_11595,N_9174,N_7747);
and U11596 (N_11596,N_6572,N_9911);
nor U11597 (N_11597,N_7064,N_7319);
xnor U11598 (N_11598,N_8103,N_9926);
or U11599 (N_11599,N_9752,N_5499);
nor U11600 (N_11600,N_8750,N_9982);
nand U11601 (N_11601,N_9572,N_6107);
nand U11602 (N_11602,N_7011,N_9364);
nand U11603 (N_11603,N_8626,N_8631);
and U11604 (N_11604,N_5174,N_7486);
xor U11605 (N_11605,N_7328,N_8256);
nand U11606 (N_11606,N_5266,N_6553);
nand U11607 (N_11607,N_5792,N_7339);
or U11608 (N_11608,N_8523,N_9823);
nor U11609 (N_11609,N_6994,N_7085);
xor U11610 (N_11610,N_6605,N_5572);
nand U11611 (N_11611,N_5368,N_7717);
or U11612 (N_11612,N_8444,N_5401);
nand U11613 (N_11613,N_6796,N_7217);
xor U11614 (N_11614,N_8102,N_7017);
nand U11615 (N_11615,N_6831,N_7764);
or U11616 (N_11616,N_6181,N_5359);
and U11617 (N_11617,N_8758,N_5986);
xnor U11618 (N_11618,N_9724,N_7824);
xor U11619 (N_11619,N_5201,N_8308);
xor U11620 (N_11620,N_7195,N_6256);
or U11621 (N_11621,N_5507,N_9494);
or U11622 (N_11622,N_6336,N_5954);
or U11623 (N_11623,N_6452,N_5933);
and U11624 (N_11624,N_7701,N_8806);
nor U11625 (N_11625,N_7572,N_6599);
or U11626 (N_11626,N_5354,N_6273);
xnor U11627 (N_11627,N_9504,N_7917);
nand U11628 (N_11628,N_5551,N_9178);
and U11629 (N_11629,N_5241,N_9855);
nand U11630 (N_11630,N_5026,N_9402);
nand U11631 (N_11631,N_9403,N_9734);
or U11632 (N_11632,N_7522,N_5358);
and U11633 (N_11633,N_7761,N_6932);
nor U11634 (N_11634,N_6292,N_6467);
xnor U11635 (N_11635,N_7506,N_9352);
nand U11636 (N_11636,N_7148,N_5620);
xnor U11637 (N_11637,N_5279,N_7725);
nand U11638 (N_11638,N_8766,N_8097);
xnor U11639 (N_11639,N_5504,N_6937);
and U11640 (N_11640,N_8658,N_6365);
and U11641 (N_11641,N_7613,N_5770);
or U11642 (N_11642,N_5450,N_7341);
nor U11643 (N_11643,N_8789,N_9214);
and U11644 (N_11644,N_8733,N_5117);
and U11645 (N_11645,N_5537,N_8351);
nand U11646 (N_11646,N_7920,N_5591);
nor U11647 (N_11647,N_5198,N_7373);
and U11648 (N_11648,N_8176,N_7032);
nor U11649 (N_11649,N_9212,N_5734);
xnor U11650 (N_11650,N_8838,N_5480);
or U11651 (N_11651,N_9202,N_5835);
nor U11652 (N_11652,N_5562,N_5525);
nor U11653 (N_11653,N_9704,N_7196);
nand U11654 (N_11654,N_5865,N_5822);
xor U11655 (N_11655,N_9014,N_6208);
or U11656 (N_11656,N_8338,N_7563);
nand U11657 (N_11657,N_7491,N_6328);
xnor U11658 (N_11658,N_8871,N_8217);
or U11659 (N_11659,N_6657,N_6888);
nor U11660 (N_11660,N_9141,N_9474);
nand U11661 (N_11661,N_6925,N_6548);
nand U11662 (N_11662,N_6265,N_6851);
or U11663 (N_11663,N_7115,N_9748);
xor U11664 (N_11664,N_9184,N_9371);
nor U11665 (N_11665,N_6033,N_8349);
nor U11666 (N_11666,N_9677,N_9932);
and U11667 (N_11667,N_9064,N_6696);
and U11668 (N_11668,N_5162,N_8311);
or U11669 (N_11669,N_6245,N_7693);
nand U11670 (N_11670,N_8652,N_9834);
and U11671 (N_11671,N_6129,N_9496);
xor U11672 (N_11672,N_5165,N_6239);
xnor U11673 (N_11673,N_6911,N_9538);
nor U11674 (N_11674,N_7632,N_5423);
nand U11675 (N_11675,N_5592,N_8125);
xnor U11676 (N_11676,N_9344,N_5147);
and U11677 (N_11677,N_8299,N_6644);
nand U11678 (N_11678,N_5508,N_6723);
nand U11679 (N_11679,N_6339,N_7228);
and U11680 (N_11680,N_9194,N_8513);
nor U11681 (N_11681,N_8841,N_7803);
xnor U11682 (N_11682,N_6736,N_6445);
nand U11683 (N_11683,N_7918,N_8015);
and U11684 (N_11684,N_7479,N_9703);
xor U11685 (N_11685,N_7586,N_7374);
nor U11686 (N_11686,N_5602,N_5842);
nand U11687 (N_11687,N_6852,N_8644);
xor U11688 (N_11688,N_9548,N_8901);
nand U11689 (N_11689,N_5300,N_6295);
xor U11690 (N_11690,N_6547,N_8747);
xnor U11691 (N_11691,N_7985,N_8012);
xnor U11692 (N_11692,N_9077,N_9542);
and U11693 (N_11693,N_7366,N_7069);
or U11694 (N_11694,N_9892,N_5078);
nor U11695 (N_11695,N_5479,N_6299);
or U11696 (N_11696,N_9122,N_7633);
xor U11697 (N_11697,N_9068,N_9683);
nand U11698 (N_11698,N_6583,N_7376);
nand U11699 (N_11699,N_5852,N_5975);
nor U11700 (N_11700,N_5227,N_5502);
or U11701 (N_11701,N_6049,N_9207);
nor U11702 (N_11702,N_5307,N_9689);
xnor U11703 (N_11703,N_7870,N_7360);
nor U11704 (N_11704,N_8345,N_6427);
nand U11705 (N_11705,N_6383,N_5115);
or U11706 (N_11706,N_5679,N_8000);
and U11707 (N_11707,N_9881,N_6013);
nor U11708 (N_11708,N_8374,N_7293);
or U11709 (N_11709,N_8497,N_5203);
and U11710 (N_11710,N_7595,N_6377);
nand U11711 (N_11711,N_6828,N_5473);
and U11712 (N_11712,N_8884,N_6773);
nor U11713 (N_11713,N_5311,N_8654);
xor U11714 (N_11714,N_9913,N_5398);
xnor U11715 (N_11715,N_8305,N_9557);
or U11716 (N_11716,N_8897,N_7886);
or U11717 (N_11717,N_8745,N_7783);
or U11718 (N_11718,N_6155,N_7021);
or U11719 (N_11719,N_7324,N_6322);
nor U11720 (N_11720,N_8169,N_5790);
and U11721 (N_11721,N_7734,N_7815);
nor U11722 (N_11722,N_7785,N_7891);
or U11723 (N_11723,N_6359,N_6042);
nand U11724 (N_11724,N_8211,N_6601);
xnor U11725 (N_11725,N_9120,N_9785);
nand U11726 (N_11726,N_8490,N_8534);
and U11727 (N_11727,N_9980,N_5730);
nand U11728 (N_11728,N_7451,N_8144);
xor U11729 (N_11729,N_6071,N_6158);
or U11730 (N_11730,N_9225,N_9825);
or U11731 (N_11731,N_7456,N_7709);
or U11732 (N_11732,N_5980,N_9705);
xor U11733 (N_11733,N_8876,N_8852);
nand U11734 (N_11734,N_5936,N_6887);
xnor U11735 (N_11735,N_7146,N_9617);
and U11736 (N_11736,N_7465,N_6041);
nand U11737 (N_11737,N_7471,N_9762);
nor U11738 (N_11738,N_8822,N_8983);
and U11739 (N_11739,N_7896,N_5623);
nand U11740 (N_11740,N_5478,N_7317);
nor U11741 (N_11741,N_6508,N_6970);
xnor U11742 (N_11742,N_9904,N_9851);
and U11743 (N_11743,N_5530,N_6419);
nor U11744 (N_11744,N_8707,N_9224);
nor U11745 (N_11745,N_9772,N_6628);
nor U11746 (N_11746,N_5891,N_8700);
or U11747 (N_11747,N_5433,N_9597);
nor U11748 (N_11748,N_5764,N_5997);
nor U11749 (N_11749,N_5652,N_8966);
xnor U11750 (N_11750,N_9299,N_9743);
or U11751 (N_11751,N_6411,N_8428);
and U11752 (N_11752,N_8388,N_9935);
nand U11753 (N_11753,N_6454,N_9231);
nor U11754 (N_11754,N_5364,N_6492);
nor U11755 (N_11755,N_6085,N_8661);
or U11756 (N_11756,N_5028,N_7571);
or U11757 (N_11757,N_8496,N_6622);
nor U11758 (N_11758,N_8826,N_7934);
xor U11759 (N_11759,N_7159,N_6406);
nand U11760 (N_11760,N_8242,N_9669);
and U11761 (N_11761,N_7201,N_5191);
and U11762 (N_11762,N_6936,N_5454);
and U11763 (N_11763,N_6230,N_9409);
nor U11764 (N_11764,N_9143,N_8486);
and U11765 (N_11765,N_7378,N_5708);
nor U11766 (N_11766,N_6801,N_8375);
or U11767 (N_11767,N_7866,N_9844);
nor U11768 (N_11768,N_9775,N_6413);
nor U11769 (N_11769,N_8787,N_5661);
xor U11770 (N_11770,N_6758,N_9107);
or U11771 (N_11771,N_9975,N_7847);
nor U11772 (N_11772,N_7499,N_6528);
and U11773 (N_11773,N_7042,N_8142);
nand U11774 (N_11774,N_9158,N_6006);
xnor U11775 (N_11775,N_5314,N_7696);
nor U11776 (N_11776,N_9697,N_7816);
nor U11777 (N_11777,N_5100,N_7565);
xnor U11778 (N_11778,N_9103,N_9072);
nand U11779 (N_11779,N_8068,N_8923);
xor U11780 (N_11780,N_9974,N_7832);
nor U11781 (N_11781,N_8790,N_6930);
and U11782 (N_11782,N_6297,N_7914);
and U11783 (N_11783,N_8556,N_6731);
and U11784 (N_11784,N_6401,N_8836);
and U11785 (N_11785,N_6068,N_7906);
nor U11786 (N_11786,N_7493,N_8199);
nand U11787 (N_11787,N_8040,N_5329);
or U11788 (N_11788,N_9351,N_6302);
or U11789 (N_11789,N_5780,N_8027);
nor U11790 (N_11790,N_8060,N_9936);
xnor U11791 (N_11791,N_7677,N_5706);
nand U11792 (N_11792,N_8997,N_8767);
nor U11793 (N_11793,N_6349,N_5895);
nor U11794 (N_11794,N_5880,N_9429);
and U11795 (N_11795,N_8557,N_7167);
and U11796 (N_11796,N_6253,N_9009);
and U11797 (N_11797,N_5704,N_6873);
xor U11798 (N_11798,N_6103,N_6371);
xnor U11799 (N_11799,N_7013,N_5415);
nand U11800 (N_11800,N_7862,N_9730);
nor U11801 (N_11801,N_5036,N_7147);
nand U11802 (N_11802,N_6645,N_8891);
nor U11803 (N_11803,N_9537,N_6104);
and U11804 (N_11804,N_9101,N_9970);
xor U11805 (N_11805,N_5858,N_8867);
nand U11806 (N_11806,N_6496,N_7192);
or U11807 (N_11807,N_5905,N_7394);
xor U11808 (N_11808,N_8937,N_7999);
nand U11809 (N_11809,N_8756,N_6701);
nand U11810 (N_11810,N_6161,N_5557);
nor U11811 (N_11811,N_9714,N_5666);
nand U11812 (N_11812,N_9593,N_8373);
nor U11813 (N_11813,N_7452,N_8030);
and U11814 (N_11814,N_9234,N_5465);
xor U11815 (N_11815,N_7460,N_7787);
xor U11816 (N_11816,N_9787,N_8090);
xnor U11817 (N_11817,N_8823,N_9808);
and U11818 (N_11818,N_6204,N_7260);
and U11819 (N_11819,N_7885,N_6093);
and U11820 (N_11820,N_9407,N_5158);
and U11821 (N_11821,N_6757,N_9342);
xnor U11822 (N_11822,N_6466,N_5302);
nand U11823 (N_11823,N_6769,N_6510);
and U11824 (N_11824,N_7370,N_5664);
and U11825 (N_11825,N_6106,N_5308);
nand U11826 (N_11826,N_5053,N_5343);
or U11827 (N_11827,N_5546,N_7600);
and U11828 (N_11828,N_7967,N_7765);
nor U11829 (N_11829,N_9220,N_5041);
nor U11830 (N_11830,N_8653,N_7023);
nand U11831 (N_11831,N_7921,N_7091);
nor U11832 (N_11832,N_7003,N_9284);
xor U11833 (N_11833,N_9801,N_9208);
and U11834 (N_11834,N_8013,N_5700);
xnor U11835 (N_11835,N_9296,N_8804);
xnor U11836 (N_11836,N_7568,N_6931);
and U11837 (N_11837,N_5340,N_6416);
xnor U11838 (N_11838,N_9763,N_6784);
xor U11839 (N_11839,N_5768,N_9672);
nand U11840 (N_11840,N_7994,N_9942);
xor U11841 (N_11841,N_5645,N_6691);
nand U11842 (N_11842,N_7728,N_7960);
nor U11843 (N_11843,N_5095,N_7007);
or U11844 (N_11844,N_6077,N_9901);
nor U11845 (N_11845,N_7098,N_9145);
and U11846 (N_11846,N_7443,N_9478);
nor U11847 (N_11847,N_7490,N_9747);
nand U11848 (N_11848,N_5292,N_7830);
nor U11849 (N_11849,N_8686,N_9441);
and U11850 (N_11850,N_8773,N_5680);
and U11851 (N_11851,N_9067,N_5282);
or U11852 (N_11852,N_9613,N_6559);
and U11853 (N_11853,N_9161,N_6354);
or U11854 (N_11854,N_9715,N_6065);
nand U11855 (N_11855,N_9857,N_5125);
and U11856 (N_11856,N_8207,N_5618);
nor U11857 (N_11857,N_9049,N_8072);
or U11858 (N_11858,N_8675,N_6690);
nor U11859 (N_11859,N_9195,N_6215);
xnor U11860 (N_11860,N_9007,N_7603);
or U11861 (N_11861,N_9720,N_5397);
or U11862 (N_11862,N_6188,N_7552);
xor U11863 (N_11863,N_7294,N_5875);
xnor U11864 (N_11864,N_5999,N_8412);
and U11865 (N_11865,N_8768,N_6910);
and U11866 (N_11866,N_9943,N_5049);
and U11867 (N_11867,N_9362,N_5293);
and U11868 (N_11868,N_9028,N_5250);
and U11869 (N_11869,N_9646,N_8334);
nand U11870 (N_11870,N_9095,N_9240);
nor U11871 (N_11871,N_9947,N_6313);
xor U11872 (N_11872,N_5072,N_9547);
or U11873 (N_11873,N_8208,N_5069);
xor U11874 (N_11874,N_9215,N_7397);
or U11875 (N_11875,N_8327,N_7583);
xor U11876 (N_11876,N_6266,N_5939);
nor U11877 (N_11877,N_8360,N_6673);
nor U11878 (N_11878,N_7186,N_9800);
and U11879 (N_11879,N_8569,N_9112);
nand U11880 (N_11880,N_8537,N_5267);
nand U11881 (N_11881,N_5848,N_7570);
and U11882 (N_11882,N_5682,N_6933);
nor U11883 (N_11883,N_5873,N_5883);
nor U11884 (N_11884,N_9596,N_8300);
and U11885 (N_11885,N_6818,N_7542);
and U11886 (N_11886,N_8025,N_6133);
nand U11887 (N_11887,N_9994,N_5099);
nor U11888 (N_11888,N_6836,N_9922);
and U11889 (N_11889,N_7819,N_9690);
nand U11890 (N_11890,N_8205,N_9977);
nor U11891 (N_11891,N_8655,N_9771);
or U11892 (N_11892,N_6145,N_9245);
nand U11893 (N_11893,N_6856,N_5949);
nand U11894 (N_11894,N_8989,N_5245);
and U11895 (N_11895,N_7152,N_9255);
nor U11896 (N_11896,N_9395,N_9506);
or U11897 (N_11897,N_5254,N_8156);
nand U11898 (N_11898,N_8936,N_9873);
nor U11899 (N_11899,N_6185,N_6603);
nand U11900 (N_11900,N_7368,N_7111);
xor U11901 (N_11901,N_5769,N_5837);
xnor U11902 (N_11902,N_7301,N_8229);
or U11903 (N_11903,N_9484,N_8730);
nand U11904 (N_11904,N_8065,N_7119);
or U11905 (N_11905,N_5260,N_8101);
and U11906 (N_11906,N_6610,N_5363);
xor U11907 (N_11907,N_5157,N_7863);
xor U11908 (N_11908,N_6301,N_9757);
or U11909 (N_11909,N_7400,N_6099);
and U11910 (N_11910,N_9600,N_6849);
xor U11911 (N_11911,N_5392,N_8245);
or U11912 (N_11912,N_9446,N_6530);
nand U11913 (N_11913,N_8900,N_9831);
nand U11914 (N_11914,N_5183,N_8267);
xnor U11915 (N_11915,N_5470,N_7238);
and U11916 (N_11916,N_8347,N_8445);
and U11917 (N_11917,N_6491,N_7692);
xnor U11918 (N_11918,N_6632,N_8682);
xor U11919 (N_11919,N_8610,N_6480);
and U11920 (N_11920,N_6403,N_5068);
or U11921 (N_11921,N_6028,N_5548);
xnor U11922 (N_11922,N_5092,N_9096);
xor U11923 (N_11923,N_5422,N_5560);
nand U11924 (N_11924,N_7405,N_9173);
and U11925 (N_11925,N_8198,N_9258);
and U11926 (N_11926,N_8056,N_9976);
or U11927 (N_11927,N_7972,N_8446);
and U11928 (N_11928,N_5317,N_8524);
and U11929 (N_11929,N_7322,N_8814);
xor U11930 (N_11930,N_9741,N_5747);
xnor U11931 (N_11931,N_8269,N_7355);
or U11932 (N_11932,N_6703,N_8280);
xnor U11933 (N_11933,N_5385,N_7822);
nand U11934 (N_11934,N_8849,N_8266);
nand U11935 (N_11935,N_5288,N_9029);
or U11936 (N_11936,N_6053,N_6000);
xnor U11937 (N_11937,N_9965,N_6683);
xnor U11938 (N_11938,N_6412,N_5721);
nor U11939 (N_11939,N_5335,N_9653);
nand U11940 (N_11940,N_9711,N_6800);
nand U11941 (N_11941,N_9725,N_9167);
nand U11942 (N_11942,N_5610,N_5137);
nor U11943 (N_11943,N_9756,N_5538);
xnor U11944 (N_11944,N_8914,N_8634);
nand U11945 (N_11945,N_7894,N_7674);
or U11946 (N_11946,N_6238,N_6338);
nor U11947 (N_11947,N_7237,N_5968);
nor U11948 (N_11948,N_6922,N_5925);
or U11949 (N_11949,N_8827,N_9444);
nand U11950 (N_11950,N_5985,N_9041);
nor U11951 (N_11951,N_6117,N_5646);
nor U11952 (N_11952,N_8692,N_7313);
nand U11953 (N_11953,N_8944,N_8409);
and U11954 (N_11954,N_5677,N_6410);
xnor U11955 (N_11955,N_5221,N_5940);
or U11956 (N_11956,N_8817,N_5286);
xnor U11957 (N_11957,N_6421,N_5776);
xor U11958 (N_11958,N_6175,N_8985);
nand U11959 (N_11959,N_9927,N_5932);
and U11960 (N_11960,N_8529,N_9657);
and U11961 (N_11961,N_5897,N_6096);
or U11962 (N_11962,N_9784,N_7793);
nor U11963 (N_11963,N_9408,N_6938);
xnor U11964 (N_11964,N_5642,N_9490);
nor U11965 (N_11965,N_6483,N_9272);
nor U11966 (N_11966,N_8738,N_5584);
or U11967 (N_11967,N_5367,N_8505);
nor U11968 (N_11968,N_8218,N_7093);
or U11969 (N_11969,N_7484,N_7422);
and U11970 (N_11970,N_8212,N_7420);
nor U11971 (N_11971,N_6498,N_7878);
nor U11972 (N_11972,N_6739,N_9841);
nand U11973 (N_11973,N_9481,N_5148);
and U11974 (N_11974,N_9529,N_9505);
or U11975 (N_11975,N_5913,N_5561);
xnor U11976 (N_11976,N_5395,N_6308);
and U11977 (N_11977,N_7312,N_7288);
xor U11978 (N_11978,N_8710,N_8075);
nor U11979 (N_11979,N_6832,N_5637);
nand U11980 (N_11980,N_7266,N_9437);
nor U11981 (N_11981,N_8184,N_6536);
xnor U11982 (N_11982,N_5406,N_5996);
and U11983 (N_11983,N_5298,N_7434);
or U11984 (N_11984,N_9654,N_5924);
and U11985 (N_11985,N_9458,N_9384);
or U11986 (N_11986,N_9565,N_9180);
and U11987 (N_11987,N_6976,N_9447);
xor U11988 (N_11988,N_8630,N_6765);
nor U11989 (N_11989,N_5767,N_5155);
nor U11990 (N_11990,N_7871,N_6814);
or U11991 (N_11991,N_5184,N_6284);
and U11992 (N_11992,N_9582,N_5866);
and U11993 (N_11993,N_7253,N_5615);
nand U11994 (N_11994,N_8099,N_6920);
or U11995 (N_11995,N_7473,N_7525);
xor U11996 (N_11996,N_5608,N_7745);
nor U11997 (N_11997,N_8036,N_6195);
nand U11998 (N_11998,N_5634,N_7695);
nor U11999 (N_11999,N_6274,N_7574);
nand U12000 (N_12000,N_7944,N_7198);
and U12001 (N_12001,N_6702,N_5042);
xor U12002 (N_12002,N_5500,N_9113);
and U12003 (N_12003,N_6450,N_6835);
nor U12004 (N_12004,N_5404,N_5570);
nor U12005 (N_12005,N_7442,N_9154);
and U12006 (N_12006,N_9124,N_9155);
nor U12007 (N_12007,N_7395,N_5503);
or U12008 (N_12008,N_8741,N_5594);
and U12009 (N_12009,N_6296,N_8458);
xor U12010 (N_12010,N_5823,N_7387);
nor U12011 (N_12011,N_9233,N_7730);
nand U12012 (N_12012,N_6756,N_8325);
and U12013 (N_12013,N_6337,N_7134);
and U12014 (N_12014,N_6658,N_5231);
nand U12015 (N_12015,N_8045,N_7184);
and U12016 (N_12016,N_8893,N_5732);
nor U12017 (N_12017,N_5816,N_5037);
nor U12018 (N_12018,N_6267,N_9944);
nand U12019 (N_12019,N_9971,N_8024);
xnor U12020 (N_12020,N_7782,N_8005);
or U12021 (N_12021,N_8500,N_9647);
and U12022 (N_12022,N_7161,N_7978);
or U12023 (N_12023,N_8259,N_9584);
xnor U12024 (N_12024,N_9423,N_5813);
nand U12025 (N_12025,N_5671,N_5420);
xor U12026 (N_12026,N_8571,N_8816);
xnor U12027 (N_12027,N_7504,N_5547);
nand U12028 (N_12028,N_8291,N_7591);
xnor U12029 (N_12029,N_7996,N_5310);
nor U12030 (N_12030,N_5501,N_7426);
or U12031 (N_12031,N_5098,N_7412);
and U12032 (N_12032,N_7664,N_6458);
nor U12033 (N_12033,N_5381,N_6653);
nor U12034 (N_12034,N_9242,N_9830);
nor U12035 (N_12035,N_6909,N_8683);
nor U12036 (N_12036,N_6819,N_5339);
nand U12037 (N_12037,N_7762,N_6241);
or U12038 (N_12038,N_7295,N_8140);
nand U12039 (N_12039,N_5482,N_7448);
or U12040 (N_12040,N_6863,N_9008);
nand U12041 (N_12041,N_6511,N_9183);
nand U12042 (N_12042,N_6081,N_6415);
and U12043 (N_12043,N_6543,N_9327);
xnor U12044 (N_12044,N_9780,N_8053);
xor U12045 (N_12045,N_7379,N_5909);
or U12046 (N_12046,N_6446,N_8306);
or U12047 (N_12047,N_5017,N_9699);
nand U12048 (N_12048,N_9074,N_5519);
and U12049 (N_12049,N_7749,N_7684);
xor U12050 (N_12050,N_8530,N_8154);
and U12051 (N_12051,N_9945,N_9164);
nand U12052 (N_12052,N_9866,N_8039);
xnor U12053 (N_12053,N_8196,N_6043);
and U12054 (N_12054,N_7869,N_8323);
and U12055 (N_12055,N_8678,N_7182);
nor U12056 (N_12056,N_6250,N_9827);
xor U12057 (N_12057,N_5108,N_6634);
nand U12058 (N_12058,N_8765,N_7351);
and U12059 (N_12059,N_9722,N_7437);
nor U12060 (N_12060,N_9172,N_8454);
nand U12061 (N_12061,N_5543,N_9349);
nor U12062 (N_12062,N_5871,N_6380);
nand U12063 (N_12063,N_9383,N_9503);
nand U12064 (N_12064,N_6616,N_7240);
or U12065 (N_12065,N_8504,N_5235);
xnor U12066 (N_12066,N_7205,N_5523);
xnor U12067 (N_12067,N_7163,N_6351);
and U12068 (N_12068,N_9025,N_7320);
and U12069 (N_12069,N_6358,N_9915);
or U12070 (N_12070,N_8362,N_7231);
xor U12071 (N_12071,N_5457,N_7215);
xor U12072 (N_12072,N_6899,N_8436);
nand U12073 (N_12073,N_9235,N_6957);
or U12074 (N_12074,N_5045,N_7330);
and U12075 (N_12075,N_8417,N_7365);
nand U12076 (N_12076,N_9885,N_9219);
and U12077 (N_12077,N_5444,N_6759);
nor U12078 (N_12078,N_9802,N_5515);
nand U12079 (N_12079,N_5831,N_8503);
nor U12080 (N_12080,N_7173,N_7478);
and U12081 (N_12081,N_8197,N_8302);
nand U12082 (N_12082,N_6120,N_9434);
nor U12083 (N_12083,N_5841,N_8255);
xor U12084 (N_12084,N_8627,N_6040);
nor U12085 (N_12085,N_7333,N_5362);
or U12086 (N_12086,N_9820,N_6705);
and U12087 (N_12087,N_5344,N_9501);
and U12088 (N_12088,N_8071,N_6646);
nor U12089 (N_12089,N_9266,N_7180);
xnor U12090 (N_12090,N_9439,N_9626);
or U12091 (N_12091,N_9045,N_8190);
xnor U12092 (N_12092,N_8739,N_9917);
and U12093 (N_12093,N_7557,N_6193);
nor U12094 (N_12094,N_7890,N_8595);
xor U12095 (N_12095,N_9745,N_7089);
nor U12096 (N_12096,N_5202,N_6733);
and U12097 (N_12097,N_7199,N_9348);
nand U12098 (N_12098,N_6281,N_6647);
nor U12099 (N_12099,N_9968,N_9253);
nand U12100 (N_12100,N_5283,N_7547);
nor U12101 (N_12101,N_7606,N_7990);
and U12102 (N_12102,N_7354,N_5990);
nor U12103 (N_12103,N_8181,N_5341);
nand U12104 (N_12104,N_7353,N_9493);
or U12105 (N_12105,N_6214,N_9614);
nand U12106 (N_12106,N_8023,N_6981);
and U12107 (N_12107,N_9104,N_8544);
nand U12108 (N_12108,N_7427,N_8461);
xor U12109 (N_12109,N_6240,N_6173);
or U12110 (N_12110,N_8802,N_5113);
xor U12111 (N_12111,N_9991,N_9908);
xor U12112 (N_12112,N_8577,N_5243);
xnor U12113 (N_12113,N_9424,N_6623);
nand U12114 (N_12114,N_7447,N_7975);
nor U12115 (N_12115,N_8546,N_9136);
nor U12116 (N_12116,N_7037,N_5569);
nor U12117 (N_12117,N_9055,N_6191);
and U12118 (N_12118,N_5299,N_7088);
xnor U12119 (N_12119,N_7149,N_6187);
nand U12120 (N_12120,N_5498,N_6812);
and U12121 (N_12121,N_7646,N_8632);
and U12122 (N_12122,N_9350,N_6912);
or U12123 (N_12123,N_8124,N_6487);
and U12124 (N_12124,N_7590,N_8121);
nor U12125 (N_12125,N_7156,N_9973);
nand U12126 (N_12126,N_8404,N_7143);
xnor U12127 (N_12127,N_6321,N_7962);
and U12128 (N_12128,N_5319,N_7817);
nand U12129 (N_12129,N_6176,N_9709);
nor U12130 (N_12130,N_7105,N_9583);
or U12131 (N_12131,N_8865,N_9325);
xnor U12132 (N_12132,N_9793,N_5908);
or U12133 (N_12133,N_6092,N_8938);
nand U12134 (N_12134,N_7271,N_7553);
nand U12135 (N_12135,N_7800,N_6168);
and U12136 (N_12136,N_7731,N_5687);
nor U12137 (N_12137,N_6034,N_5901);
nor U12138 (N_12138,N_9102,N_8018);
nor U12139 (N_12139,N_7766,N_8732);
nand U12140 (N_12140,N_8237,N_7336);
xor U12141 (N_12141,N_5440,N_9768);
and U12142 (N_12142,N_6119,N_9471);
xnor U12143 (N_12143,N_9078,N_6417);
or U12144 (N_12144,N_5614,N_7703);
nand U12145 (N_12145,N_5558,N_7038);
and U12146 (N_12146,N_8846,N_6720);
or U12147 (N_12147,N_5641,N_6786);
nor U12148 (N_12148,N_8927,N_6640);
nand U12149 (N_12149,N_5309,N_5607);
nand U12150 (N_12150,N_6978,N_6447);
and U12151 (N_12151,N_8147,N_5083);
xnor U12152 (N_12152,N_8294,N_7110);
nor U12153 (N_12153,N_9530,N_8685);
nor U12154 (N_12154,N_9540,N_9087);
nand U12155 (N_12155,N_5889,N_8501);
and U12156 (N_12156,N_6561,N_5196);
nor U12157 (N_12157,N_7502,N_8377);
xnor U12158 (N_12158,N_6984,N_9146);
and U12159 (N_12159,N_5971,N_8724);
nand U12160 (N_12160,N_9330,N_6485);
xor U12161 (N_12161,N_9132,N_5590);
or U12162 (N_12162,N_6069,N_6070);
and U12163 (N_12163,N_5289,N_6824);
and U12164 (N_12164,N_5593,N_6091);
nor U12165 (N_12165,N_6182,N_7710);
xor U12166 (N_12166,N_9569,N_5375);
or U12167 (N_12167,N_9431,N_5526);
or U12168 (N_12168,N_9149,N_8590);
or U12169 (N_12169,N_7083,N_7645);
nor U12170 (N_12170,N_7061,N_7900);
nor U12171 (N_12171,N_8479,N_6600);
xor U12172 (N_12172,N_6361,N_6234);
xnor U12173 (N_12173,N_8452,N_7588);
and U12174 (N_12174,N_5428,N_7587);
xnor U12175 (N_12175,N_7516,N_8583);
nand U12176 (N_12176,N_7076,N_5132);
or U12177 (N_12177,N_9573,N_6754);
and U12178 (N_12178,N_9570,N_5713);
or U12179 (N_12179,N_7548,N_7194);
nand U12180 (N_12180,N_7063,N_7000);
and U12181 (N_12181,N_9628,N_8538);
or U12182 (N_12182,N_8611,N_6500);
or U12183 (N_12183,N_7383,N_7039);
and U12184 (N_12184,N_7604,N_8669);
and U12185 (N_12185,N_5667,N_6056);
or U12186 (N_12186,N_9955,N_8607);
nand U12187 (N_12187,N_8689,N_6207);
nand U12188 (N_12188,N_8066,N_9358);
and U12189 (N_12189,N_9685,N_7086);
or U12190 (N_12190,N_7923,N_5210);
or U12191 (N_12191,N_9895,N_5622);
nand U12192 (N_12192,N_9400,N_8430);
and U12193 (N_12193,N_5093,N_5963);
or U12194 (N_12194,N_7431,N_5063);
nor U12195 (N_12195,N_5915,N_7008);
xor U12196 (N_12196,N_6560,N_5225);
nor U12197 (N_12197,N_5074,N_9332);
nor U12198 (N_12198,N_5073,N_5751);
xnor U12199 (N_12199,N_5427,N_8899);
nand U12200 (N_12200,N_8257,N_8645);
nand U12201 (N_12201,N_5944,N_5847);
and U12202 (N_12202,N_7270,N_9343);
nor U12203 (N_12203,N_5651,N_5360);
xnor U12204 (N_12204,N_7804,N_9116);
nand U12205 (N_12205,N_6438,N_5239);
and U12206 (N_12206,N_8096,N_6669);
nor U12207 (N_12207,N_7028,N_9410);
xnor U12208 (N_12208,N_7255,N_8801);
and U12209 (N_12209,N_6364,N_6977);
nor U12210 (N_12210,N_7045,N_9621);
xor U12211 (N_12211,N_7300,N_5845);
xnor U12212 (N_12212,N_7594,N_5598);
xor U12213 (N_12213,N_7283,N_9309);
or U12214 (N_12214,N_9086,N_6876);
and U12215 (N_12215,N_9521,N_7101);
and U12216 (N_12216,N_6465,N_5934);
nand U12217 (N_12217,N_8705,N_7888);
or U12218 (N_12218,N_5793,N_9323);
and U12219 (N_12219,N_9462,N_6805);
nand U12220 (N_12220,N_5318,N_6532);
and U12221 (N_12221,N_9897,N_7342);
nor U12222 (N_12222,N_7788,N_6558);
nand U12223 (N_12223,N_5754,N_7582);
xnor U12224 (N_12224,N_6728,N_9803);
and U12225 (N_12225,N_6606,N_6855);
nor U12226 (N_12226,N_7940,N_5448);
or U12227 (N_12227,N_7455,N_5207);
xnor U12228 (N_12228,N_8807,N_9363);
or U12229 (N_12229,N_8825,N_9930);
or U12230 (N_12230,N_9789,N_5259);
nor U12231 (N_12231,N_7415,N_8353);
nand U12232 (N_12232,N_5199,N_6388);
nand U12233 (N_12233,N_7842,N_7200);
xnor U12234 (N_12234,N_8372,N_5567);
nor U12235 (N_12235,N_7937,N_6153);
nand U12236 (N_12236,N_8770,N_9094);
or U12237 (N_12237,N_5857,N_8432);
nand U12238 (N_12238,N_9204,N_6178);
or U12239 (N_12239,N_7673,N_6573);
xnor U12240 (N_12240,N_8536,N_9499);
and U12241 (N_12241,N_9526,N_6522);
or U12242 (N_12242,N_6031,N_5575);
nor U12243 (N_12243,N_5785,N_9997);
nor U12244 (N_12244,N_8657,N_9986);
or U12245 (N_12245,N_9411,N_6382);
nand U12246 (N_12246,N_6992,N_9487);
nor U12247 (N_12247,N_6286,N_7853);
or U12248 (N_12248,N_9592,N_7829);
xor U12249 (N_12249,N_5424,N_5442);
xor U12250 (N_12250,N_8894,N_9681);
or U12251 (N_12251,N_9528,N_5799);
and U12252 (N_12252,N_6169,N_6945);
and U12253 (N_12253,N_7576,N_9637);
or U12254 (N_12254,N_8254,N_7154);
and U12255 (N_12255,N_6317,N_5212);
nor U12256 (N_12256,N_7055,N_7108);
or U12257 (N_12257,N_8141,N_6456);
nand U12258 (N_12258,N_7723,N_5740);
nor U12259 (N_12259,N_9190,N_7770);
or U12260 (N_12260,N_5836,N_8965);
and U12261 (N_12261,N_9249,N_5247);
nor U12262 (N_12262,N_7116,N_8037);
or U12263 (N_12263,N_7639,N_9753);
nor U12264 (N_12264,N_5938,N_7185);
or U12265 (N_12265,N_7569,N_6098);
or U12266 (N_12266,N_6192,N_6816);
nor U12267 (N_12267,N_9463,N_9388);
nor U12268 (N_12268,N_9508,N_9417);
xnor U12269 (N_12269,N_9151,N_5091);
nand U12270 (N_12270,N_5124,N_6998);
and U12271 (N_12271,N_7867,N_8179);
nor U12272 (N_12272,N_8133,N_7382);
nand U12273 (N_12273,N_9338,N_6326);
nor U12274 (N_12274,N_6115,N_7020);
or U12275 (N_12275,N_6650,N_6542);
xnor U12276 (N_12276,N_7797,N_6063);
nand U12277 (N_12277,N_6959,N_6597);
or U12278 (N_12278,N_6122,N_9812);
nand U12279 (N_12279,N_9182,N_5150);
nor U12280 (N_12280,N_6386,N_5251);
xnor U12281 (N_12281,N_7965,N_7262);
nor U12282 (N_12282,N_5469,N_6269);
xor U12283 (N_12283,N_6067,N_7034);
nand U12284 (N_12284,N_7369,N_9612);
or U12285 (N_12285,N_9177,N_8991);
xor U12286 (N_12286,N_7658,N_5919);
and U12287 (N_12287,N_6320,N_5660);
xnor U12288 (N_12288,N_8956,N_9815);
or U12289 (N_12289,N_9558,N_8623);
nand U12290 (N_12290,N_9912,N_8262);
nor U12291 (N_12291,N_5965,N_7081);
nand U12292 (N_12292,N_7549,N_7697);
nor U12293 (N_12293,N_7840,N_9941);
nand U12294 (N_12294,N_7950,N_8922);
nand U12295 (N_12295,N_7424,N_9469);
nand U12296 (N_12296,N_5703,N_9485);
and U12297 (N_12297,N_5070,N_7475);
and U12298 (N_12298,N_6568,N_6329);
xor U12299 (N_12299,N_8250,N_6983);
and U12300 (N_12300,N_8548,N_5619);
nor U12301 (N_12301,N_5007,N_7509);
nor U12302 (N_12302,N_9928,N_9361);
xnor U12303 (N_12303,N_7269,N_9594);
xor U12304 (N_12304,N_7230,N_7450);
or U12305 (N_12305,N_8842,N_9137);
nor U12306 (N_12306,N_7019,N_8494);
xnor U12307 (N_12307,N_6137,N_8407);
nor U12308 (N_12308,N_5606,N_5559);
and U12309 (N_12309,N_9585,N_6293);
nor U12310 (N_12310,N_9751,N_7943);
nand U12311 (N_12311,N_8980,N_9588);
and U12312 (N_12312,N_6853,N_6448);
nand U12313 (N_12313,N_8493,N_7476);
xnor U12314 (N_12314,N_7241,N_7433);
and U12315 (N_12315,N_9015,N_8222);
nand U12316 (N_12316,N_7018,N_6046);
and U12317 (N_12317,N_8420,N_5055);
xnor U12318 (N_12318,N_7092,N_9051);
or U12319 (N_12319,N_7090,N_6262);
xnor U12320 (N_12320,N_7598,N_8671);
xor U12321 (N_12321,N_5088,N_8704);
nand U12322 (N_12322,N_9674,N_5485);
or U12323 (N_12323,N_9482,N_6113);
nor U12324 (N_12324,N_8889,N_6662);
xor U12325 (N_12325,N_6283,N_7203);
xnor U12326 (N_12326,N_6044,N_6949);
nor U12327 (N_12327,N_8378,N_5846);
or U12328 (N_12328,N_6791,N_7047);
or U12329 (N_12329,N_8052,N_5205);
and U12330 (N_12330,N_5727,N_9111);
nand U12331 (N_12331,N_5009,N_7413);
nand U12332 (N_12332,N_5782,N_7082);
and U12333 (N_12333,N_7459,N_9638);
and U12334 (N_12334,N_9673,N_6741);
and U12335 (N_12335,N_6499,N_8742);
xor U12336 (N_12336,N_9282,N_6390);
nor U12337 (N_12337,N_9886,N_8390);
nand U12338 (N_12338,N_9842,N_5929);
xor U12339 (N_12339,N_9972,N_6142);
xnor U12340 (N_12340,N_8916,N_7072);
or U12341 (N_12341,N_5067,N_8426);
nand U12342 (N_12342,N_8435,N_5684);
xor U12343 (N_12343,N_6379,N_7014);
nand U12344 (N_12344,N_6700,N_8368);
nor U12345 (N_12345,N_9054,N_8717);
nand U12346 (N_12346,N_7612,N_6872);
xnor U12347 (N_12347,N_7640,N_8882);
and U12348 (N_12348,N_6052,N_8038);
nor U12349 (N_12349,N_5039,N_5967);
and U12350 (N_12350,N_9044,N_5758);
nor U12351 (N_12351,N_5912,N_9687);
nand U12352 (N_12352,N_7279,N_8518);
xnor U12353 (N_12353,N_5630,N_8593);
xor U12354 (N_12354,N_8975,N_5605);
or U12355 (N_12355,N_9285,N_8911);
or U12356 (N_12356,N_6740,N_8067);
or U12357 (N_12357,N_7982,N_5829);
and U12358 (N_12358,N_8749,N_5244);
nand U12359 (N_12359,N_6711,N_8462);
nand U12360 (N_12360,N_8007,N_8276);
nor U12361 (N_12361,N_8236,N_9835);
nand U12362 (N_12362,N_7291,N_5596);
nand U12363 (N_12363,N_9134,N_6607);
nor U12364 (N_12364,N_7432,N_6841);
or U12365 (N_12365,N_9513,N_7540);
xor U12366 (N_12366,N_7786,N_7040);
and U12367 (N_12367,N_9502,N_5211);
or U12368 (N_12368,N_8563,N_7927);
and U12369 (N_12369,N_6212,N_8559);
nor U12370 (N_12370,N_6525,N_5886);
nor U12371 (N_12371,N_9228,N_5079);
or U12372 (N_12372,N_6862,N_5313);
nand U12373 (N_12373,N_5016,N_8031);
and U12374 (N_12374,N_5694,N_6396);
nor U12375 (N_12375,N_9004,N_8410);
xor U12376 (N_12376,N_9902,N_5617);
nor U12377 (N_12377,N_5084,N_6259);
xor U12378 (N_12378,N_7607,N_8274);
and U12379 (N_12379,N_7672,N_8111);
xor U12380 (N_12380,N_7036,N_7991);
nand U12381 (N_12381,N_8085,N_8945);
nand U12382 (N_12382,N_7621,N_9900);
and U12383 (N_12383,N_9728,N_8457);
or U12384 (N_12384,N_6627,N_6834);
xor U12385 (N_12385,N_9805,N_8551);
and U12386 (N_12386,N_9440,N_5935);
or U12387 (N_12387,N_7705,N_8064);
or U12388 (N_12388,N_6101,N_5556);
and U12389 (N_12389,N_8226,N_8161);
nor U12390 (N_12390,N_9742,N_6538);
nor U12391 (N_12391,N_9270,N_7733);
xnor U12392 (N_12392,N_5983,N_8459);
xnor U12393 (N_12393,N_7503,N_6400);
nand U12394 (N_12394,N_5514,N_5521);
and U12395 (N_12395,N_6174,N_5449);
xor U12396 (N_12396,N_7409,N_7439);
or U12397 (N_12397,N_6629,N_6324);
nand U12398 (N_12398,N_9205,N_8993);
and U12399 (N_12399,N_8456,N_5096);
or U12400 (N_12400,N_7754,N_7128);
or U12401 (N_12401,N_6626,N_5926);
xor U12402 (N_12402,N_7857,N_5624);
xnor U12403 (N_12403,N_8082,N_5802);
xnor U12404 (N_12404,N_7248,N_9457);
nor U12405 (N_12405,N_9016,N_8895);
nor U12406 (N_12406,N_9551,N_7630);
xor U12407 (N_12407,N_6649,N_5182);
nand U12408 (N_12408,N_5918,N_8782);
nor U12409 (N_12409,N_7483,N_6541);
and U12410 (N_12410,N_7882,N_7367);
nand U12411 (N_12411,N_7404,N_5535);
nor U12412 (N_12412,N_6112,N_8178);
nor U12413 (N_12413,N_8419,N_7401);
and U12414 (N_12414,N_8862,N_5006);
and U12415 (N_12415,N_8087,N_6384);
xor U12416 (N_12416,N_7904,N_7211);
xnor U12417 (N_12417,N_5275,N_7179);
xor U12418 (N_12418,N_5903,N_5378);
and U12419 (N_12419,N_6464,N_5760);
nand U12420 (N_12420,N_5403,N_8761);
nor U12421 (N_12421,N_8239,N_7868);
nor U12422 (N_12422,N_9794,N_9571);
nand U12423 (N_12423,N_8416,N_9397);
xnor U12424 (N_12424,N_5900,N_5089);
nor U12425 (N_12425,N_8112,N_5613);
or U12426 (N_12426,N_8998,N_6418);
nand U12427 (N_12427,N_8840,N_6674);
or U12428 (N_12428,N_9156,N_9489);
nand U12429 (N_12429,N_6282,N_5186);
xnor U12430 (N_12430,N_7227,N_8074);
or U12431 (N_12431,N_6440,N_6346);
and U12432 (N_12432,N_9257,N_6940);
nor U12433 (N_12433,N_9810,N_9716);
and U12434 (N_12434,N_6048,N_8543);
nor U12435 (N_12435,N_5071,N_9684);
nor U12436 (N_12436,N_6821,N_5322);
xnor U12437 (N_12437,N_5008,N_5549);
or U12438 (N_12438,N_5722,N_8107);
nand U12439 (N_12439,N_6393,N_6058);
and U12440 (N_12440,N_6005,N_7907);
nor U12441 (N_12441,N_8909,N_9454);
nand U12442 (N_12442,N_9736,N_7743);
and U12443 (N_12443,N_6254,N_6902);
nor U12444 (N_12444,N_6236,N_5922);
and U12445 (N_12445,N_7631,N_7029);
and U12446 (N_12446,N_9845,N_7095);
nor U12447 (N_12447,N_7094,N_5246);
nand U12448 (N_12448,N_6578,N_5338);
nand U12449 (N_12449,N_7399,N_7106);
and U12450 (N_12450,N_8722,N_8960);
or U12451 (N_12451,N_7798,N_5209);
and U12452 (N_12452,N_7794,N_6592);
and U12453 (N_12453,N_6201,N_6776);
xnor U12454 (N_12454,N_6094,N_7137);
and U12455 (N_12455,N_6655,N_9949);
and U12456 (N_12456,N_8641,N_8674);
nor U12457 (N_12457,N_6309,N_8346);
nor U12458 (N_12458,N_5094,N_6567);
xor U12459 (N_12459,N_7191,N_6859);
or U12460 (N_12460,N_9665,N_5195);
nand U12461 (N_12461,N_6854,N_6035);
nor U12462 (N_12462,N_5827,N_8371);
nor U12463 (N_12463,N_7877,N_5779);
nand U12464 (N_12464,N_7292,N_6277);
nor U12465 (N_12465,N_9153,N_6848);
or U12466 (N_12466,N_7718,N_8429);
nor U12467 (N_12467,N_5024,N_5121);
xnor U12468 (N_12468,N_9652,N_5082);
nor U12469 (N_12469,N_7663,N_8174);
and U12470 (N_12470,N_7964,N_8057);
nand U12471 (N_12471,N_8736,N_8581);
nand U12472 (N_12472,N_6179,N_8834);
nor U12473 (N_12473,N_7234,N_5506);
nand U12474 (N_12474,N_5729,N_5943);
and U12475 (N_12475,N_7214,N_5455);
or U12476 (N_12476,N_8449,N_9632);
or U12477 (N_12477,N_8575,N_5386);
or U12478 (N_12478,N_9467,N_5812);
nand U12479 (N_12479,N_7454,N_9197);
or U12480 (N_12480,N_9848,N_5826);
or U12481 (N_12481,N_8489,N_5552);
and U12482 (N_12482,N_7276,N_9083);
or U12483 (N_12483,N_9544,N_9071);
nand U12484 (N_12484,N_6715,N_6060);
and U12485 (N_12485,N_5665,N_7911);
xor U12486 (N_12486,N_8084,N_6602);
nor U12487 (N_12487,N_7418,N_8340);
xor U12488 (N_12488,N_5797,N_7533);
or U12489 (N_12489,N_8809,N_8639);
xnor U12490 (N_12490,N_7642,N_6062);
nand U12491 (N_12491,N_8100,N_5541);
or U12492 (N_12492,N_8131,N_5304);
xor U12493 (N_12493,N_5657,N_5803);
nand U12494 (N_12494,N_5577,N_6946);
nor U12495 (N_12495,N_7356,N_5077);
nor U12496 (N_12496,N_7051,N_8727);
or U12497 (N_12497,N_7599,N_5236);
nand U12498 (N_12498,N_6648,N_9821);
nand U12499 (N_12499,N_5013,N_6124);
and U12500 (N_12500,N_6243,N_8202);
nor U12501 (N_12501,N_5089,N_6828);
nor U12502 (N_12502,N_6157,N_7497);
nand U12503 (N_12503,N_8306,N_6259);
and U12504 (N_12504,N_6761,N_6408);
and U12505 (N_12505,N_5679,N_7007);
nor U12506 (N_12506,N_8340,N_7157);
nand U12507 (N_12507,N_5401,N_5855);
nor U12508 (N_12508,N_9950,N_6340);
nor U12509 (N_12509,N_5756,N_9917);
nor U12510 (N_12510,N_9180,N_5222);
xor U12511 (N_12511,N_6660,N_7642);
nand U12512 (N_12512,N_5913,N_9144);
or U12513 (N_12513,N_5782,N_7445);
xor U12514 (N_12514,N_9672,N_8569);
or U12515 (N_12515,N_5214,N_9158);
and U12516 (N_12516,N_5828,N_5148);
or U12517 (N_12517,N_7419,N_9536);
nor U12518 (N_12518,N_7574,N_7600);
and U12519 (N_12519,N_8518,N_9684);
nor U12520 (N_12520,N_7375,N_5725);
nand U12521 (N_12521,N_5697,N_9812);
nor U12522 (N_12522,N_8097,N_8275);
or U12523 (N_12523,N_8333,N_8057);
nor U12524 (N_12524,N_6315,N_9449);
xnor U12525 (N_12525,N_7095,N_5335);
nand U12526 (N_12526,N_5925,N_5678);
xnor U12527 (N_12527,N_7023,N_6577);
xor U12528 (N_12528,N_6396,N_8377);
xnor U12529 (N_12529,N_6968,N_6521);
xor U12530 (N_12530,N_8443,N_6566);
nor U12531 (N_12531,N_9968,N_8899);
nand U12532 (N_12532,N_5857,N_5635);
and U12533 (N_12533,N_7133,N_8347);
nand U12534 (N_12534,N_6450,N_5808);
nand U12535 (N_12535,N_7685,N_8749);
nor U12536 (N_12536,N_9261,N_9729);
nor U12537 (N_12537,N_8138,N_5132);
nand U12538 (N_12538,N_8312,N_8263);
xor U12539 (N_12539,N_6471,N_8307);
nand U12540 (N_12540,N_8341,N_8761);
nor U12541 (N_12541,N_7193,N_9820);
nand U12542 (N_12542,N_6311,N_5861);
or U12543 (N_12543,N_8439,N_9464);
nand U12544 (N_12544,N_6051,N_9674);
nor U12545 (N_12545,N_7303,N_9625);
and U12546 (N_12546,N_9141,N_6404);
nor U12547 (N_12547,N_7911,N_9522);
xor U12548 (N_12548,N_5439,N_9832);
and U12549 (N_12549,N_9729,N_7858);
nand U12550 (N_12550,N_7496,N_9577);
nand U12551 (N_12551,N_8406,N_7455);
nand U12552 (N_12552,N_6331,N_7030);
nor U12553 (N_12553,N_8532,N_5163);
and U12554 (N_12554,N_7855,N_5689);
nor U12555 (N_12555,N_5208,N_8782);
or U12556 (N_12556,N_9838,N_9511);
and U12557 (N_12557,N_9174,N_7441);
or U12558 (N_12558,N_8241,N_8479);
and U12559 (N_12559,N_7269,N_7610);
nand U12560 (N_12560,N_7076,N_8783);
or U12561 (N_12561,N_8223,N_9965);
xnor U12562 (N_12562,N_9093,N_5965);
xor U12563 (N_12563,N_7829,N_9923);
or U12564 (N_12564,N_8171,N_5883);
nand U12565 (N_12565,N_8757,N_7863);
xor U12566 (N_12566,N_6444,N_5916);
or U12567 (N_12567,N_5821,N_9973);
nor U12568 (N_12568,N_6009,N_5915);
and U12569 (N_12569,N_5126,N_5805);
xnor U12570 (N_12570,N_8489,N_5794);
or U12571 (N_12571,N_9458,N_7789);
and U12572 (N_12572,N_8511,N_6880);
nor U12573 (N_12573,N_7819,N_9722);
and U12574 (N_12574,N_7784,N_5874);
xor U12575 (N_12575,N_7876,N_6497);
and U12576 (N_12576,N_9812,N_6929);
or U12577 (N_12577,N_6246,N_5060);
and U12578 (N_12578,N_9371,N_9962);
xor U12579 (N_12579,N_8185,N_7761);
nand U12580 (N_12580,N_9508,N_8907);
and U12581 (N_12581,N_7205,N_6038);
xor U12582 (N_12582,N_9880,N_9183);
or U12583 (N_12583,N_9844,N_7591);
or U12584 (N_12584,N_5492,N_7906);
xor U12585 (N_12585,N_5611,N_6545);
or U12586 (N_12586,N_6538,N_5705);
and U12587 (N_12587,N_5250,N_6860);
xnor U12588 (N_12588,N_7097,N_6361);
and U12589 (N_12589,N_8651,N_9673);
nand U12590 (N_12590,N_8638,N_7437);
xor U12591 (N_12591,N_6813,N_9602);
xnor U12592 (N_12592,N_9997,N_5443);
nand U12593 (N_12593,N_5352,N_9487);
xnor U12594 (N_12594,N_9808,N_7868);
nor U12595 (N_12595,N_9839,N_9116);
nand U12596 (N_12596,N_7734,N_7473);
nor U12597 (N_12597,N_9694,N_7859);
or U12598 (N_12598,N_5415,N_8580);
or U12599 (N_12599,N_8762,N_6282);
and U12600 (N_12600,N_6601,N_5627);
nor U12601 (N_12601,N_9139,N_7439);
nor U12602 (N_12602,N_5131,N_5924);
or U12603 (N_12603,N_5183,N_7602);
or U12604 (N_12604,N_5450,N_5932);
nand U12605 (N_12605,N_8286,N_6452);
or U12606 (N_12606,N_6514,N_7227);
xor U12607 (N_12607,N_5292,N_7506);
nor U12608 (N_12608,N_6929,N_6253);
nor U12609 (N_12609,N_5617,N_7687);
and U12610 (N_12610,N_9378,N_6589);
and U12611 (N_12611,N_6815,N_6585);
and U12612 (N_12612,N_7261,N_9636);
nand U12613 (N_12613,N_8030,N_9706);
or U12614 (N_12614,N_5230,N_6869);
xor U12615 (N_12615,N_8931,N_5985);
nor U12616 (N_12616,N_5241,N_9712);
xnor U12617 (N_12617,N_6179,N_6726);
nand U12618 (N_12618,N_9230,N_6855);
xor U12619 (N_12619,N_6950,N_5316);
xor U12620 (N_12620,N_5671,N_8353);
xor U12621 (N_12621,N_6713,N_8632);
nor U12622 (N_12622,N_7643,N_8984);
nand U12623 (N_12623,N_8032,N_9849);
and U12624 (N_12624,N_7590,N_8573);
nor U12625 (N_12625,N_8704,N_7851);
or U12626 (N_12626,N_9604,N_9572);
nand U12627 (N_12627,N_5130,N_5081);
nand U12628 (N_12628,N_8343,N_8122);
nand U12629 (N_12629,N_5779,N_8971);
xnor U12630 (N_12630,N_7488,N_5818);
nand U12631 (N_12631,N_8905,N_9858);
xor U12632 (N_12632,N_9641,N_7110);
or U12633 (N_12633,N_6922,N_7354);
xnor U12634 (N_12634,N_9763,N_7734);
nand U12635 (N_12635,N_5248,N_5500);
nor U12636 (N_12636,N_8136,N_8945);
nor U12637 (N_12637,N_6972,N_9073);
nand U12638 (N_12638,N_8019,N_7877);
nand U12639 (N_12639,N_6864,N_9852);
and U12640 (N_12640,N_6558,N_7858);
nand U12641 (N_12641,N_8605,N_7231);
xnor U12642 (N_12642,N_5249,N_8969);
nor U12643 (N_12643,N_9683,N_7239);
nor U12644 (N_12644,N_8671,N_8323);
nor U12645 (N_12645,N_9893,N_5905);
xnor U12646 (N_12646,N_9417,N_6850);
and U12647 (N_12647,N_8281,N_9242);
xnor U12648 (N_12648,N_7909,N_6243);
or U12649 (N_12649,N_9587,N_8939);
and U12650 (N_12650,N_8032,N_8297);
nand U12651 (N_12651,N_8451,N_8620);
and U12652 (N_12652,N_6752,N_9947);
xnor U12653 (N_12653,N_9735,N_8525);
nor U12654 (N_12654,N_5536,N_9586);
nand U12655 (N_12655,N_6445,N_7847);
or U12656 (N_12656,N_9633,N_9012);
and U12657 (N_12657,N_9650,N_8956);
nand U12658 (N_12658,N_8913,N_7866);
nor U12659 (N_12659,N_6780,N_9477);
or U12660 (N_12660,N_9509,N_7083);
nor U12661 (N_12661,N_5350,N_9359);
xor U12662 (N_12662,N_9559,N_8442);
nor U12663 (N_12663,N_8339,N_7430);
or U12664 (N_12664,N_5720,N_6320);
or U12665 (N_12665,N_7396,N_8387);
or U12666 (N_12666,N_9430,N_5740);
xnor U12667 (N_12667,N_6018,N_6111);
or U12668 (N_12668,N_8006,N_5503);
and U12669 (N_12669,N_5369,N_8351);
xor U12670 (N_12670,N_6669,N_9222);
nor U12671 (N_12671,N_7163,N_8386);
and U12672 (N_12672,N_8890,N_8203);
xor U12673 (N_12673,N_8029,N_6334);
nand U12674 (N_12674,N_5783,N_8053);
and U12675 (N_12675,N_6036,N_5570);
xor U12676 (N_12676,N_5557,N_5072);
xor U12677 (N_12677,N_9463,N_8643);
xnor U12678 (N_12678,N_8707,N_5254);
and U12679 (N_12679,N_7358,N_9220);
xnor U12680 (N_12680,N_7093,N_9083);
or U12681 (N_12681,N_8545,N_6976);
nor U12682 (N_12682,N_8620,N_6444);
xnor U12683 (N_12683,N_9104,N_5607);
xor U12684 (N_12684,N_6997,N_6871);
or U12685 (N_12685,N_9827,N_7383);
or U12686 (N_12686,N_9922,N_7971);
nand U12687 (N_12687,N_8562,N_8631);
xnor U12688 (N_12688,N_5362,N_5386);
nor U12689 (N_12689,N_8648,N_6410);
or U12690 (N_12690,N_9220,N_9518);
nand U12691 (N_12691,N_7923,N_9730);
xnor U12692 (N_12692,N_5004,N_9992);
and U12693 (N_12693,N_6344,N_7666);
nor U12694 (N_12694,N_5541,N_5586);
and U12695 (N_12695,N_9025,N_9634);
xor U12696 (N_12696,N_8750,N_7583);
nor U12697 (N_12697,N_8217,N_9368);
xor U12698 (N_12698,N_9026,N_8112);
nor U12699 (N_12699,N_9846,N_8104);
or U12700 (N_12700,N_8116,N_9190);
or U12701 (N_12701,N_7475,N_5531);
xor U12702 (N_12702,N_8139,N_7995);
xnor U12703 (N_12703,N_6054,N_5987);
xor U12704 (N_12704,N_6954,N_5611);
nor U12705 (N_12705,N_5069,N_6459);
nand U12706 (N_12706,N_6682,N_8476);
or U12707 (N_12707,N_9227,N_5843);
nand U12708 (N_12708,N_6123,N_8448);
and U12709 (N_12709,N_9227,N_6778);
or U12710 (N_12710,N_8510,N_6117);
nand U12711 (N_12711,N_6762,N_7905);
and U12712 (N_12712,N_7901,N_5335);
xor U12713 (N_12713,N_6285,N_9498);
xor U12714 (N_12714,N_6176,N_6102);
or U12715 (N_12715,N_9537,N_7598);
nand U12716 (N_12716,N_8328,N_7949);
or U12717 (N_12717,N_6200,N_6367);
and U12718 (N_12718,N_5613,N_7675);
or U12719 (N_12719,N_8284,N_5419);
and U12720 (N_12720,N_8622,N_7833);
xor U12721 (N_12721,N_7613,N_5535);
nor U12722 (N_12722,N_6193,N_6254);
nor U12723 (N_12723,N_5768,N_8191);
and U12724 (N_12724,N_9394,N_6498);
and U12725 (N_12725,N_9956,N_5405);
xor U12726 (N_12726,N_6563,N_6997);
nand U12727 (N_12727,N_5208,N_6251);
nand U12728 (N_12728,N_6495,N_6423);
nor U12729 (N_12729,N_9709,N_7900);
and U12730 (N_12730,N_9015,N_8460);
nor U12731 (N_12731,N_7865,N_8790);
and U12732 (N_12732,N_5233,N_5435);
nand U12733 (N_12733,N_8635,N_8463);
nor U12734 (N_12734,N_6492,N_5246);
xnor U12735 (N_12735,N_9637,N_6029);
xor U12736 (N_12736,N_7079,N_5044);
and U12737 (N_12737,N_6206,N_8612);
and U12738 (N_12738,N_7431,N_8652);
and U12739 (N_12739,N_6409,N_6207);
nand U12740 (N_12740,N_6172,N_7863);
nand U12741 (N_12741,N_6393,N_8137);
and U12742 (N_12742,N_6770,N_6889);
nor U12743 (N_12743,N_9404,N_6135);
or U12744 (N_12744,N_9104,N_6852);
nand U12745 (N_12745,N_9857,N_8443);
nor U12746 (N_12746,N_6190,N_6821);
nand U12747 (N_12747,N_9710,N_7221);
xnor U12748 (N_12748,N_5681,N_7727);
and U12749 (N_12749,N_5319,N_6477);
and U12750 (N_12750,N_5466,N_8538);
nand U12751 (N_12751,N_6131,N_8685);
or U12752 (N_12752,N_7466,N_7990);
nor U12753 (N_12753,N_8943,N_6876);
or U12754 (N_12754,N_9606,N_7981);
nor U12755 (N_12755,N_7254,N_6962);
or U12756 (N_12756,N_6511,N_9422);
or U12757 (N_12757,N_6206,N_9471);
xnor U12758 (N_12758,N_9393,N_8363);
and U12759 (N_12759,N_5361,N_7557);
and U12760 (N_12760,N_5971,N_6660);
nand U12761 (N_12761,N_9410,N_5959);
nor U12762 (N_12762,N_7937,N_7327);
nand U12763 (N_12763,N_7389,N_8707);
xnor U12764 (N_12764,N_9190,N_9159);
nor U12765 (N_12765,N_9533,N_8705);
xnor U12766 (N_12766,N_7093,N_5005);
nand U12767 (N_12767,N_5228,N_9913);
nand U12768 (N_12768,N_8449,N_8658);
xnor U12769 (N_12769,N_5020,N_6092);
and U12770 (N_12770,N_6589,N_9521);
nand U12771 (N_12771,N_7333,N_7314);
nand U12772 (N_12772,N_9040,N_5340);
or U12773 (N_12773,N_9094,N_7063);
nand U12774 (N_12774,N_8537,N_8688);
nand U12775 (N_12775,N_9345,N_9435);
nand U12776 (N_12776,N_6603,N_7765);
and U12777 (N_12777,N_9776,N_6451);
or U12778 (N_12778,N_7315,N_8619);
or U12779 (N_12779,N_7888,N_9497);
and U12780 (N_12780,N_8444,N_8172);
or U12781 (N_12781,N_7512,N_8745);
and U12782 (N_12782,N_9708,N_5397);
or U12783 (N_12783,N_6056,N_6834);
or U12784 (N_12784,N_6822,N_9879);
nor U12785 (N_12785,N_9254,N_5691);
and U12786 (N_12786,N_9000,N_8066);
nor U12787 (N_12787,N_7524,N_9141);
nand U12788 (N_12788,N_6210,N_5003);
nor U12789 (N_12789,N_7699,N_8089);
nand U12790 (N_12790,N_7211,N_8632);
and U12791 (N_12791,N_8390,N_8683);
or U12792 (N_12792,N_9974,N_8515);
and U12793 (N_12793,N_5366,N_9277);
xor U12794 (N_12794,N_5419,N_5303);
or U12795 (N_12795,N_7521,N_7509);
or U12796 (N_12796,N_6196,N_6979);
nand U12797 (N_12797,N_9517,N_7646);
xnor U12798 (N_12798,N_5816,N_9879);
xor U12799 (N_12799,N_7426,N_7184);
nand U12800 (N_12800,N_7846,N_9338);
or U12801 (N_12801,N_6111,N_7130);
and U12802 (N_12802,N_9331,N_8637);
and U12803 (N_12803,N_7647,N_8370);
and U12804 (N_12804,N_5025,N_8513);
nor U12805 (N_12805,N_7279,N_5049);
xor U12806 (N_12806,N_7289,N_7180);
xnor U12807 (N_12807,N_9750,N_9245);
nand U12808 (N_12808,N_9218,N_7215);
nand U12809 (N_12809,N_8496,N_9394);
and U12810 (N_12810,N_5204,N_8130);
and U12811 (N_12811,N_5426,N_8482);
xor U12812 (N_12812,N_9159,N_6110);
nor U12813 (N_12813,N_6447,N_9360);
xor U12814 (N_12814,N_7835,N_6039);
and U12815 (N_12815,N_8374,N_8162);
xor U12816 (N_12816,N_7493,N_9836);
nand U12817 (N_12817,N_5404,N_8075);
nand U12818 (N_12818,N_9696,N_9727);
xnor U12819 (N_12819,N_7240,N_5013);
xor U12820 (N_12820,N_6248,N_8172);
xor U12821 (N_12821,N_8225,N_7296);
and U12822 (N_12822,N_9934,N_6176);
and U12823 (N_12823,N_8931,N_9886);
nor U12824 (N_12824,N_9347,N_8133);
xor U12825 (N_12825,N_6152,N_9093);
and U12826 (N_12826,N_7409,N_7872);
and U12827 (N_12827,N_9160,N_5162);
and U12828 (N_12828,N_5193,N_8998);
nand U12829 (N_12829,N_7468,N_8536);
and U12830 (N_12830,N_9284,N_8044);
or U12831 (N_12831,N_7673,N_6267);
nand U12832 (N_12832,N_6662,N_5882);
nor U12833 (N_12833,N_6653,N_9537);
nand U12834 (N_12834,N_7492,N_8557);
xor U12835 (N_12835,N_7354,N_9695);
or U12836 (N_12836,N_5975,N_6704);
xor U12837 (N_12837,N_5180,N_8852);
nand U12838 (N_12838,N_6113,N_7304);
nor U12839 (N_12839,N_5681,N_7391);
nor U12840 (N_12840,N_9781,N_8307);
or U12841 (N_12841,N_8860,N_7608);
nand U12842 (N_12842,N_5825,N_7430);
nor U12843 (N_12843,N_9911,N_6051);
nor U12844 (N_12844,N_8465,N_8400);
xnor U12845 (N_12845,N_8002,N_7647);
xor U12846 (N_12846,N_7722,N_9046);
xnor U12847 (N_12847,N_9042,N_8762);
or U12848 (N_12848,N_7699,N_5043);
and U12849 (N_12849,N_7416,N_6032);
nand U12850 (N_12850,N_7215,N_9636);
or U12851 (N_12851,N_6637,N_7796);
or U12852 (N_12852,N_7166,N_5735);
nor U12853 (N_12853,N_5965,N_9007);
nand U12854 (N_12854,N_9277,N_6975);
nand U12855 (N_12855,N_9903,N_5302);
or U12856 (N_12856,N_6296,N_7097);
xor U12857 (N_12857,N_6204,N_7415);
nor U12858 (N_12858,N_7050,N_8481);
nor U12859 (N_12859,N_9984,N_7977);
xor U12860 (N_12860,N_5185,N_9973);
or U12861 (N_12861,N_6681,N_6982);
nand U12862 (N_12862,N_7219,N_6942);
xor U12863 (N_12863,N_9438,N_8060);
nor U12864 (N_12864,N_7588,N_8034);
nand U12865 (N_12865,N_5353,N_7049);
or U12866 (N_12866,N_6568,N_9420);
and U12867 (N_12867,N_7117,N_7781);
or U12868 (N_12868,N_8942,N_6336);
nor U12869 (N_12869,N_6444,N_8899);
or U12870 (N_12870,N_8984,N_6653);
nor U12871 (N_12871,N_7257,N_8256);
xor U12872 (N_12872,N_6343,N_6419);
nand U12873 (N_12873,N_5686,N_7043);
nand U12874 (N_12874,N_7909,N_5694);
and U12875 (N_12875,N_8482,N_8559);
xnor U12876 (N_12876,N_8414,N_7576);
nand U12877 (N_12877,N_6623,N_5871);
nor U12878 (N_12878,N_8376,N_6298);
nand U12879 (N_12879,N_8684,N_8740);
nor U12880 (N_12880,N_6558,N_6587);
and U12881 (N_12881,N_6877,N_6408);
or U12882 (N_12882,N_8273,N_9169);
xor U12883 (N_12883,N_6981,N_9127);
nor U12884 (N_12884,N_6647,N_6093);
xor U12885 (N_12885,N_7269,N_6613);
or U12886 (N_12886,N_8597,N_8541);
nor U12887 (N_12887,N_7448,N_7159);
nor U12888 (N_12888,N_9255,N_5786);
nor U12889 (N_12889,N_7136,N_8472);
or U12890 (N_12890,N_5760,N_9787);
or U12891 (N_12891,N_5197,N_7825);
nor U12892 (N_12892,N_5059,N_9712);
nor U12893 (N_12893,N_9742,N_6197);
nand U12894 (N_12894,N_5170,N_9492);
nor U12895 (N_12895,N_7440,N_9399);
or U12896 (N_12896,N_7856,N_5275);
xnor U12897 (N_12897,N_5339,N_8514);
nand U12898 (N_12898,N_5417,N_6774);
xor U12899 (N_12899,N_8867,N_6648);
nor U12900 (N_12900,N_6595,N_8978);
xor U12901 (N_12901,N_5859,N_7963);
and U12902 (N_12902,N_8141,N_6810);
nor U12903 (N_12903,N_7746,N_9938);
and U12904 (N_12904,N_5922,N_8068);
xor U12905 (N_12905,N_5939,N_8331);
and U12906 (N_12906,N_7651,N_6591);
and U12907 (N_12907,N_6649,N_5099);
or U12908 (N_12908,N_7160,N_8753);
nand U12909 (N_12909,N_6209,N_9558);
nor U12910 (N_12910,N_8811,N_7215);
nor U12911 (N_12911,N_7621,N_6731);
or U12912 (N_12912,N_8711,N_8862);
and U12913 (N_12913,N_9403,N_9314);
nand U12914 (N_12914,N_6807,N_7442);
and U12915 (N_12915,N_7280,N_9643);
xor U12916 (N_12916,N_6865,N_7366);
nor U12917 (N_12917,N_5336,N_7073);
nand U12918 (N_12918,N_7526,N_5054);
nor U12919 (N_12919,N_6973,N_9306);
nand U12920 (N_12920,N_8026,N_9443);
or U12921 (N_12921,N_9147,N_6215);
nand U12922 (N_12922,N_6653,N_5344);
nand U12923 (N_12923,N_6625,N_7085);
and U12924 (N_12924,N_8231,N_7911);
or U12925 (N_12925,N_9556,N_9002);
nor U12926 (N_12926,N_9601,N_6159);
or U12927 (N_12927,N_5137,N_5053);
nor U12928 (N_12928,N_7348,N_6408);
xor U12929 (N_12929,N_5344,N_6431);
xor U12930 (N_12930,N_6478,N_5122);
nand U12931 (N_12931,N_5609,N_6639);
xor U12932 (N_12932,N_7284,N_7360);
and U12933 (N_12933,N_5221,N_8069);
nand U12934 (N_12934,N_9977,N_8184);
nor U12935 (N_12935,N_8009,N_8948);
or U12936 (N_12936,N_8039,N_8491);
or U12937 (N_12937,N_6075,N_6719);
nor U12938 (N_12938,N_5487,N_5769);
xnor U12939 (N_12939,N_8316,N_7150);
xnor U12940 (N_12940,N_8126,N_8972);
or U12941 (N_12941,N_9669,N_8230);
nor U12942 (N_12942,N_8047,N_5002);
nand U12943 (N_12943,N_7590,N_5747);
nand U12944 (N_12944,N_9497,N_8065);
or U12945 (N_12945,N_6460,N_9681);
or U12946 (N_12946,N_7002,N_8227);
or U12947 (N_12947,N_8540,N_7520);
or U12948 (N_12948,N_7367,N_6432);
or U12949 (N_12949,N_5147,N_9756);
and U12950 (N_12950,N_7022,N_8380);
and U12951 (N_12951,N_7269,N_6076);
or U12952 (N_12952,N_8749,N_8706);
xor U12953 (N_12953,N_5395,N_9971);
nor U12954 (N_12954,N_8152,N_6428);
xor U12955 (N_12955,N_8227,N_8722);
and U12956 (N_12956,N_7513,N_8288);
nand U12957 (N_12957,N_7964,N_6916);
nor U12958 (N_12958,N_7143,N_9317);
nor U12959 (N_12959,N_7251,N_5584);
or U12960 (N_12960,N_6796,N_6366);
or U12961 (N_12961,N_9433,N_6381);
or U12962 (N_12962,N_8820,N_9457);
and U12963 (N_12963,N_7452,N_6630);
nand U12964 (N_12964,N_5297,N_9095);
nor U12965 (N_12965,N_6161,N_7833);
xor U12966 (N_12966,N_8048,N_5339);
and U12967 (N_12967,N_5146,N_9137);
xnor U12968 (N_12968,N_9380,N_6363);
and U12969 (N_12969,N_5771,N_6921);
nor U12970 (N_12970,N_7405,N_8765);
xor U12971 (N_12971,N_8027,N_8611);
nor U12972 (N_12972,N_7860,N_6427);
or U12973 (N_12973,N_9478,N_5448);
nor U12974 (N_12974,N_5531,N_7029);
nand U12975 (N_12975,N_5162,N_7044);
xnor U12976 (N_12976,N_6791,N_7791);
or U12977 (N_12977,N_5232,N_7953);
nand U12978 (N_12978,N_7234,N_9655);
xor U12979 (N_12979,N_8371,N_8904);
nand U12980 (N_12980,N_7972,N_5877);
xor U12981 (N_12981,N_6592,N_5672);
or U12982 (N_12982,N_9133,N_6201);
nand U12983 (N_12983,N_8534,N_6594);
and U12984 (N_12984,N_9668,N_6713);
or U12985 (N_12985,N_8292,N_7490);
nor U12986 (N_12986,N_9656,N_7025);
nand U12987 (N_12987,N_8948,N_8283);
and U12988 (N_12988,N_6529,N_9750);
nand U12989 (N_12989,N_7283,N_5864);
nand U12990 (N_12990,N_5578,N_5428);
xnor U12991 (N_12991,N_8305,N_6312);
nand U12992 (N_12992,N_8249,N_7753);
nor U12993 (N_12993,N_6946,N_8742);
nand U12994 (N_12994,N_6895,N_9698);
or U12995 (N_12995,N_7652,N_7525);
and U12996 (N_12996,N_8123,N_5203);
or U12997 (N_12997,N_8993,N_8412);
or U12998 (N_12998,N_6298,N_9334);
xnor U12999 (N_12999,N_7954,N_7574);
nor U13000 (N_13000,N_9456,N_5408);
and U13001 (N_13001,N_8417,N_5407);
xnor U13002 (N_13002,N_8002,N_9694);
and U13003 (N_13003,N_5395,N_9344);
nand U13004 (N_13004,N_6517,N_9140);
and U13005 (N_13005,N_7934,N_7588);
nand U13006 (N_13006,N_7910,N_7979);
and U13007 (N_13007,N_9064,N_8646);
xnor U13008 (N_13008,N_8675,N_8147);
nor U13009 (N_13009,N_5589,N_9051);
or U13010 (N_13010,N_9523,N_5328);
and U13011 (N_13011,N_6754,N_9514);
or U13012 (N_13012,N_6408,N_5808);
nand U13013 (N_13013,N_9339,N_7457);
and U13014 (N_13014,N_9086,N_6517);
and U13015 (N_13015,N_7021,N_8084);
or U13016 (N_13016,N_6966,N_9340);
nand U13017 (N_13017,N_5144,N_5553);
or U13018 (N_13018,N_7023,N_5089);
and U13019 (N_13019,N_5216,N_6830);
nand U13020 (N_13020,N_7416,N_5424);
nor U13021 (N_13021,N_9939,N_5196);
xnor U13022 (N_13022,N_8592,N_5128);
nor U13023 (N_13023,N_9156,N_6856);
or U13024 (N_13024,N_5893,N_7717);
nand U13025 (N_13025,N_7069,N_5516);
xnor U13026 (N_13026,N_7936,N_8164);
and U13027 (N_13027,N_8239,N_8269);
xnor U13028 (N_13028,N_5155,N_6312);
nor U13029 (N_13029,N_6221,N_8999);
nor U13030 (N_13030,N_9253,N_6047);
nor U13031 (N_13031,N_6739,N_9524);
or U13032 (N_13032,N_6716,N_9446);
or U13033 (N_13033,N_7650,N_5633);
nor U13034 (N_13034,N_9960,N_8427);
or U13035 (N_13035,N_5148,N_9066);
nand U13036 (N_13036,N_5919,N_9203);
nor U13037 (N_13037,N_8461,N_9978);
nand U13038 (N_13038,N_7660,N_7976);
xor U13039 (N_13039,N_6579,N_8775);
and U13040 (N_13040,N_7802,N_8253);
nand U13041 (N_13041,N_6504,N_9557);
xnor U13042 (N_13042,N_8870,N_8693);
and U13043 (N_13043,N_7645,N_8363);
nor U13044 (N_13044,N_6456,N_7590);
nand U13045 (N_13045,N_6693,N_8141);
xnor U13046 (N_13046,N_6044,N_9961);
nand U13047 (N_13047,N_8749,N_9912);
nor U13048 (N_13048,N_8887,N_9048);
nand U13049 (N_13049,N_8639,N_6379);
nand U13050 (N_13050,N_6090,N_9137);
and U13051 (N_13051,N_5403,N_7856);
xnor U13052 (N_13052,N_5248,N_8148);
and U13053 (N_13053,N_9740,N_9868);
nor U13054 (N_13054,N_6687,N_9418);
nor U13055 (N_13055,N_9420,N_7114);
or U13056 (N_13056,N_8837,N_5076);
xnor U13057 (N_13057,N_9919,N_6655);
and U13058 (N_13058,N_5115,N_8774);
nor U13059 (N_13059,N_5024,N_7292);
nand U13060 (N_13060,N_5376,N_9726);
xor U13061 (N_13061,N_6440,N_8675);
nand U13062 (N_13062,N_9791,N_8064);
nor U13063 (N_13063,N_8834,N_9927);
and U13064 (N_13064,N_6439,N_7117);
and U13065 (N_13065,N_7288,N_8168);
or U13066 (N_13066,N_8171,N_6089);
or U13067 (N_13067,N_8361,N_7705);
or U13068 (N_13068,N_7254,N_6509);
or U13069 (N_13069,N_7479,N_8931);
nor U13070 (N_13070,N_7276,N_7588);
or U13071 (N_13071,N_5924,N_7449);
or U13072 (N_13072,N_6738,N_7877);
or U13073 (N_13073,N_6805,N_8674);
or U13074 (N_13074,N_9054,N_7300);
nor U13075 (N_13075,N_5404,N_9202);
nor U13076 (N_13076,N_6293,N_8286);
and U13077 (N_13077,N_8702,N_8817);
xnor U13078 (N_13078,N_5943,N_7273);
nand U13079 (N_13079,N_7237,N_5185);
xnor U13080 (N_13080,N_6127,N_8844);
nor U13081 (N_13081,N_6688,N_9749);
nand U13082 (N_13082,N_8500,N_8327);
nor U13083 (N_13083,N_7340,N_5709);
and U13084 (N_13084,N_9012,N_9227);
and U13085 (N_13085,N_7515,N_7209);
and U13086 (N_13086,N_8408,N_7707);
xor U13087 (N_13087,N_6394,N_7036);
and U13088 (N_13088,N_5470,N_8246);
xor U13089 (N_13089,N_8047,N_9974);
xnor U13090 (N_13090,N_9346,N_5589);
or U13091 (N_13091,N_7970,N_5525);
nand U13092 (N_13092,N_7349,N_6805);
or U13093 (N_13093,N_6981,N_6257);
or U13094 (N_13094,N_8332,N_6904);
nand U13095 (N_13095,N_8058,N_9650);
and U13096 (N_13096,N_6640,N_5517);
xnor U13097 (N_13097,N_7874,N_9186);
and U13098 (N_13098,N_5171,N_5174);
and U13099 (N_13099,N_6309,N_9574);
and U13100 (N_13100,N_6981,N_9660);
nand U13101 (N_13101,N_6519,N_5262);
xnor U13102 (N_13102,N_5927,N_7945);
xnor U13103 (N_13103,N_8944,N_5212);
xnor U13104 (N_13104,N_8603,N_5451);
and U13105 (N_13105,N_8280,N_9471);
and U13106 (N_13106,N_8366,N_6105);
nand U13107 (N_13107,N_9099,N_5591);
xnor U13108 (N_13108,N_6978,N_6718);
xor U13109 (N_13109,N_6196,N_6028);
or U13110 (N_13110,N_8026,N_8212);
nand U13111 (N_13111,N_7739,N_8108);
nand U13112 (N_13112,N_8543,N_8425);
nand U13113 (N_13113,N_8310,N_6951);
nor U13114 (N_13114,N_7843,N_5309);
or U13115 (N_13115,N_6052,N_6881);
xor U13116 (N_13116,N_9885,N_7452);
nand U13117 (N_13117,N_8785,N_5429);
xnor U13118 (N_13118,N_7712,N_5501);
nor U13119 (N_13119,N_5967,N_6626);
nor U13120 (N_13120,N_7364,N_9581);
nand U13121 (N_13121,N_9685,N_7879);
or U13122 (N_13122,N_7673,N_8995);
and U13123 (N_13123,N_7106,N_6739);
nor U13124 (N_13124,N_8896,N_9987);
nor U13125 (N_13125,N_9863,N_5323);
or U13126 (N_13126,N_6572,N_6482);
xnor U13127 (N_13127,N_8564,N_9206);
xor U13128 (N_13128,N_9460,N_5137);
nand U13129 (N_13129,N_5679,N_6160);
xor U13130 (N_13130,N_6818,N_6453);
nand U13131 (N_13131,N_5024,N_9002);
and U13132 (N_13132,N_5829,N_7872);
xnor U13133 (N_13133,N_8774,N_9558);
nor U13134 (N_13134,N_9930,N_6266);
nor U13135 (N_13135,N_5151,N_9464);
and U13136 (N_13136,N_9712,N_9168);
or U13137 (N_13137,N_6796,N_8532);
or U13138 (N_13138,N_5493,N_7893);
and U13139 (N_13139,N_7778,N_9030);
and U13140 (N_13140,N_7893,N_9579);
and U13141 (N_13141,N_6656,N_5886);
nand U13142 (N_13142,N_9428,N_9206);
or U13143 (N_13143,N_9354,N_9432);
or U13144 (N_13144,N_9631,N_6553);
xnor U13145 (N_13145,N_9031,N_9671);
and U13146 (N_13146,N_7175,N_8083);
or U13147 (N_13147,N_6181,N_5226);
nor U13148 (N_13148,N_9354,N_6543);
nor U13149 (N_13149,N_9806,N_6698);
and U13150 (N_13150,N_7113,N_8475);
nor U13151 (N_13151,N_8154,N_9924);
xor U13152 (N_13152,N_5580,N_9547);
and U13153 (N_13153,N_8860,N_6101);
or U13154 (N_13154,N_5642,N_8322);
nand U13155 (N_13155,N_8406,N_6751);
or U13156 (N_13156,N_7306,N_6042);
nor U13157 (N_13157,N_7677,N_6380);
or U13158 (N_13158,N_6886,N_9413);
xor U13159 (N_13159,N_6038,N_9437);
nand U13160 (N_13160,N_5908,N_6268);
nor U13161 (N_13161,N_7293,N_7465);
xnor U13162 (N_13162,N_5922,N_5152);
xor U13163 (N_13163,N_7847,N_8445);
or U13164 (N_13164,N_9020,N_6034);
xnor U13165 (N_13165,N_7419,N_7862);
nor U13166 (N_13166,N_9416,N_9059);
nor U13167 (N_13167,N_7030,N_8904);
nand U13168 (N_13168,N_7537,N_5822);
xor U13169 (N_13169,N_8722,N_5671);
or U13170 (N_13170,N_8809,N_8007);
and U13171 (N_13171,N_7514,N_9538);
xnor U13172 (N_13172,N_8669,N_5596);
or U13173 (N_13173,N_6645,N_6630);
nor U13174 (N_13174,N_5610,N_5513);
nand U13175 (N_13175,N_6410,N_7325);
xor U13176 (N_13176,N_5913,N_8956);
nand U13177 (N_13177,N_5826,N_9034);
xor U13178 (N_13178,N_7044,N_9796);
nor U13179 (N_13179,N_8394,N_6541);
xnor U13180 (N_13180,N_8617,N_8494);
or U13181 (N_13181,N_7331,N_7285);
or U13182 (N_13182,N_9329,N_6723);
and U13183 (N_13183,N_6348,N_6924);
or U13184 (N_13184,N_5908,N_6489);
nand U13185 (N_13185,N_5519,N_7478);
nor U13186 (N_13186,N_9974,N_7130);
nor U13187 (N_13187,N_5318,N_9980);
xnor U13188 (N_13188,N_7704,N_8963);
or U13189 (N_13189,N_8000,N_8543);
or U13190 (N_13190,N_6761,N_6718);
and U13191 (N_13191,N_6859,N_8288);
nand U13192 (N_13192,N_9202,N_9728);
or U13193 (N_13193,N_8005,N_6719);
xor U13194 (N_13194,N_7775,N_7311);
nand U13195 (N_13195,N_8806,N_9723);
xor U13196 (N_13196,N_8784,N_7645);
xor U13197 (N_13197,N_9307,N_9667);
nor U13198 (N_13198,N_5541,N_6284);
xor U13199 (N_13199,N_9954,N_9993);
nor U13200 (N_13200,N_6579,N_7986);
xnor U13201 (N_13201,N_5816,N_9221);
xnor U13202 (N_13202,N_9664,N_6821);
nor U13203 (N_13203,N_6309,N_5259);
and U13204 (N_13204,N_5457,N_8965);
or U13205 (N_13205,N_6301,N_9469);
xor U13206 (N_13206,N_9248,N_7862);
nor U13207 (N_13207,N_6145,N_9694);
nor U13208 (N_13208,N_7441,N_6522);
and U13209 (N_13209,N_6206,N_8149);
xor U13210 (N_13210,N_8349,N_7704);
or U13211 (N_13211,N_8093,N_8631);
or U13212 (N_13212,N_9000,N_8760);
xnor U13213 (N_13213,N_6968,N_5924);
nand U13214 (N_13214,N_6341,N_5326);
or U13215 (N_13215,N_6782,N_8107);
nor U13216 (N_13216,N_9405,N_7883);
or U13217 (N_13217,N_5322,N_7752);
nand U13218 (N_13218,N_8142,N_9277);
and U13219 (N_13219,N_5954,N_6354);
or U13220 (N_13220,N_5100,N_5153);
xnor U13221 (N_13221,N_5752,N_5482);
and U13222 (N_13222,N_5400,N_8058);
nand U13223 (N_13223,N_5936,N_5491);
or U13224 (N_13224,N_9391,N_5509);
nand U13225 (N_13225,N_8086,N_9276);
nor U13226 (N_13226,N_9974,N_5814);
or U13227 (N_13227,N_9277,N_8771);
and U13228 (N_13228,N_6873,N_8348);
and U13229 (N_13229,N_6335,N_5197);
nand U13230 (N_13230,N_6243,N_9035);
xnor U13231 (N_13231,N_5390,N_7764);
or U13232 (N_13232,N_7313,N_7515);
nand U13233 (N_13233,N_5648,N_5412);
nor U13234 (N_13234,N_5949,N_5857);
and U13235 (N_13235,N_6367,N_7934);
xor U13236 (N_13236,N_9419,N_6497);
nor U13237 (N_13237,N_9295,N_6026);
or U13238 (N_13238,N_8616,N_8853);
nor U13239 (N_13239,N_8813,N_7388);
nand U13240 (N_13240,N_6315,N_9181);
or U13241 (N_13241,N_7736,N_6047);
xnor U13242 (N_13242,N_6075,N_9375);
or U13243 (N_13243,N_8138,N_8318);
and U13244 (N_13244,N_8835,N_9574);
or U13245 (N_13245,N_5519,N_5058);
xor U13246 (N_13246,N_7123,N_7347);
nor U13247 (N_13247,N_7974,N_7251);
nand U13248 (N_13248,N_5607,N_7865);
nor U13249 (N_13249,N_6736,N_8867);
xnor U13250 (N_13250,N_9738,N_5756);
xor U13251 (N_13251,N_6255,N_5876);
nand U13252 (N_13252,N_5582,N_9570);
nand U13253 (N_13253,N_8530,N_7251);
nand U13254 (N_13254,N_5455,N_8876);
nand U13255 (N_13255,N_7684,N_9306);
xnor U13256 (N_13256,N_8992,N_8007);
nand U13257 (N_13257,N_8431,N_5029);
xor U13258 (N_13258,N_7818,N_9756);
nand U13259 (N_13259,N_9954,N_6454);
nand U13260 (N_13260,N_9467,N_9605);
and U13261 (N_13261,N_7198,N_9137);
nand U13262 (N_13262,N_7551,N_5434);
xnor U13263 (N_13263,N_8112,N_6998);
nand U13264 (N_13264,N_8781,N_8169);
xnor U13265 (N_13265,N_9187,N_5266);
xor U13266 (N_13266,N_5925,N_5001);
nor U13267 (N_13267,N_6348,N_9201);
nand U13268 (N_13268,N_6566,N_7574);
or U13269 (N_13269,N_9741,N_5585);
xor U13270 (N_13270,N_6068,N_8037);
nor U13271 (N_13271,N_9342,N_7402);
nand U13272 (N_13272,N_9331,N_5012);
nor U13273 (N_13273,N_7568,N_9525);
xnor U13274 (N_13274,N_5943,N_5228);
nor U13275 (N_13275,N_8919,N_6331);
xnor U13276 (N_13276,N_5659,N_6878);
xnor U13277 (N_13277,N_9378,N_7997);
nand U13278 (N_13278,N_5799,N_7976);
and U13279 (N_13279,N_7077,N_9692);
nand U13280 (N_13280,N_5306,N_9431);
and U13281 (N_13281,N_8086,N_9917);
nor U13282 (N_13282,N_6982,N_6432);
nor U13283 (N_13283,N_5714,N_9890);
or U13284 (N_13284,N_7928,N_8124);
and U13285 (N_13285,N_9943,N_8862);
or U13286 (N_13286,N_6060,N_5989);
or U13287 (N_13287,N_9407,N_7211);
nor U13288 (N_13288,N_7800,N_9025);
nand U13289 (N_13289,N_9028,N_9264);
nand U13290 (N_13290,N_5218,N_9152);
or U13291 (N_13291,N_5301,N_8932);
nor U13292 (N_13292,N_6100,N_8023);
and U13293 (N_13293,N_6091,N_5124);
xnor U13294 (N_13294,N_7309,N_5138);
xnor U13295 (N_13295,N_8502,N_6788);
nand U13296 (N_13296,N_8513,N_7524);
nand U13297 (N_13297,N_8510,N_6905);
nor U13298 (N_13298,N_5701,N_6505);
xnor U13299 (N_13299,N_7319,N_6084);
nand U13300 (N_13300,N_8979,N_7899);
xnor U13301 (N_13301,N_8452,N_5718);
xor U13302 (N_13302,N_5146,N_8177);
nand U13303 (N_13303,N_9717,N_9485);
xnor U13304 (N_13304,N_6905,N_5011);
and U13305 (N_13305,N_8638,N_8699);
or U13306 (N_13306,N_7780,N_8004);
and U13307 (N_13307,N_7402,N_9912);
nor U13308 (N_13308,N_6274,N_5369);
and U13309 (N_13309,N_9483,N_8967);
nor U13310 (N_13310,N_5871,N_9038);
and U13311 (N_13311,N_9822,N_8271);
or U13312 (N_13312,N_7235,N_5342);
or U13313 (N_13313,N_6047,N_8544);
nand U13314 (N_13314,N_9984,N_5603);
or U13315 (N_13315,N_7918,N_9670);
and U13316 (N_13316,N_9971,N_6950);
nor U13317 (N_13317,N_5928,N_6587);
nand U13318 (N_13318,N_8439,N_6993);
and U13319 (N_13319,N_7854,N_9835);
nor U13320 (N_13320,N_5101,N_6672);
or U13321 (N_13321,N_9699,N_8361);
nor U13322 (N_13322,N_7402,N_5690);
nand U13323 (N_13323,N_9813,N_6335);
or U13324 (N_13324,N_9177,N_5804);
and U13325 (N_13325,N_7463,N_6913);
and U13326 (N_13326,N_5085,N_8456);
xnor U13327 (N_13327,N_7832,N_8443);
or U13328 (N_13328,N_6332,N_9217);
nand U13329 (N_13329,N_6607,N_9124);
or U13330 (N_13330,N_8713,N_8610);
xor U13331 (N_13331,N_5805,N_7794);
nor U13332 (N_13332,N_5526,N_7109);
and U13333 (N_13333,N_8139,N_9976);
xor U13334 (N_13334,N_5076,N_5410);
and U13335 (N_13335,N_6222,N_6672);
xor U13336 (N_13336,N_5189,N_5276);
nand U13337 (N_13337,N_5341,N_8340);
and U13338 (N_13338,N_7444,N_7874);
nor U13339 (N_13339,N_7051,N_9815);
nor U13340 (N_13340,N_7817,N_5304);
and U13341 (N_13341,N_9840,N_8496);
or U13342 (N_13342,N_7303,N_9349);
xnor U13343 (N_13343,N_5946,N_9988);
and U13344 (N_13344,N_5399,N_6726);
nand U13345 (N_13345,N_7845,N_6158);
nor U13346 (N_13346,N_6086,N_9457);
and U13347 (N_13347,N_9649,N_5121);
nand U13348 (N_13348,N_7486,N_6342);
xor U13349 (N_13349,N_8084,N_5332);
and U13350 (N_13350,N_5941,N_5472);
nor U13351 (N_13351,N_8892,N_6586);
xor U13352 (N_13352,N_8189,N_7627);
xor U13353 (N_13353,N_7332,N_7655);
xor U13354 (N_13354,N_5340,N_5557);
xnor U13355 (N_13355,N_6001,N_6490);
or U13356 (N_13356,N_9500,N_9602);
or U13357 (N_13357,N_8584,N_7497);
or U13358 (N_13358,N_8875,N_6140);
or U13359 (N_13359,N_8833,N_6823);
nand U13360 (N_13360,N_7742,N_7402);
nand U13361 (N_13361,N_7103,N_7860);
nand U13362 (N_13362,N_9021,N_8059);
or U13363 (N_13363,N_7660,N_8199);
and U13364 (N_13364,N_7895,N_5823);
nand U13365 (N_13365,N_8626,N_8717);
or U13366 (N_13366,N_6082,N_8868);
nor U13367 (N_13367,N_7573,N_5853);
nor U13368 (N_13368,N_8840,N_8878);
or U13369 (N_13369,N_5693,N_8895);
and U13370 (N_13370,N_7853,N_7188);
nor U13371 (N_13371,N_9694,N_6180);
or U13372 (N_13372,N_9776,N_7008);
and U13373 (N_13373,N_6535,N_8587);
xor U13374 (N_13374,N_6218,N_5663);
xnor U13375 (N_13375,N_6579,N_9787);
and U13376 (N_13376,N_9582,N_8788);
or U13377 (N_13377,N_8353,N_6827);
nor U13378 (N_13378,N_9360,N_9653);
xor U13379 (N_13379,N_9028,N_9143);
xnor U13380 (N_13380,N_9506,N_9297);
or U13381 (N_13381,N_7832,N_8892);
nor U13382 (N_13382,N_9243,N_9080);
and U13383 (N_13383,N_6465,N_5521);
xnor U13384 (N_13384,N_9615,N_7949);
nand U13385 (N_13385,N_5637,N_5961);
and U13386 (N_13386,N_9628,N_7107);
nor U13387 (N_13387,N_9607,N_5722);
nand U13388 (N_13388,N_5934,N_5666);
xnor U13389 (N_13389,N_9404,N_6884);
nand U13390 (N_13390,N_5428,N_9825);
nand U13391 (N_13391,N_9117,N_5010);
nand U13392 (N_13392,N_7260,N_6469);
nand U13393 (N_13393,N_7952,N_7845);
nor U13394 (N_13394,N_6849,N_9431);
nand U13395 (N_13395,N_7437,N_6362);
nor U13396 (N_13396,N_8404,N_8840);
nand U13397 (N_13397,N_6901,N_9838);
nand U13398 (N_13398,N_7283,N_6454);
or U13399 (N_13399,N_7473,N_6449);
and U13400 (N_13400,N_5419,N_6823);
or U13401 (N_13401,N_9684,N_8614);
nand U13402 (N_13402,N_8331,N_9656);
and U13403 (N_13403,N_9721,N_8880);
and U13404 (N_13404,N_5545,N_5355);
nand U13405 (N_13405,N_8479,N_6381);
nand U13406 (N_13406,N_7270,N_8295);
or U13407 (N_13407,N_7144,N_9820);
nor U13408 (N_13408,N_6736,N_9450);
and U13409 (N_13409,N_7094,N_5851);
or U13410 (N_13410,N_9510,N_6807);
nand U13411 (N_13411,N_5073,N_9932);
or U13412 (N_13412,N_5291,N_8981);
nand U13413 (N_13413,N_8653,N_7538);
or U13414 (N_13414,N_7680,N_8913);
nor U13415 (N_13415,N_5313,N_8288);
xnor U13416 (N_13416,N_6200,N_9191);
nor U13417 (N_13417,N_9413,N_7145);
nand U13418 (N_13418,N_5492,N_9060);
and U13419 (N_13419,N_7194,N_8619);
xor U13420 (N_13420,N_9886,N_5015);
or U13421 (N_13421,N_9162,N_6009);
nand U13422 (N_13422,N_5107,N_8361);
nand U13423 (N_13423,N_8915,N_9416);
nor U13424 (N_13424,N_8974,N_8905);
and U13425 (N_13425,N_9436,N_6391);
xor U13426 (N_13426,N_9462,N_5359);
xnor U13427 (N_13427,N_7325,N_9878);
nor U13428 (N_13428,N_8382,N_8273);
xnor U13429 (N_13429,N_6532,N_8815);
and U13430 (N_13430,N_7356,N_5216);
nand U13431 (N_13431,N_8560,N_9431);
and U13432 (N_13432,N_9774,N_8832);
nor U13433 (N_13433,N_6757,N_8888);
and U13434 (N_13434,N_7829,N_8018);
or U13435 (N_13435,N_9807,N_9282);
or U13436 (N_13436,N_7817,N_5861);
nor U13437 (N_13437,N_6101,N_6994);
nor U13438 (N_13438,N_5966,N_8451);
nand U13439 (N_13439,N_5847,N_9790);
xor U13440 (N_13440,N_7248,N_9983);
nor U13441 (N_13441,N_6778,N_9137);
xor U13442 (N_13442,N_9558,N_8864);
nand U13443 (N_13443,N_7000,N_7578);
nand U13444 (N_13444,N_9075,N_5858);
nand U13445 (N_13445,N_7040,N_6040);
and U13446 (N_13446,N_9638,N_7652);
or U13447 (N_13447,N_7105,N_5816);
or U13448 (N_13448,N_8295,N_5662);
nor U13449 (N_13449,N_5767,N_7812);
nor U13450 (N_13450,N_8645,N_8583);
nor U13451 (N_13451,N_6425,N_6103);
nand U13452 (N_13452,N_7826,N_5498);
and U13453 (N_13453,N_8478,N_6261);
and U13454 (N_13454,N_8995,N_6856);
xnor U13455 (N_13455,N_6391,N_6511);
and U13456 (N_13456,N_5673,N_7073);
or U13457 (N_13457,N_5013,N_9185);
nor U13458 (N_13458,N_8536,N_8446);
or U13459 (N_13459,N_8146,N_6976);
nor U13460 (N_13460,N_5045,N_5251);
or U13461 (N_13461,N_6816,N_5477);
nor U13462 (N_13462,N_6798,N_7142);
nor U13463 (N_13463,N_7376,N_9115);
or U13464 (N_13464,N_5204,N_6294);
xnor U13465 (N_13465,N_7072,N_5063);
or U13466 (N_13466,N_6772,N_8718);
nand U13467 (N_13467,N_8546,N_8475);
nor U13468 (N_13468,N_8684,N_8213);
xnor U13469 (N_13469,N_7977,N_9556);
nor U13470 (N_13470,N_6466,N_5002);
nand U13471 (N_13471,N_8603,N_6549);
nand U13472 (N_13472,N_7031,N_9127);
nor U13473 (N_13473,N_8239,N_7280);
and U13474 (N_13474,N_6650,N_6500);
xor U13475 (N_13475,N_6798,N_6945);
xor U13476 (N_13476,N_8742,N_5675);
or U13477 (N_13477,N_6109,N_7001);
nand U13478 (N_13478,N_8668,N_9688);
and U13479 (N_13479,N_5585,N_8014);
and U13480 (N_13480,N_8247,N_6510);
or U13481 (N_13481,N_5777,N_9869);
or U13482 (N_13482,N_6608,N_5553);
or U13483 (N_13483,N_6565,N_7635);
and U13484 (N_13484,N_8826,N_6426);
or U13485 (N_13485,N_9223,N_8268);
nand U13486 (N_13486,N_8829,N_5245);
nand U13487 (N_13487,N_8980,N_8161);
and U13488 (N_13488,N_7834,N_9680);
or U13489 (N_13489,N_7724,N_9308);
nand U13490 (N_13490,N_8462,N_9272);
nand U13491 (N_13491,N_8415,N_9805);
or U13492 (N_13492,N_6089,N_8498);
nand U13493 (N_13493,N_8905,N_8512);
xnor U13494 (N_13494,N_6524,N_9202);
or U13495 (N_13495,N_8938,N_5723);
or U13496 (N_13496,N_5205,N_7914);
and U13497 (N_13497,N_6966,N_9930);
nor U13498 (N_13498,N_5727,N_5587);
and U13499 (N_13499,N_8794,N_7054);
nor U13500 (N_13500,N_8597,N_8997);
or U13501 (N_13501,N_8704,N_8944);
nor U13502 (N_13502,N_9647,N_6119);
nand U13503 (N_13503,N_9146,N_9167);
or U13504 (N_13504,N_7536,N_5524);
nor U13505 (N_13505,N_7076,N_6479);
nor U13506 (N_13506,N_9939,N_7758);
nand U13507 (N_13507,N_8043,N_7658);
or U13508 (N_13508,N_5526,N_9932);
nand U13509 (N_13509,N_9113,N_8545);
nor U13510 (N_13510,N_9951,N_6407);
or U13511 (N_13511,N_9047,N_7784);
xor U13512 (N_13512,N_5528,N_5643);
nor U13513 (N_13513,N_6242,N_6065);
or U13514 (N_13514,N_8508,N_9877);
nand U13515 (N_13515,N_9028,N_8459);
nor U13516 (N_13516,N_9788,N_5410);
and U13517 (N_13517,N_9182,N_7676);
and U13518 (N_13518,N_9956,N_5753);
nor U13519 (N_13519,N_5863,N_6519);
xor U13520 (N_13520,N_6791,N_8484);
or U13521 (N_13521,N_8266,N_9884);
or U13522 (N_13522,N_5106,N_6606);
nor U13523 (N_13523,N_9909,N_7377);
or U13524 (N_13524,N_9774,N_7722);
nor U13525 (N_13525,N_6616,N_6962);
nand U13526 (N_13526,N_7150,N_6016);
and U13527 (N_13527,N_9462,N_5660);
or U13528 (N_13528,N_5255,N_5909);
or U13529 (N_13529,N_5628,N_8611);
xor U13530 (N_13530,N_6385,N_8353);
nand U13531 (N_13531,N_8715,N_5514);
or U13532 (N_13532,N_5281,N_5020);
xor U13533 (N_13533,N_9127,N_6314);
xor U13534 (N_13534,N_9667,N_9201);
xor U13535 (N_13535,N_6155,N_6210);
nor U13536 (N_13536,N_6092,N_6030);
nor U13537 (N_13537,N_7994,N_5092);
and U13538 (N_13538,N_9532,N_7994);
or U13539 (N_13539,N_5705,N_7689);
nor U13540 (N_13540,N_6319,N_6619);
and U13541 (N_13541,N_7776,N_5433);
or U13542 (N_13542,N_5559,N_7993);
xnor U13543 (N_13543,N_7718,N_5472);
xor U13544 (N_13544,N_6217,N_5781);
or U13545 (N_13545,N_8612,N_5388);
nor U13546 (N_13546,N_5850,N_6585);
nand U13547 (N_13547,N_9341,N_7820);
nand U13548 (N_13548,N_5374,N_8276);
or U13549 (N_13549,N_9228,N_6111);
or U13550 (N_13550,N_9635,N_7742);
nor U13551 (N_13551,N_6057,N_9523);
and U13552 (N_13552,N_5685,N_6450);
and U13553 (N_13553,N_9173,N_9786);
or U13554 (N_13554,N_6321,N_7222);
and U13555 (N_13555,N_5943,N_9023);
nand U13556 (N_13556,N_9087,N_9810);
xor U13557 (N_13557,N_8245,N_8795);
or U13558 (N_13558,N_7225,N_9510);
nor U13559 (N_13559,N_7781,N_5730);
xor U13560 (N_13560,N_6642,N_8935);
nand U13561 (N_13561,N_7520,N_9639);
nand U13562 (N_13562,N_6140,N_7753);
and U13563 (N_13563,N_5465,N_9727);
nand U13564 (N_13564,N_9677,N_6842);
nand U13565 (N_13565,N_5740,N_9670);
nand U13566 (N_13566,N_5438,N_5852);
or U13567 (N_13567,N_7466,N_8880);
nor U13568 (N_13568,N_7136,N_6110);
nand U13569 (N_13569,N_6806,N_7698);
nor U13570 (N_13570,N_9409,N_5498);
nand U13571 (N_13571,N_8486,N_9217);
nor U13572 (N_13572,N_8707,N_5676);
and U13573 (N_13573,N_9055,N_9083);
nor U13574 (N_13574,N_9204,N_6293);
xor U13575 (N_13575,N_9094,N_9751);
or U13576 (N_13576,N_7371,N_8978);
nand U13577 (N_13577,N_9002,N_9159);
or U13578 (N_13578,N_8395,N_7782);
nor U13579 (N_13579,N_6683,N_9195);
nand U13580 (N_13580,N_5343,N_8562);
nand U13581 (N_13581,N_9959,N_9056);
or U13582 (N_13582,N_5829,N_7861);
nand U13583 (N_13583,N_7537,N_5514);
or U13584 (N_13584,N_7710,N_6183);
xnor U13585 (N_13585,N_6707,N_9335);
xnor U13586 (N_13586,N_9287,N_6470);
nand U13587 (N_13587,N_5105,N_8405);
or U13588 (N_13588,N_5443,N_5796);
and U13589 (N_13589,N_9362,N_9920);
nand U13590 (N_13590,N_9491,N_9199);
xnor U13591 (N_13591,N_5623,N_8013);
and U13592 (N_13592,N_9033,N_7680);
nand U13593 (N_13593,N_5847,N_7989);
or U13594 (N_13594,N_9687,N_9192);
or U13595 (N_13595,N_9894,N_5455);
nand U13596 (N_13596,N_5984,N_7668);
nor U13597 (N_13597,N_8705,N_9772);
xor U13598 (N_13598,N_7440,N_5030);
xor U13599 (N_13599,N_7226,N_6797);
or U13600 (N_13600,N_9201,N_5956);
or U13601 (N_13601,N_8438,N_8551);
xor U13602 (N_13602,N_6553,N_9953);
or U13603 (N_13603,N_7832,N_7171);
nand U13604 (N_13604,N_5891,N_8231);
and U13605 (N_13605,N_7529,N_8919);
nor U13606 (N_13606,N_9304,N_7912);
and U13607 (N_13607,N_7901,N_8277);
or U13608 (N_13608,N_7959,N_7708);
nor U13609 (N_13609,N_6512,N_6584);
xnor U13610 (N_13610,N_8086,N_6683);
nor U13611 (N_13611,N_7468,N_8708);
or U13612 (N_13612,N_8171,N_7165);
nand U13613 (N_13613,N_7620,N_9703);
nor U13614 (N_13614,N_5866,N_7503);
xor U13615 (N_13615,N_9452,N_6499);
and U13616 (N_13616,N_9062,N_7388);
nor U13617 (N_13617,N_7313,N_7777);
and U13618 (N_13618,N_8869,N_8781);
nor U13619 (N_13619,N_6827,N_6472);
nor U13620 (N_13620,N_8073,N_6329);
and U13621 (N_13621,N_8121,N_8909);
and U13622 (N_13622,N_5940,N_5027);
nor U13623 (N_13623,N_8461,N_9897);
nand U13624 (N_13624,N_6796,N_6248);
nor U13625 (N_13625,N_6436,N_6320);
nor U13626 (N_13626,N_7459,N_5287);
nor U13627 (N_13627,N_7095,N_9546);
or U13628 (N_13628,N_7863,N_9242);
and U13629 (N_13629,N_8574,N_8114);
nor U13630 (N_13630,N_8875,N_7576);
and U13631 (N_13631,N_9050,N_6274);
nor U13632 (N_13632,N_7536,N_7476);
and U13633 (N_13633,N_7256,N_5717);
or U13634 (N_13634,N_9980,N_6209);
nor U13635 (N_13635,N_6624,N_8978);
xor U13636 (N_13636,N_6002,N_9065);
nor U13637 (N_13637,N_7758,N_8010);
and U13638 (N_13638,N_7896,N_6562);
nand U13639 (N_13639,N_8671,N_5475);
nor U13640 (N_13640,N_8681,N_7735);
or U13641 (N_13641,N_6195,N_6863);
or U13642 (N_13642,N_9678,N_6327);
and U13643 (N_13643,N_7028,N_8153);
xnor U13644 (N_13644,N_5042,N_7569);
or U13645 (N_13645,N_9789,N_9314);
and U13646 (N_13646,N_8826,N_8078);
xor U13647 (N_13647,N_6264,N_5141);
xor U13648 (N_13648,N_5371,N_6691);
or U13649 (N_13649,N_6145,N_6400);
and U13650 (N_13650,N_9400,N_6695);
and U13651 (N_13651,N_7731,N_5802);
nor U13652 (N_13652,N_6636,N_9636);
and U13653 (N_13653,N_9370,N_7660);
or U13654 (N_13654,N_6030,N_9422);
or U13655 (N_13655,N_8676,N_8990);
xnor U13656 (N_13656,N_9047,N_9934);
and U13657 (N_13657,N_8618,N_7946);
or U13658 (N_13658,N_6845,N_8349);
or U13659 (N_13659,N_9312,N_6775);
and U13660 (N_13660,N_5139,N_5717);
and U13661 (N_13661,N_8186,N_6762);
nor U13662 (N_13662,N_6188,N_5951);
and U13663 (N_13663,N_8027,N_6708);
and U13664 (N_13664,N_7048,N_6310);
xor U13665 (N_13665,N_8672,N_9164);
xnor U13666 (N_13666,N_9880,N_8607);
nor U13667 (N_13667,N_5767,N_8059);
nor U13668 (N_13668,N_6421,N_5153);
or U13669 (N_13669,N_9512,N_5483);
xnor U13670 (N_13670,N_5438,N_6941);
nor U13671 (N_13671,N_9503,N_9772);
or U13672 (N_13672,N_7459,N_7207);
xnor U13673 (N_13673,N_7234,N_6743);
nor U13674 (N_13674,N_7166,N_5073);
nand U13675 (N_13675,N_7878,N_6738);
xor U13676 (N_13676,N_8723,N_9952);
or U13677 (N_13677,N_8346,N_9074);
or U13678 (N_13678,N_8575,N_5631);
and U13679 (N_13679,N_8247,N_8554);
nor U13680 (N_13680,N_5050,N_5240);
nor U13681 (N_13681,N_7317,N_6744);
xnor U13682 (N_13682,N_6174,N_7881);
and U13683 (N_13683,N_8988,N_7481);
and U13684 (N_13684,N_5590,N_6997);
or U13685 (N_13685,N_8093,N_9585);
xor U13686 (N_13686,N_6361,N_6967);
nand U13687 (N_13687,N_8346,N_9503);
xor U13688 (N_13688,N_6162,N_9849);
nor U13689 (N_13689,N_5693,N_7335);
xnor U13690 (N_13690,N_5025,N_5394);
xnor U13691 (N_13691,N_6322,N_8439);
or U13692 (N_13692,N_8341,N_5268);
nor U13693 (N_13693,N_6755,N_8463);
nand U13694 (N_13694,N_8985,N_7056);
or U13695 (N_13695,N_7679,N_9808);
nand U13696 (N_13696,N_8962,N_5626);
or U13697 (N_13697,N_9181,N_9117);
or U13698 (N_13698,N_6103,N_6636);
nor U13699 (N_13699,N_8849,N_9795);
nand U13700 (N_13700,N_5952,N_8287);
or U13701 (N_13701,N_9293,N_6027);
xnor U13702 (N_13702,N_6292,N_9459);
xnor U13703 (N_13703,N_8151,N_8673);
nand U13704 (N_13704,N_9782,N_6069);
nand U13705 (N_13705,N_7225,N_5509);
xnor U13706 (N_13706,N_5869,N_7451);
nor U13707 (N_13707,N_6748,N_7016);
nor U13708 (N_13708,N_5841,N_5006);
nor U13709 (N_13709,N_8747,N_7473);
nand U13710 (N_13710,N_7669,N_8008);
or U13711 (N_13711,N_8374,N_8390);
xnor U13712 (N_13712,N_5550,N_5321);
and U13713 (N_13713,N_9267,N_5717);
xnor U13714 (N_13714,N_7765,N_9264);
or U13715 (N_13715,N_7826,N_6906);
nand U13716 (N_13716,N_5931,N_7417);
nand U13717 (N_13717,N_9849,N_9083);
xor U13718 (N_13718,N_5059,N_5586);
nand U13719 (N_13719,N_7952,N_7915);
nand U13720 (N_13720,N_8844,N_8920);
xor U13721 (N_13721,N_8840,N_6797);
nor U13722 (N_13722,N_7480,N_5367);
and U13723 (N_13723,N_7279,N_8228);
nand U13724 (N_13724,N_7673,N_9529);
or U13725 (N_13725,N_7038,N_7316);
xnor U13726 (N_13726,N_8549,N_9865);
and U13727 (N_13727,N_6274,N_6439);
or U13728 (N_13728,N_6163,N_6530);
or U13729 (N_13729,N_6262,N_5492);
and U13730 (N_13730,N_6721,N_5631);
and U13731 (N_13731,N_6479,N_8578);
nand U13732 (N_13732,N_7228,N_7557);
nor U13733 (N_13733,N_6294,N_6057);
nand U13734 (N_13734,N_9100,N_8413);
or U13735 (N_13735,N_9500,N_7927);
or U13736 (N_13736,N_8752,N_6340);
nand U13737 (N_13737,N_6767,N_7110);
or U13738 (N_13738,N_8167,N_5256);
nor U13739 (N_13739,N_9481,N_7987);
nor U13740 (N_13740,N_9745,N_9789);
or U13741 (N_13741,N_9912,N_8184);
and U13742 (N_13742,N_7770,N_9314);
xor U13743 (N_13743,N_6758,N_9058);
or U13744 (N_13744,N_6392,N_6616);
xnor U13745 (N_13745,N_5956,N_7201);
xnor U13746 (N_13746,N_7419,N_8374);
nand U13747 (N_13747,N_7597,N_5923);
nor U13748 (N_13748,N_5643,N_8633);
nand U13749 (N_13749,N_7562,N_8448);
and U13750 (N_13750,N_7078,N_5099);
or U13751 (N_13751,N_9594,N_6489);
and U13752 (N_13752,N_9454,N_7300);
nand U13753 (N_13753,N_7632,N_8296);
nor U13754 (N_13754,N_9833,N_7137);
or U13755 (N_13755,N_9130,N_8052);
xor U13756 (N_13756,N_8267,N_7280);
xor U13757 (N_13757,N_7701,N_8562);
and U13758 (N_13758,N_6315,N_8429);
nand U13759 (N_13759,N_9461,N_7194);
nand U13760 (N_13760,N_9288,N_8291);
nand U13761 (N_13761,N_9788,N_8004);
nor U13762 (N_13762,N_8864,N_5513);
nor U13763 (N_13763,N_7750,N_5750);
or U13764 (N_13764,N_9867,N_6945);
nand U13765 (N_13765,N_9291,N_6899);
xnor U13766 (N_13766,N_7772,N_7403);
nand U13767 (N_13767,N_5899,N_8338);
and U13768 (N_13768,N_9265,N_7465);
nand U13769 (N_13769,N_9343,N_8841);
nor U13770 (N_13770,N_9136,N_5838);
or U13771 (N_13771,N_5521,N_8863);
xor U13772 (N_13772,N_6047,N_9603);
nand U13773 (N_13773,N_6322,N_5711);
nand U13774 (N_13774,N_7002,N_9132);
nand U13775 (N_13775,N_6740,N_9361);
or U13776 (N_13776,N_7267,N_9055);
or U13777 (N_13777,N_8136,N_8096);
and U13778 (N_13778,N_5580,N_7182);
nor U13779 (N_13779,N_6555,N_8637);
and U13780 (N_13780,N_8306,N_7231);
nand U13781 (N_13781,N_7300,N_5501);
nor U13782 (N_13782,N_9713,N_9784);
xnor U13783 (N_13783,N_5943,N_8993);
or U13784 (N_13784,N_6852,N_6778);
and U13785 (N_13785,N_6512,N_6051);
xnor U13786 (N_13786,N_6186,N_5824);
xnor U13787 (N_13787,N_6820,N_5845);
or U13788 (N_13788,N_9278,N_6297);
or U13789 (N_13789,N_9845,N_5405);
nand U13790 (N_13790,N_7146,N_8184);
nor U13791 (N_13791,N_8244,N_6212);
and U13792 (N_13792,N_5246,N_9880);
nor U13793 (N_13793,N_9269,N_8278);
and U13794 (N_13794,N_7098,N_9623);
and U13795 (N_13795,N_9835,N_5236);
nor U13796 (N_13796,N_8639,N_7170);
and U13797 (N_13797,N_6328,N_6047);
nand U13798 (N_13798,N_7670,N_7829);
xnor U13799 (N_13799,N_8595,N_9273);
xnor U13800 (N_13800,N_6319,N_9461);
nor U13801 (N_13801,N_7561,N_8646);
or U13802 (N_13802,N_8756,N_9559);
or U13803 (N_13803,N_6176,N_5993);
and U13804 (N_13804,N_7339,N_9516);
xnor U13805 (N_13805,N_8957,N_6515);
xor U13806 (N_13806,N_6189,N_6135);
nor U13807 (N_13807,N_6757,N_6191);
nor U13808 (N_13808,N_8834,N_6960);
and U13809 (N_13809,N_8899,N_8759);
nand U13810 (N_13810,N_8229,N_9293);
nand U13811 (N_13811,N_6913,N_8835);
or U13812 (N_13812,N_7799,N_7714);
or U13813 (N_13813,N_7408,N_7000);
and U13814 (N_13814,N_9194,N_8914);
and U13815 (N_13815,N_8148,N_6738);
xnor U13816 (N_13816,N_7097,N_5917);
nand U13817 (N_13817,N_9163,N_7148);
nand U13818 (N_13818,N_7171,N_7791);
xnor U13819 (N_13819,N_5574,N_7596);
and U13820 (N_13820,N_8590,N_7194);
and U13821 (N_13821,N_8405,N_5634);
xor U13822 (N_13822,N_8456,N_7752);
and U13823 (N_13823,N_5373,N_5153);
nand U13824 (N_13824,N_9638,N_5369);
nor U13825 (N_13825,N_7252,N_8283);
nand U13826 (N_13826,N_6545,N_9994);
xnor U13827 (N_13827,N_8493,N_5865);
and U13828 (N_13828,N_5904,N_9706);
nand U13829 (N_13829,N_9203,N_7656);
or U13830 (N_13830,N_9439,N_8940);
nor U13831 (N_13831,N_7327,N_9615);
or U13832 (N_13832,N_8017,N_8108);
nand U13833 (N_13833,N_9653,N_9730);
nand U13834 (N_13834,N_7844,N_5730);
and U13835 (N_13835,N_6777,N_9643);
nand U13836 (N_13836,N_6068,N_8781);
xor U13837 (N_13837,N_8457,N_6422);
nand U13838 (N_13838,N_5616,N_8944);
xnor U13839 (N_13839,N_6489,N_5099);
nor U13840 (N_13840,N_7856,N_6213);
nand U13841 (N_13841,N_7871,N_8930);
nand U13842 (N_13842,N_7191,N_8444);
nor U13843 (N_13843,N_7888,N_6414);
nand U13844 (N_13844,N_7283,N_8294);
nand U13845 (N_13845,N_7810,N_5836);
nand U13846 (N_13846,N_7353,N_7478);
xor U13847 (N_13847,N_9503,N_5251);
and U13848 (N_13848,N_7094,N_7348);
or U13849 (N_13849,N_7103,N_7276);
xor U13850 (N_13850,N_9799,N_7791);
nor U13851 (N_13851,N_8375,N_5695);
nand U13852 (N_13852,N_7537,N_6995);
nand U13853 (N_13853,N_5538,N_5124);
or U13854 (N_13854,N_9885,N_5380);
nor U13855 (N_13855,N_8006,N_6955);
nand U13856 (N_13856,N_7593,N_6161);
nand U13857 (N_13857,N_6459,N_5690);
xnor U13858 (N_13858,N_5679,N_9091);
and U13859 (N_13859,N_6106,N_8141);
nor U13860 (N_13860,N_8075,N_9448);
nor U13861 (N_13861,N_9337,N_7943);
and U13862 (N_13862,N_7895,N_6307);
nand U13863 (N_13863,N_5021,N_5689);
or U13864 (N_13864,N_5267,N_9267);
nand U13865 (N_13865,N_9394,N_8096);
nor U13866 (N_13866,N_5644,N_9681);
nor U13867 (N_13867,N_7180,N_5535);
nand U13868 (N_13868,N_5748,N_5149);
or U13869 (N_13869,N_5839,N_9885);
or U13870 (N_13870,N_6490,N_7930);
and U13871 (N_13871,N_9036,N_7977);
or U13872 (N_13872,N_8397,N_5637);
and U13873 (N_13873,N_9190,N_7094);
or U13874 (N_13874,N_6349,N_8338);
or U13875 (N_13875,N_7398,N_9289);
or U13876 (N_13876,N_8527,N_9539);
nor U13877 (N_13877,N_5013,N_7864);
and U13878 (N_13878,N_6262,N_8898);
or U13879 (N_13879,N_8049,N_6988);
nor U13880 (N_13880,N_6323,N_8358);
xor U13881 (N_13881,N_5775,N_8132);
and U13882 (N_13882,N_8589,N_8747);
or U13883 (N_13883,N_6558,N_6601);
nand U13884 (N_13884,N_7562,N_6940);
xor U13885 (N_13885,N_5394,N_8626);
xnor U13886 (N_13886,N_6084,N_8921);
xor U13887 (N_13887,N_8585,N_5404);
xor U13888 (N_13888,N_5002,N_5650);
nor U13889 (N_13889,N_9200,N_8646);
nor U13890 (N_13890,N_5049,N_9026);
xor U13891 (N_13891,N_5188,N_5585);
nand U13892 (N_13892,N_8754,N_8299);
xor U13893 (N_13893,N_6277,N_9866);
or U13894 (N_13894,N_8530,N_8196);
or U13895 (N_13895,N_6894,N_7066);
nand U13896 (N_13896,N_8370,N_9380);
nor U13897 (N_13897,N_5655,N_6852);
or U13898 (N_13898,N_7362,N_6936);
nor U13899 (N_13899,N_9574,N_8848);
or U13900 (N_13900,N_7338,N_9209);
nor U13901 (N_13901,N_8584,N_5260);
xnor U13902 (N_13902,N_5082,N_8150);
and U13903 (N_13903,N_9466,N_6197);
xnor U13904 (N_13904,N_8959,N_9082);
nor U13905 (N_13905,N_7841,N_8924);
xnor U13906 (N_13906,N_9009,N_5571);
xor U13907 (N_13907,N_7858,N_8715);
nor U13908 (N_13908,N_7075,N_9446);
or U13909 (N_13909,N_8446,N_7592);
nor U13910 (N_13910,N_6532,N_6213);
xor U13911 (N_13911,N_6885,N_7204);
and U13912 (N_13912,N_8032,N_5648);
or U13913 (N_13913,N_5543,N_6844);
nor U13914 (N_13914,N_7691,N_9834);
nand U13915 (N_13915,N_8401,N_7259);
and U13916 (N_13916,N_6960,N_8585);
xor U13917 (N_13917,N_8662,N_9359);
nor U13918 (N_13918,N_8420,N_6687);
xnor U13919 (N_13919,N_9796,N_6548);
nand U13920 (N_13920,N_9613,N_6112);
nor U13921 (N_13921,N_9225,N_7843);
xnor U13922 (N_13922,N_7552,N_9720);
xnor U13923 (N_13923,N_5130,N_5327);
xor U13924 (N_13924,N_5592,N_8728);
xnor U13925 (N_13925,N_7779,N_9835);
or U13926 (N_13926,N_5832,N_7446);
or U13927 (N_13927,N_8136,N_6616);
nand U13928 (N_13928,N_9673,N_5225);
nand U13929 (N_13929,N_7263,N_8830);
or U13930 (N_13930,N_8457,N_6442);
xor U13931 (N_13931,N_7306,N_8174);
xnor U13932 (N_13932,N_6206,N_7626);
xnor U13933 (N_13933,N_7916,N_8243);
nor U13934 (N_13934,N_9236,N_7269);
and U13935 (N_13935,N_7455,N_5758);
and U13936 (N_13936,N_5707,N_6421);
and U13937 (N_13937,N_7454,N_9356);
or U13938 (N_13938,N_7202,N_7283);
and U13939 (N_13939,N_7732,N_9042);
or U13940 (N_13940,N_6626,N_9780);
and U13941 (N_13941,N_8613,N_5107);
nand U13942 (N_13942,N_9873,N_5126);
xnor U13943 (N_13943,N_8701,N_9997);
xor U13944 (N_13944,N_7793,N_8227);
nor U13945 (N_13945,N_9608,N_5370);
and U13946 (N_13946,N_7952,N_8305);
and U13947 (N_13947,N_9023,N_9646);
nor U13948 (N_13948,N_8940,N_8934);
xor U13949 (N_13949,N_8805,N_6361);
nand U13950 (N_13950,N_6851,N_5574);
nor U13951 (N_13951,N_7152,N_8619);
nand U13952 (N_13952,N_8405,N_5313);
xnor U13953 (N_13953,N_7016,N_8305);
or U13954 (N_13954,N_6903,N_9447);
and U13955 (N_13955,N_9786,N_9534);
and U13956 (N_13956,N_6109,N_7836);
or U13957 (N_13957,N_6401,N_7952);
and U13958 (N_13958,N_8357,N_8907);
nor U13959 (N_13959,N_8434,N_7251);
or U13960 (N_13960,N_7951,N_9128);
xor U13961 (N_13961,N_5051,N_5143);
nand U13962 (N_13962,N_6645,N_6936);
and U13963 (N_13963,N_8077,N_9676);
or U13964 (N_13964,N_8794,N_8136);
nand U13965 (N_13965,N_7456,N_5188);
and U13966 (N_13966,N_6821,N_6390);
nor U13967 (N_13967,N_8602,N_6810);
or U13968 (N_13968,N_7731,N_8513);
or U13969 (N_13969,N_5466,N_7308);
or U13970 (N_13970,N_6889,N_5735);
xor U13971 (N_13971,N_5353,N_5466);
nor U13972 (N_13972,N_9262,N_7615);
nor U13973 (N_13973,N_6906,N_5584);
or U13974 (N_13974,N_7652,N_8727);
nand U13975 (N_13975,N_8064,N_6847);
or U13976 (N_13976,N_8930,N_9359);
nand U13977 (N_13977,N_7644,N_9151);
nor U13978 (N_13978,N_8313,N_5174);
nand U13979 (N_13979,N_6661,N_5862);
nor U13980 (N_13980,N_5338,N_9390);
nand U13981 (N_13981,N_9405,N_6491);
nor U13982 (N_13982,N_5457,N_9322);
nand U13983 (N_13983,N_9870,N_8414);
or U13984 (N_13984,N_8238,N_8510);
nor U13985 (N_13985,N_7119,N_5151);
nor U13986 (N_13986,N_8028,N_8452);
nor U13987 (N_13987,N_6921,N_8319);
or U13988 (N_13988,N_9445,N_7448);
nor U13989 (N_13989,N_7628,N_8879);
or U13990 (N_13990,N_8516,N_6185);
and U13991 (N_13991,N_6954,N_6830);
nor U13992 (N_13992,N_7695,N_6628);
xor U13993 (N_13993,N_6184,N_8711);
and U13994 (N_13994,N_6660,N_7136);
nor U13995 (N_13995,N_5520,N_8298);
and U13996 (N_13996,N_8471,N_5495);
and U13997 (N_13997,N_8579,N_9292);
nand U13998 (N_13998,N_7465,N_9327);
and U13999 (N_13999,N_5452,N_5121);
or U14000 (N_14000,N_6158,N_7450);
xnor U14001 (N_14001,N_5687,N_7551);
and U14002 (N_14002,N_9316,N_9978);
nor U14003 (N_14003,N_5530,N_8251);
xnor U14004 (N_14004,N_5801,N_7751);
and U14005 (N_14005,N_9613,N_8606);
nand U14006 (N_14006,N_8021,N_9136);
xnor U14007 (N_14007,N_5378,N_8476);
nand U14008 (N_14008,N_5511,N_6855);
nand U14009 (N_14009,N_8829,N_6616);
nand U14010 (N_14010,N_5446,N_8095);
or U14011 (N_14011,N_6784,N_7364);
nor U14012 (N_14012,N_5520,N_7637);
xnor U14013 (N_14013,N_5290,N_7213);
xor U14014 (N_14014,N_8308,N_6349);
or U14015 (N_14015,N_7316,N_5432);
and U14016 (N_14016,N_9130,N_9265);
or U14017 (N_14017,N_5038,N_6290);
nor U14018 (N_14018,N_5613,N_6703);
and U14019 (N_14019,N_9991,N_9517);
and U14020 (N_14020,N_6101,N_9196);
or U14021 (N_14021,N_6668,N_7724);
or U14022 (N_14022,N_8252,N_5971);
or U14023 (N_14023,N_6854,N_6510);
xor U14024 (N_14024,N_6984,N_7637);
nand U14025 (N_14025,N_8677,N_6026);
or U14026 (N_14026,N_9152,N_5403);
or U14027 (N_14027,N_7655,N_5627);
and U14028 (N_14028,N_7519,N_7890);
nand U14029 (N_14029,N_9258,N_9908);
nor U14030 (N_14030,N_8705,N_7558);
nor U14031 (N_14031,N_5421,N_6180);
or U14032 (N_14032,N_8959,N_6726);
or U14033 (N_14033,N_6436,N_6634);
and U14034 (N_14034,N_9180,N_6729);
or U14035 (N_14035,N_7977,N_9683);
nor U14036 (N_14036,N_5292,N_7376);
nand U14037 (N_14037,N_5244,N_6770);
and U14038 (N_14038,N_8976,N_5781);
or U14039 (N_14039,N_7335,N_5591);
xnor U14040 (N_14040,N_7306,N_6671);
nand U14041 (N_14041,N_9347,N_5419);
nand U14042 (N_14042,N_5482,N_6270);
and U14043 (N_14043,N_6105,N_9784);
nor U14044 (N_14044,N_9470,N_6151);
and U14045 (N_14045,N_6155,N_8754);
or U14046 (N_14046,N_6080,N_6828);
nor U14047 (N_14047,N_6565,N_6228);
nand U14048 (N_14048,N_5941,N_5713);
and U14049 (N_14049,N_9062,N_7087);
xor U14050 (N_14050,N_9998,N_5513);
nand U14051 (N_14051,N_7643,N_8293);
nor U14052 (N_14052,N_8071,N_8797);
and U14053 (N_14053,N_5985,N_9797);
or U14054 (N_14054,N_8392,N_6271);
nor U14055 (N_14055,N_8932,N_8795);
nand U14056 (N_14056,N_5671,N_8622);
nand U14057 (N_14057,N_5434,N_5279);
and U14058 (N_14058,N_9018,N_8082);
nand U14059 (N_14059,N_5487,N_6901);
nor U14060 (N_14060,N_5103,N_9871);
nand U14061 (N_14061,N_8140,N_6991);
xor U14062 (N_14062,N_5015,N_9173);
nor U14063 (N_14063,N_6035,N_6568);
and U14064 (N_14064,N_5437,N_7992);
nand U14065 (N_14065,N_8592,N_5521);
nor U14066 (N_14066,N_6724,N_7398);
or U14067 (N_14067,N_5745,N_7098);
or U14068 (N_14068,N_6596,N_5949);
nand U14069 (N_14069,N_7724,N_5767);
nand U14070 (N_14070,N_7232,N_8119);
nand U14071 (N_14071,N_9496,N_5491);
or U14072 (N_14072,N_8540,N_9799);
xnor U14073 (N_14073,N_6645,N_9193);
xor U14074 (N_14074,N_9919,N_6007);
nor U14075 (N_14075,N_6025,N_9410);
nand U14076 (N_14076,N_6357,N_6820);
and U14077 (N_14077,N_5205,N_8902);
xnor U14078 (N_14078,N_6899,N_8597);
and U14079 (N_14079,N_6422,N_8471);
nand U14080 (N_14080,N_7476,N_6116);
or U14081 (N_14081,N_7958,N_8403);
nand U14082 (N_14082,N_6306,N_8204);
xnor U14083 (N_14083,N_8104,N_8348);
xor U14084 (N_14084,N_5636,N_7080);
and U14085 (N_14085,N_7524,N_8672);
and U14086 (N_14086,N_8253,N_6984);
or U14087 (N_14087,N_6218,N_6106);
and U14088 (N_14088,N_9984,N_5760);
and U14089 (N_14089,N_6364,N_9790);
and U14090 (N_14090,N_9558,N_5049);
or U14091 (N_14091,N_7747,N_7128);
nor U14092 (N_14092,N_5049,N_5167);
or U14093 (N_14093,N_5673,N_8254);
nand U14094 (N_14094,N_6273,N_9747);
xnor U14095 (N_14095,N_6114,N_6461);
nor U14096 (N_14096,N_5470,N_6887);
or U14097 (N_14097,N_5296,N_8925);
nor U14098 (N_14098,N_7444,N_9843);
nand U14099 (N_14099,N_6095,N_6720);
nand U14100 (N_14100,N_6887,N_6982);
or U14101 (N_14101,N_6909,N_7975);
nor U14102 (N_14102,N_8155,N_5900);
nor U14103 (N_14103,N_9711,N_7205);
or U14104 (N_14104,N_5390,N_9856);
or U14105 (N_14105,N_6783,N_7295);
and U14106 (N_14106,N_5761,N_7789);
and U14107 (N_14107,N_5179,N_9150);
nand U14108 (N_14108,N_7736,N_6543);
and U14109 (N_14109,N_7139,N_7073);
xnor U14110 (N_14110,N_7113,N_9666);
nor U14111 (N_14111,N_6090,N_9019);
or U14112 (N_14112,N_7842,N_8767);
nor U14113 (N_14113,N_5573,N_8338);
nor U14114 (N_14114,N_5687,N_7178);
and U14115 (N_14115,N_8907,N_6267);
nor U14116 (N_14116,N_7071,N_6571);
nor U14117 (N_14117,N_8197,N_8847);
nand U14118 (N_14118,N_7662,N_6349);
nor U14119 (N_14119,N_6180,N_9679);
nand U14120 (N_14120,N_5815,N_8804);
and U14121 (N_14121,N_9310,N_9443);
and U14122 (N_14122,N_5796,N_7757);
nor U14123 (N_14123,N_8044,N_7937);
xor U14124 (N_14124,N_6472,N_9660);
or U14125 (N_14125,N_8300,N_8571);
or U14126 (N_14126,N_5509,N_5302);
nor U14127 (N_14127,N_6097,N_6980);
and U14128 (N_14128,N_9930,N_7698);
nor U14129 (N_14129,N_5164,N_8678);
nand U14130 (N_14130,N_9331,N_9055);
nor U14131 (N_14131,N_7006,N_6374);
or U14132 (N_14132,N_7867,N_6625);
nand U14133 (N_14133,N_5928,N_5165);
and U14134 (N_14134,N_8457,N_6234);
and U14135 (N_14135,N_8181,N_6056);
nor U14136 (N_14136,N_9284,N_6785);
xnor U14137 (N_14137,N_6087,N_8671);
nor U14138 (N_14138,N_8592,N_7489);
and U14139 (N_14139,N_9444,N_5728);
xor U14140 (N_14140,N_6060,N_8674);
or U14141 (N_14141,N_6340,N_6161);
xnor U14142 (N_14142,N_8092,N_8853);
or U14143 (N_14143,N_7039,N_5434);
and U14144 (N_14144,N_5131,N_9039);
xnor U14145 (N_14145,N_8420,N_5132);
and U14146 (N_14146,N_6260,N_7364);
nor U14147 (N_14147,N_5579,N_8989);
or U14148 (N_14148,N_5055,N_9927);
xnor U14149 (N_14149,N_7663,N_7579);
or U14150 (N_14150,N_7538,N_9840);
and U14151 (N_14151,N_8585,N_9896);
nor U14152 (N_14152,N_7613,N_7327);
or U14153 (N_14153,N_5220,N_8144);
or U14154 (N_14154,N_6534,N_5713);
and U14155 (N_14155,N_5133,N_6001);
or U14156 (N_14156,N_7129,N_5957);
or U14157 (N_14157,N_6195,N_7026);
and U14158 (N_14158,N_5662,N_5713);
xor U14159 (N_14159,N_6649,N_5729);
or U14160 (N_14160,N_6928,N_8570);
xnor U14161 (N_14161,N_8140,N_9108);
nor U14162 (N_14162,N_6227,N_7013);
or U14163 (N_14163,N_5121,N_6037);
xor U14164 (N_14164,N_6792,N_7159);
or U14165 (N_14165,N_7481,N_8400);
and U14166 (N_14166,N_6473,N_8060);
nor U14167 (N_14167,N_7060,N_9555);
and U14168 (N_14168,N_7867,N_7152);
nor U14169 (N_14169,N_5868,N_6779);
nor U14170 (N_14170,N_7812,N_5352);
xor U14171 (N_14171,N_7097,N_5776);
xor U14172 (N_14172,N_8969,N_8469);
nand U14173 (N_14173,N_8158,N_8719);
nand U14174 (N_14174,N_6768,N_8493);
xnor U14175 (N_14175,N_8900,N_8216);
xnor U14176 (N_14176,N_5931,N_8652);
xor U14177 (N_14177,N_8278,N_9260);
and U14178 (N_14178,N_7415,N_7935);
nor U14179 (N_14179,N_5667,N_9372);
and U14180 (N_14180,N_7988,N_6972);
nor U14181 (N_14181,N_8389,N_6590);
nor U14182 (N_14182,N_7061,N_8011);
xnor U14183 (N_14183,N_7230,N_7606);
and U14184 (N_14184,N_9435,N_5017);
nor U14185 (N_14185,N_6229,N_5127);
and U14186 (N_14186,N_9816,N_7666);
nor U14187 (N_14187,N_9204,N_9922);
xnor U14188 (N_14188,N_6120,N_7007);
nor U14189 (N_14189,N_8892,N_9996);
nand U14190 (N_14190,N_9240,N_7166);
and U14191 (N_14191,N_9565,N_8744);
nor U14192 (N_14192,N_6332,N_9851);
xnor U14193 (N_14193,N_5897,N_5915);
or U14194 (N_14194,N_8425,N_7088);
xor U14195 (N_14195,N_5088,N_7859);
xnor U14196 (N_14196,N_8056,N_9057);
nor U14197 (N_14197,N_9907,N_9593);
xor U14198 (N_14198,N_9905,N_5986);
xor U14199 (N_14199,N_9043,N_7994);
or U14200 (N_14200,N_9975,N_9297);
nand U14201 (N_14201,N_5931,N_8341);
xor U14202 (N_14202,N_6217,N_7635);
and U14203 (N_14203,N_5755,N_9406);
nor U14204 (N_14204,N_9394,N_9688);
or U14205 (N_14205,N_6487,N_6525);
nand U14206 (N_14206,N_5303,N_9702);
or U14207 (N_14207,N_7998,N_7256);
and U14208 (N_14208,N_6081,N_8154);
or U14209 (N_14209,N_6819,N_9033);
nor U14210 (N_14210,N_7223,N_8152);
nand U14211 (N_14211,N_9809,N_9157);
or U14212 (N_14212,N_7369,N_6003);
and U14213 (N_14213,N_9247,N_6357);
and U14214 (N_14214,N_7970,N_9682);
or U14215 (N_14215,N_6044,N_8952);
nor U14216 (N_14216,N_8605,N_6669);
nor U14217 (N_14217,N_7009,N_6676);
xnor U14218 (N_14218,N_5140,N_5847);
or U14219 (N_14219,N_5899,N_7287);
and U14220 (N_14220,N_9058,N_6330);
nor U14221 (N_14221,N_7747,N_5667);
or U14222 (N_14222,N_6151,N_7593);
nand U14223 (N_14223,N_7712,N_7373);
xor U14224 (N_14224,N_7879,N_6574);
xor U14225 (N_14225,N_8251,N_8434);
and U14226 (N_14226,N_5791,N_5207);
and U14227 (N_14227,N_6546,N_7258);
nand U14228 (N_14228,N_7304,N_6320);
nand U14229 (N_14229,N_8469,N_6035);
xnor U14230 (N_14230,N_8069,N_6812);
or U14231 (N_14231,N_9797,N_6868);
nand U14232 (N_14232,N_6725,N_9965);
nor U14233 (N_14233,N_5125,N_6834);
or U14234 (N_14234,N_6657,N_9974);
or U14235 (N_14235,N_9305,N_8694);
nor U14236 (N_14236,N_6008,N_5930);
or U14237 (N_14237,N_8780,N_9263);
and U14238 (N_14238,N_8182,N_7525);
xnor U14239 (N_14239,N_9079,N_7960);
nand U14240 (N_14240,N_7103,N_9367);
and U14241 (N_14241,N_8985,N_5707);
nand U14242 (N_14242,N_9299,N_7015);
nand U14243 (N_14243,N_7054,N_7295);
nor U14244 (N_14244,N_6715,N_9897);
nor U14245 (N_14245,N_5533,N_5306);
nand U14246 (N_14246,N_5130,N_8664);
nand U14247 (N_14247,N_7663,N_7648);
and U14248 (N_14248,N_8915,N_7533);
and U14249 (N_14249,N_7976,N_9353);
nand U14250 (N_14250,N_6239,N_9595);
xor U14251 (N_14251,N_9346,N_9448);
nand U14252 (N_14252,N_9682,N_8450);
or U14253 (N_14253,N_9055,N_7515);
and U14254 (N_14254,N_5252,N_5774);
and U14255 (N_14255,N_8970,N_8934);
nor U14256 (N_14256,N_7952,N_7585);
nor U14257 (N_14257,N_5464,N_5243);
nor U14258 (N_14258,N_7414,N_6985);
nand U14259 (N_14259,N_5675,N_9377);
nor U14260 (N_14260,N_7444,N_5598);
and U14261 (N_14261,N_6503,N_8547);
and U14262 (N_14262,N_6514,N_6730);
nor U14263 (N_14263,N_8410,N_5002);
xnor U14264 (N_14264,N_5673,N_5680);
or U14265 (N_14265,N_6429,N_5771);
or U14266 (N_14266,N_6800,N_9053);
nand U14267 (N_14267,N_9224,N_8251);
and U14268 (N_14268,N_6095,N_5639);
nor U14269 (N_14269,N_8782,N_9277);
and U14270 (N_14270,N_5993,N_6700);
nand U14271 (N_14271,N_6062,N_6908);
xor U14272 (N_14272,N_8332,N_8370);
nand U14273 (N_14273,N_5120,N_7650);
nor U14274 (N_14274,N_7427,N_7348);
or U14275 (N_14275,N_7143,N_7651);
xnor U14276 (N_14276,N_7015,N_8301);
nand U14277 (N_14277,N_9094,N_5250);
nand U14278 (N_14278,N_6175,N_7789);
and U14279 (N_14279,N_9361,N_5040);
nand U14280 (N_14280,N_5011,N_8398);
nor U14281 (N_14281,N_6290,N_9679);
nor U14282 (N_14282,N_5649,N_7634);
xnor U14283 (N_14283,N_9334,N_9984);
and U14284 (N_14284,N_9497,N_6202);
or U14285 (N_14285,N_5382,N_6976);
xnor U14286 (N_14286,N_5546,N_5528);
xnor U14287 (N_14287,N_9148,N_8191);
xor U14288 (N_14288,N_9446,N_7635);
or U14289 (N_14289,N_8271,N_8247);
xnor U14290 (N_14290,N_5725,N_8025);
and U14291 (N_14291,N_9278,N_9039);
and U14292 (N_14292,N_6084,N_7828);
nand U14293 (N_14293,N_9831,N_8171);
xnor U14294 (N_14294,N_9060,N_9499);
or U14295 (N_14295,N_6403,N_7050);
xnor U14296 (N_14296,N_8532,N_8699);
nand U14297 (N_14297,N_9643,N_8660);
nand U14298 (N_14298,N_9504,N_9376);
or U14299 (N_14299,N_7202,N_9738);
or U14300 (N_14300,N_5431,N_5215);
and U14301 (N_14301,N_7599,N_9596);
xor U14302 (N_14302,N_9747,N_8850);
xor U14303 (N_14303,N_9102,N_7214);
nor U14304 (N_14304,N_6109,N_9408);
and U14305 (N_14305,N_9994,N_7268);
nor U14306 (N_14306,N_6246,N_9128);
nand U14307 (N_14307,N_6058,N_7225);
xor U14308 (N_14308,N_7566,N_8426);
and U14309 (N_14309,N_6105,N_9188);
or U14310 (N_14310,N_5579,N_6990);
or U14311 (N_14311,N_7604,N_6312);
nor U14312 (N_14312,N_6075,N_5403);
xnor U14313 (N_14313,N_5548,N_8826);
and U14314 (N_14314,N_6138,N_9767);
or U14315 (N_14315,N_5937,N_5041);
nor U14316 (N_14316,N_9382,N_7560);
and U14317 (N_14317,N_7156,N_6472);
nand U14318 (N_14318,N_5630,N_8512);
or U14319 (N_14319,N_7246,N_8425);
nand U14320 (N_14320,N_6118,N_8178);
nand U14321 (N_14321,N_5786,N_8803);
and U14322 (N_14322,N_6932,N_6236);
and U14323 (N_14323,N_5711,N_6972);
and U14324 (N_14324,N_8209,N_9187);
or U14325 (N_14325,N_6906,N_9425);
and U14326 (N_14326,N_6626,N_7256);
nand U14327 (N_14327,N_6603,N_6077);
nand U14328 (N_14328,N_9090,N_7785);
and U14329 (N_14329,N_6929,N_8957);
and U14330 (N_14330,N_7355,N_8250);
or U14331 (N_14331,N_6290,N_7259);
nand U14332 (N_14332,N_5777,N_5945);
nand U14333 (N_14333,N_7763,N_7164);
and U14334 (N_14334,N_5120,N_7250);
or U14335 (N_14335,N_6900,N_9058);
nand U14336 (N_14336,N_8196,N_7757);
and U14337 (N_14337,N_8466,N_9563);
xor U14338 (N_14338,N_6451,N_6829);
xnor U14339 (N_14339,N_6361,N_7054);
and U14340 (N_14340,N_5975,N_8158);
xnor U14341 (N_14341,N_6888,N_8132);
and U14342 (N_14342,N_6669,N_8645);
or U14343 (N_14343,N_8944,N_9047);
nor U14344 (N_14344,N_6381,N_5401);
nor U14345 (N_14345,N_9458,N_6859);
or U14346 (N_14346,N_8477,N_6133);
nor U14347 (N_14347,N_5033,N_9604);
nor U14348 (N_14348,N_5891,N_6349);
nor U14349 (N_14349,N_9867,N_9557);
and U14350 (N_14350,N_6313,N_8995);
and U14351 (N_14351,N_6938,N_5102);
xnor U14352 (N_14352,N_6090,N_5848);
xnor U14353 (N_14353,N_7084,N_9107);
or U14354 (N_14354,N_8643,N_7620);
nor U14355 (N_14355,N_8473,N_6902);
nand U14356 (N_14356,N_8145,N_8508);
and U14357 (N_14357,N_6361,N_6499);
or U14358 (N_14358,N_7628,N_7316);
nor U14359 (N_14359,N_6889,N_5257);
and U14360 (N_14360,N_9790,N_8657);
xnor U14361 (N_14361,N_8582,N_7909);
nor U14362 (N_14362,N_8266,N_9158);
and U14363 (N_14363,N_6792,N_8680);
nor U14364 (N_14364,N_5821,N_6714);
nand U14365 (N_14365,N_9933,N_7549);
xor U14366 (N_14366,N_9864,N_5282);
xor U14367 (N_14367,N_6050,N_8091);
xor U14368 (N_14368,N_5972,N_9029);
xor U14369 (N_14369,N_6107,N_5386);
nand U14370 (N_14370,N_8453,N_9943);
nor U14371 (N_14371,N_6426,N_6021);
xnor U14372 (N_14372,N_9887,N_7756);
xor U14373 (N_14373,N_7213,N_6675);
xor U14374 (N_14374,N_9437,N_7523);
and U14375 (N_14375,N_8489,N_7404);
nor U14376 (N_14376,N_6342,N_5632);
xnor U14377 (N_14377,N_8581,N_7252);
nand U14378 (N_14378,N_5927,N_9744);
or U14379 (N_14379,N_9384,N_9273);
nand U14380 (N_14380,N_7576,N_5050);
nand U14381 (N_14381,N_9590,N_8118);
nor U14382 (N_14382,N_7113,N_8270);
or U14383 (N_14383,N_5871,N_5374);
xor U14384 (N_14384,N_5342,N_8403);
nor U14385 (N_14385,N_6432,N_8859);
nand U14386 (N_14386,N_7212,N_7285);
and U14387 (N_14387,N_9157,N_9193);
or U14388 (N_14388,N_6934,N_9786);
nor U14389 (N_14389,N_7705,N_9530);
or U14390 (N_14390,N_9972,N_9980);
or U14391 (N_14391,N_6140,N_8932);
nand U14392 (N_14392,N_5232,N_8292);
or U14393 (N_14393,N_6097,N_9354);
nand U14394 (N_14394,N_5614,N_8609);
or U14395 (N_14395,N_8342,N_8971);
nor U14396 (N_14396,N_6145,N_8874);
xnor U14397 (N_14397,N_6884,N_8253);
xnor U14398 (N_14398,N_5136,N_7696);
or U14399 (N_14399,N_7940,N_9936);
xnor U14400 (N_14400,N_6343,N_5004);
nor U14401 (N_14401,N_9054,N_7849);
or U14402 (N_14402,N_5329,N_8179);
xor U14403 (N_14403,N_9522,N_5794);
and U14404 (N_14404,N_8610,N_5351);
and U14405 (N_14405,N_5966,N_6996);
nor U14406 (N_14406,N_5407,N_8492);
and U14407 (N_14407,N_6068,N_9174);
or U14408 (N_14408,N_9688,N_5774);
nor U14409 (N_14409,N_6014,N_6016);
nor U14410 (N_14410,N_6757,N_8740);
or U14411 (N_14411,N_9786,N_9990);
nor U14412 (N_14412,N_5644,N_7776);
and U14413 (N_14413,N_8385,N_8787);
nor U14414 (N_14414,N_5655,N_9358);
nand U14415 (N_14415,N_9146,N_9814);
and U14416 (N_14416,N_8495,N_7639);
or U14417 (N_14417,N_9621,N_9689);
nand U14418 (N_14418,N_6278,N_9974);
or U14419 (N_14419,N_7380,N_6957);
nand U14420 (N_14420,N_9517,N_7869);
nor U14421 (N_14421,N_6210,N_8575);
nand U14422 (N_14422,N_7843,N_9082);
or U14423 (N_14423,N_6726,N_6694);
xnor U14424 (N_14424,N_5665,N_5681);
and U14425 (N_14425,N_6263,N_8818);
nand U14426 (N_14426,N_8036,N_7960);
nor U14427 (N_14427,N_7709,N_6144);
or U14428 (N_14428,N_8478,N_5996);
xor U14429 (N_14429,N_6238,N_7616);
nor U14430 (N_14430,N_5669,N_6317);
nor U14431 (N_14431,N_5351,N_6020);
or U14432 (N_14432,N_8319,N_9195);
or U14433 (N_14433,N_6545,N_6709);
or U14434 (N_14434,N_9893,N_7334);
and U14435 (N_14435,N_8612,N_5431);
xor U14436 (N_14436,N_7818,N_6627);
nand U14437 (N_14437,N_9015,N_5287);
nand U14438 (N_14438,N_8232,N_9451);
and U14439 (N_14439,N_5360,N_8757);
or U14440 (N_14440,N_6236,N_5987);
or U14441 (N_14441,N_5158,N_5643);
or U14442 (N_14442,N_6561,N_8013);
and U14443 (N_14443,N_9309,N_9077);
nand U14444 (N_14444,N_9189,N_7044);
nand U14445 (N_14445,N_5165,N_6052);
or U14446 (N_14446,N_8801,N_7872);
nor U14447 (N_14447,N_8549,N_5502);
nand U14448 (N_14448,N_8632,N_7919);
nor U14449 (N_14449,N_7709,N_9084);
nor U14450 (N_14450,N_6792,N_6992);
xnor U14451 (N_14451,N_8162,N_9578);
and U14452 (N_14452,N_5771,N_6332);
nand U14453 (N_14453,N_5610,N_6904);
nor U14454 (N_14454,N_5298,N_8001);
and U14455 (N_14455,N_9732,N_6956);
and U14456 (N_14456,N_5646,N_5418);
nor U14457 (N_14457,N_8867,N_5319);
and U14458 (N_14458,N_6677,N_8315);
nor U14459 (N_14459,N_7526,N_8125);
and U14460 (N_14460,N_8488,N_8859);
and U14461 (N_14461,N_7112,N_7738);
xor U14462 (N_14462,N_8075,N_9347);
xnor U14463 (N_14463,N_9166,N_7739);
nand U14464 (N_14464,N_9498,N_8859);
and U14465 (N_14465,N_8065,N_7633);
xnor U14466 (N_14466,N_7226,N_6421);
xnor U14467 (N_14467,N_8150,N_8483);
and U14468 (N_14468,N_5491,N_8425);
nor U14469 (N_14469,N_5489,N_6250);
and U14470 (N_14470,N_7405,N_6095);
or U14471 (N_14471,N_8454,N_8720);
and U14472 (N_14472,N_8406,N_9834);
or U14473 (N_14473,N_8321,N_5418);
or U14474 (N_14474,N_7386,N_9723);
nand U14475 (N_14475,N_6055,N_6336);
or U14476 (N_14476,N_7705,N_6341);
nand U14477 (N_14477,N_9743,N_5273);
and U14478 (N_14478,N_9343,N_6047);
nor U14479 (N_14479,N_9009,N_7907);
nand U14480 (N_14480,N_8794,N_5266);
and U14481 (N_14481,N_9275,N_5106);
nor U14482 (N_14482,N_7091,N_8077);
nand U14483 (N_14483,N_9074,N_9607);
nor U14484 (N_14484,N_7364,N_5639);
nand U14485 (N_14485,N_6853,N_7415);
or U14486 (N_14486,N_7391,N_7258);
and U14487 (N_14487,N_7337,N_9739);
and U14488 (N_14488,N_9738,N_8372);
nand U14489 (N_14489,N_6218,N_8987);
nor U14490 (N_14490,N_7311,N_9937);
nor U14491 (N_14491,N_5865,N_6452);
nand U14492 (N_14492,N_6062,N_5130);
and U14493 (N_14493,N_5380,N_9012);
or U14494 (N_14494,N_5828,N_8400);
nand U14495 (N_14495,N_8177,N_6806);
xnor U14496 (N_14496,N_5099,N_8361);
nand U14497 (N_14497,N_6363,N_7660);
nand U14498 (N_14498,N_7561,N_6455);
xor U14499 (N_14499,N_9720,N_7854);
or U14500 (N_14500,N_7495,N_8196);
nand U14501 (N_14501,N_6038,N_7577);
nand U14502 (N_14502,N_7532,N_9527);
nor U14503 (N_14503,N_7615,N_9530);
and U14504 (N_14504,N_6342,N_5139);
nor U14505 (N_14505,N_9878,N_5780);
or U14506 (N_14506,N_9080,N_5929);
nor U14507 (N_14507,N_8505,N_5594);
and U14508 (N_14508,N_5796,N_8705);
nand U14509 (N_14509,N_5465,N_8906);
xor U14510 (N_14510,N_8807,N_6317);
or U14511 (N_14511,N_6915,N_9909);
or U14512 (N_14512,N_7696,N_8015);
xnor U14513 (N_14513,N_7022,N_7380);
and U14514 (N_14514,N_5948,N_9828);
nand U14515 (N_14515,N_6726,N_5168);
or U14516 (N_14516,N_6810,N_7844);
nand U14517 (N_14517,N_6849,N_9825);
nand U14518 (N_14518,N_6260,N_5130);
or U14519 (N_14519,N_6980,N_6271);
and U14520 (N_14520,N_9221,N_8897);
nor U14521 (N_14521,N_5149,N_9043);
xor U14522 (N_14522,N_6515,N_5257);
xor U14523 (N_14523,N_8047,N_9052);
or U14524 (N_14524,N_8822,N_6689);
nand U14525 (N_14525,N_7614,N_8155);
nand U14526 (N_14526,N_7391,N_7405);
nand U14527 (N_14527,N_9903,N_9893);
xnor U14528 (N_14528,N_7599,N_9966);
nand U14529 (N_14529,N_6672,N_6378);
nand U14530 (N_14530,N_5232,N_6934);
xnor U14531 (N_14531,N_9818,N_5247);
xor U14532 (N_14532,N_8376,N_7344);
nand U14533 (N_14533,N_9561,N_6114);
and U14534 (N_14534,N_7890,N_5624);
nand U14535 (N_14535,N_6096,N_5408);
nor U14536 (N_14536,N_5378,N_6350);
xnor U14537 (N_14537,N_6584,N_7526);
xor U14538 (N_14538,N_6649,N_5177);
and U14539 (N_14539,N_9826,N_6099);
nand U14540 (N_14540,N_5627,N_7406);
nor U14541 (N_14541,N_6552,N_9875);
nand U14542 (N_14542,N_9397,N_8367);
or U14543 (N_14543,N_6794,N_5937);
nor U14544 (N_14544,N_7217,N_5759);
nand U14545 (N_14545,N_8906,N_8535);
or U14546 (N_14546,N_7713,N_7290);
nand U14547 (N_14547,N_7304,N_9016);
nand U14548 (N_14548,N_7869,N_5643);
and U14549 (N_14549,N_9386,N_9421);
xnor U14550 (N_14550,N_5177,N_9900);
or U14551 (N_14551,N_9230,N_7685);
nand U14552 (N_14552,N_9626,N_6390);
xor U14553 (N_14553,N_6942,N_6382);
or U14554 (N_14554,N_7649,N_8863);
xor U14555 (N_14555,N_9324,N_7293);
and U14556 (N_14556,N_7659,N_5821);
or U14557 (N_14557,N_5420,N_9192);
and U14558 (N_14558,N_6869,N_9929);
nand U14559 (N_14559,N_8774,N_8996);
nor U14560 (N_14560,N_8069,N_6904);
nor U14561 (N_14561,N_9444,N_9397);
or U14562 (N_14562,N_8279,N_6521);
or U14563 (N_14563,N_6685,N_6048);
nand U14564 (N_14564,N_7749,N_7842);
or U14565 (N_14565,N_6655,N_8683);
and U14566 (N_14566,N_9390,N_5673);
and U14567 (N_14567,N_8460,N_6487);
and U14568 (N_14568,N_7856,N_5962);
xor U14569 (N_14569,N_7214,N_9080);
or U14570 (N_14570,N_8175,N_8942);
and U14571 (N_14571,N_8712,N_8083);
and U14572 (N_14572,N_6483,N_9302);
nand U14573 (N_14573,N_9762,N_9317);
nand U14574 (N_14574,N_8226,N_6582);
or U14575 (N_14575,N_8034,N_9993);
xor U14576 (N_14576,N_9317,N_7185);
nor U14577 (N_14577,N_5452,N_8774);
xor U14578 (N_14578,N_9205,N_8412);
nand U14579 (N_14579,N_9266,N_6844);
nor U14580 (N_14580,N_8940,N_7190);
nor U14581 (N_14581,N_7049,N_9473);
and U14582 (N_14582,N_9621,N_8125);
nand U14583 (N_14583,N_5188,N_6900);
or U14584 (N_14584,N_5183,N_8949);
nor U14585 (N_14585,N_9344,N_8400);
nor U14586 (N_14586,N_6068,N_9698);
or U14587 (N_14587,N_9591,N_6472);
nor U14588 (N_14588,N_7266,N_9913);
nor U14589 (N_14589,N_9487,N_5040);
nor U14590 (N_14590,N_8611,N_8572);
and U14591 (N_14591,N_6465,N_7230);
or U14592 (N_14592,N_5906,N_8512);
or U14593 (N_14593,N_8184,N_7679);
xnor U14594 (N_14594,N_7805,N_7437);
or U14595 (N_14595,N_5940,N_6347);
nor U14596 (N_14596,N_9937,N_7710);
nor U14597 (N_14597,N_8892,N_5562);
or U14598 (N_14598,N_6647,N_8161);
nand U14599 (N_14599,N_5337,N_7584);
xor U14600 (N_14600,N_9121,N_6781);
and U14601 (N_14601,N_7378,N_5165);
nand U14602 (N_14602,N_7630,N_6555);
and U14603 (N_14603,N_9824,N_8964);
xnor U14604 (N_14604,N_8132,N_9099);
and U14605 (N_14605,N_9050,N_9156);
or U14606 (N_14606,N_8573,N_5749);
xor U14607 (N_14607,N_9294,N_9223);
xnor U14608 (N_14608,N_8879,N_5506);
nor U14609 (N_14609,N_7741,N_9180);
and U14610 (N_14610,N_8361,N_6701);
nor U14611 (N_14611,N_5516,N_8712);
nor U14612 (N_14612,N_8396,N_6263);
or U14613 (N_14613,N_5850,N_8028);
or U14614 (N_14614,N_7249,N_8819);
and U14615 (N_14615,N_6806,N_9995);
or U14616 (N_14616,N_6154,N_5634);
nor U14617 (N_14617,N_9455,N_5877);
or U14618 (N_14618,N_8279,N_8312);
and U14619 (N_14619,N_7952,N_7249);
nor U14620 (N_14620,N_8802,N_9214);
nor U14621 (N_14621,N_7550,N_8546);
or U14622 (N_14622,N_7582,N_7178);
or U14623 (N_14623,N_6073,N_5062);
xnor U14624 (N_14624,N_9482,N_9307);
and U14625 (N_14625,N_7399,N_6447);
nand U14626 (N_14626,N_6535,N_8404);
xor U14627 (N_14627,N_9368,N_6526);
nor U14628 (N_14628,N_8342,N_6277);
nor U14629 (N_14629,N_6657,N_9306);
or U14630 (N_14630,N_6012,N_6526);
xnor U14631 (N_14631,N_5166,N_9137);
xor U14632 (N_14632,N_9823,N_5867);
xor U14633 (N_14633,N_9675,N_5671);
nor U14634 (N_14634,N_6979,N_7667);
and U14635 (N_14635,N_5645,N_5397);
xor U14636 (N_14636,N_5833,N_6234);
nor U14637 (N_14637,N_8405,N_5523);
nor U14638 (N_14638,N_6613,N_7272);
nor U14639 (N_14639,N_9835,N_7010);
nand U14640 (N_14640,N_8446,N_8101);
nand U14641 (N_14641,N_8103,N_5681);
or U14642 (N_14642,N_7966,N_9865);
and U14643 (N_14643,N_6896,N_9374);
or U14644 (N_14644,N_8244,N_8743);
or U14645 (N_14645,N_9006,N_9329);
nand U14646 (N_14646,N_6515,N_9410);
or U14647 (N_14647,N_5207,N_6869);
nor U14648 (N_14648,N_6559,N_9232);
or U14649 (N_14649,N_9068,N_9900);
and U14650 (N_14650,N_7448,N_5614);
nor U14651 (N_14651,N_6848,N_5561);
nor U14652 (N_14652,N_7781,N_9423);
nor U14653 (N_14653,N_8027,N_9121);
nor U14654 (N_14654,N_9244,N_6899);
xnor U14655 (N_14655,N_8218,N_9991);
or U14656 (N_14656,N_6548,N_7648);
nor U14657 (N_14657,N_8338,N_9909);
or U14658 (N_14658,N_5277,N_6588);
xnor U14659 (N_14659,N_9503,N_9324);
xnor U14660 (N_14660,N_9458,N_8267);
and U14661 (N_14661,N_5701,N_9325);
and U14662 (N_14662,N_9048,N_7019);
nand U14663 (N_14663,N_7330,N_7557);
nor U14664 (N_14664,N_7216,N_7053);
or U14665 (N_14665,N_6715,N_6181);
xnor U14666 (N_14666,N_7863,N_7403);
or U14667 (N_14667,N_5117,N_7147);
xnor U14668 (N_14668,N_9473,N_6105);
nor U14669 (N_14669,N_9758,N_9654);
and U14670 (N_14670,N_5012,N_8972);
or U14671 (N_14671,N_6505,N_9064);
and U14672 (N_14672,N_6613,N_6595);
and U14673 (N_14673,N_7558,N_5149);
xor U14674 (N_14674,N_6777,N_5268);
and U14675 (N_14675,N_5801,N_9718);
nor U14676 (N_14676,N_9942,N_5036);
and U14677 (N_14677,N_5856,N_6215);
nand U14678 (N_14678,N_5130,N_5999);
nand U14679 (N_14679,N_9572,N_8210);
or U14680 (N_14680,N_7936,N_7784);
nor U14681 (N_14681,N_6556,N_7057);
and U14682 (N_14682,N_5222,N_9686);
or U14683 (N_14683,N_8170,N_5619);
and U14684 (N_14684,N_8596,N_7228);
and U14685 (N_14685,N_5438,N_8333);
nand U14686 (N_14686,N_7435,N_9244);
and U14687 (N_14687,N_8009,N_5954);
xor U14688 (N_14688,N_9605,N_5613);
or U14689 (N_14689,N_9528,N_7344);
nand U14690 (N_14690,N_6453,N_7424);
or U14691 (N_14691,N_7930,N_5673);
nor U14692 (N_14692,N_5410,N_9304);
nor U14693 (N_14693,N_9372,N_6052);
xor U14694 (N_14694,N_9902,N_5516);
nor U14695 (N_14695,N_8190,N_6696);
nand U14696 (N_14696,N_9131,N_5456);
nand U14697 (N_14697,N_7946,N_7037);
and U14698 (N_14698,N_7738,N_6345);
nor U14699 (N_14699,N_6255,N_8528);
nor U14700 (N_14700,N_9500,N_9105);
nor U14701 (N_14701,N_8561,N_6711);
and U14702 (N_14702,N_7431,N_9602);
nor U14703 (N_14703,N_9958,N_5283);
nand U14704 (N_14704,N_6019,N_6341);
nand U14705 (N_14705,N_8437,N_9007);
or U14706 (N_14706,N_6300,N_7961);
nand U14707 (N_14707,N_6746,N_7264);
nand U14708 (N_14708,N_8681,N_5778);
nor U14709 (N_14709,N_8057,N_8569);
nand U14710 (N_14710,N_9909,N_7468);
nand U14711 (N_14711,N_5133,N_9380);
nand U14712 (N_14712,N_7440,N_9640);
xor U14713 (N_14713,N_9811,N_9739);
and U14714 (N_14714,N_8044,N_9628);
xnor U14715 (N_14715,N_9409,N_7188);
and U14716 (N_14716,N_9676,N_7525);
and U14717 (N_14717,N_9580,N_8578);
or U14718 (N_14718,N_9540,N_7009);
and U14719 (N_14719,N_6391,N_8423);
xor U14720 (N_14720,N_6312,N_8214);
or U14721 (N_14721,N_8340,N_5988);
and U14722 (N_14722,N_7575,N_7104);
and U14723 (N_14723,N_7890,N_8940);
and U14724 (N_14724,N_8453,N_6074);
and U14725 (N_14725,N_5675,N_6470);
and U14726 (N_14726,N_9991,N_8720);
and U14727 (N_14727,N_9465,N_7026);
nand U14728 (N_14728,N_5735,N_7364);
or U14729 (N_14729,N_8653,N_6228);
nor U14730 (N_14730,N_9571,N_7548);
xnor U14731 (N_14731,N_5797,N_9513);
nor U14732 (N_14732,N_5944,N_7102);
and U14733 (N_14733,N_7086,N_8891);
nand U14734 (N_14734,N_6405,N_8230);
xor U14735 (N_14735,N_6835,N_8901);
xnor U14736 (N_14736,N_9775,N_6290);
nor U14737 (N_14737,N_7856,N_9001);
or U14738 (N_14738,N_8648,N_7629);
or U14739 (N_14739,N_5220,N_7362);
or U14740 (N_14740,N_8315,N_5304);
xor U14741 (N_14741,N_9187,N_9857);
and U14742 (N_14742,N_8592,N_8525);
nor U14743 (N_14743,N_5780,N_5103);
nand U14744 (N_14744,N_5661,N_8865);
nand U14745 (N_14745,N_7753,N_7290);
xor U14746 (N_14746,N_7172,N_9951);
nor U14747 (N_14747,N_5041,N_5046);
nand U14748 (N_14748,N_6393,N_6448);
nor U14749 (N_14749,N_6960,N_8024);
xor U14750 (N_14750,N_6947,N_7741);
or U14751 (N_14751,N_8727,N_7429);
or U14752 (N_14752,N_5772,N_6295);
nor U14753 (N_14753,N_5196,N_6642);
or U14754 (N_14754,N_9591,N_9262);
nand U14755 (N_14755,N_9438,N_7562);
nand U14756 (N_14756,N_7373,N_8280);
nor U14757 (N_14757,N_8144,N_5424);
or U14758 (N_14758,N_9668,N_8079);
or U14759 (N_14759,N_7396,N_5716);
or U14760 (N_14760,N_7513,N_6727);
and U14761 (N_14761,N_8352,N_8392);
xor U14762 (N_14762,N_6902,N_9452);
nand U14763 (N_14763,N_5962,N_7913);
and U14764 (N_14764,N_5200,N_9840);
xor U14765 (N_14765,N_7053,N_6925);
and U14766 (N_14766,N_7574,N_8803);
or U14767 (N_14767,N_5364,N_6929);
xor U14768 (N_14768,N_8169,N_7976);
nor U14769 (N_14769,N_6781,N_7443);
nor U14770 (N_14770,N_5309,N_8340);
nor U14771 (N_14771,N_5128,N_5352);
and U14772 (N_14772,N_6386,N_7975);
nor U14773 (N_14773,N_7564,N_9189);
and U14774 (N_14774,N_5427,N_8811);
and U14775 (N_14775,N_6614,N_7465);
or U14776 (N_14776,N_6925,N_8212);
and U14777 (N_14777,N_6637,N_5635);
nor U14778 (N_14778,N_9985,N_7493);
and U14779 (N_14779,N_5440,N_5060);
nand U14780 (N_14780,N_6379,N_8483);
or U14781 (N_14781,N_9261,N_8355);
and U14782 (N_14782,N_7170,N_8326);
and U14783 (N_14783,N_5037,N_6579);
xnor U14784 (N_14784,N_5198,N_6478);
xnor U14785 (N_14785,N_6570,N_5565);
xor U14786 (N_14786,N_6602,N_5861);
nor U14787 (N_14787,N_6461,N_8977);
xor U14788 (N_14788,N_8116,N_8082);
nand U14789 (N_14789,N_5022,N_6350);
nand U14790 (N_14790,N_8148,N_9392);
or U14791 (N_14791,N_5435,N_9959);
nor U14792 (N_14792,N_7459,N_8095);
nor U14793 (N_14793,N_8977,N_9678);
xor U14794 (N_14794,N_5405,N_7087);
nor U14795 (N_14795,N_5775,N_6220);
xor U14796 (N_14796,N_6455,N_9301);
nor U14797 (N_14797,N_5083,N_6791);
nor U14798 (N_14798,N_7263,N_9901);
xnor U14799 (N_14799,N_7860,N_8500);
nand U14800 (N_14800,N_8667,N_9623);
or U14801 (N_14801,N_8746,N_8721);
nand U14802 (N_14802,N_8654,N_9292);
nor U14803 (N_14803,N_6969,N_5047);
nor U14804 (N_14804,N_6224,N_6979);
xor U14805 (N_14805,N_8929,N_9580);
or U14806 (N_14806,N_7633,N_7468);
nand U14807 (N_14807,N_5646,N_5199);
xnor U14808 (N_14808,N_7620,N_7926);
nand U14809 (N_14809,N_9255,N_6336);
nand U14810 (N_14810,N_9841,N_6234);
nand U14811 (N_14811,N_6283,N_7587);
or U14812 (N_14812,N_6549,N_7163);
and U14813 (N_14813,N_5461,N_7542);
nor U14814 (N_14814,N_9933,N_6888);
nor U14815 (N_14815,N_6244,N_5768);
xnor U14816 (N_14816,N_7549,N_6642);
nor U14817 (N_14817,N_5663,N_7561);
nand U14818 (N_14818,N_6009,N_8583);
nor U14819 (N_14819,N_8154,N_8834);
nor U14820 (N_14820,N_5557,N_7368);
nor U14821 (N_14821,N_9036,N_7914);
nand U14822 (N_14822,N_5892,N_8216);
nand U14823 (N_14823,N_5687,N_6676);
nand U14824 (N_14824,N_5743,N_9643);
xnor U14825 (N_14825,N_8197,N_6882);
or U14826 (N_14826,N_9517,N_8921);
and U14827 (N_14827,N_8102,N_6428);
nand U14828 (N_14828,N_5232,N_9407);
nor U14829 (N_14829,N_8882,N_9330);
nand U14830 (N_14830,N_7618,N_8234);
nor U14831 (N_14831,N_5588,N_9758);
or U14832 (N_14832,N_9168,N_5056);
xor U14833 (N_14833,N_8187,N_7049);
nor U14834 (N_14834,N_8306,N_6180);
xor U14835 (N_14835,N_6832,N_9328);
or U14836 (N_14836,N_8225,N_5010);
nor U14837 (N_14837,N_6056,N_5123);
xor U14838 (N_14838,N_9357,N_5016);
and U14839 (N_14839,N_8555,N_8745);
xnor U14840 (N_14840,N_8867,N_8300);
xnor U14841 (N_14841,N_7445,N_7877);
or U14842 (N_14842,N_6852,N_7759);
nor U14843 (N_14843,N_5238,N_8910);
nand U14844 (N_14844,N_6565,N_9977);
or U14845 (N_14845,N_8884,N_7416);
or U14846 (N_14846,N_6381,N_5849);
or U14847 (N_14847,N_6713,N_7473);
xnor U14848 (N_14848,N_8007,N_5994);
nand U14849 (N_14849,N_7473,N_5598);
or U14850 (N_14850,N_7221,N_6493);
nor U14851 (N_14851,N_7528,N_5271);
or U14852 (N_14852,N_8316,N_6237);
xor U14853 (N_14853,N_7090,N_7021);
and U14854 (N_14854,N_5583,N_6627);
nand U14855 (N_14855,N_8982,N_8897);
nor U14856 (N_14856,N_5157,N_7017);
nor U14857 (N_14857,N_6842,N_8922);
nand U14858 (N_14858,N_8056,N_6709);
nand U14859 (N_14859,N_7371,N_5246);
and U14860 (N_14860,N_7852,N_6083);
nor U14861 (N_14861,N_5484,N_8000);
and U14862 (N_14862,N_9346,N_7408);
nand U14863 (N_14863,N_8931,N_7104);
xnor U14864 (N_14864,N_8530,N_7906);
and U14865 (N_14865,N_8842,N_5701);
nand U14866 (N_14866,N_8127,N_9958);
xnor U14867 (N_14867,N_9463,N_6877);
xor U14868 (N_14868,N_5917,N_8311);
xnor U14869 (N_14869,N_6990,N_7343);
nand U14870 (N_14870,N_6906,N_9675);
xor U14871 (N_14871,N_7273,N_9775);
or U14872 (N_14872,N_6890,N_6807);
nand U14873 (N_14873,N_5221,N_6197);
nand U14874 (N_14874,N_8381,N_6947);
or U14875 (N_14875,N_5170,N_7246);
or U14876 (N_14876,N_7908,N_9486);
or U14877 (N_14877,N_7991,N_6183);
nand U14878 (N_14878,N_8065,N_9527);
xor U14879 (N_14879,N_8557,N_5678);
nor U14880 (N_14880,N_8247,N_6202);
and U14881 (N_14881,N_8169,N_9661);
and U14882 (N_14882,N_6482,N_6604);
or U14883 (N_14883,N_9230,N_9085);
nor U14884 (N_14884,N_8370,N_9930);
or U14885 (N_14885,N_6803,N_5737);
and U14886 (N_14886,N_7264,N_9437);
nor U14887 (N_14887,N_6033,N_5493);
xnor U14888 (N_14888,N_5764,N_8232);
or U14889 (N_14889,N_9531,N_7848);
nand U14890 (N_14890,N_5242,N_7759);
or U14891 (N_14891,N_7235,N_9168);
nand U14892 (N_14892,N_8356,N_7680);
and U14893 (N_14893,N_7045,N_5288);
or U14894 (N_14894,N_5652,N_9003);
and U14895 (N_14895,N_8463,N_6865);
nand U14896 (N_14896,N_6692,N_9048);
xor U14897 (N_14897,N_7222,N_6675);
and U14898 (N_14898,N_7414,N_5399);
or U14899 (N_14899,N_7712,N_7688);
and U14900 (N_14900,N_6112,N_8008);
and U14901 (N_14901,N_6453,N_9390);
nor U14902 (N_14902,N_5637,N_7631);
or U14903 (N_14903,N_9600,N_5266);
nor U14904 (N_14904,N_6183,N_9749);
xor U14905 (N_14905,N_9173,N_5765);
xor U14906 (N_14906,N_5789,N_8029);
or U14907 (N_14907,N_5836,N_8725);
nand U14908 (N_14908,N_5477,N_7974);
and U14909 (N_14909,N_6850,N_5908);
xor U14910 (N_14910,N_7962,N_9433);
nand U14911 (N_14911,N_7332,N_7323);
nor U14912 (N_14912,N_8145,N_5976);
and U14913 (N_14913,N_5011,N_9022);
nand U14914 (N_14914,N_7000,N_5804);
xor U14915 (N_14915,N_8933,N_6166);
nand U14916 (N_14916,N_9616,N_7295);
xnor U14917 (N_14917,N_7589,N_9651);
nand U14918 (N_14918,N_9900,N_8912);
or U14919 (N_14919,N_8458,N_7606);
nor U14920 (N_14920,N_8748,N_8874);
nand U14921 (N_14921,N_7811,N_9008);
xor U14922 (N_14922,N_8399,N_5616);
nor U14923 (N_14923,N_5734,N_9836);
nor U14924 (N_14924,N_8031,N_7717);
nor U14925 (N_14925,N_6446,N_8952);
and U14926 (N_14926,N_5301,N_7583);
nand U14927 (N_14927,N_9450,N_7853);
and U14928 (N_14928,N_5034,N_7414);
xor U14929 (N_14929,N_7307,N_5809);
and U14930 (N_14930,N_7578,N_6261);
or U14931 (N_14931,N_9199,N_6521);
nor U14932 (N_14932,N_7445,N_5022);
nor U14933 (N_14933,N_7017,N_8072);
nor U14934 (N_14934,N_5388,N_8101);
xnor U14935 (N_14935,N_8362,N_5438);
and U14936 (N_14936,N_9666,N_8496);
nor U14937 (N_14937,N_9459,N_7060);
nand U14938 (N_14938,N_8255,N_8537);
or U14939 (N_14939,N_6385,N_5533);
nand U14940 (N_14940,N_9905,N_6681);
nor U14941 (N_14941,N_8909,N_5433);
nand U14942 (N_14942,N_7525,N_9771);
nand U14943 (N_14943,N_8207,N_5776);
or U14944 (N_14944,N_7871,N_9967);
nor U14945 (N_14945,N_7184,N_5569);
nor U14946 (N_14946,N_6020,N_8503);
xor U14947 (N_14947,N_8693,N_5069);
nor U14948 (N_14948,N_9849,N_9041);
nand U14949 (N_14949,N_8031,N_7607);
nand U14950 (N_14950,N_9341,N_7452);
and U14951 (N_14951,N_6284,N_8802);
xnor U14952 (N_14952,N_6909,N_5718);
and U14953 (N_14953,N_7424,N_8690);
nand U14954 (N_14954,N_9672,N_7206);
xnor U14955 (N_14955,N_8422,N_8177);
nor U14956 (N_14956,N_5283,N_5053);
nor U14957 (N_14957,N_7168,N_7622);
or U14958 (N_14958,N_9237,N_6826);
nand U14959 (N_14959,N_8695,N_9626);
xor U14960 (N_14960,N_5707,N_7569);
nand U14961 (N_14961,N_5739,N_6459);
or U14962 (N_14962,N_6398,N_6967);
xnor U14963 (N_14963,N_5894,N_5244);
nor U14964 (N_14964,N_9553,N_5605);
and U14965 (N_14965,N_7000,N_7361);
or U14966 (N_14966,N_8115,N_7199);
and U14967 (N_14967,N_9280,N_6127);
nor U14968 (N_14968,N_5926,N_9144);
and U14969 (N_14969,N_8664,N_9751);
or U14970 (N_14970,N_6066,N_8188);
nor U14971 (N_14971,N_7659,N_8576);
or U14972 (N_14972,N_5189,N_6577);
nand U14973 (N_14973,N_8238,N_8160);
or U14974 (N_14974,N_5150,N_6374);
and U14975 (N_14975,N_8724,N_9433);
nor U14976 (N_14976,N_9620,N_7050);
nand U14977 (N_14977,N_6218,N_7735);
or U14978 (N_14978,N_7381,N_7408);
and U14979 (N_14979,N_6158,N_7344);
nor U14980 (N_14980,N_6456,N_6135);
or U14981 (N_14981,N_8777,N_8336);
nor U14982 (N_14982,N_8089,N_8681);
or U14983 (N_14983,N_8566,N_8775);
or U14984 (N_14984,N_8956,N_7408);
xnor U14985 (N_14985,N_5066,N_5557);
and U14986 (N_14986,N_8407,N_5857);
and U14987 (N_14987,N_7148,N_5710);
nand U14988 (N_14988,N_6247,N_7336);
nand U14989 (N_14989,N_7058,N_6691);
xor U14990 (N_14990,N_9249,N_6467);
nand U14991 (N_14991,N_7448,N_6482);
xnor U14992 (N_14992,N_7637,N_7812);
nand U14993 (N_14993,N_5391,N_9947);
xnor U14994 (N_14994,N_6676,N_6339);
and U14995 (N_14995,N_6967,N_9188);
or U14996 (N_14996,N_7845,N_6259);
nor U14997 (N_14997,N_9344,N_6040);
and U14998 (N_14998,N_6516,N_6717);
nor U14999 (N_14999,N_9273,N_5265);
xnor UO_0 (O_0,N_14530,N_12327);
xnor UO_1 (O_1,N_11996,N_11050);
nor UO_2 (O_2,N_13503,N_12713);
nand UO_3 (O_3,N_11049,N_10664);
and UO_4 (O_4,N_12503,N_13092);
or UO_5 (O_5,N_13230,N_13740);
and UO_6 (O_6,N_13269,N_14215);
xor UO_7 (O_7,N_13594,N_13150);
nand UO_8 (O_8,N_10954,N_11091);
xnor UO_9 (O_9,N_10724,N_11337);
nand UO_10 (O_10,N_13001,N_12818);
nor UO_11 (O_11,N_10304,N_11123);
or UO_12 (O_12,N_10593,N_12069);
or UO_13 (O_13,N_10982,N_10950);
nor UO_14 (O_14,N_14421,N_13499);
xnor UO_15 (O_15,N_13517,N_13931);
nand UO_16 (O_16,N_13577,N_13544);
xor UO_17 (O_17,N_10101,N_10678);
nor UO_18 (O_18,N_11006,N_11412);
xor UO_19 (O_19,N_11712,N_10334);
and UO_20 (O_20,N_14265,N_14484);
xnor UO_21 (O_21,N_11113,N_12320);
or UO_22 (O_22,N_12902,N_12598);
nand UO_23 (O_23,N_14678,N_13134);
and UO_24 (O_24,N_13378,N_11786);
nor UO_25 (O_25,N_14982,N_14953);
nand UO_26 (O_26,N_14842,N_13601);
nor UO_27 (O_27,N_14791,N_14451);
and UO_28 (O_28,N_14980,N_10415);
xnor UO_29 (O_29,N_12367,N_14622);
and UO_30 (O_30,N_10327,N_11731);
nor UO_31 (O_31,N_12502,N_14985);
xor UO_32 (O_32,N_12858,N_14337);
nand UO_33 (O_33,N_12872,N_12197);
or UO_34 (O_34,N_10467,N_14814);
and UO_35 (O_35,N_14464,N_11410);
xor UO_36 (O_36,N_11755,N_12315);
xor UO_37 (O_37,N_11235,N_12224);
or UO_38 (O_38,N_11945,N_11707);
nand UO_39 (O_39,N_12838,N_14684);
nor UO_40 (O_40,N_10994,N_12391);
or UO_41 (O_41,N_11082,N_12664);
xor UO_42 (O_42,N_14778,N_13535);
nand UO_43 (O_43,N_14359,N_14685);
and UO_44 (O_44,N_11210,N_11851);
nand UO_45 (O_45,N_12677,N_11704);
or UO_46 (O_46,N_11879,N_11663);
and UO_47 (O_47,N_11402,N_13272);
and UO_48 (O_48,N_14015,N_14206);
and UO_49 (O_49,N_11703,N_10707);
nand UO_50 (O_50,N_13438,N_10516);
and UO_51 (O_51,N_13158,N_14368);
or UO_52 (O_52,N_14094,N_13864);
or UO_53 (O_53,N_10591,N_11459);
nand UO_54 (O_54,N_14029,N_11368);
xnor UO_55 (O_55,N_13971,N_11422);
xor UO_56 (O_56,N_13338,N_10661);
nor UO_57 (O_57,N_11333,N_14146);
nor UO_58 (O_58,N_11365,N_14793);
xnor UO_59 (O_59,N_10945,N_14382);
and UO_60 (O_60,N_14351,N_10603);
nand UO_61 (O_61,N_12030,N_13953);
nor UO_62 (O_62,N_12336,N_12715);
or UO_63 (O_63,N_11407,N_11685);
nor UO_64 (O_64,N_14097,N_13390);
and UO_65 (O_65,N_12341,N_10692);
or UO_66 (O_66,N_14922,N_10976);
nor UO_67 (O_67,N_10372,N_10310);
nor UO_68 (O_68,N_13321,N_11386);
nand UO_69 (O_69,N_10790,N_10818);
nand UO_70 (O_70,N_13500,N_14560);
or UO_71 (O_71,N_14873,N_10739);
xor UO_72 (O_72,N_13729,N_11285);
nor UO_73 (O_73,N_10071,N_11668);
nand UO_74 (O_74,N_14396,N_11093);
nand UO_75 (O_75,N_13606,N_14690);
or UO_76 (O_76,N_11983,N_12092);
nor UO_77 (O_77,N_12509,N_11366);
nor UO_78 (O_78,N_13944,N_13485);
xor UO_79 (O_79,N_11022,N_11071);
and UO_80 (O_80,N_13682,N_13068);
nor UO_81 (O_81,N_10972,N_13524);
nor UO_82 (O_82,N_14027,N_13016);
or UO_83 (O_83,N_10640,N_12692);
xnor UO_84 (O_84,N_10674,N_13012);
or UO_85 (O_85,N_12082,N_12089);
nor UO_86 (O_86,N_13827,N_12255);
nand UO_87 (O_87,N_13198,N_12786);
or UO_88 (O_88,N_14978,N_11261);
and UO_89 (O_89,N_13803,N_10180);
and UO_90 (O_90,N_10620,N_11315);
and UO_91 (O_91,N_13849,N_10051);
xnor UO_92 (O_92,N_11832,N_11721);
xor UO_93 (O_93,N_12409,N_10813);
and UO_94 (O_94,N_11545,N_10480);
xnor UO_95 (O_95,N_13315,N_10019);
or UO_96 (O_96,N_11000,N_14118);
nand UO_97 (O_97,N_12694,N_11966);
and UO_98 (O_98,N_12100,N_13916);
xor UO_99 (O_99,N_13200,N_11438);
nand UO_100 (O_100,N_11608,N_11310);
or UO_101 (O_101,N_12987,N_12157);
xnor UO_102 (O_102,N_13534,N_11468);
nor UO_103 (O_103,N_11498,N_12569);
nand UO_104 (O_104,N_10965,N_12526);
and UO_105 (O_105,N_11259,N_14030);
or UO_106 (O_106,N_11530,N_13239);
and UO_107 (O_107,N_10733,N_13800);
and UO_108 (O_108,N_10748,N_13954);
or UO_109 (O_109,N_10393,N_13723);
xor UO_110 (O_110,N_10219,N_10424);
xor UO_111 (O_111,N_10884,N_11348);
and UO_112 (O_112,N_10123,N_11487);
nor UO_113 (O_113,N_14525,N_11859);
and UO_114 (O_114,N_11393,N_11780);
nand UO_115 (O_115,N_14649,N_14944);
nand UO_116 (O_116,N_14743,N_12477);
nor UO_117 (O_117,N_10951,N_11497);
or UO_118 (O_118,N_11409,N_13402);
or UO_119 (O_119,N_13757,N_14531);
and UO_120 (O_120,N_13293,N_12777);
and UO_121 (O_121,N_13764,N_12400);
xor UO_122 (O_122,N_14967,N_14420);
nor UO_123 (O_123,N_10969,N_14900);
nand UO_124 (O_124,N_14458,N_11522);
nand UO_125 (O_125,N_10249,N_13069);
and UO_126 (O_126,N_10187,N_11566);
nor UO_127 (O_127,N_12175,N_11757);
nor UO_128 (O_128,N_12994,N_14223);
and UO_129 (O_129,N_11930,N_14557);
xnor UO_130 (O_130,N_11538,N_11650);
xor UO_131 (O_131,N_13486,N_12669);
and UO_132 (O_132,N_11248,N_10611);
nor UO_133 (O_133,N_10040,N_14954);
xnor UO_134 (O_134,N_14467,N_14833);
nor UO_135 (O_135,N_13103,N_12107);
and UO_136 (O_136,N_12035,N_11100);
and UO_137 (O_137,N_12130,N_12771);
or UO_138 (O_138,N_14772,N_14960);
nor UO_139 (O_139,N_12024,N_13368);
xor UO_140 (O_140,N_10181,N_14958);
nand UO_141 (O_141,N_10117,N_13162);
nor UO_142 (O_142,N_14492,N_14242);
or UO_143 (O_143,N_10490,N_14611);
or UO_144 (O_144,N_13060,N_10523);
xnor UO_145 (O_145,N_12889,N_14164);
nor UO_146 (O_146,N_10358,N_10789);
or UO_147 (O_147,N_14241,N_14113);
nand UO_148 (O_148,N_14911,N_11536);
nor UO_149 (O_149,N_13000,N_14823);
or UO_150 (O_150,N_12769,N_13354);
and UO_151 (O_151,N_12155,N_13648);
or UO_152 (O_152,N_13874,N_12952);
xnor UO_153 (O_153,N_10229,N_12439);
nor UO_154 (O_154,N_13169,N_14133);
nor UO_155 (O_155,N_10518,N_10094);
xor UO_156 (O_156,N_13733,N_13192);
and UO_157 (O_157,N_12856,N_13151);
and UO_158 (O_158,N_10305,N_13048);
and UO_159 (O_159,N_13624,N_14219);
xnor UO_160 (O_160,N_14719,N_12532);
xnor UO_161 (O_161,N_13231,N_14427);
and UO_162 (O_162,N_11234,N_14835);
nand UO_163 (O_163,N_13703,N_14295);
or UO_164 (O_164,N_12279,N_12547);
nand UO_165 (O_165,N_11787,N_11576);
xnor UO_166 (O_166,N_12448,N_14274);
nand UO_167 (O_167,N_13718,N_13867);
and UO_168 (O_168,N_10171,N_14992);
and UO_169 (O_169,N_12198,N_12955);
nor UO_170 (O_170,N_11766,N_12142);
or UO_171 (O_171,N_11301,N_13223);
and UO_172 (O_172,N_13132,N_10000);
xor UO_173 (O_173,N_11726,N_14808);
nor UO_174 (O_174,N_14091,N_11958);
xnor UO_175 (O_175,N_11687,N_14800);
and UO_176 (O_176,N_13118,N_11026);
xnor UO_177 (O_177,N_11299,N_12621);
nor UO_178 (O_178,N_10909,N_10460);
xor UO_179 (O_179,N_13090,N_13398);
nand UO_180 (O_180,N_11223,N_14306);
nand UO_181 (O_181,N_11122,N_13545);
and UO_182 (O_182,N_14312,N_14682);
nor UO_183 (O_183,N_10957,N_10793);
or UO_184 (O_184,N_11702,N_13256);
nand UO_185 (O_185,N_14576,N_14618);
nand UO_186 (O_186,N_13879,N_13082);
or UO_187 (O_187,N_11451,N_10428);
nor UO_188 (O_188,N_10411,N_14613);
nand UO_189 (O_189,N_11253,N_14184);
nor UO_190 (O_190,N_13114,N_13769);
or UO_191 (O_191,N_11225,N_14775);
and UO_192 (O_192,N_13309,N_13749);
nor UO_193 (O_193,N_13843,N_11920);
nor UO_194 (O_194,N_10588,N_10336);
xor UO_195 (O_195,N_14086,N_10226);
nor UO_196 (O_196,N_10092,N_11985);
nor UO_197 (O_197,N_11676,N_14018);
xor UO_198 (O_198,N_12779,N_12529);
nand UO_199 (O_199,N_10551,N_11053);
nor UO_200 (O_200,N_12938,N_14756);
nor UO_201 (O_201,N_13014,N_10289);
and UO_202 (O_202,N_10996,N_14986);
and UO_203 (O_203,N_14709,N_14154);
xor UO_204 (O_204,N_10183,N_13887);
nor UO_205 (O_205,N_13586,N_13182);
xor UO_206 (O_206,N_14221,N_10010);
or UO_207 (O_207,N_11743,N_11723);
or UO_208 (O_208,N_13728,N_14783);
xnor UO_209 (O_209,N_12049,N_10280);
xor UO_210 (O_210,N_14822,N_11471);
nand UO_211 (O_211,N_13033,N_13999);
nor UO_212 (O_212,N_13685,N_11079);
or UO_213 (O_213,N_14324,N_12654);
nor UO_214 (O_214,N_12438,N_12873);
nor UO_215 (O_215,N_14140,N_11021);
nor UO_216 (O_216,N_12304,N_12071);
nor UO_217 (O_217,N_14616,N_14742);
nor UO_218 (O_218,N_10462,N_10434);
nor UO_219 (O_219,N_12234,N_13777);
xor UO_220 (O_220,N_10447,N_11326);
nand UO_221 (O_221,N_11830,N_11914);
nor UO_222 (O_222,N_13659,N_11441);
nand UO_223 (O_223,N_14872,N_13570);
or UO_224 (O_224,N_10152,N_13616);
or UO_225 (O_225,N_14928,N_13066);
xor UO_226 (O_226,N_13208,N_11233);
nand UO_227 (O_227,N_10690,N_10385);
or UO_228 (O_228,N_14705,N_12498);
xnor UO_229 (O_229,N_10989,N_12080);
or UO_230 (O_230,N_11466,N_12523);
xnor UO_231 (O_231,N_11774,N_14995);
and UO_232 (O_232,N_12445,N_10778);
nor UO_233 (O_233,N_14383,N_14089);
nor UO_234 (O_234,N_14731,N_14138);
nor UO_235 (O_235,N_10938,N_14385);
and UO_236 (O_236,N_13125,N_10819);
xnor UO_237 (O_237,N_11265,N_10242);
and UO_238 (O_238,N_14250,N_12842);
or UO_239 (O_239,N_11925,N_14232);
and UO_240 (O_240,N_13765,N_12762);
xnor UO_241 (O_241,N_13666,N_11291);
xor UO_242 (O_242,N_12874,N_13582);
or UO_243 (O_243,N_11257,N_10743);
nor UO_244 (O_244,N_11841,N_12580);
or UO_245 (O_245,N_14264,N_13113);
or UO_246 (O_246,N_10556,N_10536);
nor UO_247 (O_247,N_12256,N_14212);
nor UO_248 (O_248,N_10799,N_10643);
and UO_249 (O_249,N_12454,N_10064);
or UO_250 (O_250,N_11917,N_10437);
or UO_251 (O_251,N_12225,N_12741);
and UO_252 (O_252,N_11105,N_10512);
and UO_253 (O_253,N_11311,N_13343);
or UO_254 (O_254,N_11309,N_14201);
nand UO_255 (O_255,N_10711,N_12330);
nor UO_256 (O_256,N_12728,N_11847);
and UO_257 (O_257,N_10355,N_10083);
or UO_258 (O_258,N_12368,N_13583);
nor UO_259 (O_259,N_12824,N_12346);
or UO_260 (O_260,N_11708,N_12956);
or UO_261 (O_261,N_12572,N_14857);
nand UO_262 (O_262,N_12505,N_14096);
and UO_263 (O_263,N_13865,N_11488);
nand UO_264 (O_264,N_14165,N_11806);
or UO_265 (O_265,N_14887,N_10286);
nand UO_266 (O_266,N_11955,N_11031);
xnor UO_267 (O_267,N_11264,N_12174);
xnor UO_268 (O_268,N_10855,N_12193);
and UO_269 (O_269,N_14660,N_13549);
and UO_270 (O_270,N_13919,N_10436);
nor UO_271 (O_271,N_10344,N_14378);
xor UO_272 (O_272,N_10189,N_10543);
and UO_273 (O_273,N_10205,N_11725);
nand UO_274 (O_274,N_13417,N_13716);
nor UO_275 (O_275,N_12002,N_11646);
or UO_276 (O_276,N_12846,N_12806);
or UO_277 (O_277,N_13504,N_10208);
nand UO_278 (O_278,N_10433,N_13339);
xnor UO_279 (O_279,N_14147,N_12209);
nand UO_280 (O_280,N_12273,N_12831);
nor UO_281 (O_281,N_11308,N_12906);
or UO_282 (O_282,N_12133,N_13021);
xor UO_283 (O_283,N_13667,N_12784);
xnor UO_284 (O_284,N_12007,N_10314);
or UO_285 (O_285,N_13751,N_11621);
or UO_286 (O_286,N_10315,N_14794);
xor UO_287 (O_287,N_10768,N_12959);
nor UO_288 (O_288,N_11502,N_13376);
xnor UO_289 (O_289,N_13056,N_13079);
nand UO_290 (O_290,N_13473,N_10176);
xnor UO_291 (O_291,N_13319,N_11164);
nand UO_292 (O_292,N_10560,N_14507);
and UO_293 (O_293,N_10857,N_11426);
xor UO_294 (O_294,N_13469,N_13799);
nor UO_295 (O_295,N_12251,N_10851);
nor UO_296 (O_296,N_12504,N_10617);
nand UO_297 (O_297,N_11720,N_13185);
and UO_298 (O_298,N_12283,N_13225);
xor UO_299 (O_299,N_14869,N_10666);
nor UO_300 (O_300,N_13392,N_11697);
or UO_301 (O_301,N_14361,N_14127);
xor UO_302 (O_302,N_12984,N_14667);
xor UO_303 (O_303,N_13389,N_10874);
and UO_304 (O_304,N_11295,N_11331);
nor UO_305 (O_305,N_11273,N_12849);
xor UO_306 (O_306,N_12474,N_10856);
or UO_307 (O_307,N_14514,N_11396);
nand UO_308 (O_308,N_14784,N_13929);
nand UO_309 (O_309,N_10257,N_12268);
and UO_310 (O_310,N_14327,N_11912);
nor UO_311 (O_311,N_11959,N_14653);
and UO_312 (O_312,N_11298,N_12396);
or UO_313 (O_313,N_14290,N_10339);
or UO_314 (O_314,N_14797,N_11777);
and UO_315 (O_315,N_11012,N_14879);
nand UO_316 (O_316,N_12099,N_12708);
and UO_317 (O_317,N_11963,N_13160);
and UO_318 (O_318,N_10839,N_14190);
and UO_319 (O_319,N_13318,N_12663);
or UO_320 (O_320,N_10243,N_13797);
and UO_321 (O_321,N_10861,N_13394);
nor UO_322 (O_322,N_12941,N_11988);
or UO_323 (O_323,N_11605,N_11927);
xor UO_324 (O_324,N_10862,N_11457);
xor UO_325 (O_325,N_11700,N_10489);
or UO_326 (O_326,N_10721,N_11373);
or UO_327 (O_327,N_11472,N_13420);
xor UO_328 (O_328,N_10641,N_13128);
xnor UO_329 (O_329,N_11679,N_11729);
nor UO_330 (O_330,N_12781,N_13801);
nor UO_331 (O_331,N_11736,N_13934);
and UO_332 (O_332,N_14213,N_13030);
and UO_333 (O_333,N_13434,N_13527);
nor UO_334 (O_334,N_10416,N_14374);
xnor UO_335 (O_335,N_12292,N_11816);
xor UO_336 (O_336,N_13708,N_10323);
nand UO_337 (O_337,N_14100,N_11599);
or UO_338 (O_338,N_13566,N_13706);
or UO_339 (O_339,N_12684,N_14905);
nand UO_340 (O_340,N_10514,N_12465);
nand UO_341 (O_341,N_11099,N_13928);
nand UO_342 (O_342,N_13140,N_12834);
and UO_343 (O_343,N_14384,N_10598);
and UO_344 (O_344,N_13176,N_14651);
nor UO_345 (O_345,N_13631,N_10853);
or UO_346 (O_346,N_14395,N_13671);
nand UO_347 (O_347,N_13579,N_12429);
and UO_348 (O_348,N_10241,N_11358);
nor UO_349 (O_349,N_14647,N_10740);
nor UO_350 (O_350,N_10747,N_13575);
xnor UO_351 (O_351,N_14406,N_10378);
xnor UO_352 (O_352,N_13896,N_10899);
xor UO_353 (O_353,N_13004,N_11589);
nand UO_354 (O_354,N_14575,N_11886);
or UO_355 (O_355,N_13107,N_11761);
or UO_356 (O_356,N_14693,N_11825);
and UO_357 (O_357,N_10133,N_10066);
nand UO_358 (O_358,N_14081,N_11212);
and UO_359 (O_359,N_12001,N_12607);
or UO_360 (O_360,N_14319,N_10594);
xor UO_361 (O_361,N_14227,N_14391);
and UO_362 (O_362,N_11652,N_12323);
nor UO_363 (O_363,N_14292,N_14897);
nand UO_364 (O_364,N_12709,N_12690);
nor UO_365 (O_365,N_13205,N_12086);
and UO_366 (O_366,N_13036,N_13796);
xnor UO_367 (O_367,N_10933,N_12507);
xnor UO_368 (O_368,N_11790,N_13657);
or UO_369 (O_369,N_10354,N_10476);
nand UO_370 (O_370,N_14988,N_10233);
nand UO_371 (O_371,N_10614,N_12020);
and UO_372 (O_372,N_12468,N_13687);
xor UO_373 (O_373,N_12073,N_11889);
xor UO_374 (O_374,N_10439,N_13951);
nor UO_375 (O_375,N_12931,N_14275);
or UO_376 (O_376,N_13353,N_13083);
or UO_377 (O_377,N_10455,N_11518);
nand UO_378 (O_378,N_11829,N_10231);
nor UO_379 (O_379,N_14826,N_12188);
nor UO_380 (O_380,N_12508,N_13977);
or UO_381 (O_381,N_12845,N_12372);
nand UO_382 (O_382,N_13869,N_10624);
nor UO_383 (O_383,N_14883,N_10332);
xnor UO_384 (O_384,N_13304,N_10026);
or UO_385 (O_385,N_11572,N_11684);
and UO_386 (O_386,N_10113,N_13755);
nand UO_387 (O_387,N_12672,N_14855);
or UO_388 (O_388,N_12434,N_10601);
nand UO_389 (O_389,N_10492,N_11905);
nand UO_390 (O_390,N_10595,N_12312);
nor UO_391 (O_391,N_12308,N_12156);
or UO_392 (O_392,N_14448,N_14811);
or UO_393 (O_393,N_13640,N_13171);
xnor UO_394 (O_394,N_10118,N_13110);
xor UO_395 (O_395,N_10256,N_12294);
xnor UO_396 (O_396,N_14832,N_14952);
nand UO_397 (O_397,N_13308,N_12929);
nand UO_398 (O_398,N_11217,N_11427);
xor UO_399 (O_399,N_10665,N_12643);
xor UO_400 (O_400,N_12550,N_14973);
xor UO_401 (O_401,N_11199,N_13581);
and UO_402 (O_402,N_12926,N_13320);
and UO_403 (O_403,N_14457,N_13446);
or UO_404 (O_404,N_10764,N_10932);
and UO_405 (O_405,N_11982,N_10824);
nand UO_406 (O_406,N_13739,N_11376);
nand UO_407 (O_407,N_14529,N_13399);
or UO_408 (O_408,N_14913,N_11296);
or UO_409 (O_409,N_10902,N_10074);
and UO_410 (O_410,N_13555,N_12334);
xnor UO_411 (O_411,N_13258,N_10268);
xnor UO_412 (O_412,N_10279,N_14544);
or UO_413 (O_413,N_13771,N_13493);
nand UO_414 (O_414,N_11208,N_11686);
and UO_415 (O_415,N_14204,N_10426);
nand UO_416 (O_416,N_11906,N_13266);
xnor UO_417 (O_417,N_10088,N_12676);
and UO_418 (O_418,N_13760,N_13988);
nor UO_419 (O_419,N_11741,N_10458);
xnor UO_420 (O_420,N_14701,N_11878);
nand UO_421 (O_421,N_13508,N_14191);
xnor UO_422 (O_422,N_13040,N_12940);
xnor UO_423 (O_423,N_11035,N_14652);
and UO_424 (O_424,N_10502,N_14158);
nor UO_425 (O_425,N_11013,N_12836);
or UO_426 (O_426,N_11595,N_14067);
nand UO_427 (O_427,N_12245,N_10469);
and UO_428 (O_428,N_12287,N_12366);
xnor UO_429 (O_429,N_10767,N_12881);
and UO_430 (O_430,N_12094,N_11585);
nand UO_431 (O_431,N_14802,N_13959);
or UO_432 (O_432,N_10124,N_12964);
nor UO_433 (O_433,N_10410,N_10169);
and UO_434 (O_434,N_13778,N_11633);
nand UO_435 (O_435,N_12339,N_11342);
xnor UO_436 (O_436,N_10986,N_11718);
or UO_437 (O_437,N_11092,N_14237);
nor UO_438 (O_438,N_14901,N_12190);
nand UO_439 (O_439,N_10662,N_10816);
or UO_440 (O_440,N_11915,N_14442);
or UO_441 (O_441,N_11060,N_10225);
nand UO_442 (O_442,N_10686,N_12267);
nand UO_443 (O_443,N_13121,N_12093);
nor UO_444 (O_444,N_12785,N_11961);
xor UO_445 (O_445,N_10255,N_11397);
or UO_446 (O_446,N_11689,N_11857);
xnor UO_447 (O_447,N_13122,N_11424);
and UO_448 (O_448,N_13271,N_12860);
xnor UO_449 (O_449,N_14444,N_13976);
xnor UO_450 (O_450,N_13761,N_13857);
xnor UO_451 (O_451,N_12973,N_13673);
nand UO_452 (O_452,N_10604,N_13567);
nand UO_453 (O_453,N_13448,N_13249);
nor UO_454 (O_454,N_12618,N_10081);
xor UO_455 (O_455,N_14418,N_10251);
nor UO_456 (O_456,N_12577,N_10043);
xor UO_457 (O_457,N_12571,N_13780);
nand UO_458 (O_458,N_12921,N_14942);
nor UO_459 (O_459,N_10377,N_14931);
or UO_460 (O_460,N_12564,N_10277);
and UO_461 (O_461,N_13522,N_13554);
nand UO_462 (O_462,N_14139,N_10559);
nand UO_463 (O_463,N_10600,N_13404);
or UO_464 (O_464,N_12172,N_14740);
nor UO_465 (O_465,N_14281,N_10836);
xor UO_466 (O_466,N_11270,N_12866);
nor UO_467 (O_467,N_10049,N_12309);
and UO_468 (O_468,N_14485,N_10947);
xor UO_469 (O_469,N_12631,N_12970);
xnor UO_470 (O_470,N_10090,N_11797);
xnor UO_471 (O_471,N_10186,N_11903);
xnor UO_472 (O_472,N_13525,N_11144);
and UO_473 (O_473,N_14640,N_13495);
or UO_474 (O_474,N_11696,N_10712);
nand UO_475 (O_475,N_10347,N_12586);
nor UO_476 (O_476,N_12844,N_14052);
nor UO_477 (O_477,N_12295,N_11484);
and UO_478 (O_478,N_12306,N_13585);
nor UO_479 (O_479,N_10901,N_11362);
or UO_480 (O_480,N_11462,N_12742);
nor UO_481 (O_481,N_10448,N_10878);
and UO_482 (O_482,N_13984,N_14581);
or UO_483 (O_483,N_11068,N_13351);
xor UO_484 (O_484,N_13773,N_11429);
xor UO_485 (O_485,N_13732,N_12021);
and UO_486 (O_486,N_14925,N_11737);
nor UO_487 (O_487,N_13155,N_10503);
or UO_488 (O_488,N_14160,N_12296);
nand UO_489 (O_489,N_10002,N_11789);
xnor UO_490 (O_490,N_12935,N_10346);
and UO_491 (O_491,N_11128,N_11478);
and UO_492 (O_492,N_14523,N_11182);
and UO_493 (O_493,N_10528,N_11918);
or UO_494 (O_494,N_14548,N_10449);
xnor UO_495 (O_495,N_13693,N_11503);
or UO_496 (O_496,N_10779,N_12271);
xor UO_497 (O_497,N_13428,N_11984);
or UO_498 (O_498,N_14328,N_14129);
nor UO_499 (O_499,N_14856,N_10917);
or UO_500 (O_500,N_13297,N_12318);
nand UO_501 (O_501,N_11486,N_14600);
nor UO_502 (O_502,N_12488,N_13476);
nand UO_503 (O_503,N_10524,N_10285);
and UO_504 (O_504,N_10540,N_13507);
xnor UO_505 (O_505,N_13106,N_11660);
or UO_506 (O_506,N_11683,N_14592);
or UO_507 (O_507,N_12096,N_11330);
or UO_508 (O_508,N_11453,N_14430);
nor UO_509 (O_509,N_12297,N_14720);
and UO_510 (O_510,N_10655,N_10405);
xor UO_511 (O_511,N_10894,N_12992);
nor UO_512 (O_512,N_13099,N_11335);
and UO_513 (O_513,N_11442,N_13430);
or UO_514 (O_514,N_11623,N_14716);
nor UO_515 (O_515,N_10960,N_13994);
or UO_516 (O_516,N_12408,N_14666);
nor UO_517 (O_517,N_11615,N_10589);
nor UO_518 (O_518,N_11106,N_14261);
or UO_519 (O_519,N_14612,N_11287);
nor UO_520 (O_520,N_14689,N_11944);
nand UO_521 (O_521,N_14211,N_14637);
and UO_522 (O_522,N_12032,N_14659);
nand UO_523 (O_523,N_13049,N_10833);
nand UO_524 (O_524,N_10261,N_14224);
xnor UO_525 (O_525,N_11166,N_12835);
or UO_526 (O_526,N_12619,N_11379);
nor UO_527 (O_527,N_10499,N_13387);
and UO_528 (O_528,N_13287,N_13444);
nor UO_529 (O_529,N_12958,N_11874);
nand UO_530 (O_530,N_12658,N_14379);
and UO_531 (O_531,N_11549,N_11559);
nand UO_532 (O_532,N_11962,N_12919);
nand UO_533 (O_533,N_10105,N_10511);
or UO_534 (O_534,N_13301,N_11692);
or UO_535 (O_535,N_12937,N_12026);
and UO_536 (O_536,N_14589,N_11413);
and UO_537 (O_537,N_11746,N_10422);
nand UO_538 (O_538,N_12972,N_10333);
nor UO_539 (O_539,N_10207,N_12905);
and UO_540 (O_540,N_10659,N_12591);
nand UO_541 (O_541,N_10693,N_12351);
nor UO_542 (O_542,N_13913,N_13441);
nand UO_543 (O_543,N_11266,N_10995);
nand UO_544 (O_544,N_12207,N_12424);
nand UO_545 (O_545,N_11483,N_10754);
nor UO_546 (O_546,N_13250,N_10039);
nand UO_547 (O_547,N_14917,N_10209);
nor UO_548 (O_548,N_14607,N_10897);
xor UO_549 (O_549,N_14508,N_10991);
xnor UO_550 (O_550,N_10263,N_10457);
nand UO_551 (O_551,N_12679,N_12893);
nor UO_552 (O_552,N_14696,N_13449);
nor UO_553 (O_553,N_11445,N_11821);
and UO_554 (O_554,N_13597,N_13904);
and UO_555 (O_555,N_12702,N_12269);
and UO_556 (O_556,N_14515,N_13602);
nand UO_557 (O_557,N_11455,N_13625);
nor UO_558 (O_558,N_11583,N_12119);
nand UO_559 (O_559,N_11801,N_13280);
nand UO_560 (O_560,N_12971,N_10014);
xnor UO_561 (O_561,N_12943,N_11688);
or UO_562 (O_562,N_12622,N_12496);
and UO_563 (O_563,N_11117,N_11016);
and UO_564 (O_564,N_13480,N_12531);
nand UO_565 (O_565,N_13550,N_12208);
xnor UO_566 (O_566,N_13413,N_12122);
nand UO_567 (O_567,N_12756,N_10657);
and UO_568 (O_568,N_12652,N_13491);
xnor UO_569 (O_569,N_14584,N_13414);
and UO_570 (O_570,N_12442,N_10599);
nor UO_571 (O_571,N_10046,N_11942);
nor UO_572 (O_572,N_12173,N_12803);
xnor UO_573 (O_573,N_12395,N_12333);
nand UO_574 (O_574,N_14195,N_12854);
or UO_575 (O_575,N_12410,N_11070);
and UO_576 (O_576,N_14977,N_11389);
nand UO_577 (O_577,N_12361,N_12981);
xnor UO_578 (O_578,N_11228,N_13375);
nor UO_579 (O_579,N_11074,N_11193);
nand UO_580 (O_580,N_12534,N_13829);
and UO_581 (O_581,N_13870,N_12891);
xor UO_582 (O_582,N_12440,N_13199);
and UO_583 (O_583,N_12750,N_13047);
or UO_584 (O_584,N_11404,N_11714);
or UO_585 (O_585,N_11854,N_12775);
nor UO_586 (O_586,N_14362,N_11476);
or UO_587 (O_587,N_10041,N_12832);
and UO_588 (O_588,N_13759,N_11227);
xnor UO_589 (O_589,N_13993,N_12484);
and UO_590 (O_590,N_12298,N_10926);
nor UO_591 (O_591,N_14178,N_11246);
or UO_592 (O_592,N_12584,N_11170);
nor UO_593 (O_593,N_11856,N_11065);
or UO_594 (O_594,N_14538,N_13405);
nor UO_595 (O_595,N_10267,N_11511);
or UO_596 (O_596,N_10296,N_13653);
xnor UO_597 (O_597,N_13034,N_13005);
or UO_598 (O_598,N_10485,N_14326);
and UO_599 (O_599,N_10681,N_12678);
and UO_600 (O_600,N_14363,N_10783);
nand UO_601 (O_601,N_12597,N_11994);
and UO_602 (O_602,N_14321,N_11738);
nor UO_603 (O_603,N_12557,N_12210);
and UO_604 (O_604,N_14907,N_14512);
nand UO_605 (O_605,N_13029,N_10220);
or UO_606 (O_606,N_13006,N_12732);
xnor UO_607 (O_607,N_11400,N_11709);
nor UO_608 (O_608,N_12220,N_13807);
or UO_609 (O_609,N_14408,N_10224);
and UO_610 (O_610,N_14183,N_11140);
or UO_611 (O_611,N_12079,N_14884);
or UO_612 (O_612,N_11072,N_14805);
and UO_613 (O_613,N_14574,N_12403);
and UO_614 (O_614,N_11051,N_10825);
and UO_615 (O_615,N_11431,N_12384);
nand UO_616 (O_616,N_12614,N_13483);
xnor UO_617 (O_617,N_13720,N_11173);
nor UO_618 (O_618,N_12514,N_13812);
and UO_619 (O_619,N_12851,N_11802);
nand UO_620 (O_620,N_14425,N_14017);
or UO_621 (O_621,N_12281,N_12978);
and UO_622 (O_622,N_10359,N_14381);
xor UO_623 (O_623,N_10919,N_12491);
nand UO_624 (O_624,N_14170,N_13860);
and UO_625 (O_625,N_14565,N_13333);
and UO_626 (O_626,N_10924,N_14606);
and UO_627 (O_627,N_13770,N_13241);
and UO_628 (O_628,N_14573,N_13274);
or UO_629 (O_629,N_10179,N_14028);
nor UO_630 (O_630,N_12650,N_11220);
nand UO_631 (O_631,N_10885,N_10629);
nand UO_632 (O_632,N_10806,N_13835);
and UO_633 (O_633,N_11527,N_12149);
xnor UO_634 (O_634,N_12112,N_14344);
xnor UO_635 (O_635,N_12212,N_12138);
or UO_636 (O_636,N_11627,N_12880);
nand UO_637 (O_637,N_10274,N_13337);
nand UO_638 (O_638,N_10953,N_13725);
nand UO_639 (O_639,N_10639,N_14434);
xor UO_640 (O_640,N_10342,N_14179);
nor UO_641 (O_641,N_11577,N_10203);
nor UO_642 (O_642,N_14866,N_13377);
nand UO_643 (O_643,N_12413,N_12033);
nor UO_644 (O_644,N_13850,N_13146);
and UO_645 (O_645,N_12057,N_12483);
xnor UO_646 (O_646,N_14777,N_12913);
xnor UO_647 (O_647,N_10784,N_12321);
nand UO_648 (O_648,N_12261,N_13805);
or UO_649 (O_649,N_14131,N_12065);
nor UO_650 (O_650,N_14282,N_12387);
xnor UO_651 (O_651,N_13661,N_13498);
nand UO_652 (O_652,N_10076,N_11262);
xnor UO_653 (O_653,N_14143,N_11949);
and UO_654 (O_654,N_11710,N_13163);
nand UO_655 (O_655,N_11807,N_14587);
nand UO_656 (O_656,N_12977,N_13932);
nor UO_657 (O_657,N_12160,N_10774);
and UO_658 (O_658,N_11109,N_13785);
nand UO_659 (O_659,N_13683,N_11313);
and UO_660 (O_660,N_14024,N_10196);
xnor UO_661 (O_661,N_14994,N_12812);
and UO_662 (O_662,N_14598,N_13939);
nand UO_663 (O_663,N_14608,N_11165);
xnor UO_664 (O_664,N_11657,N_11575);
nor UO_665 (O_665,N_11919,N_14750);
and UO_666 (O_666,N_13822,N_10401);
nand UO_667 (O_667,N_10916,N_11867);
or UO_668 (O_668,N_14825,N_13123);
xnor UO_669 (O_669,N_12512,N_12329);
nor UO_670 (O_670,N_12538,N_14339);
xnor UO_671 (O_671,N_14423,N_10802);
nand UO_672 (O_672,N_11586,N_11473);
and UO_673 (O_673,N_12217,N_11048);
xor UO_674 (O_674,N_13943,N_14697);
nor UO_675 (O_675,N_13911,N_10755);
nand UO_676 (O_676,N_14631,N_14710);
and UO_677 (O_677,N_14516,N_11606);
nor UO_678 (O_678,N_10345,N_13331);
nand UO_679 (O_679,N_10312,N_10510);
and UO_680 (O_680,N_11659,N_14435);
nor UO_681 (O_681,N_14506,N_10412);
and UO_682 (O_682,N_13753,N_14460);
nand UO_683 (O_683,N_11382,N_13591);
or UO_684 (O_684,N_14012,N_12660);
and UO_685 (O_685,N_13334,N_14120);
and UO_686 (O_686,N_14661,N_10365);
and UO_687 (O_687,N_12249,N_10442);
xor UO_688 (O_688,N_14727,N_10098);
nor UO_689 (O_689,N_12415,N_14177);
or UO_690 (O_690,N_11177,N_11464);
xnor UO_691 (O_691,N_13855,N_10998);
nor UO_692 (O_692,N_13306,N_14671);
nor UO_693 (O_693,N_11493,N_12667);
xor UO_694 (O_694,N_10148,N_13116);
or UO_695 (O_695,N_14534,N_11045);
nand UO_696 (O_696,N_12282,N_13455);
and UO_697 (O_697,N_14472,N_11809);
nor UO_698 (O_698,N_14632,N_14056);
nor UO_699 (O_699,N_12238,N_12983);
nand UO_700 (O_700,N_10077,N_10319);
or UO_701 (O_701,N_11184,N_14828);
or UO_702 (O_702,N_10282,N_10987);
and UO_703 (O_703,N_12171,N_13881);
or UO_704 (O_704,N_10759,N_13813);
xnor UO_705 (O_705,N_12359,N_12725);
or UO_706 (O_706,N_11661,N_12303);
xor UO_707 (O_707,N_12179,N_13696);
and UO_708 (O_708,N_11791,N_12452);
or UO_709 (O_709,N_11334,N_12003);
or UO_710 (O_710,N_13262,N_12882);
or UO_711 (O_711,N_14715,N_13009);
or UO_712 (O_712,N_10929,N_12863);
nor UO_713 (O_713,N_13057,N_13639);
nand UO_714 (O_714,N_11805,N_12604);
or UO_715 (O_715,N_13310,N_10718);
nor UO_716 (O_716,N_11634,N_12229);
nor UO_717 (O_717,N_14914,N_14711);
nor UO_718 (O_718,N_11869,N_14517);
xnor UO_719 (O_719,N_11800,N_12839);
nand UO_720 (O_720,N_12888,N_10505);
or UO_721 (O_721,N_11747,N_14034);
and UO_722 (O_722,N_13431,N_12034);
nor UO_723 (O_723,N_12894,N_12219);
and UO_724 (O_724,N_13593,N_12807);
and UO_725 (O_725,N_12945,N_11926);
and UO_726 (O_726,N_11353,N_14466);
and UO_727 (O_727,N_11190,N_11813);
xor UO_728 (O_728,N_13384,N_10920);
and UO_729 (O_729,N_13344,N_12134);
nor UO_730 (O_730,N_14122,N_13622);
and UO_731 (O_731,N_14604,N_10873);
xor UO_732 (O_732,N_13823,N_14289);
and UO_733 (O_733,N_11271,N_10621);
or UO_734 (O_734,N_11171,N_10238);
nand UO_735 (O_735,N_13152,N_10165);
and UO_736 (O_736,N_11254,N_12521);
nand UO_737 (O_737,N_10992,N_12470);
or UO_738 (O_738,N_12284,N_12516);
nor UO_739 (O_739,N_11244,N_10730);
or UO_740 (O_740,N_14533,N_14555);
or UO_741 (O_741,N_14624,N_14005);
nand UO_742 (O_742,N_10637,N_14022);
or UO_743 (O_743,N_10567,N_10544);
or UO_744 (O_744,N_10970,N_10038);
nand UO_745 (O_745,N_10881,N_10357);
or UO_746 (O_746,N_10968,N_12291);
xor UO_747 (O_747,N_14104,N_10495);
and UO_748 (O_748,N_10999,N_12852);
or UO_749 (O_749,N_11209,N_13349);
and UO_750 (O_750,N_12482,N_12635);
xnor UO_751 (O_751,N_13336,N_13917);
and UO_752 (O_752,N_12879,N_13628);
and UO_753 (O_753,N_14733,N_10394);
or UO_754 (O_754,N_12867,N_12432);
and UO_755 (O_755,N_13427,N_13681);
nand UO_756 (O_756,N_14657,N_12443);
xnor UO_757 (O_757,N_10099,N_11649);
nor UO_758 (O_758,N_12562,N_10635);
and UO_759 (O_759,N_13302,N_10752);
and UO_760 (O_760,N_10111,N_14915);
nor UO_761 (O_761,N_13370,N_14735);
nor UO_762 (O_762,N_13435,N_11232);
or UO_763 (O_763,N_10018,N_10150);
nor UO_764 (O_764,N_10468,N_14405);
nor UO_765 (O_765,N_13292,N_13073);
nand UO_766 (O_766,N_11179,N_13573);
or UO_767 (O_767,N_11990,N_14683);
nand UO_768 (O_768,N_13665,N_13873);
xnor UO_769 (O_769,N_14130,N_13179);
or UO_770 (O_770,N_10121,N_14550);
nor UO_771 (O_771,N_10299,N_10780);
nand UO_772 (O_772,N_11341,N_14817);
and UO_773 (O_773,N_12989,N_10302);
nor UO_774 (O_774,N_14042,N_10823);
or UO_775 (O_775,N_14257,N_12045);
nand UO_776 (O_776,N_11428,N_13425);
xor UO_777 (O_777,N_12783,N_10529);
nor UO_778 (O_778,N_13261,N_14782);
nor UO_779 (O_779,N_13101,N_10284);
nand UO_780 (O_780,N_13089,N_14103);
nor UO_781 (O_781,N_10407,N_14044);
or UO_782 (O_782,N_12078,N_13966);
xor UO_783 (O_783,N_13015,N_10736);
xor UO_784 (O_784,N_12227,N_12567);
or UO_785 (O_785,N_14882,N_13011);
or UO_786 (O_786,N_12319,N_12936);
or UO_787 (O_787,N_11881,N_11052);
or UO_788 (O_788,N_10444,N_11514);
nor UO_789 (O_789,N_10837,N_11767);
xnor UO_790 (O_790,N_13969,N_11669);
and UO_791 (O_791,N_14675,N_13027);
xor UO_792 (O_792,N_11302,N_13551);
xnor UO_793 (O_793,N_11862,N_14590);
xor UO_794 (O_794,N_11345,N_14965);
and UO_795 (O_795,N_13561,N_14043);
xnor UO_796 (O_796,N_13195,N_13008);
xnor UO_797 (O_797,N_10147,N_12602);
xnor UO_798 (O_798,N_14233,N_10673);
and UO_799 (O_799,N_11758,N_11643);
or UO_800 (O_800,N_11443,N_10218);
nor UO_801 (O_801,N_13833,N_13051);
nor UO_802 (O_802,N_14424,N_12814);
or UO_803 (O_803,N_12640,N_10497);
nor UO_804 (O_804,N_12383,N_13906);
xor UO_805 (O_805,N_12611,N_10934);
nand UO_806 (O_806,N_11195,N_13180);
xnor UO_807 (O_807,N_12734,N_13590);
or UO_808 (O_808,N_14572,N_10979);
and UO_809 (O_809,N_13898,N_10520);
xor UO_810 (O_810,N_12800,N_12206);
nor UO_811 (O_811,N_13875,N_11826);
nor UO_812 (O_812,N_14745,N_13768);
nor UO_813 (O_813,N_11019,N_11896);
nand UO_814 (O_814,N_10138,N_13492);
nand UO_815 (O_815,N_12698,N_13861);
nor UO_816 (O_816,N_14989,N_10652);
nor UO_817 (O_817,N_12561,N_13960);
xor UO_818 (O_818,N_10791,N_13868);
nand UO_819 (O_819,N_12923,N_11059);
nand UO_820 (O_820,N_11937,N_11936);
nand UO_821 (O_821,N_12588,N_10091);
nand UO_822 (O_822,N_10977,N_13157);
and UO_823 (O_823,N_14345,N_13406);
or UO_824 (O_824,N_12402,N_14990);
or UO_825 (O_825,N_12605,N_10212);
and UO_826 (O_826,N_12975,N_14433);
nand UO_827 (O_827,N_10723,N_10230);
or UO_828 (O_828,N_13830,N_11971);
and UO_829 (O_829,N_12075,N_10796);
and UO_830 (O_830,N_11768,N_10847);
nor UO_831 (O_831,N_13002,N_10496);
nor UO_832 (O_832,N_12405,N_14670);
nand UO_833 (O_833,N_10648,N_13364);
xnor UO_834 (O_834,N_14724,N_11260);
nor UO_835 (O_835,N_12641,N_14192);
xor UO_836 (O_836,N_12090,N_14862);
nand UO_837 (O_837,N_10921,N_14541);
or UO_838 (O_838,N_10131,N_13202);
xnor UO_839 (O_839,N_10997,N_11977);
xor UO_840 (O_840,N_10705,N_10928);
nor UO_841 (O_841,N_13126,N_14956);
nor UO_842 (O_842,N_10308,N_14526);
nand UO_843 (O_843,N_14074,N_14700);
xnor UO_844 (O_844,N_12363,N_11319);
and UO_845 (O_845,N_13885,N_13041);
nor UO_846 (O_846,N_11524,N_14375);
xor UO_847 (O_847,N_13281,N_12453);
or UO_848 (O_848,N_12124,N_11943);
and UO_849 (O_849,N_12960,N_12996);
nand UO_850 (O_850,N_12645,N_10057);
xor UO_851 (O_851,N_14203,N_10055);
nand UO_852 (O_852,N_11406,N_12671);
xor UO_853 (O_853,N_14524,N_14059);
or UO_854 (O_854,N_11561,N_14908);
nor UO_855 (O_855,N_14930,N_14248);
and UO_856 (O_856,N_11148,N_13747);
xor UO_857 (O_857,N_14730,N_13745);
xor UO_858 (O_858,N_14315,N_12951);
nor UO_859 (O_859,N_11224,N_10036);
nor UO_860 (O_860,N_13980,N_14528);
xor UO_861 (O_861,N_11213,N_14940);
or UO_862 (O_862,N_14149,N_12299);
nand UO_863 (O_863,N_14767,N_11913);
xor UO_864 (O_864,N_13788,N_11808);
nand UO_865 (O_865,N_12129,N_10773);
or UO_866 (O_866,N_10808,N_13145);
and UO_867 (O_867,N_12928,N_12144);
or UO_868 (O_868,N_11003,N_13750);
and UO_869 (O_869,N_10785,N_12419);
nor UO_870 (O_870,N_14920,N_13743);
xor UO_871 (O_871,N_13265,N_13188);
nor UO_872 (O_872,N_10262,N_12162);
nor UO_873 (O_873,N_14283,N_12182);
or UO_874 (O_874,N_13997,N_11965);
nor UO_875 (O_875,N_11374,N_11573);
or UO_876 (O_876,N_14539,N_11207);
nor UO_877 (O_877,N_13731,N_12260);
xor UO_878 (O_878,N_11203,N_14176);
xnor UO_879 (O_879,N_14049,N_10908);
nor UO_880 (O_880,N_13286,N_14747);
xor UO_881 (O_881,N_13704,N_11934);
nor UO_882 (O_882,N_10893,N_14957);
nand UO_883 (O_883,N_11694,N_12720);
nor UO_884 (O_884,N_11900,N_11238);
or UO_885 (O_885,N_13046,N_10763);
nand UO_886 (O_886,N_14809,N_11978);
and UO_887 (O_887,N_12695,N_13903);
xor UO_888 (O_888,N_10311,N_10223);
xor UO_889 (O_889,N_11836,N_14360);
or UO_890 (O_890,N_12993,N_11508);
xor UO_891 (O_891,N_13902,N_10406);
nor UO_892 (O_892,N_12322,N_13397);
xnor UO_893 (O_893,N_13936,N_11756);
xor UO_894 (O_894,N_14205,N_10638);
xor UO_895 (O_895,N_11546,N_14634);
nand UO_896 (O_896,N_10840,N_10821);
and UO_897 (O_897,N_14329,N_13806);
and UO_898 (O_898,N_10826,N_13894);
and UO_899 (O_899,N_12216,N_10777);
nand UO_900 (O_900,N_10031,N_13978);
nor UO_901 (O_901,N_12651,N_14934);
and UO_902 (O_902,N_13248,N_14501);
or UO_903 (O_903,N_11088,N_11763);
or UO_904 (O_904,N_10573,N_12106);
or UO_905 (O_905,N_11432,N_14836);
or UO_906 (O_906,N_13093,N_12656);
and UO_907 (O_907,N_13986,N_11492);
and UO_908 (O_908,N_10163,N_14235);
and UO_909 (O_909,N_10050,N_10167);
nand UO_910 (O_910,N_13466,N_10035);
and UO_911 (O_911,N_12091,N_13316);
nor UO_912 (O_912,N_11294,N_13727);
nand UO_913 (O_913,N_12084,N_11975);
nand UO_914 (O_914,N_12004,N_12884);
nand UO_915 (O_915,N_10860,N_14753);
xnor UO_916 (O_916,N_13595,N_10431);
nand UO_917 (O_917,N_11064,N_11998);
xor UO_918 (O_918,N_13096,N_11027);
nand UO_919 (O_919,N_13558,N_14868);
or UO_920 (O_920,N_11760,N_11286);
xor UO_921 (O_921,N_14803,N_14085);
and UO_922 (O_922,N_12527,N_11258);
or UO_923 (O_923,N_10338,N_10488);
nor UO_924 (O_924,N_11292,N_11654);
or UO_925 (O_925,N_14629,N_10575);
xnor UO_926 (O_926,N_10466,N_10606);
xnor UO_927 (O_927,N_10197,N_11121);
and UO_928 (O_928,N_14046,N_10024);
nor UO_929 (O_929,N_12204,N_11976);
nor UO_930 (O_930,N_11054,N_11845);
and UO_931 (O_931,N_13819,N_13721);
or UO_932 (O_932,N_12345,N_12105);
nand UO_933 (O_933,N_11844,N_10832);
or UO_934 (O_934,N_12653,N_10025);
nand UO_935 (O_935,N_11640,N_14331);
xor UO_936 (O_936,N_10605,N_11619);
nor UO_937 (O_937,N_11705,N_13224);
xor UO_938 (O_938,N_14037,N_11550);
or UO_939 (O_939,N_10876,N_11873);
and UO_940 (O_940,N_12401,N_14801);
nor UO_941 (O_941,N_13838,N_13372);
xnor UO_942 (O_942,N_12871,N_11784);
and UO_943 (O_943,N_11202,N_11517);
or UO_944 (O_944,N_12612,N_14112);
nor UO_945 (O_945,N_14937,N_14741);
and UO_946 (O_946,N_14487,N_11631);
xor UO_947 (O_947,N_11485,N_14737);
and UO_948 (O_948,N_11876,N_13232);
nor UO_949 (O_949,N_12196,N_11765);
or UO_950 (O_950,N_11329,N_12925);
xnor UO_951 (O_951,N_13763,N_10786);
xor UO_952 (O_952,N_12311,N_10214);
nand UO_953 (O_953,N_12444,N_14157);
xor UO_954 (O_954,N_14999,N_12120);
nand UO_955 (O_955,N_10271,N_11570);
nand UO_956 (O_956,N_10380,N_12480);
and UO_957 (O_957,N_10482,N_10470);
and UO_958 (O_958,N_10443,N_11534);
and UO_959 (O_959,N_11058,N_10656);
nand UO_960 (O_960,N_13445,N_13705);
xor UO_961 (O_961,N_11811,N_12390);
or UO_962 (O_962,N_14365,N_11097);
nor UO_963 (O_963,N_14676,N_12592);
nand UO_964 (O_964,N_11317,N_12051);
nand UO_965 (O_965,N_12773,N_14414);
nand UO_966 (O_966,N_14546,N_14503);
nand UO_967 (O_967,N_14732,N_13910);
xor UO_968 (O_968,N_14121,N_12965);
nor UO_969 (O_969,N_13587,N_10384);
and UO_970 (O_970,N_13407,N_14062);
xnor UO_971 (O_971,N_11745,N_10362);
and UO_972 (O_972,N_13111,N_11423);
nor UO_973 (O_973,N_14304,N_12109);
nand UO_974 (O_974,N_12525,N_10070);
nor UO_975 (O_975,N_13183,N_12553);
nor UO_976 (O_976,N_10891,N_12853);
nor UO_977 (O_977,N_11263,N_11617);
nor UO_978 (O_978,N_13235,N_14209);
xor UO_979 (O_979,N_11138,N_13854);
or UO_980 (O_980,N_13598,N_14297);
and UO_981 (O_981,N_14692,N_12335);
nand UO_982 (O_982,N_13259,N_12447);
nor UO_983 (O_983,N_12822,N_14603);
nand UO_984 (O_984,N_10340,N_11742);
xnor UO_985 (O_985,N_11467,N_13120);
nor UO_986 (O_986,N_11728,N_10918);
and UO_987 (O_987,N_10725,N_10479);
or UO_988 (O_988,N_14725,N_10585);
or UO_989 (O_989,N_11594,N_10658);
nand UO_990 (O_990,N_12542,N_11899);
nand UO_991 (O_991,N_14267,N_13452);
and UO_992 (O_992,N_10100,N_10550);
xnor UO_993 (O_993,N_13307,N_12780);
nor UO_994 (O_994,N_12481,N_13276);
xor UO_995 (O_995,N_11935,N_10766);
and UO_996 (O_996,N_10925,N_13804);
nand UO_997 (O_997,N_11507,N_12214);
or UO_998 (O_998,N_13285,N_13828);
or UO_999 (O_999,N_12776,N_13694);
or UO_1000 (O_1000,N_10590,N_13713);
nand UO_1001 (O_1001,N_10134,N_14633);
nand UO_1002 (O_1002,N_13355,N_10735);
and UO_1003 (O_1003,N_11474,N_12378);
nor UO_1004 (O_1004,N_14366,N_12898);
and UO_1005 (O_1005,N_14446,N_14686);
and UO_1006 (O_1006,N_10265,N_12670);
nand UO_1007 (O_1007,N_11460,N_13512);
nor UO_1008 (O_1008,N_14827,N_10143);
nand UO_1009 (O_1009,N_11842,N_13691);
xnor UO_1010 (O_1010,N_10596,N_14938);
nor UO_1011 (O_1011,N_13629,N_13626);
or UO_1012 (O_1012,N_11675,N_12163);
xnor UO_1013 (O_1013,N_11229,N_13085);
nand UO_1014 (O_1014,N_13357,N_11370);
or UO_1015 (O_1015,N_11119,N_13494);
and UO_1016 (O_1016,N_13408,N_12587);
nor UO_1017 (O_1017,N_11794,N_11590);
nand UO_1018 (O_1018,N_12520,N_13141);
or UO_1019 (O_1019,N_14107,N_14619);
nand UO_1020 (O_1020,N_10574,N_14780);
nand UO_1021 (O_1021,N_10464,N_11602);
xor UO_1022 (O_1022,N_11997,N_13139);
xnor UO_1023 (O_1023,N_13484,N_14202);
nor UO_1024 (O_1024,N_14933,N_12192);
nor UO_1025 (O_1025,N_13792,N_10830);
xnor UO_1026 (O_1026,N_11018,N_13065);
or UO_1027 (O_1027,N_13536,N_12787);
nor UO_1028 (O_1028,N_13359,N_12680);
and UO_1029 (O_1029,N_14198,N_12275);
and UO_1030 (O_1030,N_12280,N_11610);
nand UO_1031 (O_1031,N_11469,N_13356);
nor UO_1032 (O_1032,N_13559,N_13095);
nor UO_1033 (O_1033,N_13824,N_12878);
xor UO_1034 (O_1034,N_14646,N_12450);
nor UO_1035 (O_1035,N_14688,N_12371);
nor UO_1036 (O_1036,N_10102,N_10454);
nor UO_1037 (O_1037,N_12342,N_12633);
nor UO_1038 (O_1038,N_13516,N_11540);
nand UO_1039 (O_1039,N_11864,N_12761);
and UO_1040 (O_1040,N_12747,N_11584);
and UO_1041 (O_1041,N_10072,N_11205);
nor UO_1042 (O_1042,N_12223,N_11005);
and UO_1043 (O_1043,N_10063,N_14975);
nor UO_1044 (O_1044,N_14371,N_13013);
nand UO_1045 (O_1045,N_12263,N_13670);
nand UO_1046 (O_1046,N_13736,N_11846);
nand UO_1047 (O_1047,N_10452,N_11837);
nor UO_1048 (O_1048,N_12535,N_10771);
nor UO_1049 (O_1049,N_12017,N_14736);
or UO_1050 (O_1050,N_10576,N_12897);
nand UO_1051 (O_1051,N_14478,N_14163);
nor UO_1052 (O_1052,N_11416,N_13724);
nand UO_1053 (O_1053,N_10349,N_11461);
nand UO_1054 (O_1054,N_10126,N_13211);
nor UO_1055 (O_1055,N_13381,N_13323);
or UO_1056 (O_1056,N_14599,N_12127);
nor UO_1057 (O_1057,N_10409,N_10260);
nor UO_1058 (O_1058,N_10719,N_13138);
nand UO_1059 (O_1059,N_12539,N_12437);
or UO_1060 (O_1060,N_10688,N_10110);
nand UO_1061 (O_1061,N_12682,N_13519);
nor UO_1062 (O_1062,N_13837,N_13643);
xor UO_1063 (O_1063,N_10569,N_14256);
or UO_1064 (O_1064,N_14038,N_13938);
and UO_1065 (O_1065,N_14496,N_11355);
xnor UO_1066 (O_1066,N_11383,N_12540);
nor UO_1067 (O_1067,N_11569,N_13710);
or UO_1068 (O_1068,N_10939,N_11197);
or UO_1069 (O_1069,N_13147,N_14076);
or UO_1070 (O_1070,N_12847,N_11277);
and UO_1071 (O_1071,N_10642,N_12168);
nand UO_1072 (O_1072,N_14247,N_10967);
xor UO_1073 (O_1073,N_14053,N_11770);
nand UO_1074 (O_1074,N_13599,N_11762);
nand UO_1075 (O_1075,N_11637,N_10335);
and UO_1076 (O_1076,N_11750,N_10671);
or UO_1077 (O_1077,N_11029,N_13553);
nand UO_1078 (O_1078,N_12215,N_11436);
and UO_1079 (O_1079,N_13254,N_10952);
or UO_1080 (O_1080,N_14861,N_10337);
or UO_1081 (O_1081,N_10246,N_12548);
nor UO_1082 (O_1082,N_12301,N_13070);
nor UO_1083 (O_1083,N_12203,N_12486);
xor UO_1084 (O_1084,N_12037,N_12820);
xnor UO_1085 (O_1085,N_10389,N_10615);
and UO_1086 (O_1086,N_14323,N_12043);
xnor UO_1087 (O_1087,N_12050,N_11448);
xnor UO_1088 (O_1088,N_14852,N_14230);
nand UO_1089 (O_1089,N_12235,N_10361);
or UO_1090 (O_1090,N_14033,N_12354);
or UO_1091 (O_1091,N_10259,N_12999);
or UO_1092 (O_1092,N_10376,N_12809);
nand UO_1093 (O_1093,N_14276,N_13291);
nor UO_1094 (O_1094,N_13895,N_10142);
nor UO_1095 (O_1095,N_10751,N_12950);
or UO_1096 (O_1096,N_11648,N_10198);
or UO_1097 (O_1097,N_10364,N_12524);
and UO_1098 (O_1098,N_10669,N_13680);
and UO_1099 (O_1099,N_10890,N_12374);
nand UO_1100 (O_1100,N_10494,N_10419);
xor UO_1101 (O_1101,N_11154,N_11491);
nor UO_1102 (O_1102,N_12685,N_10616);
and UO_1103 (O_1103,N_11480,N_11979);
and UO_1104 (O_1104,N_11162,N_11759);
or UO_1105 (O_1105,N_13809,N_13078);
nand UO_1106 (O_1106,N_14841,N_12752);
or UO_1107 (O_1107,N_14450,N_14481);
nor UO_1108 (O_1108,N_11752,N_13518);
nand UO_1109 (O_1109,N_12111,N_12751);
nand UO_1110 (O_1110,N_11773,N_14309);
xnor UO_1111 (O_1111,N_11456,N_13858);
and UO_1112 (O_1112,N_13196,N_14310);
nand UO_1113 (O_1113,N_13299,N_14563);
xor UO_1114 (O_1114,N_12058,N_14948);
or UO_1115 (O_1115,N_11954,N_10331);
or UO_1116 (O_1116,N_13312,N_12338);
xor UO_1117 (O_1117,N_11641,N_13831);
nor UO_1118 (O_1118,N_12537,N_11630);
and UO_1119 (O_1119,N_12862,N_12136);
nand UO_1120 (O_1120,N_13229,N_13915);
nand UO_1121 (O_1121,N_11458,N_13131);
xnor UO_1122 (O_1122,N_14906,N_13490);
and UO_1123 (O_1123,N_10772,N_11901);
xor UO_1124 (O_1124,N_10222,N_10155);
and UO_1125 (O_1125,N_10403,N_10122);
or UO_1126 (O_1126,N_12435,N_14432);
nor UO_1127 (O_1127,N_14311,N_12054);
nor UO_1128 (O_1128,N_10770,N_14040);
and UO_1129 (O_1129,N_10697,N_10670);
nor UO_1130 (O_1130,N_14511,N_14456);
or UO_1131 (O_1131,N_10519,N_12185);
and UO_1132 (O_1132,N_11421,N_10158);
and UO_1133 (O_1133,N_10896,N_13238);
nor UO_1134 (O_1134,N_11717,N_12890);
xor UO_1135 (O_1135,N_11603,N_11894);
xnor UO_1136 (O_1136,N_12982,N_12735);
nor UO_1137 (O_1137,N_13949,N_11133);
nand UO_1138 (O_1138,N_14586,N_14032);
nand UO_1139 (O_1139,N_10966,N_10776);
and UO_1140 (O_1140,N_10971,N_12013);
and UO_1141 (O_1141,N_13412,N_10264);
and UO_1142 (O_1142,N_13421,N_14302);
nand UO_1143 (O_1143,N_11967,N_12270);
xnor UO_1144 (O_1144,N_14291,N_10498);
nand UO_1145 (O_1145,N_14820,N_13613);
nor UO_1146 (O_1146,N_14483,N_11588);
nand UO_1147 (O_1147,N_13655,N_14000);
or UO_1148 (O_1148,N_11168,N_10788);
and UO_1149 (O_1149,N_11499,N_10045);
nor UO_1150 (O_1150,N_11446,N_12169);
nand UO_1151 (O_1151,N_11433,N_12264);
and UO_1152 (O_1152,N_14781,N_12608);
and UO_1153 (O_1153,N_10441,N_12759);
nand UO_1154 (O_1154,N_13656,N_13294);
or UO_1155 (O_1155,N_14639,N_10157);
and UO_1156 (O_1156,N_11678,N_11611);
nand UO_1157 (O_1157,N_12146,N_14870);
xor UO_1158 (O_1158,N_12826,N_13956);
nor UO_1159 (O_1159,N_13242,N_13373);
or UO_1160 (O_1160,N_13841,N_12417);
nand UO_1161 (O_1161,N_13863,N_11147);
or UO_1162 (O_1162,N_12115,N_11875);
nand UO_1163 (O_1163,N_12064,N_12148);
nor UO_1164 (O_1164,N_12724,N_13300);
and UO_1165 (O_1165,N_11403,N_11108);
or UO_1166 (O_1166,N_14057,N_13290);
nand UO_1167 (O_1167,N_13808,N_11609);
and UO_1168 (O_1168,N_12147,N_14626);
and UO_1169 (O_1169,N_13632,N_10204);
and UO_1170 (O_1170,N_12675,N_14243);
or UO_1171 (O_1171,N_10103,N_12056);
xnor UO_1172 (O_1172,N_14812,N_13081);
and UO_1173 (O_1173,N_10613,N_12770);
nand UO_1174 (O_1174,N_12549,N_12620);
and UO_1175 (O_1175,N_10195,N_11009);
or UO_1176 (O_1176,N_14403,N_10650);
nand UO_1177 (O_1177,N_13091,N_14376);
nand UO_1178 (O_1178,N_14695,N_10852);
nor UO_1179 (O_1179,N_10481,N_11470);
and UO_1180 (O_1180,N_12805,N_14482);
nand UO_1181 (O_1181,N_14352,N_11490);
xnor UO_1182 (O_1182,N_12012,N_12536);
and UO_1183 (O_1183,N_10703,N_13352);
and UO_1184 (O_1184,N_14099,N_11798);
nor UO_1185 (O_1185,N_11084,N_13514);
nor UO_1186 (O_1186,N_14278,N_12326);
nand UO_1187 (O_1187,N_13964,N_12451);
and UO_1188 (O_1188,N_11504,N_14815);
nor UO_1189 (O_1189,N_13877,N_13450);
and UO_1190 (O_1190,N_13365,N_11354);
or UO_1191 (O_1191,N_11895,N_13112);
nand UO_1192 (O_1192,N_13962,N_10351);
nand UO_1193 (O_1193,N_11835,N_12272);
nor UO_1194 (O_1194,N_12825,N_14899);
nand UO_1195 (O_1195,N_10128,N_14810);
nor UO_1196 (O_1196,N_10843,N_10627);
xnor UO_1197 (O_1197,N_10429,N_13530);
nor UO_1198 (O_1198,N_12038,N_14537);
nor UO_1199 (O_1199,N_10914,N_11336);
nor UO_1200 (O_1200,N_12864,N_10396);
or UO_1201 (O_1201,N_14798,N_11247);
nor UO_1202 (O_1202,N_11434,N_10558);
or UO_1203 (O_1203,N_13513,N_14969);
or UO_1204 (O_1204,N_14674,N_14650);
nand UO_1205 (O_1205,N_10834,N_10581);
and UO_1206 (O_1206,N_14325,N_14703);
and UO_1207 (O_1207,N_10554,N_11186);
and UO_1208 (O_1208,N_12025,N_12868);
nand UO_1209 (O_1209,N_13909,N_12039);
and UO_1210 (O_1210,N_12494,N_10234);
xor UO_1211 (O_1211,N_10782,N_10708);
and UO_1212 (O_1212,N_13509,N_11230);
or UO_1213 (O_1213,N_14706,N_12665);
and UO_1214 (O_1214,N_11241,N_11897);
xor UO_1215 (O_1215,N_13995,N_11535);
and UO_1216 (O_1216,N_13010,N_13654);
nand UO_1217 (O_1217,N_14014,N_11435);
nor UO_1218 (O_1218,N_14518,N_12022);
xnor UO_1219 (O_1219,N_12717,N_13634);
nor UO_1220 (O_1220,N_12358,N_10484);
and UO_1221 (O_1221,N_11043,N_12638);
nand UO_1222 (O_1222,N_14497,N_11343);
xnor UO_1223 (O_1223,N_14010,N_13965);
xor UO_1224 (O_1224,N_13063,N_11810);
xor UO_1225 (O_1225,N_11553,N_14077);
or UO_1226 (O_1226,N_14171,N_12242);
and UO_1227 (O_1227,N_11776,N_11924);
nand UO_1228 (O_1228,N_12317,N_14465);
nand UO_1229 (O_1229,N_14218,N_14876);
or UO_1230 (O_1230,N_11548,N_10020);
xor UO_1231 (O_1231,N_11613,N_14388);
nor UO_1232 (O_1232,N_12953,N_13635);
xor UO_1233 (O_1233,N_10807,N_13538);
xor UO_1234 (O_1234,N_10898,N_11276);
nand UO_1235 (O_1235,N_11506,N_10021);
and UO_1236 (O_1236,N_10168,N_13596);
and UO_1237 (O_1237,N_14285,N_10154);
nor UO_1238 (O_1238,N_12355,N_12596);
nor UO_1239 (O_1239,N_13779,N_14349);
xnor UO_1240 (O_1240,N_12792,N_14079);
nor UO_1241 (O_1241,N_12855,N_13037);
xor UO_1242 (O_1242,N_10413,N_12221);
xnor UO_1243 (O_1243,N_10961,N_14889);
nand UO_1244 (O_1244,N_13914,N_14026);
and UO_1245 (O_1245,N_14638,N_14335);
nor UO_1246 (O_1246,N_13216,N_13968);
or UO_1247 (O_1247,N_14712,N_10622);
or UO_1248 (O_1248,N_12154,N_10463);
or UO_1249 (O_1249,N_14357,N_13022);
or UO_1250 (O_1250,N_12760,N_13234);
nor UO_1251 (O_1251,N_13071,N_13275);
nor UO_1252 (O_1252,N_12828,N_10698);
nand UO_1253 (O_1253,N_13342,N_11107);
nor UO_1254 (O_1254,N_10445,N_11078);
nand UO_1255 (O_1255,N_11030,N_12714);
nor UO_1256 (O_1256,N_11598,N_12313);
nand UO_1257 (O_1257,N_10129,N_10521);
or UO_1258 (O_1258,N_14417,N_10988);
nand UO_1259 (O_1259,N_10749,N_13062);
nor UO_1260 (O_1260,N_13707,N_13026);
or UO_1261 (O_1261,N_12963,N_10432);
or UO_1262 (O_1262,N_14840,N_11555);
and UO_1263 (O_1263,N_12246,N_13711);
and UO_1264 (O_1264,N_12519,N_13578);
nand UO_1265 (O_1265,N_13820,N_10201);
and UO_1266 (O_1266,N_11156,N_11189);
and UO_1267 (O_1267,N_12886,N_10145);
nand UO_1268 (O_1268,N_10316,N_11387);
nor UO_1269 (O_1269,N_11131,N_10539);
nand UO_1270 (O_1270,N_12909,N_12916);
or UO_1271 (O_1271,N_11629,N_11596);
xor UO_1272 (O_1272,N_10211,N_13892);
nand UO_1273 (O_1273,N_14754,N_13987);
nand UO_1274 (O_1274,N_12011,N_10533);
nor UO_1275 (O_1275,N_13053,N_10879);
and UO_1276 (O_1276,N_14003,N_11381);
or UO_1277 (O_1277,N_12949,N_12924);
nand UO_1278 (O_1278,N_11563,N_12394);
xnor UO_1279 (O_1279,N_12681,N_12513);
or UO_1280 (O_1280,N_11116,N_11479);
xnor UO_1281 (O_1281,N_14597,N_12609);
nand UO_1282 (O_1282,N_12422,N_12991);
nand UO_1283 (O_1283,N_10281,N_10525);
nor UO_1284 (O_1284,N_10160,N_13174);
nor UO_1285 (O_1285,N_14509,N_10292);
or UO_1286 (O_1286,N_13233,N_12857);
nor UO_1287 (O_1287,N_14462,N_14134);
and UO_1288 (O_1288,N_11155,N_10630);
nand UO_1289 (O_1289,N_10164,N_14924);
or UO_1290 (O_1290,N_13423,N_13094);
and UO_1291 (O_1291,N_12616,N_13277);
and UO_1292 (O_1292,N_10287,N_12141);
nor UO_1293 (O_1293,N_11822,N_12347);
nor UO_1294 (O_1294,N_12573,N_13883);
and UO_1295 (O_1295,N_14308,N_14390);
or UO_1296 (O_1296,N_11855,N_11834);
or UO_1297 (O_1297,N_14594,N_14571);
nand UO_1298 (O_1298,N_11564,N_11547);
and UO_1299 (O_1299,N_13630,N_11868);
xnor UO_1300 (O_1300,N_11638,N_11880);
or UO_1301 (O_1301,N_14367,N_13611);
nand UO_1302 (O_1302,N_11500,N_10727);
or UO_1303 (O_1303,N_12691,N_12455);
and UO_1304 (O_1304,N_11681,N_11713);
or UO_1305 (O_1305,N_12758,N_10676);
nand UO_1306 (O_1306,N_10023,N_12276);
and UO_1307 (O_1307,N_10247,N_14255);
xnor UO_1308 (O_1308,N_13226,N_10235);
xor UO_1309 (O_1309,N_12729,N_12661);
nand UO_1310 (O_1310,N_14672,N_10350);
or UO_1311 (O_1311,N_10417,N_13470);
and UO_1312 (O_1312,N_12887,N_12472);
nand UO_1313 (O_1313,N_11840,N_11946);
nand UO_1314 (O_1314,N_11715,N_11948);
nor UO_1315 (O_1315,N_13975,N_12819);
nand UO_1316 (O_1316,N_13871,N_11284);
nor UO_1317 (O_1317,N_10188,N_12930);
and UO_1318 (O_1318,N_11929,N_13646);
xor UO_1319 (O_1319,N_12132,N_12005);
nand UO_1320 (O_1320,N_11194,N_10958);
nand UO_1321 (O_1321,N_12574,N_11706);
or UO_1322 (O_1322,N_11993,N_10317);
and UO_1323 (O_1323,N_10112,N_12988);
nand UO_1324 (O_1324,N_14253,N_10461);
or UO_1325 (O_1325,N_14455,N_11519);
and UO_1326 (O_1326,N_12036,N_13719);
nor UO_1327 (O_1327,N_13983,N_10870);
and UO_1328 (O_1328,N_11980,N_14871);
and UO_1329 (O_1329,N_11325,N_11032);
nand UO_1330 (O_1330,N_12473,N_11267);
xnor UO_1331 (O_1331,N_12088,N_13609);
and UO_1332 (O_1332,N_14779,N_12551);
xor UO_1333 (O_1333,N_10955,N_13783);
nor UO_1334 (O_1334,N_13497,N_13638);
xnor UO_1335 (O_1335,N_11020,N_13166);
nor UO_1336 (O_1336,N_14155,N_11034);
and UO_1337 (O_1337,N_10963,N_11632);
nand UO_1338 (O_1338,N_12460,N_12915);
or UO_1339 (O_1339,N_10863,N_12362);
xor UO_1340 (O_1340,N_11923,N_10135);
xor UO_1341 (O_1341,N_12420,N_10526);
nor UO_1342 (O_1342,N_12430,N_12293);
and UO_1343 (O_1343,N_13193,N_12199);
nand UO_1344 (O_1344,N_13059,N_11653);
nand UO_1345 (O_1345,N_12565,N_13961);
and UO_1346 (O_1346,N_14239,N_14115);
and UO_1347 (O_1347,N_11531,N_14976);
and UO_1348 (O_1348,N_10486,N_13844);
xor UO_1349 (O_1349,N_13737,N_10326);
xnor UO_1350 (O_1350,N_12948,N_14168);
nor UO_1351 (O_1351,N_13564,N_11293);
nor UO_1352 (O_1352,N_12974,N_13781);
nand UO_1353 (O_1353,N_11160,N_10848);
and UO_1354 (O_1354,N_12563,N_10003);
xor UO_1355 (O_1355,N_11159,N_14947);
or UO_1356 (O_1356,N_10877,N_13479);
nor UO_1357 (O_1357,N_14343,N_10273);
nand UO_1358 (O_1358,N_11297,N_10423);
and UO_1359 (O_1359,N_13818,N_10115);
nand UO_1360 (O_1360,N_11062,N_14713);
nand UO_1361 (O_1361,N_10803,N_10085);
nand UO_1362 (O_1362,N_14578,N_11970);
and UO_1363 (O_1363,N_12774,N_12583);
nor UO_1364 (O_1364,N_14041,N_10858);
xnor UO_1365 (O_1365,N_12240,N_13528);
nor UO_1366 (O_1366,N_13617,N_14058);
xnor UO_1367 (O_1367,N_12375,N_12493);
nand UO_1368 (O_1368,N_11909,N_10200);
or UO_1369 (O_1369,N_13967,N_12289);
or UO_1370 (O_1370,N_14020,N_14910);
and UO_1371 (O_1371,N_13542,N_11089);
and UO_1372 (O_1372,N_14843,N_13927);
or UO_1373 (O_1373,N_14141,N_13204);
xnor UO_1374 (O_1374,N_14231,N_12407);
nor UO_1375 (O_1375,N_11290,N_10557);
and UO_1376 (O_1376,N_13998,N_12546);
nor UO_1377 (O_1377,N_10942,N_13035);
or UO_1378 (O_1378,N_13897,N_13409);
nand UO_1379 (O_1379,N_10383,N_12060);
nand UO_1380 (O_1380,N_12490,N_10911);
and UO_1381 (O_1381,N_10527,N_10438);
xor UO_1382 (O_1382,N_11866,N_12176);
and UO_1383 (O_1383,N_11796,N_11328);
nand UO_1384 (O_1384,N_13164,N_12125);
and UO_1385 (O_1385,N_11157,N_10800);
nor UO_1386 (O_1386,N_10975,N_12377);
and UO_1387 (O_1387,N_13360,N_12166);
nor UO_1388 (O_1388,N_10912,N_13537);
xor UO_1389 (O_1389,N_11622,N_10069);
or UO_1390 (O_1390,N_13496,N_11340);
nor UO_1391 (O_1391,N_12944,N_14124);
and UO_1392 (O_1392,N_10297,N_10949);
nand UO_1393 (O_1393,N_10959,N_11240);
xor UO_1394 (O_1394,N_13722,N_14623);
nand UO_1395 (O_1395,N_13651,N_14313);
nor UO_1396 (O_1396,N_13100,N_11785);
or UO_1397 (O_1397,N_10728,N_12063);
xnor UO_1398 (O_1398,N_14585,N_10835);
nand UO_1399 (O_1399,N_10571,N_14847);
or UO_1400 (O_1400,N_11356,N_13464);
nand UO_1401 (O_1401,N_14898,N_12161);
nor UO_1402 (O_1402,N_12870,N_12290);
and UO_1403 (O_1403,N_10374,N_10555);
xor UO_1404 (O_1404,N_13649,N_11670);
nand UO_1405 (O_1405,N_10797,N_11574);
nand UO_1406 (O_1406,N_10139,N_13926);
and UO_1407 (O_1407,N_10300,N_13018);
nor UO_1408 (O_1408,N_12755,N_13135);
xnor UO_1409 (O_1409,N_14108,N_10329);
or UO_1410 (O_1410,N_13584,N_12029);
nand UO_1411 (O_1411,N_11995,N_14562);
nor UO_1412 (O_1412,N_13295,N_14152);
nand UO_1413 (O_1413,N_10565,N_11693);
nand UO_1414 (O_1414,N_10653,N_14955);
nor UO_1415 (O_1415,N_14090,N_14355);
xor UO_1416 (O_1416,N_14443,N_12042);
or UO_1417 (O_1417,N_11411,N_10079);
and UO_1418 (O_1418,N_13563,N_10753);
and UO_1419 (O_1419,N_10679,N_11711);
nor UO_1420 (O_1420,N_14480,N_14520);
or UO_1421 (O_1421,N_10517,N_14919);
or UO_1422 (O_1422,N_14818,N_11371);
or UO_1423 (O_1423,N_13912,N_10116);
nor UO_1424 (O_1424,N_11999,N_13474);
xor UO_1425 (O_1425,N_12511,N_14926);
and UO_1426 (O_1426,N_12610,N_10553);
and UO_1427 (O_1427,N_10397,N_13627);
or UO_1428 (O_1428,N_10704,N_12019);
and UO_1429 (O_1429,N_12441,N_14927);
nand UO_1430 (O_1430,N_13784,N_13767);
nor UO_1431 (O_1431,N_14932,N_13437);
or UO_1432 (O_1432,N_12464,N_10244);
or UO_1433 (O_1433,N_11614,N_10325);
nor UO_1434 (O_1434,N_10258,N_14389);
nor UO_1435 (O_1435,N_13385,N_13025);
nand UO_1436 (O_1436,N_10420,N_10880);
or UO_1437 (O_1437,N_11180,N_13623);
or UO_1438 (O_1438,N_14474,N_11792);
or UO_1439 (O_1439,N_11312,N_10093);
or UO_1440 (O_1440,N_10140,N_13794);
xnor UO_1441 (O_1441,N_10610,N_12976);
nor UO_1442 (O_1442,N_10106,N_13371);
xnor UO_1443 (O_1443,N_11537,N_13689);
and UO_1444 (O_1444,N_11814,N_10983);
nor UO_1445 (O_1445,N_14317,N_13674);
nand UO_1446 (O_1446,N_14259,N_12883);
xnor UO_1447 (O_1447,N_14216,N_11185);
xor UO_1448 (O_1448,N_12181,N_10228);
nor UO_1449 (O_1449,N_12159,N_10015);
or UO_1450 (O_1450,N_10618,N_12258);
nor UO_1451 (O_1451,N_11231,N_12392);
and UO_1452 (O_1452,N_11094,N_14386);
nor UO_1453 (O_1453,N_14886,N_13612);
or UO_1454 (O_1454,N_14132,N_11593);
nand UO_1455 (O_1455,N_11067,N_14595);
nor UO_1456 (O_1456,N_14807,N_11541);
and UO_1457 (O_1457,N_10321,N_14760);
xor UO_1458 (O_1458,N_12576,N_10844);
nand UO_1459 (O_1459,N_11871,N_14251);
nand UO_1460 (O_1460,N_13278,N_12637);
and UO_1461 (O_1461,N_13348,N_13756);
nand UO_1462 (O_1462,N_12875,N_10232);
nand UO_1463 (O_1463,N_12097,N_10948);
or UO_1464 (O_1464,N_14263,N_13853);
nand UO_1465 (O_1465,N_14126,N_13859);
or UO_1466 (O_1466,N_12968,N_11275);
nand UO_1467 (O_1467,N_14117,N_11183);
nand UO_1468 (O_1468,N_11513,N_12232);
xnor UO_1469 (O_1469,N_11691,N_11044);
xor UO_1470 (O_1470,N_12425,N_14439);
nor UO_1471 (O_1471,N_13505,N_11114);
or UO_1472 (O_1472,N_14095,N_10801);
nand UO_1473 (O_1473,N_12393,N_13955);
nand UO_1474 (O_1474,N_14945,N_14238);
xnor UO_1475 (O_1475,N_13893,N_14615);
nand UO_1476 (O_1476,N_10677,N_12310);
or UO_1477 (O_1477,N_11494,N_13521);
nand UO_1478 (O_1478,N_12433,N_13482);
and UO_1479 (O_1479,N_14540,N_12731);
and UO_1480 (O_1480,N_12848,N_12841);
or UO_1481 (O_1481,N_14758,N_14072);
or UO_1482 (O_1482,N_11872,N_10645);
and UO_1483 (O_1483,N_11529,N_11974);
nand UO_1484 (O_1484,N_14272,N_14987);
nand UO_1485 (O_1485,N_13950,N_14316);
or UO_1486 (O_1486,N_13684,N_14199);
and UO_1487 (O_1487,N_13477,N_12016);
xnor UO_1488 (O_1488,N_14504,N_13679);
nor UO_1489 (O_1489,N_11788,N_12381);
or UO_1490 (O_1490,N_11161,N_14187);
or UO_1491 (O_1491,N_12031,N_14566);
xor UO_1492 (O_1492,N_14698,N_12186);
nand UO_1493 (O_1493,N_12254,N_14153);
xnor UO_1494 (O_1494,N_10668,N_14494);
nand UO_1495 (O_1495,N_14036,N_13440);
or UO_1496 (O_1496,N_14060,N_12648);
nor UO_1497 (O_1497,N_12052,N_10831);
or UO_1498 (O_1498,N_12739,N_10838);
nor UO_1499 (O_1499,N_11245,N_10850);
nand UO_1500 (O_1500,N_13186,N_14426);
or UO_1501 (O_1501,N_11014,N_10646);
nor UO_1502 (O_1502,N_11218,N_10547);
or UO_1503 (O_1503,N_14284,N_10579);
nand UO_1504 (O_1504,N_14354,N_12331);
xor UO_1505 (O_1505,N_11690,N_14471);
xor UO_1506 (O_1506,N_12189,N_12626);
nor UO_1507 (O_1507,N_13424,N_11042);
and UO_1508 (O_1508,N_14918,N_13816);
nand UO_1509 (O_1509,N_14762,N_13154);
nor UO_1510 (O_1510,N_10067,N_14150);
or UO_1511 (O_1511,N_12344,N_11888);
nor UO_1512 (O_1512,N_13695,N_14110);
nor UO_1513 (O_1513,N_14522,N_10382);
xnor UO_1514 (O_1514,N_10381,N_13221);
xnor UO_1515 (O_1515,N_14019,N_10446);
or UO_1516 (O_1516,N_12764,N_14532);
nand UO_1517 (O_1517,N_12908,N_11730);
and UO_1518 (O_1518,N_12559,N_10475);
and UO_1519 (O_1519,N_14510,N_12302);
xor UO_1520 (O_1520,N_13284,N_11134);
or UO_1521 (O_1521,N_11848,N_10859);
xor UO_1522 (O_1522,N_11405,N_11350);
nand UO_1523 (O_1523,N_11558,N_10097);
nand UO_1524 (O_1524,N_11587,N_10647);
nand UO_1525 (O_1525,N_14186,N_14644);
or UO_1526 (O_1526,N_13548,N_11439);
xnor UO_1527 (O_1527,N_13447,N_13087);
xor UO_1528 (O_1528,N_11226,N_10253);
or UO_1529 (O_1529,N_11141,N_12615);
nor UO_1530 (O_1530,N_13546,N_12349);
nand UO_1531 (O_1531,N_14776,N_11698);
and UO_1532 (O_1532,N_13489,N_11118);
nor UO_1533 (O_1533,N_10313,N_11838);
nand UO_1534 (O_1534,N_12068,N_11139);
nand UO_1535 (O_1535,N_13571,N_14123);
xor UO_1536 (O_1536,N_14536,N_14294);
nand UO_1537 (O_1537,N_10137,N_14287);
or UO_1538 (O_1538,N_10941,N_13672);
and UO_1539 (O_1539,N_13252,N_10252);
xor UO_1540 (O_1540,N_14051,N_13658);
nor UO_1541 (O_1541,N_10981,N_13592);
and UO_1542 (O_1542,N_10175,N_10820);
nor UO_1543 (O_1543,N_13836,N_14831);
and UO_1544 (O_1544,N_14893,N_11597);
and UO_1545 (O_1545,N_11673,N_13439);
or UO_1546 (O_1546,N_10577,N_13039);
or UO_1547 (O_1547,N_14751,N_11239);
or UO_1548 (O_1548,N_14004,N_13847);
or UO_1549 (O_1549,N_12830,N_13992);
or UO_1550 (O_1550,N_10125,N_13379);
or UO_1551 (O_1551,N_13774,N_10762);
nor UO_1552 (O_1552,N_10182,N_10368);
and UO_1553 (O_1553,N_13712,N_13789);
or UO_1554 (O_1554,N_14838,N_11516);
nor UO_1555 (O_1555,N_14547,N_12350);
nor UO_1556 (O_1556,N_13899,N_14845);
nor UO_1557 (O_1557,N_10086,N_12797);
and UO_1558 (O_1558,N_13531,N_12101);
xnor UO_1559 (O_1559,N_14475,N_13411);
xor UO_1560 (O_1560,N_10804,N_14723);
nor UO_1561 (O_1561,N_13846,N_10030);
or UO_1562 (O_1562,N_12492,N_10729);
nand UO_1563 (O_1563,N_14369,N_13588);
and UO_1564 (O_1564,N_10694,N_14236);
and UO_1565 (O_1565,N_13766,N_11740);
nand UO_1566 (O_1566,N_14144,N_10587);
or UO_1567 (O_1567,N_12594,N_10450);
and UO_1568 (O_1568,N_10330,N_12014);
nor UO_1569 (O_1569,N_14662,N_13247);
and UO_1570 (O_1570,N_13734,N_12325);
xor UO_1571 (O_1571,N_14016,N_11824);
and UO_1572 (O_1572,N_10414,N_13660);
xor UO_1573 (O_1573,N_12046,N_12266);
or UO_1574 (O_1574,N_14582,N_10303);
and UO_1575 (O_1575,N_10980,N_14262);
nor UO_1576 (O_1576,N_12711,N_11320);
or UO_1577 (O_1577,N_10298,N_12528);
nor UO_1578 (O_1578,N_14468,N_11465);
xnor UO_1579 (O_1579,N_12365,N_10887);
and UO_1580 (O_1580,N_11252,N_14610);
and UO_1581 (O_1581,N_14593,N_13260);
nor UO_1582 (O_1582,N_11861,N_10159);
nand UO_1583 (O_1583,N_14628,N_10109);
xor UO_1584 (O_1584,N_14799,N_12634);
nand UO_1585 (O_1585,N_12248,N_10828);
nand UO_1586 (O_1586,N_11111,N_13569);
nand UO_1587 (O_1587,N_11562,N_13589);
and UO_1588 (O_1588,N_13429,N_13511);
and UO_1589 (O_1589,N_13935,N_13317);
and UO_1590 (O_1590,N_12967,N_11363);
and UO_1591 (O_1591,N_14860,N_12668);
or UO_1592 (O_1592,N_14621,N_14114);
or UO_1593 (O_1593,N_12522,N_12957);
xor UO_1594 (O_1594,N_12625,N_13974);
and UO_1595 (O_1595,N_14963,N_12316);
nor UO_1596 (O_1596,N_10864,N_14429);
nor UO_1597 (O_1597,N_12733,N_14819);
nor UO_1598 (O_1598,N_13787,N_12061);
xor UO_1599 (O_1599,N_11642,N_11557);
or UO_1600 (O_1600,N_12772,N_12630);
xor UO_1601 (O_1601,N_14773,N_10156);
xnor UO_1602 (O_1602,N_14765,N_14996);
xor UO_1603 (O_1603,N_14093,N_10731);
nor UO_1604 (O_1604,N_14148,N_14364);
nand UO_1605 (O_1605,N_11143,N_10386);
nand UO_1606 (O_1606,N_13515,N_13206);
or UO_1607 (O_1607,N_14761,N_11249);
and UO_1608 (O_1608,N_13471,N_13621);
or UO_1609 (O_1609,N_12104,N_11719);
and UO_1610 (O_1610,N_13880,N_11318);
nand UO_1611 (O_1611,N_12411,N_10166);
or UO_1612 (O_1612,N_11656,N_11198);
and UO_1613 (O_1613,N_10250,N_10534);
nor UO_1614 (O_1614,N_12191,N_13369);
and UO_1615 (O_1615,N_13332,N_11206);
nand UO_1616 (O_1616,N_10477,N_10136);
xnor UO_1617 (O_1617,N_11151,N_11110);
and UO_1618 (O_1618,N_11677,N_12700);
and UO_1619 (O_1619,N_12356,N_12933);
nor UO_1620 (O_1620,N_13882,N_11283);
and UO_1621 (O_1621,N_13350,N_12748);
xor UO_1622 (O_1622,N_14972,N_10717);
and UO_1623 (O_1623,N_11501,N_13255);
or UO_1624 (O_1624,N_11452,N_14461);
nor UO_1625 (O_1625,N_13017,N_14240);
xnor UO_1626 (O_1626,N_11509,N_13064);
and UO_1627 (O_1627,N_12348,N_12581);
xnor UO_1628 (O_1628,N_13523,N_12899);
nor UO_1629 (O_1629,N_13675,N_10266);
nand UO_1630 (O_1630,N_13529,N_14194);
nand UO_1631 (O_1631,N_10193,N_10931);
and UO_1632 (O_1632,N_12570,N_11087);
nor UO_1633 (O_1633,N_13074,N_10532);
and UO_1634 (O_1634,N_14721,N_11204);
or UO_1635 (O_1635,N_12723,N_14449);
and UO_1636 (O_1636,N_10388,N_11102);
xor UO_1637 (O_1637,N_13996,N_10882);
or UO_1638 (O_1638,N_10216,N_14197);
nand UO_1639 (O_1639,N_10889,N_14252);
and UO_1640 (O_1640,N_13852,N_13058);
or UO_1641 (O_1641,N_12980,N_14083);
xor UO_1642 (O_1642,N_13119,N_10936);
nand UO_1643 (O_1643,N_12195,N_12901);
xnor UO_1644 (O_1644,N_11063,N_11651);
nor UO_1645 (O_1645,N_12689,N_13303);
nand UO_1646 (O_1646,N_13652,N_11175);
nand UO_1647 (O_1647,N_10978,N_10549);
xnor UO_1648 (O_1648,N_14047,N_13245);
or UO_1649 (O_1649,N_14347,N_11036);
and UO_1650 (O_1650,N_13475,N_14656);
nand UO_1651 (O_1651,N_10017,N_11391);
or UO_1652 (O_1652,N_14888,N_12517);
or UO_1653 (O_1653,N_11236,N_14909);
xor UO_1654 (O_1654,N_13786,N_10047);
xor UO_1655 (O_1655,N_14156,N_12642);
nor UO_1656 (O_1656,N_10294,N_14463);
or UO_1657 (O_1657,N_11523,N_11425);
nand UO_1658 (O_1658,N_12145,N_10685);
or UO_1659 (O_1659,N_13396,N_12428);
nor UO_1660 (O_1660,N_11489,N_11137);
or UO_1661 (O_1661,N_13758,N_13557);
and UO_1662 (O_1662,N_10538,N_12961);
and UO_1663 (O_1663,N_13191,N_12829);
and UO_1664 (O_1664,N_10435,N_13426);
or UO_1665 (O_1665,N_12353,N_14962);
and UO_1666 (O_1666,N_13165,N_11505);
nor UO_1667 (O_1667,N_10811,N_12601);
and UO_1668 (O_1668,N_10570,N_13795);
and UO_1669 (O_1669,N_14577,N_12047);
or UO_1670 (O_1670,N_10663,N_11812);
or UO_1671 (O_1671,N_14486,N_12969);
xnor UO_1672 (O_1672,N_14073,N_10631);
nand UO_1673 (O_1673,N_14277,N_14137);
nor UO_1674 (O_1674,N_14728,N_10696);
nor UO_1675 (O_1675,N_14874,N_11153);
or UO_1676 (O_1676,N_12817,N_13726);
and UO_1677 (O_1677,N_14068,N_12998);
or UO_1678 (O_1678,N_10578,N_11853);
nand UO_1679 (O_1679,N_14708,N_14891);
xor UO_1680 (O_1680,N_13636,N_11992);
xnor UO_1681 (O_1681,N_14602,N_13851);
xnor UO_1682 (O_1682,N_12794,N_10141);
xnor UO_1683 (O_1683,N_13908,N_14260);
or UO_1684 (O_1684,N_11778,N_13086);
nor UO_1685 (O_1685,N_13663,N_11314);
xnor UO_1686 (O_1686,N_11454,N_14763);
nor UO_1687 (O_1687,N_10787,N_10798);
and UO_1688 (O_1688,N_13267,N_12911);
xnor UO_1689 (O_1689,N_10984,N_11192);
or UO_1690 (O_1690,N_13080,N_10900);
or UO_1691 (O_1691,N_14098,N_10210);
xnor UO_1692 (O_1692,N_11124,N_13752);
and UO_1693 (O_1693,N_11852,N_14470);
and UO_1694 (O_1694,N_11863,N_12545);
nor UO_1695 (O_1695,N_11552,N_12416);
or UO_1696 (O_1696,N_13633,N_11542);
nor UO_1697 (O_1697,N_10387,N_11392);
nor UO_1698 (O_1698,N_12500,N_10275);
xor UO_1699 (O_1699,N_14341,N_13510);
and UO_1700 (O_1700,N_10146,N_14981);
and UO_1701 (O_1701,N_10699,N_10451);
xnor UO_1702 (O_1702,N_13762,N_13501);
xnor UO_1703 (O_1703,N_12789,N_12721);
xor UO_1704 (O_1704,N_14543,N_10702);
or UO_1705 (O_1705,N_11359,N_12152);
nand UO_1706 (O_1706,N_11344,N_12114);
or UO_1707 (O_1707,N_12222,N_13744);
xnor UO_1708 (O_1708,N_13305,N_10626);
or UO_1709 (O_1709,N_12324,N_14088);
and UO_1710 (O_1710,N_13811,N_14591);
nand UO_1711 (O_1711,N_10710,N_11481);
or UO_1712 (O_1712,N_14234,N_13776);
nand UO_1713 (O_1713,N_14642,N_13552);
and UO_1714 (O_1714,N_14307,N_10602);
xnor UO_1715 (O_1715,N_14771,N_10053);
xor UO_1716 (O_1716,N_12479,N_14894);
and UO_1717 (O_1717,N_10430,N_13130);
or UO_1718 (O_1718,N_13547,N_10507);
nor UO_1719 (O_1719,N_13821,N_11533);
nor UO_1720 (O_1720,N_12462,N_12343);
nand UO_1721 (O_1721,N_10061,N_11818);
or UO_1722 (O_1722,N_14054,N_11911);
or UO_1723 (O_1723,N_13189,N_13327);
or UO_1724 (O_1724,N_13201,N_11158);
xor UO_1725 (O_1725,N_13212,N_14066);
nor UO_1726 (O_1726,N_13142,N_11865);
nor UO_1727 (O_1727,N_14880,N_12458);
and UO_1728 (O_1728,N_14722,N_13031);
nor UO_1729 (O_1729,N_11306,N_10130);
nand UO_1730 (O_1730,N_13532,N_14867);
nand UO_1731 (O_1731,N_11125,N_12892);
nor UO_1732 (O_1732,N_14314,N_10867);
nand UO_1733 (O_1733,N_12578,N_12431);
or UO_1734 (O_1734,N_14001,N_11316);
nor UO_1735 (O_1735,N_14109,N_13775);
xnor UO_1736 (O_1736,N_12624,N_12703);
or UO_1737 (O_1737,N_11024,N_14971);
or UO_1738 (O_1738,N_13923,N_10478);
or UO_1739 (O_1739,N_12710,N_13947);
and UO_1740 (O_1740,N_12008,N_10107);
nand UO_1741 (O_1741,N_14717,N_12337);
nand UO_1742 (O_1742,N_10084,N_14946);
xnor UO_1743 (O_1743,N_10915,N_12211);
xnor UO_1744 (O_1744,N_10869,N_13156);
and UO_1745 (O_1745,N_14336,N_13210);
or UO_1746 (O_1746,N_12740,N_10078);
xor UO_1747 (O_1747,N_12510,N_12823);
or UO_1748 (O_1748,N_12070,N_11447);
or UO_1749 (O_1749,N_11565,N_13478);
nand UO_1750 (O_1750,N_13197,N_11450);
nand UO_1751 (O_1751,N_14694,N_13460);
and UO_1752 (O_1752,N_12966,N_10399);
nor UO_1753 (O_1753,N_14207,N_12153);
and UO_1754 (O_1754,N_14974,N_14553);
or UO_1755 (O_1755,N_13620,N_14437);
nor UO_1756 (O_1756,N_10632,N_10812);
nor UO_1757 (O_1757,N_14863,N_11626);
nand UO_1758 (O_1758,N_11028,N_11591);
nor UO_1759 (O_1759,N_14921,N_12554);
nand UO_1760 (O_1760,N_11551,N_11417);
nor UO_1761 (O_1761,N_13488,N_10027);
nor UO_1762 (O_1762,N_13862,N_13178);
or UO_1763 (O_1763,N_10033,N_10841);
nor UO_1764 (O_1764,N_13814,N_12595);
or UO_1765 (O_1765,N_10301,N_13097);
nor UO_1766 (O_1766,N_14569,N_11007);
xor UO_1767 (O_1767,N_11885,N_14769);
and UO_1768 (O_1768,N_12727,N_14964);
xnor UO_1769 (O_1769,N_10568,N_14495);
nor UO_1770 (O_1770,N_10745,N_12449);
nor UO_1771 (O_1771,N_12164,N_12201);
nor UO_1772 (O_1772,N_11129,N_12859);
or UO_1773 (O_1773,N_12495,N_13270);
nand UO_1774 (O_1774,N_12177,N_12544);
nor UO_1775 (O_1775,N_14635,N_10700);
xnor UO_1776 (O_1776,N_13901,N_11781);
or UO_1777 (O_1777,N_13702,N_11385);
xor UO_1778 (O_1778,N_14182,N_13190);
and UO_1779 (O_1779,N_12457,N_14142);
or UO_1780 (O_1780,N_14392,N_14266);
nor UO_1781 (O_1781,N_12942,N_10471);
nand UO_1782 (O_1782,N_12918,N_11582);
xnor UO_1783 (O_1783,N_12170,N_10562);
or UO_1784 (O_1784,N_14469,N_10236);
xor UO_1785 (O_1785,N_11037,N_10974);
nor UO_1786 (O_1786,N_13289,N_13220);
or UO_1787 (O_1787,N_13754,N_11662);
xnor UO_1788 (O_1788,N_14500,N_14070);
xnor UO_1789 (O_1789,N_10075,N_12357);
nand UO_1790 (O_1790,N_13697,N_11339);
and UO_1791 (O_1791,N_10278,N_11399);
and UO_1792 (O_1792,N_14229,N_11256);
xnor UO_1793 (O_1793,N_14961,N_10715);
or UO_1794 (O_1794,N_14013,N_14303);
nand UO_1795 (O_1795,N_11839,N_12706);
or UO_1796 (O_1796,N_13137,N_11512);
xor UO_1797 (O_1797,N_12300,N_11305);
nor UO_1798 (O_1798,N_14966,N_11870);
or UO_1799 (O_1799,N_14459,N_14502);
nor UO_1800 (O_1800,N_10504,N_12074);
xnor UO_1801 (O_1801,N_14641,N_10306);
and UO_1802 (O_1802,N_14542,N_11620);
nor UO_1803 (O_1803,N_10709,N_12241);
and UO_1804 (O_1804,N_14356,N_14348);
or UO_1805 (O_1805,N_12277,N_13388);
nand UO_1806 (O_1806,N_13236,N_11779);
and UO_1807 (O_1807,N_10962,N_12467);
and UO_1808 (O_1808,N_10854,N_10269);
or UO_1809 (O_1809,N_14959,N_13043);
nand UO_1810 (O_1810,N_12244,N_13888);
xor UO_1811 (O_1811,N_10162,N_11321);
xor UO_1812 (O_1812,N_14398,N_12497);
nand UO_1813 (O_1813,N_12466,N_11401);
nand UO_1814 (O_1814,N_14174,N_14949);
or UO_1815 (O_1815,N_14305,N_10144);
and UO_1816 (O_1816,N_12259,N_11281);
or UO_1817 (O_1817,N_14453,N_14979);
and UO_1818 (O_1818,N_14664,N_12736);
nor UO_1819 (O_1819,N_13283,N_10408);
nor UO_1820 (O_1820,N_11482,N_10343);
nand UO_1821 (O_1821,N_12766,N_10320);
nor UO_1822 (O_1822,N_10004,N_10293);
xnor UO_1823 (O_1823,N_12126,N_12228);
nand UO_1824 (O_1824,N_11219,N_11324);
nand UO_1825 (O_1825,N_10937,N_10541);
nor UO_1826 (O_1826,N_11075,N_12543);
and UO_1827 (O_1827,N_12278,N_10500);
and UO_1828 (O_1828,N_13839,N_13730);
and UO_1829 (O_1829,N_13257,N_11732);
or UO_1830 (O_1830,N_11015,N_14404);
xor UO_1831 (O_1831,N_10809,N_12763);
nand UO_1832 (O_1832,N_11085,N_12954);
and UO_1833 (O_1833,N_14755,N_10185);
nand UO_1834 (O_1834,N_11940,N_11922);
nor UO_1835 (O_1835,N_14271,N_14774);
nor UO_1836 (O_1836,N_11601,N_11987);
nand UO_1837 (O_1837,N_10270,N_10011);
nor UO_1838 (O_1838,N_10013,N_14320);
nand UO_1839 (O_1839,N_14298,N_10868);
or UO_1840 (O_1840,N_10943,N_13647);
nor UO_1841 (O_1841,N_13576,N_10845);
nor UO_1842 (O_1842,N_10307,N_12081);
xor UO_1843 (O_1843,N_12575,N_10667);
or UO_1844 (O_1844,N_12990,N_11772);
or UO_1845 (O_1845,N_13433,N_14746);
xor UO_1846 (O_1846,N_14865,N_10903);
or UO_1847 (O_1847,N_12194,N_13279);
nor UO_1848 (O_1848,N_11907,N_13419);
xor UO_1849 (O_1849,N_14691,N_13108);
nand UO_1850 (O_1850,N_13699,N_12098);
nand UO_1851 (O_1851,N_13243,N_11749);
and UO_1852 (O_1852,N_11332,N_13793);
and UO_1853 (O_1853,N_14125,N_11753);
nand UO_1854 (O_1854,N_10506,N_13454);
nand UO_1855 (O_1855,N_12385,N_12151);
and UO_1856 (O_1856,N_13981,N_12421);
nor UO_1857 (O_1857,N_11933,N_12885);
or UO_1858 (O_1858,N_11017,N_13244);
nand UO_1859 (O_1859,N_12617,N_10814);
or UO_1860 (O_1860,N_10866,N_11369);
nor UO_1861 (O_1861,N_12478,N_14214);
and UO_1862 (O_1862,N_13314,N_12239);
nand UO_1863 (O_1863,N_10095,N_14135);
or UO_1864 (O_1864,N_11004,N_14785);
nand UO_1865 (O_1865,N_10990,N_10221);
nor UO_1866 (O_1866,N_11616,N_14804);
nor UO_1867 (O_1867,N_11136,N_11221);
nor UO_1868 (O_1868,N_10895,N_13922);
nand UO_1869 (O_1869,N_11268,N_10672);
nand UO_1870 (O_1870,N_14279,N_12802);
nand UO_1871 (O_1871,N_10493,N_10757);
xor UO_1872 (O_1872,N_10871,N_12566);
nor UO_1873 (O_1873,N_11126,N_12840);
or UO_1874 (O_1874,N_10973,N_12655);
or UO_1875 (O_1875,N_10564,N_13481);
nor UO_1876 (O_1876,N_14567,N_11952);
xor UO_1877 (O_1877,N_13076,N_14286);
xnor UO_1878 (O_1878,N_13264,N_14564);
nor UO_1879 (O_1879,N_10048,N_13172);
nor UO_1880 (O_1880,N_13641,N_10625);
xor UO_1881 (O_1881,N_12095,N_12471);
or UO_1882 (O_1882,N_11989,N_11174);
and UO_1883 (O_1883,N_13990,N_11882);
or UO_1884 (O_1884,N_14473,N_13717);
nand UO_1885 (O_1885,N_11734,N_10946);
or UO_1886 (O_1886,N_11046,N_14175);
xnor UO_1887 (O_1887,N_12373,N_10744);
xnor UO_1888 (O_1888,N_14454,N_11636);
or UO_1889 (O_1889,N_10369,N_12986);
xnor UO_1890 (O_1890,N_11056,N_14605);
xor UO_1891 (O_1891,N_13298,N_13463);
and UO_1892 (O_1892,N_12628,N_11196);
nor UO_1893 (O_1893,N_13700,N_12015);
or UO_1894 (O_1894,N_12804,N_10634);
and UO_1895 (O_1895,N_13161,N_14766);
nand UO_1896 (O_1896,N_13217,N_10172);
and UO_1897 (O_1897,N_13526,N_11947);
nor UO_1898 (O_1898,N_14669,N_11916);
xnor UO_1899 (O_1899,N_12837,N_11430);
nand UO_1900 (O_1900,N_11098,N_10032);
and UO_1901 (O_1901,N_14617,N_14489);
and UO_1902 (O_1902,N_11057,N_10552);
or UO_1903 (O_1903,N_12796,N_13400);
and UO_1904 (O_1904,N_12117,N_11303);
and UO_1905 (O_1905,N_12738,N_12939);
and UO_1906 (O_1906,N_14169,N_13215);
nand UO_1907 (O_1907,N_14663,N_13815);
and UO_1908 (O_1908,N_14222,N_11346);
xnor UO_1909 (O_1909,N_13952,N_14166);
xnor UO_1910 (O_1910,N_10120,N_12352);
xor UO_1911 (O_1911,N_14851,N_14770);
or UO_1912 (O_1912,N_14065,N_13325);
nand UO_1913 (O_1913,N_10132,N_11176);
xor UO_1914 (O_1914,N_11055,N_12801);
and UO_1915 (O_1915,N_13251,N_10108);
nor UO_1916 (O_1916,N_13600,N_14441);
xnor UO_1917 (O_1917,N_12746,N_10473);
and UO_1918 (O_1918,N_10537,N_12744);
or UO_1919 (O_1919,N_14850,N_10904);
nand UO_1920 (O_1920,N_10291,N_14431);
xnor UO_1921 (O_1921,N_12233,N_13692);
xnor UO_1922 (O_1922,N_11408,N_14844);
xnor UO_1923 (O_1923,N_13989,N_13925);
and UO_1924 (O_1924,N_11289,N_11887);
and UO_1925 (O_1925,N_14419,N_14968);
xor UO_1926 (O_1926,N_12328,N_10561);
or UO_1927 (O_1927,N_14902,N_13144);
and UO_1928 (O_1928,N_12530,N_13604);
nand UO_1929 (O_1929,N_10701,N_14821);
nand UO_1930 (O_1930,N_14436,N_12066);
nor UO_1931 (O_1931,N_11860,N_12754);
nand UO_1932 (O_1932,N_10706,N_10649);
or UO_1933 (O_1933,N_12150,N_12213);
xnor UO_1934 (O_1934,N_14167,N_10295);
and UO_1935 (O_1935,N_12730,N_10623);
xor UO_1936 (O_1936,N_10865,N_10456);
nand UO_1937 (O_1937,N_12406,N_12072);
xor UO_1938 (O_1938,N_13326,N_11338);
and UO_1939 (O_1939,N_12436,N_13362);
or UO_1940 (O_1940,N_10006,N_11953);
and UO_1941 (O_1941,N_11378,N_14679);
and UO_1942 (O_1942,N_14759,N_14087);
or UO_1943 (O_1943,N_13045,N_10501);
and UO_1944 (O_1944,N_10348,N_14668);
and UO_1945 (O_1945,N_12877,N_13328);
or UO_1946 (O_1946,N_13810,N_12627);
and UO_1947 (O_1947,N_13615,N_11187);
or UO_1948 (O_1948,N_11902,N_12475);
nand UO_1949 (O_1949,N_12810,N_11237);
or UO_1950 (O_1950,N_10005,N_10586);
nand UO_1951 (O_1951,N_11908,N_10373);
and UO_1952 (O_1952,N_14846,N_14839);
nor UO_1953 (O_1953,N_14936,N_11823);
xor UO_1954 (O_1954,N_12932,N_13802);
xor UO_1955 (O_1955,N_10644,N_12370);
xor UO_1956 (O_1956,N_12743,N_10288);
nor UO_1957 (O_1957,N_13361,N_12701);
nand UO_1958 (O_1958,N_11038,N_13574);
and UO_1959 (O_1959,N_11380,N_10682);
and UO_1960 (O_1960,N_13382,N_11010);
or UO_1961 (O_1961,N_10513,N_12041);
xor UO_1962 (O_1962,N_10846,N_13686);
and UO_1963 (O_1963,N_14438,N_12113);
and UO_1964 (O_1964,N_12582,N_10756);
nor UO_1965 (O_1965,N_13367,N_13149);
nand UO_1966 (O_1966,N_14885,N_13052);
xnor UO_1967 (O_1967,N_10245,N_12404);
nor UO_1968 (O_1968,N_14554,N_12252);
or UO_1969 (O_1969,N_13177,N_14950);
and UO_1970 (O_1970,N_13924,N_14757);
nor UO_1971 (O_1971,N_11817,N_11658);
nand UO_1972 (O_1972,N_10008,N_13457);
or UO_1973 (O_1973,N_12518,N_13472);
nand UO_1974 (O_1974,N_10675,N_13109);
nor UO_1975 (O_1975,N_10792,N_13393);
and UO_1976 (O_1976,N_14895,N_12506);
or UO_1977 (O_1977,N_11672,N_14244);
nand UO_1978 (O_1978,N_12600,N_13817);
or UO_1979 (O_1979,N_11831,N_10583);
and UO_1980 (O_1980,N_14535,N_13136);
or UO_1981 (O_1981,N_14892,N_13556);
or UO_1982 (O_1982,N_10609,N_10395);
or UO_1983 (O_1983,N_12040,N_12674);
and UO_1984 (O_1984,N_10508,N_12085);
nand UO_1985 (O_1985,N_11384,N_14330);
xnor UO_1986 (O_1986,N_10044,N_14991);
or UO_1987 (O_1987,N_13442,N_12128);
nor UO_1988 (O_1988,N_10769,N_13363);
xnor UO_1989 (O_1989,N_13117,N_10060);
or UO_1990 (O_1990,N_13296,N_10612);
xor UO_1991 (O_1991,N_14288,N_11222);
nor UO_1992 (O_1992,N_14039,N_14848);
and UO_1993 (O_1993,N_14749,N_11211);
xnor UO_1994 (O_1994,N_12590,N_13366);
or UO_1995 (O_1995,N_12165,N_11804);
or UO_1996 (O_1996,N_11600,N_10545);
nand UO_1997 (O_1997,N_10425,N_11578);
nand UO_1998 (O_1998,N_10276,N_11795);
nor UO_1999 (O_1999,N_10065,N_12237);
endmodule